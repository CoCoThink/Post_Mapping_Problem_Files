module usb_phy_fast (
DataOut_i_0_,
DataOut_i_1_,
DataOut_i_2_,
DataOut_i_3_,
DataOut_i_4_,
DataOut_i_5_,
DataOut_i_6_,
DataOut_i_7_,
TxValid_i,
ispd_clk,
phy_tx_mode,
rst,
rxd,
rxdn,
rxdp,
DataIn_o_0_,
DataIn_o_1_,
DataIn_o_2_,
DataIn_o_3_,
DataIn_o_4_,
DataIn_o_5_,
DataIn_o_6_,
DataIn_o_7_,
LineState_o_0_,
LineState_o_1_,
RxActive_o,
RxError_o,
RxValid_o,
TxReady_o,
g1897_u0_o,
txdn,
txdp,
txoe,
usb_rst
);

// Start PIs
input DataOut_i_0_;
input DataOut_i_1_;
input DataOut_i_2_;
input DataOut_i_3_;
input DataOut_i_4_;
input DataOut_i_5_;
input DataOut_i_6_;
input DataOut_i_7_;
input TxValid_i;
input ispd_clk;
input phy_tx_mode;
input rst;
input rxd;
input rxdn;
input rxdp;

// Start POs
output DataIn_o_0_;
output DataIn_o_1_;
output DataIn_o_2_;
output DataIn_o_3_;
output DataIn_o_4_;
output DataIn_o_5_;
output DataIn_o_6_;
output DataIn_o_7_;
output LineState_o_0_;
output LineState_o_1_;
output RxActive_o;
output RxError_o;
output RxValid_o;
output TxReady_o;
output g1897_u0_o;
output txdn;
output txdp;
output txoe;
output usb_rst;

// Start wires
wire DataOut_i_0_;
wire DataOut_i_1_;
wire DataOut_i_2_;
wire DataOut_i_3_;
wire DataOut_i_4_;
wire DataOut_i_5_;
wire DataOut_i_6_;
wire DataOut_i_7_;
wire TxValid_i;
wire ispd_clk;
wire phy_tx_mode;
wire rst;
wire rxd;
wire rxdn;
wire rxdp;
wire DataIn_o_0_;
wire DataIn_o_1_;
wire DataIn_o_2_;
wire DataIn_o_3_;
wire DataIn_o_4_;
wire DataIn_o_5_;
wire DataIn_o_6_;
wire DataIn_o_7_;
wire LineState_o_0_;
wire LineState_o_1_;
wire RxActive_o;
wire RxError_o;
wire RxValid_o;
wire TxReady_o;
wire g1897_u0_o;
wire txdn;
wire txdp;
wire txoe;
wire usb_rst;
wire FE_RN_0_0;
wire FE_RN_1_0;
wire FE_RN_2_0;
wire g11_p;
wire g15_p;
wire g1737_p;
wire g1738_p;
wire g1739_p;
wire g1740_p;
wire g1741_p;
wire g1742_p;
wire g1743_p;
wire g1757_p;
wire TIMEBOOST_net_114;
wire g1776_db;
wire g1776_sb;
wire g1777_da;
wire g1777_db;
wire g1777_sb;
wire TIMEBOOST_net_49;
wire g1778_db;
wire g1778_sb;
wire TIMEBOOST_net_50;
wire g1779_db;
wire g1779_sb;
wire TIMEBOOST_net_69;
wire g1780_db;
wire g1780_sb;
wire TIMEBOOST_net_52;
wire g1781_db;
wire g1781_sb;
wire TIMEBOOST_net_53;
wire g1782_db;
wire g1782_sb;
wire g1855_da;
wire g1855_db;
wire g1855_sb;
wire g1857_p;
wire g1881_p;
wire g1884_p;
wire g1901_p;
wire g1923_p;
wire g1942_p;
wire g1965_p;
wire g1975_p;
wire g1980_p;
wire g2028_p;
wire g2035_p;
wire g2050_p;
wire g2057_p;
wire TIMEBOOST_net_59;
wire TIMEBOOST_net_157;
wire g2063_sb;
wire g2066_p;
wire g2067_p;
wire g2068_p;
wire g2069_p;
wire g2091_p;
wire g2103_p;
wire g2108_p;
wire g2113_p;
wire g2116_p;
wire g2128_p;
wire g2130_p;
wire g2141_p;
wire g2385_p;
wire g2412_p;
wire g2413_p;
wire g2494_p;
wire g2506_p;
wire g2651_p;
wire g2674_p;
wire g41_p;
wire i_rx_phy_bit_cnt_0_;
wire i_rx_phy_bit_cnt_2_;
wire i_rx_phy_bit_stuff_err;
wire i_rx_phy_bit_stuff_err_reg_Q;
wire i_rx_phy_byte_err;
wire i_rx_phy_byte_err_reg_Q;
wire i_rx_phy_dpll_state_0_;
wire i_rx_phy_dpll_state_1_;
wire i_rx_phy_fs_ce_r1;
wire i_rx_phy_fs_ce_r2;
wire i_rx_phy_fs_state_0_;
wire i_rx_phy_fs_state_2_;
wire i_rx_phy_one_cnt_0_;
wire i_rx_phy_one_cnt_1_;
wire i_rx_phy_one_cnt_2_;
wire i_rx_phy_rx_en;
wire i_rx_phy_rx_valid1;
wire i_rx_phy_rx_valid_r;
wire i_rx_phy_rxd_r;
wire i_rx_phy_rxd_s;
wire i_rx_phy_rxd_s0;
wire i_rx_phy_rxd_s1;
wire i_rx_phy_rxd_s1_reg_Q;
wire i_rx_phy_rxdn_s;
wire i_rx_phy_rxdn_s0;
wire i_rx_phy_rxdn_s_r;
wire i_rx_phy_rxdn_s_r_reg_Q;
wire i_rx_phy_rxdp_s;
wire i_rx_phy_rxdp_s0;
wire i_rx_phy_rxdp_s_r;
wire i_rx_phy_rxdp_s_r_reg_Q;
wire i_rx_phy_sd_nrzi;
wire i_rx_phy_sd_r;
wire i_rx_phy_se0_r;
wire i_rx_phy_se0_r_reg_Q;
wire i_rx_phy_se0_s;
wire i_rx_phy_shift_en;
wire i_rx_phy_sync_err;
wire i_rx_phy_sync_err_reg_Q;
wire i_tx_phy_append_eop;
wire i_tx_phy_append_eop_sync1;
wire i_tx_phy_append_eop_sync2;
wire i_tx_phy_append_eop_sync4;
wire i_tx_phy_bit_cnt_0_;
wire i_tx_phy_bit_cnt_1_;
wire i_tx_phy_bit_cnt_2_;
wire i_tx_phy_data_done;
wire i_tx_phy_hold_reg;
wire i_tx_phy_hold_reg_10;
wire i_tx_phy_hold_reg_4;
wire i_tx_phy_hold_reg_5;
wire i_tx_phy_hold_reg_6;
wire i_tx_phy_hold_reg_7;
wire i_tx_phy_hold_reg_8;
wire i_tx_phy_hold_reg_9;
wire i_tx_phy_hold_reg_d;
wire i_tx_phy_hold_reg_d_11;
wire i_tx_phy_hold_reg_d_12;
wire i_tx_phy_hold_reg_d_13;
wire i_tx_phy_hold_reg_d_14;
wire i_tx_phy_hold_reg_d_15;
wire i_tx_phy_hold_reg_d_17;
wire i_tx_phy_hold_reg_d_reg_1__Q;
wire i_tx_phy_hold_reg_d_reg_3__Q;
wire i_tx_phy_hold_reg_d_reg_5__Q;
wire i_tx_phy_hold_reg_d_reg_6__Q;
wire i_tx_phy_ld_data;
wire i_tx_phy_ld_data_reg_Q;
wire i_tx_phy_one_cnt_0_;
wire i_tx_phy_one_cnt_1_;
wire i_tx_phy_one_cnt_2_;
wire i_tx_phy_sd_bs_o;
wire i_tx_phy_sd_nrzi_o;
wire i_tx_phy_sd_raw_o;
wire i_tx_phy_sft_done;
wire i_tx_phy_sft_done_r;
wire i_tx_phy_state_1_;
wire i_tx_phy_state_2_;
wire i_tx_phy_tx_ip;
wire i_tx_phy_txoe_r1;
wire i_tx_phy_txoe_r2;
wire n_10;
wire n_100;
wire n_103;
wire n_105;
wire n_106;
wire n_108;
wire n_11;
wire n_111;
wire n_112;
wire n_115;
wire n_116;
wire n_118;
wire n_12;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_138;
wire n_139;
wire n_141;
wire n_142;
wire n_15;
wire n_150;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_157;
wire n_161;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_172;
wire n_175;
wire n_176;
wire n_18;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_191;
wire n_192;
wire n_193;
wire n_195;
wire n_197;
wire n_198;
wire n_201;
wire n_203;
wire n_204;
wire n_209;
wire n_21;
wire n_210;
wire n_213;
wire n_217;
wire n_22;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_235;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_248;
wire n_251;
wire n_252;
wire n_254;
wire n_255;
wire n_256;
wire TIMEBOOST_net_0;
wire n_258;
wire n_259;
wire n_263;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_27;
wire TIMEBOOST_net_44;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_28;
wire n_280;
wire n_283;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_296;
wire TIMEBOOST_net_43;
wire n_299;
wire n_300;
wire n_301;
wire TIMEBOOST_net_109;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_33;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_347;
wire n_35;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_359;
wire TIMEBOOST_net_154;
wire n_361;
wire n_362;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_37;
wire n_370;
wire n_373;
wire n_375;
wire n_377;
wire n_378;
wire n_380;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_394;
wire n_395;
wire n_400;
wire n_401;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_409;
wire TIMEBOOST_net_94;
wire n_411;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_420;
wire n_421;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_439;
wire n_440;
wire n_443;
wire n_444;
wire n_446;
wire n_447;
wire n_449;
wire n_450;
wire TIMEBOOST_net_151;
wire TIMEBOOST_net_144;
wire TIMEBOOST_net_117;
wire TIMEBOOST_net_141;
wire TIMEBOOST_net_159;
wire TIMEBOOST_net_98;
wire TIMEBOOST_net_108;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_471;
wire n_472;
wire n_479;
wire n_48;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_489;
wire n_49;
wire n_490;
wire TIMEBOOST_net_3;
wire n_493;
wire n_499;
wire n_50;
wire n_505;
wire n_506;
wire n_507;
wire n_509;
wire n_51;
wire n_511;
wire n_52;
wire n_523;
wire n_529;
wire n_53;
wire n_538;
wire n_539;
wire n_54;
wire n_540;
wire n_55;
wire n_559;
wire n_56;
wire n_567;
wire n_57;
wire n_573;
wire TIMEBOOST_net_46;
wire n_58;
wire n_583;
wire n_588;
wire n_590;
wire n_593;
wire n_598;
wire n_60;
wire n_604;
wire n_61;
wire n_628;
wire n_629;
wire n_63;
wire n_631;
wire n_632;
wire n_64;
wire n_66;
wire n_660;
wire n_661;
wire n_665;
wire n_666;
wire n_69;
wire n_697;
wire n_699;
wire n_7;
wire n_70;
wire n_700;
wire TIMEBOOST_net_158;
wire n_703;
wire n_704;
wire n_706;
wire TIMEBOOST_net_4;
wire TIMEBOOST_net_96;
wire n_709;
wire n_71;
wire TIMEBOOST_net_5;
wire n_722;
wire n_726;
wire n_727;
wire n_734;
wire n_735;
wire n_737;
wire n_74;
wire n_741;
wire n_742;
wire n_743;
wire TIMEBOOST_net_80;
wire n_749;
wire n_752;
wire n_753;
wire n_754;
wire n_755;
wire n_756;
wire n_758;
wire n_759;
wire n_763;
wire n_764;
wire n_767;
wire n_77;
wire n_782;
wire n_783;
wire n_785;
wire n_786;
wire n_788;
wire n_794;
wire n_796;
wire n_8;
wire n_800;
wire n_804;
wire n_81;
wire n_840;
wire n_841;
wire n_85;
wire n_852;
wire n_864;
wire n_873;
wire n_878;
wire n_88;
wire n_882;
wire n_884;
wire n_885;
wire n_888;
wire n_894;
wire n_9;
wire n_90;
wire n_91;
wire n_910;
wire n_911;
wire n_913;
wire n_914;
wire n_915;
wire n_916;
wire n_919;
wire n_920;
wire n_921;
wire n_922;
wire n_923;
wire n_924;
wire n_925;
wire n_926;
wire n_927;
wire n_928;
wire n_929;
wire n_930;
wire n_932;
wire n_933;
wire n_934;
wire n_935;
wire n_937;
wire n_938;
wire n_940;
wire n_941;
wire n_942;
wire n_943;
wire n_944;
wire n_945;
wire n_947;
wire n_948;
wire n_949;
wire n_951;
wire n_952;
wire n_957;
wire n_958;
wire n_959;
wire n_960;
wire n_961;
wire n_962;
wire TIMEBOOST_net_142;
wire n_965;
wire n_966;
wire n_967;
wire n_968;
wire TIMEBOOST_net_111;
wire n_97;
wire n_970;
wire n_971;
wire n_972;
wire n_974;
wire n_976;
wire n_977;
wire n_980;
wire n_981;
wire n_982;
wire n_984;
wire n_988;
wire TIMEBOOST_net_143;
wire TIMEBOOST_net_160;
wire TIMEBOOST_net_70;
wire n_992;
wire rst_cnt_0_;
wire rst_cnt_1_;
wire rst_cnt_3_;
wire rst_cnt_4_;
wire TIMEBOOST_net_126;
wire TIMEBOOST_net_8;
wire TIMEBOOST_net_148;
wire TIMEBOOST_net_155;
wire TIMEBOOST_net_11;
wire TIMEBOOST_net_12;
wire TIMEBOOST_net_13;
wire TIMEBOOST_net_14;
wire TIMEBOOST_net_15;
wire TIMEBOOST_net_137;
wire TIMEBOOST_net_55;
wire TIMEBOOST_net_156;
wire TIMEBOOST_net_93;
wire TIMEBOOST_net_95;
wire TIMEBOOST_net_21;
wire TIMEBOOST_net_22;
wire TIMEBOOST_net_23;
wire TIMEBOOST_net_24;
wire TIMEBOOST_net_25;
wire TIMEBOOST_net_26;
wire TIMEBOOST_net_27;
wire TIMEBOOST_net_54;
wire TIMEBOOST_net_29;
wire TIMEBOOST_net_30;
wire TIMEBOOST_net_162;
wire TIMEBOOST_net_32;
wire TIMEBOOST_net_135;
wire TIMEBOOST_net_34;
wire TIMEBOOST_net_35;
wire TIMEBOOST_net_36;
wire TIMEBOOST_net_145;
wire TIMEBOOST_net_38;
wire TIMEBOOST_net_45;
wire TIMEBOOST_net_40;
wire TIMEBOOST_net_147;
wire TIMEBOOST_net_140;
wire TIMEBOOST_net_152;
wire TIMEBOOST_net_161;
wire TIMEBOOST_net_163;
wire TIMEBOOST_net_146;
wire TIMEBOOST_net_149;
wire TIMEBOOST_net_153;
wire TIMEBOOST_net_164;
wire TIMEBOOST_net_165;
wire TIMEBOOST_net_166;
wire TIMEBOOST_net_167;
wire TIMEBOOST_net_168;
wire TIMEBOOST_net_169;
wire TIMEBOOST_net_170;
wire TIMEBOOST_net_171;

// Start cells
na02f02 FE_RC_0_0 ( .a(n_629), .b(FE_RN_0_0), .o(n_632) );
no02s02 FE_RC_1_0 ( .a(FE_RN_2_0), .b(FE_RN_1_0), .o(FE_RN_0_0) );
in01s02 FE_RC_2_0 ( .a(n_631), .o(FE_RN_1_0) );
in01s01 FE_RC_3_0 ( .a(rst), .o(FE_RN_2_0) );
no02s04 g10_u0 ( .a(n_911), .b(n_913), .o(n_914) );
no02s02 g11_u0 ( .a(n_980), .b(n_947), .o(g11_p) );
in01s02 g11_u1 ( .a(g11_p), .o(n_911) );
in01s08 g12_u0 ( .a(i_rx_phy_rx_en), .o(n_540) );
in01s04 g13_u0 ( .a(n_794), .o(n_913) );
no02s02 g14_u0 ( .a(n_981), .b(n_788), .o(n_604) );
na02s02 g15_u0 ( .a(n_948), .b(n_796), .o(g15_p) );
in01s01 g15_u1 ( .a(g15_p), .o(n_949) );
na02s02 TIMEBOOST_cell_16 ( .a(TIMEBOOST_net_4), .b(n_952), .o(n_930) );
in01m02 g1653_u0 ( .a(n_632), .o(n_529) );
ao12s02 g1661_u0 ( .a(FE_RN_2_0), .b(n_506), .c(n_660), .o(n_523) );
no02s02 g1680_u0 ( .a(n_386), .b(n_416), .o(n_417) );
na02s02 g1681_u0 ( .a(n_493), .b(n_440), .o(n_511) );
ao12s02 g1695_u0 ( .a(FE_RN_2_0), .b(n_704), .c(n_935), .o(n_459) );
na02s02 g1696_u0 ( .a(n_938), .b(n_480), .o(n_481) );
na02s02 g1697_u0 ( .a(n_490), .b(n_786), .o(n_506) );
in01s01 g1702_u0 ( .a(n_404), .o(n_423) );
na02s01 g1703_u0 ( .a(n_380), .b(n_269), .o(n_404) );
no02s01 g1707_u0 ( .a(n_472), .b(n_444), .o(n_499) );
ao12s02 g1709_u0 ( .a(n_370), .b(n_384), .c(rst_cnt_3_), .o(n_386) );
na02s01 TIMEBOOST_cell_431 ( .a(TIMEBOOST_net_156), .b(n_443), .o(TIMEBOOST_net_151) );
na02s04 g1717_u0 ( .a(n_916), .b(n_74), .o(n_439) );
no02s02 g1718_u0 ( .a(n_942), .b(n_916), .o(n_783) );
na02s02 g1719_u0 ( .a(n_926), .b(n_982), .o(n_480) );
na02s10 TIMEBOOST_cell_7 ( .a(i_rx_phy_rx_en), .b(i_rx_phy_rxdn_s), .o(TIMEBOOST_net_0) );
no02s01 g1725_u0 ( .a(n_385), .b(n_416), .o(n_428) );
ao12s02 g1726_u0 ( .a(n_384), .b(n_292), .c(n_256), .o(n_370) );
na02s01 TIMEBOOST_cell_83 ( .a(n_426), .b(i_rx_phy_sd_nrzi), .o(TIMEBOOST_net_38) );
ao12s01 g1729_u0 ( .a(n_961), .b(n_359), .c(n_347), .o(n_414) );
in01s01 g1731_u0 ( .a(n_754), .o(n_490) );
in01s01 g1733_u0 ( .a(n_753), .o(n_461) );
in01s01 g1734_u0 ( .a(n_753), .o(n_460) );
ao12s02 g1736_u0 ( .a(n_27), .b(n_369), .c(n_337), .o(n_411) );
na02s01 TIMEBOOST_cell_422 ( .a(n_450), .b(n_974), .o(TIMEBOOST_net_152) );
in01s01 g1737_u1 ( .a(g1737_p), .o(n_489) );
na02s01 TIMEBOOST_cell_399 ( .a(g1781_db), .b(n_974), .o(TIMEBOOST_net_145) );
in01s01 g1738_u1 ( .a(g1738_p), .o(n_487) );
na02s01 TIMEBOOST_cell_434 ( .a(n_852), .b(i_rx_phy_sd_r), .o(TIMEBOOST_net_158) );
in01s01 g1739_u1 ( .a(g1739_p), .o(n_486) );
na02s02 TIMEBOOST_cell_244 ( .a(TIMEBOOST_net_93), .b(n_511), .o(n_992) );
in01s01 g1740_u1 ( .a(g1740_p), .o(n_485) );
na02s02 TIMEBOOST_cell_295 ( .a(TIMEBOOST_net_111), .b(n_700), .o(TIMEBOOST_net_26) );
in01s01 g1741_u1 ( .a(g1741_p), .o(n_484) );
na02s02 TIMEBOOST_cell_317 ( .a(n_929), .b(n_894), .o(TIMEBOOST_net_114) );
in01s01 g1742_u1 ( .a(g1742_p), .o(n_483) );
na02s01 TIMEBOOST_cell_404 ( .a(TIMEBOOST_net_147), .b(g1777_da), .o(g1738_p) );
in01s01 g1743_u1 ( .a(g1743_p), .o(n_482) );
oa12s01 g1744_u0 ( .a(i_rx_phy_se0_r), .b(n_353), .c(i_rx_phy_bit_cnt_2_), .o(n_472) );
oa12s02 g1745_u0 ( .a(n_252), .b(n_311), .c(n_384), .o(n_380) );
in01s01 g1746_u0 ( .a(n_479), .o(n_505) );
na02s01 TIMEBOOST_cell_181 ( .a(TIMEBOOST_net_38), .b(n_248), .o(TIMEBOOST_net_69) );
oa12s01 g1748_u0 ( .a(n_447), .b(n_9), .c(n_885), .o(n_471) );
na03s02 TIMEBOOST_cell_444 ( .a(n_966), .b(TIMEBOOST_net_117), .c(n_927), .o(TIMEBOOST_net_163) );
in01s02 g1757_u1 ( .a(g1757_p), .o(n_420) );
ao12s02 g1758_u0 ( .a(n_318), .b(n_538), .c(n_539), .o(n_432) );
na02s01 g1759_u0 ( .a(n_446), .b(g2674_p), .o(n_447) );
na02s01 g1760_u0 ( .a(RxActive_o), .b(n_446), .o(n_444) );
na02s01 g1762_u0 ( .a(i_rx_phy_rx_valid_r), .b(n_446), .o(n_443) );
ao12s02 g1763_u0 ( .a(n_400), .b(n_163), .c(n_342), .o(n_388) );
na02s02 TIMEBOOST_cell_426 ( .a(n_841), .b(TIMEBOOST_net_98), .o(TIMEBOOST_net_154) );
na02s02 TIMEBOOST_cell_342 ( .a(TIMEBOOST_net_126), .b(n_278), .o(n_361) );
ao12s02 g1775_u0 ( .a(n_368), .b(n_384), .c(n_306), .o(n_385) );
in01s01 g1776_u0 ( .a(i_tx_phy_ld_data), .o(g1776_sb) );
na02s02 TIMEBOOST_cell_424 ( .a(i_tx_phy_sd_raw_o), .b(n_296), .o(TIMEBOOST_net_153) );
na02s01 g1776_u2 ( .a(i_tx_phy_ld_data), .b(i_tx_phy_hold_reg), .o(g1776_db) );
na03s02 TIMEBOOST_cell_420 ( .a(TIMEBOOST_net_151), .b(n_461), .c(n_511), .o(n_709) );
in01s01 g1777_u0 ( .a(i_tx_phy_ld_data), .o(g1777_sb) );
na02s01 g1777_u1 ( .a(DataOut_i_1_), .b(g1777_sb), .o(g1777_da) );
na02s01 g1777_u2 ( .a(i_tx_phy_ld_data), .b(i_tx_phy_hold_reg_4), .o(g1777_db) );
na02s01 TIMEBOOST_cell_124 ( .a(g1779_sb), .b(DataOut_i_3_), .o(TIMEBOOST_net_50) );
in01s01 g1778_u0 ( .a(i_tx_phy_ld_data), .o(g1778_sb) );
na02s01 TIMEBOOST_cell_437 ( .a(TIMEBOOST_net_159), .b(TIMEBOOST_net_109), .o(n_392) );
na02s01 g1778_u2 ( .a(i_tx_phy_ld_data), .b(i_tx_phy_hold_reg_5), .o(g1778_db) );
na02s02 TIMEBOOST_cell_425 ( .a(TIMEBOOST_net_153), .b(n_85), .o(TIMEBOOST_net_126) );
in01s01 g1779_u0 ( .a(i_tx_phy_ld_data), .o(g1779_sb) );
na02s01 TIMEBOOST_cell_405 ( .a(n_130), .b(g2063_sb), .o(TIMEBOOST_net_148) );
na02s01 g1779_u2 ( .a(i_tx_phy_ld_data), .b(i_tx_phy_hold_reg_6), .o(g1779_db) );
na03s03 TIMEBOOST_cell_256 ( .a(n_940), .b(n_942), .c(n_112), .o(n_943) );
in01s01 g1780_u0 ( .a(i_tx_phy_ld_data), .o(g1780_sb) );
na02s02 TIMEBOOST_cell_204 ( .a(TIMEBOOST_net_80), .b(n_938), .o(TIMEBOOST_net_32) );
na02s01 g1780_u2 ( .a(i_tx_phy_ld_data), .b(i_tx_phy_hold_reg_7), .o(g1780_db) );
na02s01 TIMEBOOST_cell_430 ( .a(n_706), .b(TIMEBOOST_net_21), .o(TIMEBOOST_net_156) );
in01s01 g1781_u0 ( .a(i_tx_phy_ld_data), .o(g1781_sb) );
na02s01 TIMEBOOST_cell_395 ( .a(g1776_db), .b(n_974), .o(TIMEBOOST_net_143) );
na02s01 g1781_u2 ( .a(i_tx_phy_ld_data), .b(i_tx_phy_hold_reg_8), .o(g1781_db) );
na02s01 TIMEBOOST_cell_433 ( .a(TIMEBOOST_net_157), .b(TIMEBOOST_net_140), .o(n_431) );
in01s01 g1782_u0 ( .a(i_tx_phy_ld_data), .o(g1782_sb) );
in01s01 TIMEBOOST_cell_114 ( .a(rst), .o(TIMEBOOST_net_43) );
na02s01 g1782_u2 ( .a(i_tx_phy_ld_data), .b(i_tx_phy_hold_reg_9), .o(g1782_db) );
in01s01 TIMEBOOST_cell_115 ( .a(TIMEBOOST_net_43), .o(TIMEBOOST_net_44) );
no02s02 g1806_u0 ( .a(n_232), .b(n_300), .o(n_369) );
na02s02 g1807_u0 ( .a(n_142), .b(n_764), .o(n_347) );
no02s02 g1808_u0 ( .a(n_307), .b(n_384), .o(n_368) );
na02s02 g1809_u0 ( .a(n_198), .b(rst_cnt_3_), .o(n_292) );
na02s01 g1810_u0 ( .a(n_197), .b(n_69), .o(n_256) );
no02s02 g1811_u0 ( .a(n_377), .b(n_400), .o(n_415) );
ao12s01 g1812_u0 ( .a(n_961), .b(n_152), .c(n_375), .o(n_427) );
na02s01 g1813_u0 ( .a(n_434), .b(DataOut_i_7_), .o(n_462) );
na02s01 g1814_u0 ( .a(i_tx_phy_ld_data), .b(i_tx_phy_hold_reg_10), .o(n_450) );
ao12s02 g1815_u0 ( .a(n_400), .b(n_154), .c(n_341), .o(n_401) );
na02s01 TIMEBOOST_cell_132 ( .a(g1782_sb), .b(DataOut_i_6_), .o(TIMEBOOST_net_54) );
no02s06 g1817_u0 ( .a(n_540), .b(n_666), .o(n_413) );
in01s01 g1819_u0 ( .a(n_426), .o(n_446) );
na02s02 g1820_u0 ( .a(n_424), .b(n_666), .o(n_426) );
ao12s01 g1821_u0 ( .a(FE_RN_2_0), .b(n_435), .c(n_389), .o(n_436) );
no02s01 g1822_u0 ( .a(n_424), .b(n_665), .o(n_425) );
na02s01 TIMEBOOST_cell_392 ( .a(TIMEBOOST_net_141), .b(TIMEBOOST_net_50), .o(g1740_p) );
in01s01 g1828_u0 ( .a(i_tx_phy_ld_data), .o(n_434) );
in01s04 g1830_u0 ( .a(i_rx_phy_rxdn_s), .o(n_424) );
ao12s01 g1837_u0 ( .a(FE_RN_2_0), .b(n_63), .c(n_968), .o(n_409) );
ao12s01 g1838_u0 ( .a(n_416), .b(n_251), .c(n_268), .o(n_367) );
ao12s02 g1840_u0 ( .a(n_322), .b(n_330), .c(n_952), .o(n_538) );
ao12s01 g1841_u0 ( .a(n_961), .b(n_355), .c(n_331), .o(n_407) );
na02s01 g1842_u0 ( .a(n_308), .b(TIMEBOOST_net_44), .o(n_366) );
ao12s02 g1843_u0 ( .a(n_400), .b(n_332), .c(n_301), .o(n_395) );
ao12s02 g1844_u0 ( .a(n_400), .b(n_344), .c(n_294), .o(n_394) );
ao12s01 g1845_u0 ( .a(n_961), .b(n_157), .c(n_352), .o(n_406) );
ao12s01 g1846_u0 ( .a(n_961), .b(n_354), .c(n_334), .o(n_405) );
ao12s01 g1848_u0 ( .a(n_400), .b(n_161), .c(n_299), .o(n_378) );
na02s02 g1849_u0 ( .a(n_340), .b(n_138), .o(n_342) );
ao12s01 g1851_u0 ( .a(FE_RN_2_0), .b(n_267), .c(RxActive_o), .o(n_365) );
na02s02 TIMEBOOST_cell_407 ( .a(n_968), .b(n_967), .o(TIMEBOOST_net_149) );
ao12s01 g1853_u0 ( .a(FE_RN_2_0), .b(n_153), .c(n_265), .o(n_364) );
oa12s01 g1854_u0 ( .a(n_133), .b(n_231), .c(i_tx_phy_hold_reg_d_13), .o(n_232) );
in01s01 g1855_u0 ( .a(n_274), .o(g1855_sb) );
na02s02 g1855_u1 ( .a(rst_cnt_4_), .b(g1855_sb), .o(g1855_da) );
na02s01 g1855_u2 ( .a(n_11), .b(n_274), .o(g1855_db) );
na02s02 g1855_u3 ( .a(g1855_da), .b(g1855_db), .o(n_311) );
ao12s02 g1856_u0 ( .a(n_339), .b(n_343), .c(i_tx_phy_bit_cnt_2_), .o(n_377) );
no02s01 g1857_u0 ( .a(n_155), .b(RxValid_o), .o(g1857_p) );
in01s01 g1857_u1 ( .a(g1857_p), .o(n_433) );
na02s01 TIMEBOOST_cell_37 ( .a(n_50), .b(g2674_p), .o(TIMEBOOST_net_15) );
ao12s02 g1859_u0 ( .a(n_391), .b(n_88), .c(n_390), .o(n_421) );
in01s01 g1860_u0 ( .a(n_197), .o(n_198) );
no02s01 g1865_u0 ( .a(n_274), .b(n_11), .o(n_275) );
na02s02 g1867_u0 ( .a(n_121), .b(n_958), .o(n_375) );
na02s02 g1868_u0 ( .a(n_340), .b(n_116), .o(n_341) );
no02s02 g1869_u0 ( .a(n_313), .b(n_416), .o(n_362) );
ao12s02 g1870_u0 ( .a(n_343), .b(n_126), .c(n_231), .o(n_339) );
na02s01 g1871_u0 ( .a(n_223), .b(i_rx_phy_rxdn_s_r), .o(n_310) );
na02s01 g1872_u0 ( .a(n_227), .b(i_rx_phy_rxdp_s_r), .o(n_309) );
na02s01 TIMEBOOST_cell_435 ( .a(TIMEBOOST_net_158), .b(TIMEBOOST_net_148), .o(n_203) );
no02s02 g1874_u0 ( .a(n_390), .b(n_389), .o(n_391) );
na02s01 TIMEBOOST_cell_67 ( .a(n_435), .b(rst), .o(TIMEBOOST_net_30) );
na02s02 TIMEBOOST_cell_442 ( .a(n_783), .b(n_176), .o(TIMEBOOST_net_162) );
ao12s02 g1877_u0 ( .a(n_228), .b(n_254), .c(i_tx_phy_bit_cnt_2_), .o(n_337) );
oa12s01 g1878_u0 ( .a(n_351), .b(n_290), .c(n_583), .o(n_387) );
ao22s01 g1879_u0 ( .a(n_225), .b(i_tx_phy_sd_nrzi_o), .c(n_873), .d(txdp), .o(n_308) );
in01s01 TIMEBOOST_cell_116 ( .a(TIMEBOOST_net_45), .o(DataIn_o_7_) );
no02s01 g1881_u0 ( .a(i_rx_phy_bit_cnt_2_), .b(n_141), .o(g1881_p) );
ao12s01 g1881_u1 ( .a(g1881_p), .b(i_rx_phy_bit_cnt_2_), .c(n_141), .o(n_142) );
ao12s02 g1882_u0 ( .a(n_230), .b(n_132), .c(n_306), .o(n_307) );
no02s01 g1884_u0 ( .a(i_tx_phy_one_cnt_2_), .b(n_51), .o(g1884_p) );
ao12s01 g1884_u1 ( .a(g1884_p), .b(i_tx_phy_one_cnt_2_), .c(n_51), .o(n_138) );
na02s01 TIMEBOOST_cell_55 ( .a(n_53), .b(g2674_p), .o(TIMEBOOST_net_24) );
no02s02 g1896_u0 ( .a(n_132), .b(n_70), .o(n_197) );
na02s01 g1897_u0 ( .a(n_764), .b(i_rx_phy_shift_en), .o(g1897_u0_o) );
no02s02 g1899_u0 ( .a(n_258), .b(n_984), .o(n_340) );
na02s02 g1900_u0 ( .a(n_764), .b(n_118), .o(n_334) );
na02s01 g1901_u0 ( .a(n_764), .b(i_rx_phy_rx_valid1), .o(g1901_p) );
in01s01 g1901_u1 ( .a(g1901_p), .o(n_373) );
na02s01 g1902_u0 ( .a(n_763), .b(i_rx_phy_bit_cnt_2_), .o(n_359) );
na02s01 TIMEBOOST_cell_128 ( .a(g1780_sb), .b(DataOut_i_4_), .o(TIMEBOOST_net_52) );
na02s01 g1904_u0 ( .a(rst), .b(n_283), .o(n_333) );
in01s01 g1905_u0 ( .a(n_416), .o(n_269) );
na02s01 g1906_u0 ( .a(n_191), .b(rst), .o(n_416) );
na02s02 g1907_u0 ( .a(n_106), .b(n_103), .o(n_268) );
no02s02 g1908_u0 ( .a(n_132), .b(n_306), .o(n_230) );
na02s02 g1913_u0 ( .a(n_343), .b(i_tx_phy_bit_cnt_0_), .o(n_332) );
na02s02 g1914_u0 ( .a(n_296), .b(n_56), .o(n_301) );
na02s02 g1915_u0 ( .a(n_343), .b(n_15), .o(n_344) );
na02s02 g1916_u0 ( .a(n_764), .b(n_37), .o(n_331) );
na02s02 g1917_u0 ( .a(n_930), .b(n_841), .o(n_330) );
na02s01 g1918_u0 ( .a(n_763), .b(n_353), .o(n_354) );
na02s01 g1919_u0 ( .a(n_763), .b(i_rx_phy_bit_cnt_0_), .o(n_355) );
no02s02 g1921_u0 ( .a(n_255), .b(i_tx_phy_bit_cnt_2_), .o(n_300) );
na02s02 g1922_u0 ( .a(n_71), .b(n_66), .o(n_274) );
no02s02 g1923_u0 ( .a(n_312), .b(n_540), .o(g1923_p) );
in01s02 g1923_u1 ( .a(g1923_p), .o(n_390) );
na02s01 TIMEBOOST_cell_57 ( .a(n_425), .b(n_175), .o(TIMEBOOST_net_25) );
na02s01 TIMEBOOST_cell_65 ( .a(i_rx_phy_dpll_state_1_), .b(n_60), .o(TIMEBOOST_net_29) );
na02s02 TIMEBOOST_cell_429 ( .a(TIMEBOOST_net_155), .b(n_942), .o(TIMEBOOST_net_80) );
na02s01 TIMEBOOST_cell_75 ( .a(n_238), .b(rst), .o(TIMEBOOST_net_34) );
oa12s01 g1928_u0 ( .a(n_131), .b(n_127), .c(i_rx_phy_rxd_s1), .o(n_229) );
na02s02 g1931_u0 ( .a(n_169), .b(n_296), .o(n_294) );
oa12s02 g1932_u0 ( .a(n_193), .b(n_97), .c(n_804), .o(n_228) );
ao22s02 g1933_u0 ( .a(n_122), .b(n_266), .c(n_150), .d(i_rx_phy_sd_nrzi), .o(n_267) );
oa12s01 g1934_u0 ( .a(n_184), .b(n_186), .c(n_48), .o(n_265) );
in01s01 g1935_u0 ( .a(n_263), .o(n_293) );
na02s01 TIMEBOOST_cell_400 ( .a(TIMEBOOST_net_145), .b(TIMEBOOST_net_49), .o(g1742_p) );
ao22s01 g1937_u0 ( .a(n_100), .b(n_885), .c(i_tx_phy_sd_nrzi_o), .d(n_873), .o(n_195) );
na02s01 g1942_u0 ( .a(i_tx_phy_data_done), .b(n_937), .o(g1942_p) );
in01s01 g1942_u1 ( .a(g1942_p), .o(n_350) );
no02s02 g1950_u0 ( .a(n_210), .b(n_882), .o(n_296) );
na02s02 g1951_u0 ( .a(n_182), .b(n_885), .o(n_343) );
in01s01 g1952_u0 ( .a(n_324), .o(n_325) );
na02s02 g1953_u0 ( .a(n_759), .b(i_rx_phy_sd_nrzi), .o(n_324) );
in01s01 g1954_u0 ( .a(n_258), .o(n_259) );
na02s02 g1955_u0 ( .a(n_182), .b(i_tx_phy_sd_raw_o), .o(n_258) );
no02s01 g1956_u0 ( .a(n_965), .b(n_929), .o(n_323) );
na02s01 TIMEBOOST_cell_432 ( .a(TIMEBOOST_net_36), .b(n_141), .o(TIMEBOOST_net_157) );
in01s02 g1959_u0 ( .a(n_573), .o(n_322) );
no02s01 g1961_u0 ( .a(n_233), .b(n_318), .o(n_320) );
no02s01 g1962_u0 ( .a(n_239), .b(n_318), .o(n_319) );
no02s01 g1963_u0 ( .a(n_318), .b(n_201), .o(n_291) );
in01s01 g1964_u0 ( .a(n_289), .o(n_290) );
na02s01 g1965_u0 ( .a(n_965), .b(n_937), .o(g1965_p) );
in01s01 g1965_u1 ( .a(g1965_p), .o(n_289) );
no02s01 g1966_u0 ( .a(n_237), .b(n_318), .o(n_317) );
no02s01 g1967_u0 ( .a(n_235), .b(FE_RN_2_0), .o(n_316) );
no02s01 g1968_u0 ( .a(n_204), .b(FE_RN_2_0), .o(n_288) );
na02s01 TIMEBOOST_cell_31 ( .a(i_rx_phy_rx_valid1), .b(rst), .o(TIMEBOOST_net_12) );
in01s01 g1974_u0 ( .a(n_226), .o(n_227) );
na02s01 g1975_u0 ( .a(i_rx_phy_rxdp_s0), .b(LineState_o_0_), .o(g1975_p) );
in01s01 g1975_u1 ( .a(g1975_p), .o(n_226) );
oa12s01 g1977_u0 ( .a(n_183), .b(n_185), .c(n_224), .o(n_225) );
oa12s02 g1978_u0 ( .a(n_927), .b(n_952), .c(n_224), .o(n_539) );
in01s01 g1979_u0 ( .a(n_222), .o(n_223) );
na02s01 g1980_u0 ( .a(i_rx_phy_rxdn_s0), .b(LineState_o_1_), .o(g1980_p) );
in01s01 g1980_u1 ( .a(g1980_p), .o(n_222) );
no02s02 g1981_u0 ( .a(LineState_o_0_), .b(LineState_o_1_), .o(n_191) );
na02s04 TIMEBOOST_cell_23 ( .a(n_894), .b(TxValid_i), .o(TIMEBOOST_net_8) );
ao12s01 g1983_u0 ( .a(n_167), .b(n_192), .c(i_tx_phy_hold_reg_d), .o(n_255) );
oa12s02 g1984_u0 ( .a(n_172), .b(i_tx_phy_hold_reg_d_15), .c(n_168), .o(n_254) );
ao12s01 g1985_u0 ( .a(n_213), .b(n_852), .c(txoe), .o(n_283) );
ao12s01 g1986_u0 ( .a(n_241), .b(n_384), .c(n_240), .o(n_313) );
na02s02 g1987_u0 ( .a(n_246), .b(n_245), .o(n_312) );
in01s02 g1991_u0 ( .a(n_66), .o(n_132) );
in01s01 g1998_u0 ( .a(n_949), .o(n_782) );
na02s01 g2000_u0 ( .a(i_rx_phy_rxd_s0), .b(n_130), .o(n_131) );
in01s01 g2003_u0 ( .a(n_982), .o(n_217) );
no02s01 g2010_u0 ( .a(n_185), .b(i_tx_phy_sd_nrzi_o), .o(n_186) );
na02s01 g2011_u0 ( .a(n_384), .b(rst_cnt_4_), .o(n_252) );
na02s01 g2012_u0 ( .a(n_224), .b(n_183), .o(n_184) );
no02s04 TIMEBOOST_cell_17 ( .a(n_929), .b(n_735), .o(TIMEBOOST_net_5) );
na02s01 g2015_u0 ( .a(n_277), .b(n_48), .o(n_280) );
na02s01 g2016_u0 ( .a(n_384), .b(n_105), .o(n_251) );
in01s01 g2020_u0 ( .a(n_759), .o(n_248) );
no02s01 g2024_u0 ( .a(i_rx_phy_rxd_s0), .b(n_130), .o(n_127) );
in01s01 g2026_u0 ( .a(n_182), .o(n_210) );
na02s04 g2027_u0 ( .a(n_55), .b(n_50), .o(n_182) );
no02s04 g2028_u0 ( .a(n_244), .b(n_243), .o(g2028_p) );
in01s02 g2028_u1 ( .a(g2028_p), .o(n_246) );
na02s02 g2029_u0 ( .a(n_244), .b(n_243), .o(n_245) );
na02s01 g2030_u0 ( .a(i_tx_phy_hold_reg_d_12), .b(n_124), .o(n_97) );
no02s01 g2035_u0 ( .a(n_125), .b(n_124), .o(g2035_p) );
in01s01 g2035_u1 ( .a(g2035_p), .o(n_126) );
na02s02 g2036_u0 ( .a(n_125), .b(n_124), .o(n_231) );
in01s01 g2038_u0 ( .a(n_604), .o(n_209) );
no02s02 g2040_u0 ( .a(n_384), .b(n_240), .o(n_241) );
in01s01 g2042_u0 ( .a(n_175), .o(n_176) );
na02s02 g2043_u0 ( .a(n_948), .b(n_794), .o(n_175) );
na02s01 g2048_u0 ( .a(n_277), .b(i_tx_phy_sd_bs_o), .o(n_278) );
no02s01 g2050_u0 ( .a(n_804), .b(n_785), .o(g2050_p) );
in01s01 g2050_u1 ( .a(g2050_p), .o(n_172) );
in01s01 g2051_u0 ( .a(n_123), .o(n_170) );
ao12s01 g2052_u0 ( .a(i_tx_phy_append_eop_sync2), .b(n_7), .c(n_48), .o(n_123) );
na02s01 g2053_u0 ( .a(n_804), .b(n_168), .o(n_169) );
no02s01 g2054_u0 ( .a(n_168), .b(i_tx_phy_hold_reg_d_11), .o(n_167) );
ao12s01 g2055_u0 ( .a(n_164), .b(n_10), .c(i_tx_phy_tx_ip), .o(n_166) );
ao12s01 g2056_u0 ( .a(n_164), .b(n_888), .c(n_737), .o(n_165) );
no02s01 g2057_u0 ( .a(i_rx_phy_sd_r), .b(n_243), .o(g2057_p) );
ao12s01 g2057_u1 ( .a(g2057_p), .b(i_rx_phy_sd_r), .c(n_243), .o(n_122) );
oa12s01 g2058_u0 ( .a(n_35), .b(i_tx_phy_sd_bs_o), .c(i_tx_phy_sd_nrzi_o), .o(n_100) );
ao22s01 g2059_u0 ( .a(i_tx_phy_tx_ip), .b(n_885), .c(n_238), .d(n_984), .o(n_239) );
ao22s01 g2060_u0 ( .a(i_tx_phy_append_eop), .b(g2674_p), .c(i_tx_phy_append_eop_sync1), .d(n_984), .o(n_237) );
ao22s01 g2061_u0 ( .a(i_tx_phy_append_eop_sync1), .b(n_885), .c(i_tx_phy_append_eop_sync2), .d(n_864), .o(n_235) );
ao22s01 g2062_u0 ( .a(i_tx_phy_append_eop_sync4), .b(n_852), .c(n_48), .d(g2674_p), .o(n_204) );
in01s01 g2063_u0 ( .a(n_852), .o(g2063_sb) );
na02s01 TIMEBOOST_cell_262 ( .a(i_tx_phy_hold_reg_d_17), .b(i_tx_phy_bit_cnt_2_), .o(TIMEBOOST_net_95) );
na02s02 TIMEBOOST_cell_443 ( .a(TIMEBOOST_net_162), .b(n_782), .o(n_493) );
na02s01 TIMEBOOST_cell_288 ( .a(n_583), .b(n_800), .o(TIMEBOOST_net_108) );
ao22s01 g2064_u0 ( .a(i_tx_phy_txoe_r2), .b(n_852), .c(i_tx_phy_txoe_r1), .d(g2674_p), .o(n_201) );
ao22s01 g2065_u0 ( .a(n_238), .b(g2674_p), .c(i_tx_phy_txoe_r1), .d(n_984), .o(n_233) );
no02s02 g2066_u0 ( .a(n_105), .b(n_240), .o(g2066_p) );
ao12s02 g2066_u1 ( .a(g2066_p), .b(n_105), .c(n_240), .o(n_106) );
no02s01 g2067_u0 ( .a(n_120), .b(i_rx_phy_one_cnt_0_), .o(g2067_p) );
ao12s02 g2067_u1 ( .a(g2067_p), .b(n_120), .c(i_rx_phy_one_cnt_0_), .o(n_121) );
no02s01 g2068_u0 ( .a(n_353), .b(i_rx_phy_bit_cnt_0_), .o(g2068_p) );
ao12s01 g2068_u1 ( .a(g2068_p), .b(n_353), .c(i_rx_phy_bit_cnt_0_), .o(n_118) );
no02s01 g2069_u0 ( .a(n_115), .b(i_tx_phy_one_cnt_0_), .o(g2069_p) );
ao12s02 g2069_u1 ( .a(g2069_p), .b(n_115), .c(i_tx_phy_one_cnt_0_), .o(n_116) );
in01s02 g2072_u0 ( .a(i_tx_phy_sft_done_r), .o(n_64) );
in01s03 g2084_u0 ( .a(i_rx_phy_rxd_r), .o(n_244) );
na02s01 g2087_u0 ( .a(i_tx_phy_one_cnt_2_), .b(n_873), .o(n_163) );
na02s01 g2088_u0 ( .a(n_873), .b(i_tx_phy_one_cnt_0_), .o(n_161) );
na02s01 g2090_u0 ( .a(i_tx_phy_append_eop), .b(n_12), .o(n_63) );
no02s01 g2091_u0 ( .a(phy_tx_mode), .b(n_984), .o(g2091_p) );
in01s01 g2091_u1 ( .a(g2091_p), .o(n_183) );
in01s02 g2092_u0 ( .a(n_111), .o(n_112) );
na02s04 g2093_u0 ( .a(n_910), .b(n_91), .o(n_111) );
in01s04 g2095_u0 ( .a(n_103), .o(n_384) );
no02s03 g2096_u0 ( .a(n_984), .b(usb_rst), .o(n_103) );
na02s02 g2099_u0 ( .a(n_57), .b(i_tx_phy_bit_cnt_0_), .o(n_168) );
na02s01 TIMEBOOST_cell_393 ( .a(g1780_db), .b(n_974), .o(TIMEBOOST_net_142) );
no02s04 g2100_u0 ( .a(RxActive_o), .b(n_878), .o(n_61) );
na02s01 g2103_u0 ( .a(n_882), .b(rst), .o(g2103_p) );
in01s01 g2103_u1 ( .a(g2103_p), .o(n_277) );
na02s01 g2104_u0 ( .a(i_rx_phy_one_cnt_0_), .b(n_873), .o(n_157) );
in01s01 g2106_u0 ( .a(n_598), .o(n_661) );
na02s01 g2108_u0 ( .a(n_882), .b(i_rx_phy_rx_valid_r), .o(g2108_p) );
in01s01 g2108_u1 ( .a(g2108_p), .o(n_155) );
na02s01 g2109_u0 ( .a(n_115), .b(n_873), .o(n_154) );
na02s02 g2111_u0 ( .a(i_tx_phy_bit_cnt_1_), .b(n_56), .o(n_804) );
in01s01 g2112_u0 ( .a(n_389), .o(n_81) );
no02s01 g2113_u0 ( .a(i_rx_phy_dpll_state_1_), .b(n_60), .o(g2113_p) );
in01s01 g2113_u1 ( .a(g2113_p), .o(n_389) );
na02s01 g2114_u0 ( .a(n_852), .b(txdn), .o(n_153) );
na02s01 g2115_u0 ( .a(n_873), .b(n_120), .o(n_152) );
na02s02 g2116_u0 ( .a(n_57), .b(n_56), .o(g2116_p) );
in01s01 g2116_u1 ( .a(g2116_p), .o(n_192) );
in01s01 g2117_u0 ( .a(n_164), .o(n_108) );
na02s01 g2118_u0 ( .a(rst), .b(TxValid_i), .o(n_164) );
in01m02 g2119_u0 ( .a(n_697), .o(n_90) );
no02s06 g2122_u0 ( .a(n_52), .b(n_28), .o(n_58) );
no02s02 g2123_u0 ( .a(n_56), .b(n_57), .o(n_125) );
no02s01 g2124_u0 ( .a(i_rx_phy_dpll_state_1_), .b(i_rx_phy_dpll_state_0_), .o(n_88) );
in01s01 g2127_u0 ( .a(n_400), .o(n_85) );
no02s02 g2128_u0 ( .a(n_27), .b(n_318), .o(g2128_p) );
in01s02 g2128_u1 ( .a(g2128_p), .o(n_400) );
in01s01 g2129_u0 ( .a(n_150), .o(n_266) );
no02s01 g2130_u0 ( .a(n_884), .b(n_509), .o(g2130_p) );
in01s01 g2130_u1 ( .a(g2130_p), .o(n_150) );
no02s02 g2131_u0 ( .a(n_70), .b(n_69), .o(n_71) );
no02s02 g2135_u0 ( .a(n_37), .b(n_18), .o(n_141) );
no02s02 g2136_u0 ( .a(n_21), .b(n_22), .o(n_66) );
no02s02 g2137_u0 ( .a(n_53), .b(n_52), .o(n_54) );
na02s01 g2138_u0 ( .a(i_tx_phy_sd_bs_o), .b(i_tx_phy_sd_nrzi_o), .o(n_35) );
no02s02 g2139_u0 ( .a(n_50), .b(n_49), .o(n_51) );
no02s04 g2140_u0 ( .a(n_49), .b(n_33), .o(n_55) );
no02s02 g2141_u0 ( .a(n_8), .b(n_984), .o(g2141_p) );
in01s01 g2141_u1 ( .a(g2141_p), .o(n_185) );
in01s01 g2145_u0 ( .a(n_559), .o(n_48) );
in01s01 g2149_u0 ( .a(n_306), .o(n_70) );
in01s01 g2152_u0 ( .a(i_rx_phy_bit_cnt_0_), .o(n_37) );
in01s04 g2155_u0 ( .a(i_tx_phy_one_cnt_0_), .o(n_50) );
in01s01 g2157_u0 ( .a(i_rx_phy_dpll_state_0_), .o(n_60) );
in01s01 g2158_u0 ( .a(phy_tx_mode), .o(n_8) );
in01s02 g2159_u0 ( .a(n_52), .o(n_120) );
in01s08 g2160_u0 ( .a(i_rx_phy_one_cnt_1_), .o(n_52) );
in01s01 g2161_u0 ( .a(i_tx_phy_append_eop_sync2), .o(n_12) );
in01s01 g2162_u0 ( .a(rst_cnt_4_), .o(n_11) );
in01s01 g2164_u0 ( .a(n_238), .o(n_27) );
in01s01 g2172_u0 ( .a(n_22), .o(n_105) );
in01s02 g2173_u0 ( .a(rst_cnt_1_), .o(n_22) );
in01s01 g2174_u0 ( .a(i_tx_phy_append_eop_sync4), .o(n_7) );
in01s01 g2178_u0 ( .a(n_56), .o(n_77) );
in01s02 g2182_u0 ( .a(i_tx_phy_bit_cnt_0_), .o(n_56) );
in01s01 g2183_u0 ( .a(n_57), .o(n_15) );
in01s02 g2186_u0 ( .a(i_tx_phy_bit_cnt_1_), .o(n_57) );
in01s02 g2190_u0 ( .a(RxActive_o), .o(n_509) );
in01s01 g2194_u0 ( .a(i_tx_phy_bit_cnt_2_), .o(n_124) );
in01s02 g2195_u0 ( .a(rst), .o(n_318) );
in01s01 g2218_u0 ( .a(n_49), .o(n_115) );
in01s04 g2219_u0 ( .a(i_tx_phy_one_cnt_1_), .o(n_49) );
in01s01 g2224_u0 ( .a(n_28), .o(n_139) );
in01s06 g2225_u0 ( .a(i_rx_phy_one_cnt_2_), .o(n_28) );
in01s02 g2226_u0 ( .a(n_91), .o(n_74) );
in01s06 g2227_u0 ( .a(n_980), .o(n_91) );
in01s01 g2251_u0 ( .a(i_tx_phy_data_done), .o(n_10) );
in01s02 g2253_u0 ( .a(n_21), .o(n_240) );
in01s02 g2254_u0 ( .a(rst_cnt_0_), .o(n_21) );
in01s02 g2257_u0 ( .a(rst_cnt_3_), .o(n_69) );
in01s01 g2258_u0 ( .a(i_rx_phy_se0_s), .o(n_9) );
in01s01 g2270_u0 ( .a(n_353), .o(n_18) );
in01s02 g2272_u0 ( .a(i_tx_phy_one_cnt_2_), .o(n_33) );
in01s01 g2273_u0 ( .a(n_243), .o(n_130) );
in01s04 g2275_u0 ( .a(i_rx_phy_rxd_s), .o(n_243) );
in01s03 g2278_u0 ( .a(i_rx_phy_one_cnt_0_), .o(n_53) );
in01s01 g22_u0 ( .a(n_852), .o(n_988) );
na02s01 g2385_u0 ( .a(n_885), .b(n_559), .o(g2385_p) );
in01s02 g2385_u1 ( .a(g2385_p), .o(n_567) );
na02s02 g2389_u0 ( .a(n_840), .b(n_567), .o(n_573) );
na02s01 TIMEBOOST_cell_182 ( .a(TIMEBOOST_net_69), .b(n_266), .o(n_479) );
no02s02 g2392_u0 ( .a(n_932), .b(n_952), .o(n_590) );
no02s02 g2397_u0 ( .a(n_952), .b(n_735), .o(n_598) );
na02s02 g23_u0 ( .a(n_604), .b(n_926), .o(n_938) );
no02m02 g2412_u0 ( .a(n_481), .b(n_628), .o(g2412_p) );
in01m02 g2412_u1 ( .a(g2412_p), .o(n_629) );
no02m02 g2413_u0 ( .a(n_727), .b(n_753), .o(g2413_p) );
in01m02 g2413_u1 ( .a(g2413_p), .o(n_628) );
na02s02 g2415_u0 ( .a(n_753), .b(n_74), .o(n_631) );
na02s02 g2431_u0 ( .a(n_749), .b(n_754), .o(n_660) );
in01s01 g2438_u0 ( .a(n_666), .o(n_665) );
in01s10 g2440_u0 ( .a(i_rx_phy_rxdp_s), .o(n_666) );
na02s08 g2459_u0 ( .a(n_980), .b(n_910), .o(n_697) );
in01m02 g2460_u0 ( .a(n_703), .o(n_704) );
na02s01 TIMEBOOST_cell_398 ( .a(TIMEBOOST_net_144), .b(TIMEBOOST_net_54), .o(g1743_p) );
na02s01 TIMEBOOST_cell_183 ( .a(i_rx_phy_shift_en), .b(n_852), .o(TIMEBOOST_net_70) );
na02s01 TIMEBOOST_cell_289 ( .a(TIMEBOOST_net_108), .b(n_350), .o(n_351) );
no02s01 g2465_u0 ( .a(n_540), .b(n_318), .o(n_706) );
na04s02 TIMEBOOST_cell_226 ( .a(n_280), .b(rst), .c(g2674_p), .d(n_170), .o(n_338) );
na02m02 g2477_u0 ( .a(n_726), .b(n_741), .o(n_727) );
no02s06 g2479_u0 ( .a(n_788), .b(n_697), .o(n_722) );
na02s01 TIMEBOOST_cell_134 ( .a(g1778_sb), .b(DataOut_i_2_), .o(TIMEBOOST_net_55) );
in01s01 g2487_u0 ( .a(n_735), .o(n_734) );
in01s02 g2491_u0 ( .a(n_735), .o(n_737) );
na02s02 g2494_u0 ( .a(n_742), .b(n_741), .o(g2494_p) );
in01s02 g2494_u1 ( .a(g2494_p), .o(n_743) );
na02s04 g2495_u0 ( .a(n_942), .b(n_914), .o(n_742) );
na02s01 TIMEBOOST_cell_440 ( .a(n_559), .b(rst), .o(TIMEBOOST_net_161) );
in01s06 g24_u0 ( .a(n_941), .o(n_942) );
ao12m02 g2501_u0 ( .a(n_318), .b(n_755), .c(n_756), .o(n_758) );
oa12m02 g2502_u0 ( .a(n_754), .b(n_944), .c(n_752), .o(n_755) );
na02s02 g2503_u0 ( .a(n_480), .b(n_742), .o(n_752) );
in01s02 g2504_u0 ( .a(n_753), .o(n_754) );
na02s01 TIMEBOOST_cell_384 ( .a(TIMEBOOST_net_137), .b(TIMEBOOST_net_35), .o(n_263) );
no02s02 g2506_u0 ( .a(n_460), .b(n_910), .o(g2506_p) );
in01s02 g2506_u1 ( .a(g2506_p), .o(n_756) );
na02s02 TIMEBOOST_cell_33 ( .a(n_593), .b(n_737), .o(TIMEBOOST_net_13) );
in01s02 g2511_u0 ( .a(n_763), .o(n_764) );
na02s04 g2512_u0 ( .a(n_759), .b(n_885), .o(n_763) );
na02s06 g2513_u0 ( .a(n_58), .b(n_53), .o(n_759) );
in01s01 g2527_u0 ( .a(n_788), .o(n_786) );
in01s01 g2537_u0 ( .a(n_965), .o(n_800) );
in01s02 g2568_u0 ( .a(n_841), .o(n_840) );
in01s02 g2573_u0 ( .a(g2674_p), .o(n_852) );
in01s01 g2584_u0 ( .a(n_885), .o(n_864) );
in01s01 g2593_u0 ( .a(n_885), .o(n_873) );
in01s02 g2595_u0 ( .a(n_885), .o(n_878) );
in01s01 g2599_u0 ( .a(n_885), .o(n_882) );
no02s04 TIMEBOOST_cell_18 ( .a(TIMEBOOST_net_5), .b(n_952), .o(n_583) );
in01s01 g2601_u0 ( .a(n_885), .o(n_884) );
in01s01 g2604_u0 ( .a(n_929), .o(n_888) );
in01s08 g2610_u0 ( .a(n_929), .o(n_894) );
no02s01 g2620_u0 ( .a(n_923), .b(n_924), .o(n_925) );
ao12s02 g2621_u0 ( .a(n_922), .b(n_915), .c(n_916), .o(n_923) );
na02s02 g2622_u0 ( .a(n_920), .b(n_921), .o(n_922) );
ao22s01 g2623_u0 ( .a(n_919), .b(n_945), .c(n_722), .d(n_916), .o(n_920) );
ao22s02 g2624_u0 ( .a(n_927), .b(n_928), .c(n_934), .d(n_929), .o(n_935) );
no02s02 g2625_u0 ( .a(n_661), .b(n_888), .o(n_927) );
no02s01 g2626_u0 ( .a(n_224), .b(n_888), .o(n_928) );
na02s02 g2627_u0 ( .a(n_930), .b(n_933), .o(n_934) );
na02s01 TIMEBOOST_cell_79 ( .a(i_rx_phy_bit_cnt_2_), .b(rst), .o(TIMEBOOST_net_36) );
na02s02 g2630_u0 ( .a(n_965), .b(n_932), .o(n_933) );
na02s03 g2632_u0 ( .a(n_64), .b(i_tx_phy_sft_done), .o(n_932) );
in01s01 g2634_u0 ( .a(n_932), .o(n_937) );
na02s02 g2635_u0 ( .a(n_938), .b(n_943), .o(n_944) );
na02s01 TIMEBOOST_cell_49 ( .a(RxActive_o), .b(rst), .o(TIMEBOOST_net_21) );
in01s01 g2637_u0 ( .a(n_794), .o(n_940) );
na02s06 g2638_u0 ( .a(n_413), .b(n_424), .o(n_941) );
no02s01 g2639_u0 ( .a(n_794), .b(n_111), .o(n_945) );
no02s02 g2640_u0 ( .a(n_980), .b(n_947), .o(n_948) );
in01s02 g2642_u0 ( .a(i_rx_phy_fs_state_2_), .o(n_947) );
in01s08 g2643_u0 ( .a(n_796), .o(n_788) );
na02s01 TIMEBOOST_cell_394 ( .a(TIMEBOOST_net_142), .b(TIMEBOOST_net_52), .o(g1741_p) );
in01s10 g2645_u0 ( .a(n_951), .o(n_952) );
in01s20 g2646_u0 ( .a(i_tx_phy_state_2_), .o(n_951) );
in01s08 g2648_u0 ( .a(i_tx_phy_state_1_), .o(n_735) );
ao12s01 g2650_u0 ( .a(n_961), .b(n_959), .c(n_960), .o(n_962) );
no02s02 g2651_u0 ( .a(n_139), .b(n_54), .o(g2651_p) );
ao12s02 g2651_u1 ( .a(g2651_p), .b(n_139), .c(n_54), .o(n_957) );
no02s04 g2652_u0 ( .a(n_324), .b(n_984), .o(n_958) );
na02s01 g2653_u0 ( .a(i_rx_phy_shift_en), .b(rst), .o(n_961) );
na02s01 TIMEBOOST_cell_290 ( .a(n_289), .b(n_165), .o(TIMEBOOST_net_109) );
oa12s02 g2655_u0 ( .a(n_965), .b(n_734), .c(n_937), .o(n_966) );
na02s01 g2656_u0 ( .a(n_583), .b(n_737), .o(n_967) );
ao12s01 g2657_u0 ( .a(n_318), .b(n_970), .c(n_974), .o(n_976) );
na02s01 g2658_u0 ( .a(n_559), .b(i_tx_phy_tx_ip), .o(n_970) );
na02s02 TIMEBOOST_cell_445 ( .a(TIMEBOOST_net_163), .b(TIMEBOOST_net_149), .o(g1757_p) );
in01s02 g2661_u0 ( .a(n_971), .o(n_972) );
na02s04 g2662_u0 ( .a(n_735), .b(n_951), .o(n_971) );
in01s02 g2664_u0 ( .a(n_974), .o(n_977) );
no02s04 g2665_u0 ( .a(n_913), .b(n_981), .o(n_982) );
in01s06 g2667_u0 ( .a(n_796), .o(n_794) );
na02s04 g2668_u0 ( .a(n_980), .b(i_rx_phy_fs_state_2_), .o(n_981) );
in01s10 g2669_u0 ( .a(i_rx_phy_fs_state_0_), .o(n_980) );
in01s10 g2670_u0 ( .a(i_rx_phy_fs_state_2_), .o(n_910) );
na02s06 TIMEBOOST_cell_14 ( .a(TIMEBOOST_net_3), .b(n_894), .o(n_841) );
na02s06 TIMEBOOST_cell_13 ( .a(n_952), .b(n_735), .o(TIMEBOOST_net_3) );
in01s02 g2674_u0 ( .a(n_984), .o(g2674_p) );
in01s06 g2676_u0 ( .a(n_885), .o(n_984) );
na02s01 TIMEBOOST_cell_401 ( .a(g1778_db), .b(n_974), .o(TIMEBOOST_net_146) );
na02s01 TIMEBOOST_cell_51 ( .a(n_112), .b(n_788), .o(TIMEBOOST_net_22) );
in01s02 g27_u0 ( .a(n_224), .o(n_559) );
na02s02 g31_u0 ( .a(n_958), .b(n_957), .o(n_959) );
na02s02 TIMEBOOST_cell_427 ( .a(TIMEBOOST_net_154), .b(n_968), .o(TIMEBOOST_net_111) );
no02s02 g33_u0 ( .a(n_929), .b(i_tx_phy_data_done), .o(n_593) );
na02s01 g34_u0 ( .a(n_139), .b(n_873), .o(n_960) );
na02m04 g35_u0 ( .a(n_926), .b(n_722), .o(n_741) );
na02m02 TIMEBOOST_cell_87 ( .a(n_90), .b(n_794), .o(TIMEBOOST_net_40) );
ao12s02 g39_u0 ( .a(n_977), .b(n_840), .c(n_567), .o(n_699) );
na02s01 TIMEBOOST_cell_142 ( .a(n_737), .b(n_108), .o(TIMEBOOST_net_59) );
no02s02 g41_u0 ( .a(n_588), .b(n_888), .o(g41_p) );
in01s02 g41_u1 ( .a(g41_p), .o(n_700) );
na02s01 TIMEBOOST_cell_77 ( .a(i_tx_phy_bit_cnt_2_), .b(n_77), .o(TIMEBOOST_net_35) );
no02s02 g44_u0 ( .a(n_971), .b(n_894), .o(n_965) );
in01s01 g51_u0 ( .a(n_583), .o(n_588) );
na02s08 TIMEBOOST_cell_8 ( .a(TIMEBOOST_net_0), .b(n_666), .o(n_916) );
in01s04 g56_u0 ( .a(n_916), .o(n_926) );
na02s02 TIMEBOOST_cell_428 ( .a(n_788), .b(n_112), .o(TIMEBOOST_net_155) );
na03s02 TIMEBOOST_cell_53 ( .a(n_919), .b(n_217), .c(n_209), .o(TIMEBOOST_net_23) );
in01s01 g61_u0 ( .a(n_942), .o(n_919) );
na02s01 g64_u0 ( .a(n_754), .b(n_509), .o(n_924) );
ms00f80 i_rx_phy_bit_cnt_reg_0__u0 ( .ck(ispd_clk), .d(n_407), .o(i_rx_phy_bit_cnt_0_) );
ms00f80 i_rx_phy_bit_cnt_reg_1__u0 ( .ck(ispd_clk), .d(n_405), .o(n_353) );
ms00f80 i_rx_phy_bit_cnt_reg_2__u0 ( .ck(ispd_clk), .d(n_414), .o(i_rx_phy_bit_cnt_2_) );
ms00f80 i_rx_phy_bit_stuff_err_reg_u0 ( .ck(ispd_clk), .d(n_505), .o(i_rx_phy_bit_stuff_err_reg_Q) );
in01s01 i_rx_phy_bit_stuff_err_reg_u1 ( .a(i_rx_phy_bit_stuff_err_reg_Q), .o(i_rx_phy_bit_stuff_err) );
ms00f80 i_rx_phy_byte_err_reg_u0 ( .ck(ispd_clk), .d(n_499), .o(i_rx_phy_byte_err_reg_Q) );
in01s01 i_rx_phy_byte_err_reg_u1 ( .a(i_rx_phy_byte_err_reg_Q), .o(i_rx_phy_byte_err) );
ms00f80 i_rx_phy_dpll_state_reg_0__u0 ( .ck(ispd_clk), .d(n_449), .o(i_rx_phy_dpll_state_0_) );
ms00f80 i_rx_phy_dpll_state_reg_1__u0 ( .ck(ispd_clk), .d(n_436), .o(i_rx_phy_dpll_state_1_) );
ms00f80 i_rx_phy_fs_ce_r1_reg_u0 ( .ck(ispd_clk), .d(n_81), .o(i_rx_phy_fs_ce_r1) );
ms00f80 i_rx_phy_fs_ce_r2_reg_u0 ( .ck(ispd_clk), .d(i_rx_phy_fs_ce_r1), .o(i_rx_phy_fs_ce_r2) );
ms00f80 i_rx_phy_fs_ce_reg_u0 ( .ck(ispd_clk), .d(i_rx_phy_fs_ce_r2), .o(n_885) );
ms00f80 i_rx_phy_fs_state_reg_0__u0 ( .ck(ispd_clk), .d(n_529), .o(i_rx_phy_fs_state_0_) );
ms00f80 i_rx_phy_fs_state_reg_1__u0 ( .ck(ispd_clk), .d(n_523), .o(n_796) );
ms00f80 i_rx_phy_fs_state_reg_2__u0 ( .ck(ispd_clk), .d(n_758), .o(i_rx_phy_fs_state_2_) );
ms00f80 i_rx_phy_hold_reg_reg_0__u0 ( .ck(ispd_clk), .d(DataIn_o_1_), .o(DataIn_o_0_) );
ms00f80 i_rx_phy_hold_reg_reg_1__u0 ( .ck(ispd_clk), .d(DataIn_o_2_), .o(DataIn_o_1_) );
ms00f80 i_rx_phy_hold_reg_reg_2__u0 ( .ck(ispd_clk), .d(DataIn_o_3_), .o(DataIn_o_2_) );
ms00f80 i_rx_phy_hold_reg_reg_3__u0 ( .ck(ispd_clk), .d(DataIn_o_4_), .o(DataIn_o_3_) );
ms00f80 i_rx_phy_hold_reg_reg_4__u0 ( .ck(ispd_clk), .d(DataIn_o_5_), .o(DataIn_o_4_) );
ms00f80 i_rx_phy_hold_reg_reg_5__u0 ( .ck(ispd_clk), .d(DataIn_o_6_), .o(DataIn_o_5_) );
ms00f80 i_rx_phy_hold_reg_reg_6__u0 ( .ck(ispd_clk), .d(DataIn_o_7_), .o(DataIn_o_6_) );
ms00f80 i_rx_phy_hold_reg_reg_7__u0 ( .ck(ispd_clk), .d(i_rx_phy_sd_nrzi), .o(TIMEBOOST_net_46) );
ms00f80 i_rx_phy_one_cnt_reg_0__u0 ( .ck(ispd_clk), .d(n_406), .o(i_rx_phy_one_cnt_0_) );
ms00f80 i_rx_phy_one_cnt_reg_1__u0 ( .ck(ispd_clk), .d(n_427), .o(i_rx_phy_one_cnt_1_) );
ms00f80 i_rx_phy_one_cnt_reg_2__u0 ( .ck(ispd_clk), .d(n_962), .o(i_rx_phy_one_cnt_2_) );
ms00f80 i_rx_phy_rx_active_reg_u0 ( .ck(ispd_clk), .d(n_709), .o(RxActive_o) );
ms00f80 i_rx_phy_rx_en_reg_u0 ( .ck(ispd_clk), .d(txoe), .o(i_rx_phy_rx_en) );
ms00f80 i_rx_phy_rx_valid1_reg_u0 ( .ck(ispd_clk), .d(n_431), .o(i_rx_phy_rx_valid1) );
ms00f80 i_rx_phy_rx_valid_r_reg_u0 ( .ck(ispd_clk), .d(n_433), .o(i_rx_phy_rx_valid_r) );
ms00f80 i_rx_phy_rx_valid_reg_u0 ( .ck(ispd_clk), .d(n_373), .o(RxValid_o) );
ms00f80 i_rx_phy_rxd_r_reg_u0 ( .ck(ispd_clk), .d(n_130), .o(i_rx_phy_rxd_r) );
ms00f80 i_rx_phy_rxd_s0_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_165), .o(i_rx_phy_rxd_s0) );
ms00f80 i_rx_phy_rxd_s1_reg_u0 ( .ck(ispd_clk), .d(i_rx_phy_rxd_s0), .o(i_rx_phy_rxd_s1_reg_Q) );
in01s01 i_rx_phy_rxd_s1_reg_u1 ( .a(i_rx_phy_rxd_s1_reg_Q), .o(i_rx_phy_rxd_s1) );
ms00f80 i_rx_phy_rxd_s_reg_u0 ( .ck(ispd_clk), .d(n_229), .o(i_rx_phy_rxd_s) );
ms00f80 i_rx_phy_rxdn_s0_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_167), .o(i_rx_phy_rxdn_s0) );
ms00f80 i_rx_phy_rxdn_s1_reg_u0 ( .ck(ispd_clk), .d(i_rx_phy_rxdn_s0), .o(LineState_o_1_) );
ms00f80 i_rx_phy_rxdn_s_r_reg_u0 ( .ck(ispd_clk), .d(n_222), .o(i_rx_phy_rxdn_s_r_reg_Q) );
in01s01 i_rx_phy_rxdn_s_r_reg_u1 ( .a(i_rx_phy_rxdn_s_r_reg_Q), .o(i_rx_phy_rxdn_s_r) );
ms00f80 i_rx_phy_rxdn_s_reg_u0 ( .ck(ispd_clk), .d(n_310), .o(i_rx_phy_rxdn_s) );
ms00f80 i_rx_phy_rxdp_s0_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_169), .o(i_rx_phy_rxdp_s0) );
ms00f80 i_rx_phy_rxdp_s1_reg_u0 ( .ck(ispd_clk), .d(i_rx_phy_rxdp_s0), .o(LineState_o_0_) );
ms00f80 i_rx_phy_rxdp_s_r_reg_u0 ( .ck(ispd_clk), .d(n_226), .o(i_rx_phy_rxdp_s_r_reg_Q) );
in01s01 i_rx_phy_rxdp_s_r_reg_u1 ( .a(i_rx_phy_rxdp_s_r_reg_Q), .o(i_rx_phy_rxdp_s_r) );
ms00f80 i_rx_phy_rxdp_s_reg_u0 ( .ck(ispd_clk), .d(n_309), .o(i_rx_phy_rxdp_s) );
ms00f80 i_rx_phy_sd_nrzi_reg_u0 ( .ck(ispd_clk), .d(n_365), .o(i_rx_phy_sd_nrzi) );
ms00f80 i_rx_phy_sd_r_reg_u0 ( .ck(ispd_clk), .d(n_203), .o(i_rx_phy_sd_r) );
ms00f80 i_rx_phy_se0_r_reg_u0 ( .ck(ispd_clk), .d(n_446), .o(i_rx_phy_se0_r_reg_Q) );
in01s01 i_rx_phy_se0_r_reg_u1 ( .a(i_rx_phy_se0_r_reg_Q), .o(i_rx_phy_se0_r) );
ms00f80 i_rx_phy_se0_s_reg_u0 ( .ck(ispd_clk), .d(n_471), .o(i_rx_phy_se0_s) );
ms00f80 i_rx_phy_shift_en_reg_u0 ( .ck(ispd_clk), .d(n_992), .o(i_rx_phy_shift_en) );
ms00f80 i_rx_phy_sync_err_reg_u0 ( .ck(ispd_clk), .d(n_925), .o(i_rx_phy_sync_err_reg_Q) );
in01s01 i_rx_phy_sync_err_reg_u1 ( .a(i_rx_phy_sync_err_reg_Q), .o(i_rx_phy_sync_err) );
ms00f80 i_tx_phy_TxReady_o_reg_u0 ( .ck(ispd_clk), .d(n_392), .o(TxReady_o) );
ms00f80 i_tx_phy_append_eop_reg_u0 ( .ck(ispd_clk), .d(n_409), .o(i_tx_phy_append_eop) );
ms00f80 i_tx_phy_append_eop_sync1_reg_u0 ( .ck(ispd_clk), .d(n_317), .o(i_tx_phy_append_eop_sync1) );
ms00f80 i_tx_phy_append_eop_sync2_reg_u0 ( .ck(ispd_clk), .d(n_316), .o(i_tx_phy_append_eop_sync2) );
ms00f80 i_tx_phy_append_eop_sync3_reg_u0 ( .ck(ispd_clk), .d(n_338), .o(n_224) );
ms00f80 i_tx_phy_append_eop_sync4_reg_u0 ( .ck(ispd_clk), .d(n_288), .o(i_tx_phy_append_eop_sync4) );
ms00f80 i_tx_phy_bit_cnt_reg_0__u0 ( .ck(ispd_clk), .d(n_395), .o(i_tx_phy_bit_cnt_0_) );
ms00f80 i_tx_phy_bit_cnt_reg_1__u0 ( .ck(ispd_clk), .d(n_394), .o(i_tx_phy_bit_cnt_1_) );
ms00f80 i_tx_phy_bit_cnt_reg_2__u0 ( .ck(ispd_clk), .d(n_415), .o(i_tx_phy_bit_cnt_2_) );
ms00f80 i_tx_phy_data_done_reg_u0 ( .ck(ispd_clk), .d(n_166), .o(i_tx_phy_data_done) );
ms00f80 i_tx_phy_hold_reg_d_reg_0__u0 ( .ck(ispd_clk), .d(i_tx_phy_hold_reg), .o(i_tx_phy_hold_reg_d) );
ms00f80 i_tx_phy_hold_reg_d_reg_1__u0 ( .ck(ispd_clk), .d(i_tx_phy_hold_reg_4), .o(i_tx_phy_hold_reg_d_reg_1__Q) );
in01s01 i_tx_phy_hold_reg_d_reg_1__u1 ( .a(i_tx_phy_hold_reg_d_reg_1__Q), .o(i_tx_phy_hold_reg_d_11) );
ms00f80 i_tx_phy_hold_reg_d_reg_2__u0 ( .ck(ispd_clk), .d(i_tx_phy_hold_reg_5), .o(i_tx_phy_hold_reg_d_12) );
ms00f80 i_tx_phy_hold_reg_d_reg_3__u0 ( .ck(ispd_clk), .d(i_tx_phy_hold_reg_6), .o(i_tx_phy_hold_reg_d_reg_3__Q) );
in01s01 i_tx_phy_hold_reg_d_reg_3__u1 ( .a(i_tx_phy_hold_reg_d_reg_3__Q), .o(i_tx_phy_hold_reg_d_13) );
ms00f80 i_tx_phy_hold_reg_d_reg_4__u0 ( .ck(ispd_clk), .d(i_tx_phy_hold_reg_7), .o(i_tx_phy_hold_reg_d_14) );
ms00f80 i_tx_phy_hold_reg_d_reg_5__u0 ( .ck(ispd_clk), .d(i_tx_phy_hold_reg_8), .o(i_tx_phy_hold_reg_d_reg_5__Q) );
in01s01 i_tx_phy_hold_reg_d_reg_5__u1 ( .a(i_tx_phy_hold_reg_d_reg_5__Q), .o(i_tx_phy_hold_reg_d_15) );
ms00f80 i_tx_phy_hold_reg_d_reg_6__u0 ( .ck(ispd_clk), .d(i_tx_phy_hold_reg_9), .o(i_tx_phy_hold_reg_d_reg_6__Q) );
in01s01 i_tx_phy_hold_reg_d_reg_6__u1 ( .a(i_tx_phy_hold_reg_d_reg_6__Q), .o(n_785) );
ms00f80 i_tx_phy_hold_reg_d_reg_7__u0 ( .ck(ispd_clk), .d(i_tx_phy_hold_reg_10), .o(i_tx_phy_hold_reg_d_17) );
ms00f80 i_tx_phy_hold_reg_reg_0__u0 ( .ck(ispd_clk), .d(n_489), .o(i_tx_phy_hold_reg) );
ms00f80 i_tx_phy_hold_reg_reg_1__u0 ( .ck(ispd_clk), .d(n_487), .o(i_tx_phy_hold_reg_4) );
ms00f80 i_tx_phy_hold_reg_reg_2__u0 ( .ck(ispd_clk), .d(n_486), .o(i_tx_phy_hold_reg_5) );
ms00f80 i_tx_phy_hold_reg_reg_3__u0 ( .ck(ispd_clk), .d(n_485), .o(i_tx_phy_hold_reg_6) );
ms00f80 i_tx_phy_hold_reg_reg_4__u0 ( .ck(ispd_clk), .d(n_484), .o(i_tx_phy_hold_reg_7) );
ms00f80 i_tx_phy_hold_reg_reg_5__u0 ( .ck(ispd_clk), .d(n_483), .o(i_tx_phy_hold_reg_8) );
ms00f80 i_tx_phy_hold_reg_reg_6__u0 ( .ck(ispd_clk), .d(n_482), .o(i_tx_phy_hold_reg_9) );
ms00f80 i_tx_phy_hold_reg_reg_7__u0 ( .ck(ispd_clk), .d(n_507), .o(i_tx_phy_hold_reg_10) );
ms00f80 i_tx_phy_ld_data_reg_u0 ( .ck(ispd_clk), .d(n_387), .o(i_tx_phy_ld_data_reg_Q) );
in01s02 i_tx_phy_ld_data_reg_u1 ( .a(i_tx_phy_ld_data_reg_Q), .o(i_tx_phy_ld_data) );
ms00f80 i_tx_phy_one_cnt_reg_0__u0 ( .ck(ispd_clk), .d(n_378), .o(i_tx_phy_one_cnt_0_) );
ms00f80 i_tx_phy_one_cnt_reg_1__u0 ( .ck(ispd_clk), .d(n_401), .o(i_tx_phy_one_cnt_1_) );
ms00f80 i_tx_phy_one_cnt_reg_2__u0 ( .ck(ispd_clk), .d(n_388), .o(i_tx_phy_one_cnt_2_) );
ms00f80 i_tx_phy_sd_bs_o_reg_u0 ( .ck(ispd_clk), .d(n_361), .o(i_tx_phy_sd_bs_o) );
ms00f80 i_tx_phy_sd_nrzi_o_reg_u0 ( .ck(ispd_clk), .d(n_276), .o(i_tx_phy_sd_nrzi_o) );
ms00f80 i_tx_phy_sd_raw_o_reg_u0 ( .ck(ispd_clk), .d(n_411), .o(i_tx_phy_sd_raw_o) );
ms00f80 i_tx_phy_sft_done_r_reg_u0 ( .ck(ispd_clk), .d(i_tx_phy_sft_done), .o(i_tx_phy_sft_done_r) );
ms00f80 i_tx_phy_sft_done_reg_u0 ( .ck(ispd_clk), .d(n_293), .o(i_tx_phy_sft_done) );
ms00f80 i_tx_phy_state_reg_0__u0 ( .ck(ispd_clk), .d(n_459), .o(n_929) );
ms00f80 i_tx_phy_state_reg_1__u0 ( .ck(ispd_clk), .d(n_420), .o(i_tx_phy_state_1_) );
ms00f80 i_tx_phy_state_reg_2__u0 ( .ck(ispd_clk), .d(n_432), .o(i_tx_phy_state_2_) );
ms00f80 i_tx_phy_tx_ip_reg_u0 ( .ck(ispd_clk), .d(n_976), .o(i_tx_phy_tx_ip) );
ms00f80 i_tx_phy_tx_ip_sync_reg_u0 ( .ck(ispd_clk), .d(n_319), .o(n_238) );
ms00f80 i_tx_phy_txdn_reg_u0 ( .ck(ispd_clk), .d(n_364), .o(txdn) );
ms00f80 i_tx_phy_txdp_reg_u0 ( .ck(ispd_clk), .d(n_366), .o(txdp) );
ms00f80 i_tx_phy_txoe_r1_reg_u0 ( .ck(ispd_clk), .d(n_320), .o(i_tx_phy_txoe_r1) );
ms00f80 i_tx_phy_txoe_r2_reg_u0 ( .ck(ispd_clk), .d(n_291), .o(i_tx_phy_txoe_r2) );
ms00f80 i_tx_phy_txoe_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_171), .o(txoe) );
ms00f80 rst_cnt_reg_0__u0 ( .ck(ispd_clk), .d(n_362), .o(rst_cnt_0_) );
ms00f80 rst_cnt_reg_1__u0 ( .ck(ispd_clk), .d(n_367), .o(rst_cnt_1_) );
ms00f80 rst_cnt_reg_2__u0 ( .ck(ispd_clk), .d(n_428), .o(n_306) );
ms00f80 rst_cnt_reg_3__u0 ( .ck(ispd_clk), .d(n_417), .o(rst_cnt_3_) );
ms00f80 rst_cnt_reg_4__u0 ( .ck(ispd_clk), .d(n_423), .o(rst_cnt_4_) );
ms00f80 usb_rst_reg_u0 ( .ck(ispd_clk), .d(n_275), .o(usb_rst) );
na02s01 TIMEBOOST_cell_29 ( .a(i_tx_phy_hold_reg_d_14), .b(i_tx_phy_bit_cnt_2_), .o(TIMEBOOST_net_11) );
na02s01 TIMEBOOST_cell_260 ( .a(i_rx_phy_bit_stuff_err), .b(i_rx_phy_byte_err), .o(TIMEBOOST_net_94) );
na02s04 TIMEBOOST_cell_24 ( .a(TIMEBOOST_net_8), .b(n_972), .o(n_974) );
na02s01 TIMEBOOST_cell_436 ( .a(n_350), .b(TIMEBOOST_net_27), .o(TIMEBOOST_net_159) );
na02s01 TIMEBOOST_cell_396 ( .a(TIMEBOOST_net_143), .b(TIMEBOOST_net_53), .o(g1737_p) );
na02s01 TIMEBOOST_cell_30 ( .a(TIMEBOOST_net_11), .b(n_192), .o(n_193) );
na02s01 TIMEBOOST_cell_32 ( .a(TIMEBOOST_net_12), .b(n_763), .o(n_767) );
na02s04 TIMEBOOST_cell_34 ( .a(n_590), .b(TIMEBOOST_net_13), .o(n_968) );
na02s02 TIMEBOOST_cell_36 ( .a(TIMEBOOST_net_14), .b(n_195), .o(n_276) );
na02s02 TIMEBOOST_cell_38 ( .a(TIMEBOOST_net_15), .b(n_259), .o(n_299) );
na03s02 TIMEBOOST_cell_438 ( .a(n_509), .b(TIMEBOOST_net_70), .c(n_988), .o(TIMEBOOST_net_160) );
na02s01 TIMEBOOST_cell_261 ( .a(TIMEBOOST_net_94), .b(i_rx_phy_sync_err), .o(RxError_o) );
na02s01 TIMEBOOST_cell_122 ( .a(g1781_sb), .b(DataOut_i_5_), .o(TIMEBOOST_net_49) );
na02s01 TIMEBOOST_cell_130 ( .a(g1776_sb), .b(DataOut_i_0_), .o(TIMEBOOST_net_53) );
na02s01 TIMEBOOST_cell_263 ( .a(TIMEBOOST_net_95), .b(n_125), .o(n_133) );
na02s04 TIMEBOOST_cell_264 ( .a(n_61), .b(n_9), .o(TIMEBOOST_net_96) );
na02s01 TIMEBOOST_cell_52 ( .a(TIMEBOOST_net_22), .b(n_919), .o(n_921) );
na02s01 TIMEBOOST_cell_54 ( .a(TIMEBOOST_net_23), .b(n_914), .o(n_915) );
na02s02 TIMEBOOST_cell_56 ( .a(TIMEBOOST_net_24), .b(n_325), .o(n_352) );
na02s01 TIMEBOOST_cell_58 ( .a(TIMEBOOST_net_25), .b(n_949), .o(n_440) );
na02m02 TIMEBOOST_cell_60 ( .a(n_699), .b(TIMEBOOST_net_26), .o(n_703) );
na02s01 TIMEBOOST_cell_441 ( .a(TIMEBOOST_net_161), .b(n_734), .o(TIMEBOOST_net_117) );
in01s01 TIMEBOOST_cell_117 ( .a(TIMEBOOST_net_46), .o(TIMEBOOST_net_45) );
na02s02 TIMEBOOST_cell_66 ( .a(TIMEBOOST_net_29), .b(n_390), .o(n_435) );
na02s01 TIMEBOOST_cell_68 ( .a(TIMEBOOST_net_30), .b(n_421), .o(n_449) );
no02s01 TIMEBOOST_cell_380 ( .a(TIMEBOOST_net_135), .b(i_tx_phy_txoe_r2), .o(n_213) );
na02s02 TIMEBOOST_cell_72 ( .a(n_743), .b(TIMEBOOST_net_32), .o(n_749) );
na02s06 TIMEBOOST_cell_265 ( .a(TIMEBOOST_net_96), .b(n_426), .o(n_753) );
na02s01 TIMEBOOST_cell_76 ( .a(TIMEBOOST_net_34), .b(i_tx_phy_txoe_r1), .o(TIMEBOOST_net_14) );
na02s01 TIMEBOOST_cell_403 ( .a(g1777_db), .b(n_974), .o(TIMEBOOST_net_147) );
in01s01 TIMEBOOST_cell_446 ( .a(rxd), .o(TIMEBOOST_net_164) );
na02s01 TIMEBOOST_cell_143 ( .a(TIMEBOOST_net_59), .b(n_323), .o(TIMEBOOST_net_27) );
na03s02 TIMEBOOST_cell_359 ( .a(n_735), .b(n_984), .c(n_929), .o(TIMEBOOST_net_4) );
na02s02 TIMEBOOST_cell_439 ( .a(TIMEBOOST_net_160), .b(n_461), .o(TIMEBOOST_net_93) );
na02m02 TIMEBOOST_cell_88 ( .a(n_439), .b(TIMEBOOST_net_40), .o(n_726) );
na02s02 TIMEBOOST_cell_318 ( .a(TIMEBOOST_net_114), .b(n_972), .o(TIMEBOOST_net_98) );
no02s01 TIMEBOOST_cell_379 ( .a(i_tx_phy_txoe_r1), .b(n_864), .o(TIMEBOOST_net_135) );
na02s01 TIMEBOOST_cell_391 ( .a(g1779_db), .b(n_974), .o(TIMEBOOST_net_141) );
na02s01 TIMEBOOST_cell_402 ( .a(TIMEBOOST_net_146), .b(TIMEBOOST_net_55), .o(g1739_p) );
na02s01 TIMEBOOST_cell_423 ( .a(TIMEBOOST_net_152), .b(n_462), .o(n_507) );
na02s01 TIMEBOOST_cell_383 ( .a(n_15), .b(n_182), .o(TIMEBOOST_net_137) );
na02s01 TIMEBOOST_cell_389 ( .a(n_767), .b(n_764), .o(TIMEBOOST_net_140) );
na02s01 TIMEBOOST_cell_397 ( .a(g1782_db), .b(n_974), .o(TIMEBOOST_net_144) );
in01s01 TIMEBOOST_cell_447 ( .a(TIMEBOOST_net_164), .o(TIMEBOOST_net_165) );
in01s01 TIMEBOOST_cell_448 ( .a(rxdn), .o(TIMEBOOST_net_166) );
in01s01 TIMEBOOST_cell_449 ( .a(TIMEBOOST_net_166), .o(TIMEBOOST_net_167) );
in01s01 TIMEBOOST_cell_450 ( .a(rxdp), .o(TIMEBOOST_net_168) );
in01s01 TIMEBOOST_cell_451 ( .a(TIMEBOOST_net_168), .o(TIMEBOOST_net_169) );
in01s01 TIMEBOOST_cell_452 ( .a(n_333), .o(TIMEBOOST_net_170) );
in01s01 TIMEBOOST_cell_453 ( .a(TIMEBOOST_net_170), .o(TIMEBOOST_net_171) );

endmodule
