module pci_bridge32_fast (
ispd_clk,
pci_ad_i_0_,
pci_ad_i_10_,
pci_ad_i_11_,
pci_ad_i_12_,
pci_ad_i_13_,
pci_ad_i_14_,
pci_ad_i_15_,
pci_ad_i_16_,
pci_ad_i_17_,
pci_ad_i_18_,
pci_ad_i_19_,
pci_ad_i_1_,
pci_ad_i_20_,
pci_ad_i_21_,
pci_ad_i_22_,
pci_ad_i_23_,
pci_ad_i_24_,
pci_ad_i_25_,
pci_ad_i_26_,
pci_ad_i_27_,
pci_ad_i_28_,
pci_ad_i_29_,
pci_ad_i_2_,
pci_ad_i_30_,
pci_ad_i_31_,
pci_ad_i_3_,
pci_ad_i_4_,
pci_ad_i_5_,
pci_ad_i_6_,
pci_ad_i_7_,
pci_ad_i_8_,
pci_ad_i_9_,
pci_cbe_i_0_,
pci_cbe_i_1_,
pci_cbe_i_2_,
pci_cbe_i_3_,
pci_devsel_i,
pci_frame_i,
pci_gnt_i,
pci_idsel_i,
pci_irdy_i,
pci_par_i,
pci_perr_i,
pci_rst_i,
pci_rst_oe_o,
pci_stop_i,
pci_trdy_i,
wb_int_i,
wbm_ack_i,
wbm_dat_i_0_,
wbm_dat_i_10_,
wbm_dat_i_11_,
wbm_dat_i_12_,
wbm_dat_i_13_,
wbm_dat_i_14_,
wbm_dat_i_15_,
wbm_dat_i_16_,
wbm_dat_i_17_,
wbm_dat_i_18_,
wbm_dat_i_19_,
wbm_dat_i_1_,
wbm_dat_i_20_,
wbm_dat_i_21_,
wbm_dat_i_22_,
wbm_dat_i_23_,
wbm_dat_i_24_,
wbm_dat_i_25_,
wbm_dat_i_26_,
wbm_dat_i_27_,
wbm_dat_i_28_,
wbm_dat_i_29_,
wbm_dat_i_2_,
wbm_dat_i_30_,
wbm_dat_i_31_,
wbm_dat_i_3_,
wbm_dat_i_4_,
wbm_dat_i_5_,
wbm_dat_i_6_,
wbm_dat_i_7_,
wbm_dat_i_8_,
wbm_dat_i_9_,
wbm_err_i,
wbm_rty_i,
wbs_adr_i_0_,
wbs_adr_i_10_,
wbs_adr_i_11_,
wbs_adr_i_12_,
wbs_adr_i_13_,
wbs_adr_i_14_,
wbs_adr_i_15_,
wbs_adr_i_16_,
wbs_adr_i_17_,
wbs_adr_i_18_,
wbs_adr_i_19_,
wbs_adr_i_1_,
wbs_adr_i_20_,
wbs_adr_i_21_,
wbs_adr_i_22_,
wbs_adr_i_23_,
wbs_adr_i_24_,
wbs_adr_i_25_,
wbs_adr_i_26_,
wbs_adr_i_27_,
wbs_adr_i_28_,
wbs_adr_i_29_,
wbs_adr_i_2_,
wbs_adr_i_30_,
wbs_adr_i_31_,
wbs_adr_i_3_,
wbs_adr_i_4_,
wbs_adr_i_5_,
wbs_adr_i_6_,
wbs_adr_i_7_,
wbs_adr_i_8_,
wbs_adr_i_9_,
wbs_bte_i_0_,
wbs_bte_i_1_,
wbs_cti_i_0_,
wbs_cti_i_1_,
wbs_cti_i_2_,
wbs_cyc_i,
wbs_dat_i_0_,
wbs_dat_i_10_,
wbs_dat_i_11_,
wbs_dat_i_12_,
wbs_dat_i_13_,
wbs_dat_i_14_,
wbs_dat_i_15_,
wbs_dat_i_16_,
wbs_dat_i_17_,
wbs_dat_i_18_,
wbs_dat_i_19_,
wbs_dat_i_1_,
wbs_dat_i_20_,
wbs_dat_i_21_,
wbs_dat_i_22_,
wbs_dat_i_23_,
wbs_dat_i_24_,
wbs_dat_i_25_,
wbs_dat_i_26_,
wbs_dat_i_27_,
wbs_dat_i_28_,
wbs_dat_i_29_,
wbs_dat_i_2_,
wbs_dat_i_30_,
wbs_dat_i_31_,
wbs_dat_i_3_,
wbs_dat_i_4_,
wbs_dat_i_5_,
wbs_dat_i_6_,
wbs_dat_i_7_,
wbs_dat_i_8_,
wbs_dat_i_9_,
wbs_sel_i_0_,
wbs_sel_i_1_,
wbs_sel_i_2_,
wbs_sel_i_3_,
wbs_stb_i,
wbs_we_i,
pci_ad_o_0_,
pci_ad_o_10_,
pci_ad_o_11_,
pci_ad_o_12_,
pci_ad_o_13_,
pci_ad_o_14_,
pci_ad_o_15_,
pci_ad_o_16_,
pci_ad_o_17_,
pci_ad_o_18_,
pci_ad_o_19_,
pci_ad_o_1_,
pci_ad_o_20_,
pci_ad_o_21_,
pci_ad_o_22_,
pci_ad_o_23_,
pci_ad_o_24_,
pci_ad_o_25_,
pci_ad_o_26_,
pci_ad_o_27_,
pci_ad_o_28_,
pci_ad_o_29_,
pci_ad_o_2_,
pci_ad_o_30_,
pci_ad_o_31_,
pci_ad_o_3_,
pci_ad_o_4_,
pci_ad_o_5_,
pci_ad_o_6_,
pci_ad_o_7_,
pci_ad_o_8_,
pci_ad_o_9_,
pci_ad_oe_o_0_,
pci_ad_oe_o_10_,
pci_ad_oe_o_11_,
pci_ad_oe_o_12_,
pci_ad_oe_o_13_,
pci_ad_oe_o_14_,
pci_ad_oe_o_15_,
pci_ad_oe_o_16_,
pci_ad_oe_o_17_,
pci_ad_oe_o_18_,
pci_ad_oe_o_19_,
pci_ad_oe_o_1_,
pci_ad_oe_o_20_,
pci_ad_oe_o_21_,
pci_ad_oe_o_22_,
pci_ad_oe_o_23_,
pci_ad_oe_o_24_,
pci_ad_oe_o_25_,
pci_ad_oe_o_26_,
pci_ad_oe_o_27_,
pci_ad_oe_o_28_,
pci_ad_oe_o_29_,
pci_ad_oe_o_2_,
pci_ad_oe_o_30_,
pci_ad_oe_o_31_,
pci_ad_oe_o_3_,
pci_ad_oe_o_4_,
pci_ad_oe_o_5_,
pci_ad_oe_o_6_,
pci_ad_oe_o_7_,
pci_ad_oe_o_8_,
pci_ad_oe_o_9_,
pci_cbe_o_0_,
pci_cbe_o_1_,
pci_cbe_o_2_,
pci_cbe_o_3_,
pci_cbe_oe_o_0_,
pci_cbe_oe_o_1_,
pci_cbe_oe_o_2_,
pci_cbe_oe_o_3_,
pci_devsel_o,
pci_devsel_oe_o,
pci_frame_o,
pci_frame_oe_o,
pci_inta_oe_o,
pci_irdy_o,
pci_irdy_oe_o,
pci_par_o,
pci_par_oe_o,
pci_perr_o,
pci_perr_oe_o,
pci_req_o,
pci_req_oe_o,
pci_serr_o,
pci_serr_oe_o,
pci_stop_o,
pci_stop_oe_o,
pci_trdy_o,
pci_trdy_oe_o,
wb_rst_o,
wbm_adr_o_0_,
wbm_adr_o_10_,
wbm_adr_o_11_,
wbm_adr_o_12_,
wbm_adr_o_13_,
wbm_adr_o_14_,
wbm_adr_o_15_,
wbm_adr_o_16_,
wbm_adr_o_17_,
wbm_adr_o_18_,
wbm_adr_o_19_,
wbm_adr_o_1_,
wbm_adr_o_20_,
wbm_adr_o_21_,
wbm_adr_o_22_,
wbm_adr_o_23_,
wbm_adr_o_24_,
wbm_adr_o_25_,
wbm_adr_o_26_,
wbm_adr_o_27_,
wbm_adr_o_28_,
wbm_adr_o_29_,
wbm_adr_o_2_,
wbm_adr_o_30_,
wbm_adr_o_31_,
wbm_adr_o_3_,
wbm_adr_o_4_,
wbm_adr_o_5_,
wbm_adr_o_6_,
wbm_adr_o_7_,
wbm_adr_o_8_,
wbm_adr_o_9_,
wbm_cti_o_0_,
wbm_cti_o_1_,
wbm_cti_o_2_,
wbm_cyc_o,
wbm_dat_o_0_,
wbm_dat_o_10_,
wbm_dat_o_11_,
wbm_dat_o_12_,
wbm_dat_o_13_,
wbm_dat_o_14_,
wbm_dat_o_15_,
wbm_dat_o_16_,
wbm_dat_o_17_,
wbm_dat_o_18_,
wbm_dat_o_19_,
wbm_dat_o_1_,
wbm_dat_o_20_,
wbm_dat_o_21_,
wbm_dat_o_22_,
wbm_dat_o_23_,
wbm_dat_o_24_,
wbm_dat_o_25_,
wbm_dat_o_26_,
wbm_dat_o_27_,
wbm_dat_o_28_,
wbm_dat_o_29_,
wbm_dat_o_2_,
wbm_dat_o_30_,
wbm_dat_o_31_,
wbm_dat_o_3_,
wbm_dat_o_4_,
wbm_dat_o_5_,
wbm_dat_o_6_,
wbm_dat_o_7_,
wbm_dat_o_8_,
wbm_dat_o_9_,
wbm_sel_o_0_,
wbm_sel_o_1_,
wbm_sel_o_2_,
wbm_sel_o_3_,
wbm_stb_o,
wbm_we_o,
wbs_ack_o,
wbs_dat_o_0_,
wbs_dat_o_10_,
wbs_dat_o_11_,
wbs_dat_o_12_,
wbs_dat_o_13_,
wbs_dat_o_14_,
wbs_dat_o_15_,
wbs_dat_o_16_,
wbs_dat_o_17_,
wbs_dat_o_18_,
wbs_dat_o_19_,
wbs_dat_o_1_,
wbs_dat_o_20_,
wbs_dat_o_21_,
wbs_dat_o_22_,
wbs_dat_o_23_,
wbs_dat_o_24_,
wbs_dat_o_25_,
wbs_dat_o_26_,
wbs_dat_o_27_,
wbs_dat_o_28_,
wbs_dat_o_29_,
wbs_dat_o_2_,
wbs_dat_o_30_,
wbs_dat_o_31_,
wbs_dat_o_3_,
wbs_dat_o_4_,
wbs_dat_o_5_,
wbs_dat_o_6_,
wbs_dat_o_7_,
wbs_dat_o_8_,
wbs_dat_o_9_,
wbs_err_o,
wbs_rty_o
);

// Start PIs
input ispd_clk;
input pci_ad_i_0_;
input pci_ad_i_10_;
input pci_ad_i_11_;
input pci_ad_i_12_;
input pci_ad_i_13_;
input pci_ad_i_14_;
input pci_ad_i_15_;
input pci_ad_i_16_;
input pci_ad_i_17_;
input pci_ad_i_18_;
input pci_ad_i_19_;
input pci_ad_i_1_;
input pci_ad_i_20_;
input pci_ad_i_21_;
input pci_ad_i_22_;
input pci_ad_i_23_;
input pci_ad_i_24_;
input pci_ad_i_25_;
input pci_ad_i_26_;
input pci_ad_i_27_;
input pci_ad_i_28_;
input pci_ad_i_29_;
input pci_ad_i_2_;
input pci_ad_i_30_;
input pci_ad_i_31_;
input pci_ad_i_3_;
input pci_ad_i_4_;
input pci_ad_i_5_;
input pci_ad_i_6_;
input pci_ad_i_7_;
input pci_ad_i_8_;
input pci_ad_i_9_;
input pci_cbe_i_0_;
input pci_cbe_i_1_;
input pci_cbe_i_2_;
input pci_cbe_i_3_;
input pci_devsel_i;
input pci_frame_i;
input pci_gnt_i;
input pci_idsel_i;
input pci_irdy_i;
input pci_par_i;
input pci_perr_i;
input pci_rst_i;
input pci_rst_oe_o;
input pci_stop_i;
input pci_trdy_i;
input wb_int_i;
input wbm_ack_i;
input wbm_dat_i_0_;
input wbm_dat_i_10_;
input wbm_dat_i_11_;
input wbm_dat_i_12_;
input wbm_dat_i_13_;
input wbm_dat_i_14_;
input wbm_dat_i_15_;
input wbm_dat_i_16_;
input wbm_dat_i_17_;
input wbm_dat_i_18_;
input wbm_dat_i_19_;
input wbm_dat_i_1_;
input wbm_dat_i_20_;
input wbm_dat_i_21_;
input wbm_dat_i_22_;
input wbm_dat_i_23_;
input wbm_dat_i_24_;
input wbm_dat_i_25_;
input wbm_dat_i_26_;
input wbm_dat_i_27_;
input wbm_dat_i_28_;
input wbm_dat_i_29_;
input wbm_dat_i_2_;
input wbm_dat_i_30_;
input wbm_dat_i_31_;
input wbm_dat_i_3_;
input wbm_dat_i_4_;
input wbm_dat_i_5_;
input wbm_dat_i_6_;
input wbm_dat_i_7_;
input wbm_dat_i_8_;
input wbm_dat_i_9_;
input wbm_err_i;
input wbm_rty_i;
input wbs_adr_i_0_;
input wbs_adr_i_10_;
input wbs_adr_i_11_;
input wbs_adr_i_12_;
input wbs_adr_i_13_;
input wbs_adr_i_14_;
input wbs_adr_i_15_;
input wbs_adr_i_16_;
input wbs_adr_i_17_;
input wbs_adr_i_18_;
input wbs_adr_i_19_;
input wbs_adr_i_1_;
input wbs_adr_i_20_;
input wbs_adr_i_21_;
input wbs_adr_i_22_;
input wbs_adr_i_23_;
input wbs_adr_i_24_;
input wbs_adr_i_25_;
input wbs_adr_i_26_;
input wbs_adr_i_27_;
input wbs_adr_i_28_;
input wbs_adr_i_29_;
input wbs_adr_i_2_;
input wbs_adr_i_30_;
input wbs_adr_i_31_;
input wbs_adr_i_3_;
input wbs_adr_i_4_;
input wbs_adr_i_5_;
input wbs_adr_i_6_;
input wbs_adr_i_7_;
input wbs_adr_i_8_;
input wbs_adr_i_9_;
input wbs_bte_i_0_;
input wbs_bte_i_1_;
input wbs_cti_i_0_;
input wbs_cti_i_1_;
input wbs_cti_i_2_;
input wbs_cyc_i;
input wbs_dat_i_0_;
input wbs_dat_i_10_;
input wbs_dat_i_11_;
input wbs_dat_i_12_;
input wbs_dat_i_13_;
input wbs_dat_i_14_;
input wbs_dat_i_15_;
input wbs_dat_i_16_;
input wbs_dat_i_17_;
input wbs_dat_i_18_;
input wbs_dat_i_19_;
input wbs_dat_i_1_;
input wbs_dat_i_20_;
input wbs_dat_i_21_;
input wbs_dat_i_22_;
input wbs_dat_i_23_;
input wbs_dat_i_24_;
input wbs_dat_i_25_;
input wbs_dat_i_26_;
input wbs_dat_i_27_;
input wbs_dat_i_28_;
input wbs_dat_i_29_;
input wbs_dat_i_2_;
input wbs_dat_i_30_;
input wbs_dat_i_31_;
input wbs_dat_i_3_;
input wbs_dat_i_4_;
input wbs_dat_i_5_;
input wbs_dat_i_6_;
input wbs_dat_i_7_;
input wbs_dat_i_8_;
input wbs_dat_i_9_;
input wbs_sel_i_0_;
input wbs_sel_i_1_;
input wbs_sel_i_2_;
input wbs_sel_i_3_;
input wbs_stb_i;
input wbs_we_i;

// Start POs
output pci_ad_o_0_;
output pci_ad_o_10_;
output pci_ad_o_11_;
output pci_ad_o_12_;
output pci_ad_o_13_;
output pci_ad_o_14_;
output pci_ad_o_15_;
output pci_ad_o_16_;
output pci_ad_o_17_;
output pci_ad_o_18_;
output pci_ad_o_19_;
output pci_ad_o_1_;
output pci_ad_o_20_;
output pci_ad_o_21_;
output pci_ad_o_22_;
output pci_ad_o_23_;
output pci_ad_o_24_;
output pci_ad_o_25_;
output pci_ad_o_26_;
output pci_ad_o_27_;
output pci_ad_o_28_;
output pci_ad_o_29_;
output pci_ad_o_2_;
output pci_ad_o_30_;
output pci_ad_o_31_;
output pci_ad_o_3_;
output pci_ad_o_4_;
output pci_ad_o_5_;
output pci_ad_o_6_;
output pci_ad_o_7_;
output pci_ad_o_8_;
output pci_ad_o_9_;
output pci_ad_oe_o_0_;
output pci_ad_oe_o_10_;
output pci_ad_oe_o_11_;
output pci_ad_oe_o_12_;
output pci_ad_oe_o_13_;
output pci_ad_oe_o_14_;
output pci_ad_oe_o_15_;
output pci_ad_oe_o_16_;
output pci_ad_oe_o_17_;
output pci_ad_oe_o_18_;
output pci_ad_oe_o_19_;
output pci_ad_oe_o_1_;
output pci_ad_oe_o_20_;
output pci_ad_oe_o_21_;
output pci_ad_oe_o_22_;
output pci_ad_oe_o_23_;
output pci_ad_oe_o_24_;
output pci_ad_oe_o_25_;
output pci_ad_oe_o_26_;
output pci_ad_oe_o_27_;
output pci_ad_oe_o_28_;
output pci_ad_oe_o_29_;
output pci_ad_oe_o_2_;
output pci_ad_oe_o_30_;
output pci_ad_oe_o_31_;
output pci_ad_oe_o_3_;
output pci_ad_oe_o_4_;
output pci_ad_oe_o_5_;
output pci_ad_oe_o_6_;
output pci_ad_oe_o_7_;
output pci_ad_oe_o_8_;
output pci_ad_oe_o_9_;
output pci_cbe_o_0_;
output pci_cbe_o_1_;
output pci_cbe_o_2_;
output pci_cbe_o_3_;
output pci_cbe_oe_o_0_;
output pci_cbe_oe_o_1_;
output pci_cbe_oe_o_2_;
output pci_cbe_oe_o_3_;
output pci_devsel_o;
output pci_devsel_oe_o;
output pci_frame_o;
output pci_frame_oe_o;
output pci_inta_oe_o;
output pci_irdy_o;
output pci_irdy_oe_o;
output pci_par_o;
output pci_par_oe_o;
output pci_perr_o;
output pci_perr_oe_o;
output pci_req_o;
output pci_req_oe_o;
output pci_serr_o;
output pci_serr_oe_o;
output pci_stop_o;
output pci_stop_oe_o;
output pci_trdy_o;
output pci_trdy_oe_o;
output wb_rst_o;
output wbm_adr_o_0_;
output wbm_adr_o_10_;
output wbm_adr_o_11_;
output wbm_adr_o_12_;
output wbm_adr_o_13_;
output wbm_adr_o_14_;
output wbm_adr_o_15_;
output wbm_adr_o_16_;
output wbm_adr_o_17_;
output wbm_adr_o_18_;
output wbm_adr_o_19_;
output wbm_adr_o_1_;
output wbm_adr_o_20_;
output wbm_adr_o_21_;
output wbm_adr_o_22_;
output wbm_adr_o_23_;
output wbm_adr_o_24_;
output wbm_adr_o_25_;
output wbm_adr_o_26_;
output wbm_adr_o_27_;
output wbm_adr_o_28_;
output wbm_adr_o_29_;
output wbm_adr_o_2_;
output wbm_adr_o_30_;
output wbm_adr_o_31_;
output wbm_adr_o_3_;
output wbm_adr_o_4_;
output wbm_adr_o_5_;
output wbm_adr_o_6_;
output wbm_adr_o_7_;
output wbm_adr_o_8_;
output wbm_adr_o_9_;
output wbm_cti_o_0_;
output wbm_cti_o_1_;
output wbm_cti_o_2_;
output wbm_cyc_o;
output wbm_dat_o_0_;
output wbm_dat_o_10_;
output wbm_dat_o_11_;
output wbm_dat_o_12_;
output wbm_dat_o_13_;
output wbm_dat_o_14_;
output wbm_dat_o_15_;
output wbm_dat_o_16_;
output wbm_dat_o_17_;
output wbm_dat_o_18_;
output wbm_dat_o_19_;
output wbm_dat_o_1_;
output wbm_dat_o_20_;
output wbm_dat_o_21_;
output wbm_dat_o_22_;
output wbm_dat_o_23_;
output wbm_dat_o_24_;
output wbm_dat_o_25_;
output wbm_dat_o_26_;
output wbm_dat_o_27_;
output wbm_dat_o_28_;
output wbm_dat_o_29_;
output wbm_dat_o_2_;
output wbm_dat_o_30_;
output wbm_dat_o_31_;
output wbm_dat_o_3_;
output wbm_dat_o_4_;
output wbm_dat_o_5_;
output wbm_dat_o_6_;
output wbm_dat_o_7_;
output wbm_dat_o_8_;
output wbm_dat_o_9_;
output wbm_sel_o_0_;
output wbm_sel_o_1_;
output wbm_sel_o_2_;
output wbm_sel_o_3_;
output wbm_stb_o;
output wbm_we_o;
output wbs_ack_o;
output wbs_dat_o_0_;
output wbs_dat_o_10_;
output wbs_dat_o_11_;
output wbs_dat_o_12_;
output wbs_dat_o_13_;
output wbs_dat_o_14_;
output wbs_dat_o_15_;
output wbs_dat_o_16_;
output wbs_dat_o_17_;
output wbs_dat_o_18_;
output wbs_dat_o_19_;
output wbs_dat_o_1_;
output wbs_dat_o_20_;
output wbs_dat_o_21_;
output wbs_dat_o_22_;
output wbs_dat_o_23_;
output wbs_dat_o_24_;
output wbs_dat_o_25_;
output wbs_dat_o_26_;
output wbs_dat_o_27_;
output wbs_dat_o_28_;
output wbs_dat_o_29_;
output wbs_dat_o_2_;
output wbs_dat_o_30_;
output wbs_dat_o_31_;
output wbs_dat_o_3_;
output wbs_dat_o_4_;
output wbs_dat_o_5_;
output wbs_dat_o_6_;
output wbs_dat_o_7_;
output wbs_dat_o_8_;
output wbs_dat_o_9_;
output wbs_err_o;
output wbs_rty_o;

// Start wires
wire ispd_clk;
wire pci_ad_i_0_;
wire pci_ad_i_10_;
wire pci_ad_i_11_;
wire pci_ad_i_12_;
wire pci_ad_i_13_;
wire pci_ad_i_14_;
wire pci_ad_i_15_;
wire pci_ad_i_16_;
wire pci_ad_i_17_;
wire pci_ad_i_18_;
wire pci_ad_i_19_;
wire pci_ad_i_1_;
wire pci_ad_i_20_;
wire pci_ad_i_21_;
wire pci_ad_i_22_;
wire pci_ad_i_23_;
wire pci_ad_i_24_;
wire pci_ad_i_25_;
wire pci_ad_i_26_;
wire pci_ad_i_27_;
wire pci_ad_i_28_;
wire pci_ad_i_29_;
wire pci_ad_i_2_;
wire pci_ad_i_30_;
wire pci_ad_i_31_;
wire pci_ad_i_3_;
wire pci_ad_i_4_;
wire pci_ad_i_5_;
wire pci_ad_i_6_;
wire pci_ad_i_7_;
wire pci_ad_i_8_;
wire pci_ad_i_9_;
wire pci_cbe_i_0_;
wire pci_cbe_i_1_;
wire pci_cbe_i_2_;
wire pci_cbe_i_3_;
wire pci_devsel_i;
wire pci_frame_i;
wire pci_gnt_i;
wire pci_idsel_i;
wire pci_irdy_i;
wire pci_par_i;
wire pci_perr_i;
wire pci_rst_i;
wire pci_rst_oe_o;
wire pci_stop_i;
wire pci_trdy_i;
wire wb_int_i;
wire wbm_ack_i;
wire wbm_dat_i_0_;
wire wbm_dat_i_10_;
wire wbm_dat_i_11_;
wire wbm_dat_i_12_;
wire wbm_dat_i_13_;
wire wbm_dat_i_14_;
wire wbm_dat_i_15_;
wire wbm_dat_i_16_;
wire wbm_dat_i_17_;
wire wbm_dat_i_18_;
wire wbm_dat_i_19_;
wire wbm_dat_i_1_;
wire wbm_dat_i_20_;
wire wbm_dat_i_21_;
wire wbm_dat_i_22_;
wire wbm_dat_i_23_;
wire wbm_dat_i_24_;
wire wbm_dat_i_25_;
wire wbm_dat_i_26_;
wire wbm_dat_i_27_;
wire wbm_dat_i_28_;
wire wbm_dat_i_29_;
wire wbm_dat_i_2_;
wire wbm_dat_i_30_;
wire wbm_dat_i_31_;
wire wbm_dat_i_3_;
wire wbm_dat_i_4_;
wire wbm_dat_i_5_;
wire wbm_dat_i_6_;
wire wbm_dat_i_7_;
wire wbm_dat_i_8_;
wire wbm_dat_i_9_;
wire wbm_err_i;
wire wbm_rty_i;
wire wbs_adr_i_0_;
wire wbs_adr_i_10_;
wire wbs_adr_i_11_;
wire wbs_adr_i_12_;
wire wbs_adr_i_13_;
wire wbs_adr_i_14_;
wire wbs_adr_i_15_;
wire wbs_adr_i_16_;
wire wbs_adr_i_17_;
wire wbs_adr_i_18_;
wire wbs_adr_i_19_;
wire wbs_adr_i_1_;
wire wbs_adr_i_20_;
wire wbs_adr_i_21_;
wire wbs_adr_i_22_;
wire wbs_adr_i_23_;
wire wbs_adr_i_24_;
wire wbs_adr_i_25_;
wire wbs_adr_i_26_;
wire wbs_adr_i_27_;
wire wbs_adr_i_28_;
wire wbs_adr_i_29_;
wire wbs_adr_i_2_;
wire wbs_adr_i_30_;
wire wbs_adr_i_31_;
wire wbs_adr_i_3_;
wire wbs_adr_i_4_;
wire wbs_adr_i_5_;
wire wbs_adr_i_6_;
wire wbs_adr_i_7_;
wire wbs_adr_i_8_;
wire wbs_adr_i_9_;
wire wbs_bte_i_0_;
wire wbs_bte_i_1_;
wire wbs_cti_i_0_;
wire wbs_cti_i_1_;
wire wbs_cti_i_2_;
wire wbs_cyc_i;
wire wbs_dat_i_0_;
wire wbs_dat_i_10_;
wire wbs_dat_i_11_;
wire wbs_dat_i_12_;
wire wbs_dat_i_13_;
wire wbs_dat_i_14_;
wire wbs_dat_i_15_;
wire wbs_dat_i_16_;
wire wbs_dat_i_17_;
wire wbs_dat_i_18_;
wire wbs_dat_i_19_;
wire wbs_dat_i_1_;
wire wbs_dat_i_20_;
wire wbs_dat_i_21_;
wire wbs_dat_i_22_;
wire wbs_dat_i_23_;
wire wbs_dat_i_24_;
wire wbs_dat_i_25_;
wire wbs_dat_i_26_;
wire wbs_dat_i_27_;
wire wbs_dat_i_28_;
wire wbs_dat_i_29_;
wire wbs_dat_i_2_;
wire wbs_dat_i_30_;
wire wbs_dat_i_31_;
wire wbs_dat_i_3_;
wire wbs_dat_i_4_;
wire wbs_dat_i_5_;
wire wbs_dat_i_6_;
wire wbs_dat_i_7_;
wire wbs_dat_i_8_;
wire wbs_dat_i_9_;
wire wbs_sel_i_0_;
wire wbs_sel_i_1_;
wire wbs_sel_i_2_;
wire wbs_sel_i_3_;
wire wbs_stb_i;
wire wbs_we_i;
wire pci_ad_o_0_;
wire pci_ad_o_10_;
wire pci_ad_o_11_;
wire pci_ad_o_12_;
wire pci_ad_o_13_;
wire pci_ad_o_14_;
wire pci_ad_o_15_;
wire pci_ad_o_16_;
wire pci_ad_o_17_;
wire pci_ad_o_18_;
wire pci_ad_o_19_;
wire pci_ad_o_1_;
wire pci_ad_o_20_;
wire pci_ad_o_21_;
wire pci_ad_o_22_;
wire pci_ad_o_23_;
wire pci_ad_o_24_;
wire pci_ad_o_25_;
wire pci_ad_o_26_;
wire pci_ad_o_27_;
wire pci_ad_o_28_;
wire pci_ad_o_29_;
wire pci_ad_o_2_;
wire pci_ad_o_30_;
wire pci_ad_o_31_;
wire pci_ad_o_3_;
wire pci_ad_o_4_;
wire pci_ad_o_5_;
wire pci_ad_o_6_;
wire pci_ad_o_7_;
wire pci_ad_o_8_;
wire pci_ad_o_9_;
wire pci_ad_oe_o_0_;
wire pci_ad_oe_o_10_;
wire pci_ad_oe_o_11_;
wire pci_ad_oe_o_12_;
wire pci_ad_oe_o_13_;
wire pci_ad_oe_o_14_;
wire pci_ad_oe_o_15_;
wire pci_ad_oe_o_16_;
wire pci_ad_oe_o_17_;
wire pci_ad_oe_o_18_;
wire pci_ad_oe_o_19_;
wire pci_ad_oe_o_1_;
wire pci_ad_oe_o_20_;
wire pci_ad_oe_o_21_;
wire pci_ad_oe_o_22_;
wire pci_ad_oe_o_23_;
wire pci_ad_oe_o_24_;
wire pci_ad_oe_o_25_;
wire pci_ad_oe_o_26_;
wire pci_ad_oe_o_27_;
wire pci_ad_oe_o_28_;
wire pci_ad_oe_o_29_;
wire pci_ad_oe_o_2_;
wire pci_ad_oe_o_30_;
wire pci_ad_oe_o_31_;
wire pci_ad_oe_o_3_;
wire pci_ad_oe_o_4_;
wire pci_ad_oe_o_5_;
wire pci_ad_oe_o_6_;
wire pci_ad_oe_o_7_;
wire pci_ad_oe_o_8_;
wire pci_ad_oe_o_9_;
wire pci_cbe_o_0_;
wire pci_cbe_o_1_;
wire pci_cbe_o_2_;
wire pci_cbe_o_3_;
wire pci_cbe_oe_o_0_;
wire pci_cbe_oe_o_1_;
wire pci_cbe_oe_o_2_;
wire pci_cbe_oe_o_3_;
wire pci_devsel_o;
wire pci_devsel_oe_o;
wire pci_frame_o;
wire pci_frame_oe_o;
wire pci_inta_oe_o;
wire pci_irdy_o;
wire pci_irdy_oe_o;
wire pci_par_o;
wire pci_par_oe_o;
wire pci_perr_o;
wire pci_perr_oe_o;
wire pci_req_o;
wire pci_req_oe_o;
wire pci_serr_o;
wire pci_serr_oe_o;
wire pci_stop_o;
wire pci_stop_oe_o;
wire pci_trdy_o;
wire pci_trdy_oe_o;
wire wb_rst_o;
wire wbm_adr_o_0_;
wire wbm_adr_o_10_;
wire wbm_adr_o_11_;
wire wbm_adr_o_12_;
wire wbm_adr_o_13_;
wire wbm_adr_o_14_;
wire wbm_adr_o_15_;
wire wbm_adr_o_16_;
wire wbm_adr_o_17_;
wire wbm_adr_o_18_;
wire wbm_adr_o_19_;
wire wbm_adr_o_1_;
wire wbm_adr_o_20_;
wire wbm_adr_o_21_;
wire wbm_adr_o_22_;
wire wbm_adr_o_23_;
wire wbm_adr_o_24_;
wire wbm_adr_o_25_;
wire wbm_adr_o_26_;
wire wbm_adr_o_27_;
wire wbm_adr_o_28_;
wire wbm_adr_o_29_;
wire wbm_adr_o_2_;
wire wbm_adr_o_30_;
wire wbm_adr_o_31_;
wire wbm_adr_o_3_;
wire wbm_adr_o_4_;
wire wbm_adr_o_5_;
wire wbm_adr_o_6_;
wire wbm_adr_o_7_;
wire wbm_adr_o_8_;
wire wbm_adr_o_9_;
wire wbm_cti_o_0_;
wire wbm_cti_o_1_;
wire wbm_cti_o_2_;
wire wbm_cyc_o;
wire wbm_dat_o_0_;
wire wbm_dat_o_10_;
wire wbm_dat_o_11_;
wire wbm_dat_o_12_;
wire wbm_dat_o_13_;
wire wbm_dat_o_14_;
wire wbm_dat_o_15_;
wire wbm_dat_o_16_;
wire wbm_dat_o_17_;
wire wbm_dat_o_18_;
wire wbm_dat_o_19_;
wire wbm_dat_o_1_;
wire wbm_dat_o_20_;
wire wbm_dat_o_21_;
wire wbm_dat_o_22_;
wire wbm_dat_o_23_;
wire wbm_dat_o_24_;
wire wbm_dat_o_25_;
wire wbm_dat_o_26_;
wire wbm_dat_o_27_;
wire wbm_dat_o_28_;
wire wbm_dat_o_29_;
wire wbm_dat_o_2_;
wire wbm_dat_o_30_;
wire wbm_dat_o_31_;
wire wbm_dat_o_3_;
wire wbm_dat_o_4_;
wire wbm_dat_o_5_;
wire wbm_dat_o_6_;
wire wbm_dat_o_7_;
wire wbm_dat_o_8_;
wire wbm_dat_o_9_;
wire wbm_sel_o_0_;
wire wbm_sel_o_1_;
wire wbm_sel_o_2_;
wire wbm_sel_o_3_;
wire wbm_stb_o;
wire wbm_we_o;
wire wbs_ack_o;
wire wbs_dat_o_0_;
wire wbs_dat_o_10_;
wire wbs_dat_o_11_;
wire wbs_dat_o_12_;
wire wbs_dat_o_13_;
wire wbs_dat_o_14_;
wire wbs_dat_o_15_;
wire wbs_dat_o_16_;
wire wbs_dat_o_17_;
wire wbs_dat_o_18_;
wire wbs_dat_o_19_;
wire wbs_dat_o_1_;
wire wbs_dat_o_20_;
wire wbs_dat_o_21_;
wire wbs_dat_o_22_;
wire wbs_dat_o_23_;
wire wbs_dat_o_24_;
wire wbs_dat_o_25_;
wire wbs_dat_o_26_;
wire wbs_dat_o_27_;
wire wbs_dat_o_28_;
wire wbs_dat_o_29_;
wire wbs_dat_o_2_;
wire wbs_dat_o_30_;
wire wbs_dat_o_31_;
wire wbs_dat_o_3_;
wire wbs_dat_o_4_;
wire wbs_dat_o_5_;
wire wbs_dat_o_6_;
wire wbs_dat_o_7_;
wire wbs_dat_o_8_;
wire wbs_dat_o_9_;
wire wbs_err_o;
wire wbs_rty_o;
wire FE_OCPN1822_n_16560;
wire FE_OCPN1823_n_16560;
wire FE_OCPN1824_n_12030;
wire FE_OCPN1825_n_12030;
wire FE_OCPN1827_n_14995;
wire FE_OCPN1831_n_16949;
wire FE_OCPN1832_n_16949;
wire FE_OCPN1833_n_11884;
wire FE_OCPN1834_n_11884;
wire FE_OCPN1835_n_16798;
wire FE_OCPN1836_n_16798;
wire FE_OCPN1837_n_1238;
wire FE_OCPN1838_n_1238;
wire FE_OCPN1839_n_1238;
wire FE_OCPN1840_n_16089;
wire FE_OCPN1841_n_16089;
wire FE_OCPN1842_n_16033;
wire FE_OCPN1843_n_16033;
wire FE_OCPN1844_n_16427;
wire FE_OCPN1845_n_16427;
wire FE_OCPN1846_n_14981;
wire FE_OCPN1847_n_14981;
wire FE_OCPN1848_n_15998;
wire FE_OCPN1849_n_15998;
wire FE_OCPN1850_n_15998;
wire FE_OCPN1851_n_16538;
wire FE_OCPN1852_n_16538;
wire FE_OCPN1853_n_2071;
wire FE_OCPN1854_n_2071;
wire FE_OCPN1855_n_2071;
wire FE_OCPN1856_FE_OFN1774_n_13800;
wire FE_OCPN1860_FE_OFN468_n_15534;
wire FE_OCPN1861_FE_OFN468_n_15534;
wire FE_OCPN1862_FE_OFN474_n_16992;
wire FE_OCPN1863_FE_OFN474_n_16992;
wire FE_OCPN1865_n_12377;
wire FE_OCPN1866_n_12377;
wire FE_OCPN1868_n_16289;
wire FE_OCPN1871_FE_OFN474_n_16992;
wire FE_OCPN1872_FE_OFN474_n_16992;
wire FE_OCPN1873_FE_OFN474_n_16992;
wire FE_OCPN1875_n_14526;
wire FE_OCPN1876_n_13903;
wire FE_OCPN1877_n_13903;
wire FE_OCPN1878_FE_OFN470_n_10588;
wire FE_OCPN1879_FE_OFN470_n_10588;
wire FE_OCPN1880_n_9991;
wire FE_OCPN1881_n_9991;
wire FE_OCPN1882_n_9991;
wire FE_OCPN1883_n_15566;
wire FE_OCPN1884_n_15566;
wire FE_OCPN1885_FE_OFN1508_n_15587;
wire FE_OCPN1886_FE_OFN1508_n_15587;
wire FE_OCPN1887_FE_OFN473_n_16992;
wire FE_OCPN1888_FE_OFN473_n_16992;
wire FE_OCPN1889_n_16553;
wire FE_OCPN1890_n_16553;
wire FE_OCPN1891_FE_OFN1727_n_9975;
wire FE_OCPN1892_FE_OFN1727_n_9975;
wire FE_OCPN1895_FE_OFN1559_n_12042;
wire FE_OCPN1897_n_3231;
wire FE_OCPN1898_n_3231;
wire FE_OCPN1899_n_16810;
wire FE_OCPN1900_n_16810;
wire FE_OCPN1901_n_16810;
wire FE_OCPN1902_FE_OFN1061_n_16720;
wire FE_OCPN1903_FE_OFN1061_n_16720;
wire FE_OCPN1904_n_8927;
wire FE_OCPN1905_n_8927;
wire FE_OCPN1907_n_11767;
wire FE_OCPN1908_n_16497;
wire FE_OCPN1909_n_16497;
wire FE_OCPN1910_FE_OFN1152_n_13249;
wire FE_OCPN1911_FE_OFN1152_n_13249;
wire FE_OCPN1912_FE_OFN1150_n_13249;
wire FE_OCPN1913_FE_OFN1150_n_13249;
wire FE_OCPN1914_FE_OFN1522_n_10892;
wire FE_OCPN1915_FE_OFN1522_n_10892;
wire FE_OCPN2014_n_10195;
wire FE_OCPN2015_n_10195;
wire FE_OCPN2217_n_13997;
wire FE_OCPN2218_n_13997;
wire FE_OCPN2219_n_13997;
wire FE_OCPUNCON1951_FE_OFN697_n_16760;
wire FE_OCPUNCON1952_FE_OFN697_n_16760;
wire FE_OCP_DRV_N1949_n_8660;
wire FE_OCP_DRV_N1950_n_8660;
wire FE_OCP_DRV_N2261_n_8660;
wire FE_OCP_DRV_N2262_n_8660;
wire FE_OCP_RBN1917_wbs_cti_i_1_;
wire FE_OCP_RBN1918_wbs_cti_i_1_;
wire FE_OCP_RBN1921_n_10273;
wire FE_OCP_RBN1922_n_10273;
wire FE_OCP_RBN1923_n_10273;
wire FE_OCP_RBN1924_n_10273;
wire FE_OCP_RBN1925_n_10259;
wire FE_OCP_RBN1926_n_10259;
wire FE_OCP_RBN1927_n_10259;
wire FE_OCP_RBN1928_n_10259;
wire FE_OCP_RBN1929_parchk_pci_trdy_reg_in;
wire FE_OCP_RBN1930_parchk_pci_trdy_reg_in;
wire FE_OCP_RBN1932_FE_OFN1515_n_10538;
wire FE_OCP_RBN1933_FE_OFN1515_n_10538;
wire FE_OCP_RBN1934_FE_OFN1515_n_10538;
wire FE_OCP_RBN1954_FE_RN_462_0;
wire FE_OCP_RBN1955_n_16981;
wire FE_OCP_RBN1956_n_16981;
wire FE_OCP_RBN1961_FE_OFN1591_n_13741;
wire FE_OCP_RBN1962_FE_OFN1591_n_13741;
wire FE_OCP_RBN1963_FE_OFN1591_n_13741;
wire FE_OCP_RBN1964_FE_OFN1591_n_13741;
wire FE_OCP_RBN1965_FE_RN_459_0;
wire FE_OCP_RBN1966_FE_RN_459_0;
wire FE_OCP_RBN1967_FE_RN_459_0;
wire FE_OCP_RBN1968_FE_OFN1532_n_10143;
wire FE_OCP_RBN1969_FE_OFN1532_n_10143;
wire FE_OCP_RBN1970_n_11767;
wire FE_OCP_RBN1971_n_11767;
wire FE_OCP_RBN1972_n_11767;
wire FE_OCP_RBN1973_n_12381;
wire FE_OCP_RBN1974_n_12381;
wire FE_OCP_RBN1975_n_12381;
wire FE_OCP_RBN1976_n_12381;
wire FE_OCP_RBN1977_n_10273;
wire FE_OCP_RBN1978_n_10273;
wire FE_OCP_RBN1979_n_10273;
wire FE_OCP_RBN1980_n_10273;
wire FE_OCP_RBN1981_FE_OFN1591_n_13741;
wire FE_OCP_RBN1983_FE_OFN1591_n_13741;
wire FE_OCP_RBN1984_FE_OFN1591_n_13741;
wire FE_OCP_RBN1985_FE_OFN1591_n_13741;
wire FE_OCP_RBN1994_n_13971;
wire FE_OCP_RBN1995_n_13971;
wire FE_OCP_RBN1996_n_13971;
wire FE_OCP_RBN1997_n_13971;
wire FE_OCP_RBN1998_n_13971;
wire FE_OCP_RBN1999_n_13971;
wire FE_OCP_RBN2000_n_1403;
wire FE_OCP_RBN2003_FE_OFN1026_n_16760;
wire FE_OCP_RBN2004_FE_OFN1026_n_16760;
wire FE_OCP_RBN2005_FE_RN_459_0;
wire FE_OCP_RBN2006_FE_RN_459_0;
wire FE_OCP_RBN2007_n_16698;
wire FE_OCP_RBN2008_n_16698;
wire FE_OCP_RBN2009_n_16698;
wire FE_OCP_RBN2010_n_16698;
wire FE_OCP_RBN2011_n_16698;
wire FE_OCP_RBN2012_n_16698;
wire FE_OCP_RBN2013_FE_OCPN1895_FE_OFN1559_n_12042;
wire FE_OCP_RBN2016_n_16970;
wire FE_OCP_RBN2017_n_16970;
wire FE_OCP_RBN2018_n_16970;
wire FE_OCP_RBN2019_n_16970;
wire FE_OCP_RBN2220_n_15347;
wire FE_OCP_RBN2221_n_15347;
wire FE_OCP_RBN2222_n_15347;
wire FE_OCP_RBN2223_n_15347;
wire FE_OCP_RBN2224_n_16322;
wire FE_OCP_RBN2225_n_16322;
wire FE_OCP_RBN2226_g75174_p;
wire FE_OCP_RBN2227_g75174_p;
wire FE_OCP_RBN2228_n_15969;
wire FE_OCP_RBN2229_n_15969;
wire FE_OCP_RBN2231_FE_RN_390_0;
wire FE_OCP_RBN2232_n_16273;
wire FE_OCP_RBN2233_n_16273;
wire FE_OCP_RBN2237_g74749_p;
wire FE_OCP_RBN2238_g74749_p;
wire FE_OCP_RBN2239_g74749_p;
wire FE_OCP_RBN2265_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_;
wire FE_OCP_RBN2269_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_;
wire FE_OCP_RBN2270_g75061_p;
wire FE_OCP_RBN2271_g75061_p;
wire FE_OCP_RBN2272_n_10268;
wire FE_OCP_RBN2273_n_10268;
wire FE_OCP_RBN2274_n_10268;
wire FE_OCP_RBN2275_n_10268;
wire FE_OCP_RBN2277_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_;
wire FE_OCP_RBN2278_n_16974;
wire FE_OCP_RBN2279_n_16974;
wire FE_OCP_RBN2280_g74996_p;
wire FE_OCP_RBN2281_g74996_p;
wire FE_OCP_RBN2282_g74996_p;
wire FE_OCP_RBN2283_g74996_p;
wire FE_OCP_RBN2284_FE_RN_494_0;
wire FE_OCP_RBN2285_FE_RN_494_0;
wire FE_OCP_RBN2286_FE_RN_494_0;
wire FE_OCP_RBN2289_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_;
wire FE_OCP_RBN2290_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_;
wire FE_OCP_RBN2291_FE_OFN1575_n_12028;
wire FE_OCP_RBN2292_FE_OFN1575_n_12028;
wire FE_OCP_RBN2293_FE_OFN1581_n_12306;
wire FE_OFN1000_n_15978;
wire FE_OFN1001_n_15978;
wire FE_OFN1002_n_2047;
wire FE_OFN1003_n_2047;
wire FE_OFN1004_n_16288;
wire FE_OFN1005_n_16288;
wire FE_OFN1006_n_16288;
wire FE_OFN1007_n_4734;
wire FE_OFN1008_n_4734;
wire FE_OFN1009_n_4734;
wire FE_OFN1010_n_4734;
wire FE_OFN1011_n_4734;
wire FE_OFN1012_n_4734;
wire FE_OFN1013_n_4734;
wire FE_OFN1014_n_2053;
wire FE_OFN1015_n_2053;
wire FE_OFN1016_n_2053;
wire FE_OFN1017_n_2053;
wire FE_OFN1018_n_11877;
wire FE_OFN1019_n_11877;
wire FE_OFN1020_n_11877;
wire FE_OFN1021_n_11877;
wire FE_OFN1022_n_11877;
wire FE_OFN1023_n_11877;
wire FE_OFN1024_n_11877;
wire FE_OFN1025_n_11877;
wire FE_OFN1026_n_16760;
wire FE_OFN1028_n_4732;
wire FE_OFN1029_n_4732;
wire FE_OFN1030_n_4732;
wire FE_OFN1031_n_4732;
wire FE_OFN1032_n_4732;
wire FE_OFN1033_n_4732;
wire FE_OFN1034_n_4732;
wire FE_OFN1035_n_4732;
wire FE_OFN1036_n_4732;
wire FE_OFN1037_n_4732;
wire FE_OFN1038_n_2037;
wire FE_OFN1039_n_2037;
wire FE_OFN1040_n_2037;
wire FE_OFN1041_n_2037;
wire FE_OFN1042_n_2037;
wire FE_OFN1043_n_2037;
wire FE_OFN1044_n_2037;
wire FE_OFN1045_n_16657;
wire FE_OFN1046_n_16657;
wire FE_OFN1047_n_16657;
wire FE_OFN1048_n_16657;
wire FE_OFN1049_n_16657;
wire FE_OFN1050_n_16657;
wire FE_OFN1051_n_16657;
wire FE_OFN1052_n_4727;
wire FE_OFN1053_n_4727;
wire FE_OFN1054_n_4727;
wire FE_OFN1055_n_4727;
wire FE_OFN1056_n_4727;
wire FE_OFN1057_n_4727;
wire FE_OFN1058_n_4727;
wire FE_OFN1059_n_4727;
wire FE_OFN1060_n_16720;
wire FE_OFN1061_n_16720;
wire FE_OFN1062_n_15808;
wire FE_OFN1063_n_15808;
wire FE_OFN1064_n_15808;
wire FE_OFN1065_n_15808;
wire FE_OFN1066_n_15808;
wire FE_OFN1067_n_15729;
wire FE_OFN1068_n_15729;
wire FE_OFN1069_n_15729;
wire FE_OFN1070_n_15729;
wire FE_OFN1071_n_15729;
wire FE_OFN1072_n_4740;
wire FE_OFN1073_n_4740;
wire FE_OFN1074_n_4740;
wire FE_OFN1075_n_4740;
wire FE_OFN1076_n_4740;
wire FE_OFN1077_n_4740;
wire FE_OFN1078_n_4778;
wire FE_OFN1079_n_4778;
wire FE_OFN1080_n_13221;
wire FE_OFN1081_n_13221;
wire FE_OFN1082_n_13221;
wire FE_OFN1083_n_13221;
wire FE_OFN1084_n_13221;
wire FE_OFN1085_n_13221;
wire FE_OFN1086_g64577_p;
wire FE_OFN1087_g64577_p;
wire FE_OFN1088_g64577_p;
wire FE_OFN1089_g64577_p;
wire FE_OFN1090_g64577_p;
wire FE_OFN1091_g64577_p;
wire FE_OFN1092_g64577_p;
wire FE_OFN1093_g64577_p;
wire FE_OFN1094_g64577_p;
wire FE_OFN1095_g64577_p;
wire FE_OFN1096_g64577_p;
wire FE_OFN1097_g64577_p;
wire FE_OFN1098_g64577_p;
wire FE_OFN1099_g64577_p;
wire FE_OFN1100_g64577_p;
wire FE_OFN1101_g64577_p;
wire FE_OFN1102_g64577_p;
wire FE_OFN1103_g64577_p;
wire FE_OFN1104_g64577_p;
wire FE_OFN1105_g64577_p;
wire FE_OFN1106_g64577_p;
wire FE_OFN1107_g64577_p;
wire FE_OFN1108_g64577_p;
wire FE_OFN1109_g64577_p;
wire FE_OFN1110_g64577_p;
wire FE_OFN1111_g64577_p;
wire FE_OFN1112_g64577_p;
wire FE_OFN1113_g64577_p;
wire FE_OFN1114_g64577_p;
wire FE_OFN1115_g64577_p;
wire FE_OFN1116_g64577_p;
wire FE_OFN1117_g64577_p;
wire FE_OFN1118_g64577_p;
wire FE_OFN1119_g64577_p;
wire FE_OFN1120_g64577_p;
wire FE_OFN1121_g64577_p;
wire FE_OFN1122_g64577_p;
wire FE_OFN1123_g64577_p;
wire FE_OFN1124_g64577_p;
wire FE_OFN1125_g64577_p;
wire FE_OFN1126_g64577_p;
wire FE_OFN1127_g64577_p;
wire FE_OFN1128_g64577_p;
wire FE_OFN1129_g64577_p;
wire FE_OFN1130_g64577_p;
wire FE_OFN1131_g64577_p;
wire FE_OFN1132_g64577_p;
wire FE_OFN1133_g64577_p;
wire FE_OFN1134_g64577_p;
wire FE_OFN1135_g64577_p;
wire FE_OFN1136_g64577_p;
wire FE_OFN1137_g64577_p;
wire FE_OFN1138_g64577_p;
wire FE_OFN1139_g64577_p;
wire FE_OFN1140_g64577_p;
wire FE_OFN1141_n_15261;
wire FE_OFN1142_n_15261;
wire FE_OFN1143_n_15261;
wire FE_OFN1144_n_15261;
wire FE_OFN1145_n_15261;
wire FE_OFN1146_n_13249;
wire FE_OFN1147_n_13249;
wire FE_OFN1148_n_13249;
wire FE_OFN1149_n_13249;
wire FE_OFN1150_n_13249;
wire FE_OFN1151_n_13249;
wire FE_OFN1152_n_13249;
wire FE_OFN1153_n_3464;
wire FE_OFN1154_n_3464;
wire FE_OFN1155_n_3464;
wire FE_OFN1156_n_7498;
wire FE_OFN1157_n_15325;
wire FE_OFN1158_n_15325;
wire FE_OFN1159_n_15325;
wire FE_OFN1160_n_5615;
wire FE_OFN1161_n_5615;
wire FE_OFN1162_n_5615;
wire FE_OFN1163_n_5615;
wire FE_OFN1164_n_5615;
wire FE_OFN1165_n_5615;
wire FE_OFN1166_n_5615;
wire FE_OFN1167_n_5592;
wire FE_OFN1168_n_5592;
wire FE_OFN1169_n_5592;
wire FE_OFN1170_n_5592;
wire FE_OFN1171_n_5592;
wire FE_OFN1172_n_5592;
wire FE_OFN1173_n_5592;
wire FE_OFN1174_n_5592;
wire FE_OFN1175_n_3476;
wire FE_OFN1176_n_3476;
wire FE_OFN1177_n_3476;
wire FE_OFN1178_n_3476;
wire FE_OFN1179_n_3476;
wire FE_OFN1180_n_3476;
wire FE_OFN1181_n_3476;
wire FE_OFN1182_n_3476;
wire FE_OFN1183_n_3476;
wire FE_OFN1184_n_3476;
wire FE_OFN1185_n_3476;
wire FE_OFN1186_n_3476;
wire FE_OFN1187_n_5742;
wire FE_OFN1188_n_5742;
wire FE_OFN1189_n_5742;
wire FE_OFN1190_n_6935;
wire FE_OFN1191_n_6935;
wire FE_OFN1192_n_6935;
wire FE_OFN1193_n_6935;
wire FE_OFN1194_n_6935;
wire FE_OFN1195_n_4090;
wire FE_OFN1196_n_4090;
wire FE_OFN1197_n_4090;
wire FE_OFN1198_n_4090;
wire FE_OFN1199_n_4090;
wire FE_OFN1200_n_4090;
wire FE_OFN1201_n_4090;
wire FE_OFN1202_n_4090;
wire FE_OFN1203_n_4090;
wire FE_OFN1204_n_4090;
wire FE_OFN1205_n_6356;
wire FE_OFN1206_n_6356;
wire FE_OFN1207_n_6356;
wire FE_OFN1208_n_6356;
wire FE_OFN1209_n_4151;
wire FE_OFN1210_n_4151;
wire FE_OFN1211_n_4151;
wire FE_OFN1212_n_4151;
wire FE_OFN1213_n_4151;
wire FE_OFN1214_n_4151;
wire FE_OFN1215_n_4151;
wire FE_OFN1216_n_4151;
wire FE_OFN1217_n_6886;
wire FE_OFN1218_n_6886;
wire FE_OFN1219_n_6886;
wire FE_OFN1220_n_6391;
wire FE_OFN1221_n_6391;
wire FE_OFN1222_n_6391;
wire FE_OFN1223_n_6391;
wire FE_OFN1224_n_6391;
wire FE_OFN1225_n_6391;
wire FE_OFN1226_n_6391;
wire FE_OFN1227_n_6391;
wire FE_OFN1228_n_6391;
wire FE_OFN1229_n_6391;
wire FE_OFN1230_n_6391;
wire FE_OFN1231_n_6391;
wire FE_OFN1232_n_6391;
wire FE_OFN1233_n_6391;
wire FE_OFN1234_n_6391;
wire FE_OFN1235_n_6391;
wire FE_OFN1236_n_6391;
wire FE_OFN1237_n_4092;
wire FE_OFN1238_n_4092;
wire FE_OFN1239_n_4092;
wire FE_OFN1240_n_4092;
wire FE_OFN1241_n_4092;
wire FE_OFN1242_n_4092;
wire FE_OFN1243_n_4092;
wire FE_OFN1244_n_4092;
wire FE_OFN1245_n_4093;
wire FE_OFN1246_n_4093;
wire FE_OFN1247_n_4093;
wire FE_OFN1248_n_4093;
wire FE_OFN1249_n_4093;
wire FE_OFN1250_n_4093;
wire FE_OFN1251_n_4143;
wire FE_OFN1252_n_4143;
wire FE_OFN1253_n_4143;
wire FE_OFN1254_n_4143;
wire FE_OFN1255_n_4143;
wire FE_OFN1256_n_4143;
wire FE_OFN1257_n_4143;
wire FE_OFN1258_n_4143;
wire FE_OFN1259_n_4143;
wire FE_OFN1260_n_4143;
wire FE_OFN1261_n_4143;
wire FE_OFN1262_n_4095;
wire FE_OFN1263_n_4095;
wire FE_OFN1264_n_4095;
wire FE_OFN1265_n_4095;
wire FE_OFN1266_n_4095;
wire FE_OFN1267_n_4095;
wire FE_OFN1268_n_4095;
wire FE_OFN1269_n_4095;
wire FE_OFN1270_n_4095;
wire FE_OFN1271_n_4096;
wire FE_OFN1272_n_4096;
wire FE_OFN1273_n_4096;
wire FE_OFN1274_n_4096;
wire FE_OFN1275_n_4096;
wire FE_OFN1276_n_4096;
wire FE_OFN1277_n_4097;
wire FE_OFN1278_n_4097;
wire FE_OFN1279_n_4097;
wire FE_OFN1280_n_4097;
wire FE_OFN1281_n_4097;
wire FE_OFN1282_n_4097;
wire FE_OFN1283_n_4097;
wire FE_OFN1284_n_4097;
wire FE_OFN1285_n_4097;
wire FE_OFN1286_n_4098;
wire FE_OFN1287_n_4098;
wire FE_OFN1288_n_4098;
wire FE_OFN1289_n_4098;
wire FE_OFN1290_n_4098;
wire FE_OFN1291_n_4098;
wire FE_OFN1292_n_4098;
wire FE_OFN1293_n_4098;
wire FE_OFN1294_n_4098;
wire FE_OFN1295_n_4098;
wire FE_OFN1296_n_5763;
wire FE_OFN1297_n_5763;
wire FE_OFN1298_n_5763;
wire FE_OFN1299_n_5763;
wire FE_OFN1300_n_5763;
wire FE_OFN1301_n_5763;
wire FE_OFN1302_n_5763;
wire FE_OFN1303_n_13124;
wire FE_OFN1304_n_13124;
wire FE_OFN1305_n_13124;
wire FE_OFN1306_n_13124;
wire FE_OFN1307_n_6624;
wire FE_OFN1308_n_6624;
wire FE_OFN1309_n_6624;
wire FE_OFN1310_n_6624;
wire FE_OFN1311_n_6624;
wire FE_OFN1312_n_6624;
wire FE_OFN1313_n_6624;
wire FE_OFN1314_n_6624;
wire FE_OFN1315_n_6624;
wire FE_OFN1316_n_6624;
wire FE_OFN1317_n_6624;
wire FE_OFN1318_n_6436;
wire FE_OFN1319_n_6436;
wire FE_OFN1320_n_6436;
wire FE_OFN1321_n_6436;
wire FE_OFN1322_n_6436;
wire FE_OFN1323_n_6436;
wire FE_OFN1324_n_13547;
wire FE_OFN1325_n_13547;
wire FE_OFN1326_n_13547;
wire FE_OFN1327_n_13547;
wire FE_OFN1328_n_13547;
wire FE_OFN1329_n_13547;
wire FE_OFN1330_n_13547;
wire FE_OFN1331_n_13547;
wire FE_OFN1332_n_13547;
wire FE_OFN1333_n_13547;
wire FE_OFN1334_n_13720;
wire FE_OFN1335_n_13720;
wire FE_OFN1336_n_16439;
wire FE_OFN1337_n_16439;
wire FE_OFN1338_n_8567;
wire FE_OFN1339_n_8567;
wire FE_OFN1340_n_8567;
wire FE_OFN1341_n_8567;
wire FE_OFN1342_n_8567;
wire FE_OFN1343_n_8567;
wire FE_OFN1344_n_8567;
wire FE_OFN1345_n_8567;
wire FE_OFN1346_n_8567;
wire FE_OFN1347_n_8567;
wire FE_OFN1348_n_8567;
wire FE_OFN1349_n_8567;
wire FE_OFN1350_n_8567;
wire FE_OFN1351_n_8567;
wire FE_OFN1352_n_8567;
wire FE_OFN1353_n_8567;
wire FE_OFN1354_n_8567;
wire FE_OFN1355_n_8567;
wire FE_OFN1356_n_8567;
wire FE_OFN1357_n_8567;
wire FE_OFN1358_n_8567;
wire FE_OFN1359_n_8567;
wire FE_OFN1360_n_8567;
wire FE_OFN1361_n_8567;
wire FE_OFN1362_n_8567;
wire FE_OFN1363_n_8567;
wire FE_OFN1364_n_8567;
wire FE_OFN1365_n_8567;
wire FE_OFN1366_n_8567;
wire FE_OFN1367_n_8567;
wire FE_OFN1368_n_8567;
wire FE_OFN1369_n_8567;
wire FE_OFN1370_n_8567;
wire FE_OFN1371_n_8567;
wire FE_OFN1372_n_8567;
wire FE_OFN1373_n_8567;
wire FE_OFN1374_n_8567;
wire FE_OFN1376_n_8567;
wire FE_OFN1377_n_8567;
wire FE_OFN1378_n_8567;
wire FE_OFN1379_n_8567;
wire FE_OFN1380_n_8567;
wire FE_OFN1381_n_8567;
wire FE_OFN1382_n_8567;
wire FE_OFN1383_n_8567;
wire FE_OFN1384_n_8567;
wire FE_OFN1385_n_8567;
wire FE_OFN1386_n_8567;
wire FE_OFN1387_n_8567;
wire FE_OFN1388_n_8567;
wire FE_OFN1389_n_8567;
wire FE_OFN1390_n_8567;
wire FE_OFN1391_n_8567;
wire FE_OFN1392_n_8567;
wire FE_OFN1394_n_8567;
wire FE_OFN1396_n_8567;
wire FE_OFN1397_n_8567;
wire FE_OFN1398_n_8567;
wire FE_OFN1399_n_8567;
wire FE_OFN1400_n_8567;
wire FE_OFN1401_n_8567;
wire FE_OFN1402_n_8567;
wire FE_OFN1403_n_8567;
wire FE_OFN1404_n_8567;
wire FE_OFN1405_n_8567;
wire FE_OFN1406_n_8567;
wire FE_OFN1407_n_8567;
wire FE_OFN1408_n_8567;
wire FE_OFN1409_n_8567;
wire FE_OFN1410_n_8567;
wire FE_OFN1411_n_8567;
wire FE_OFN1412_n_8567;
wire FE_OFN1413_n_8567;
wire FE_OFN1414_n_8567;
wire FE_OFN1415_n_8567;
wire FE_OFN1416_n_8567;
wire FE_OFN1417_n_8567;
wire FE_OFN1419_n_8567;
wire FE_OFN1420_n_8567;
wire FE_OFN1421_n_8567;
wire FE_OFN1422_n_8567;
wire FE_OFN1423_n_8567;
wire FE_OFN1424_n_8567;
wire FE_OFN1425_n_8567;
wire FE_OFN1426_n_8567;
wire FE_OFN1427_n_8567;
wire FE_OFN1428_n_8567;
wire FE_OFN1429_n_16779;
wire FE_OFN1430_n_16779;
wire FE_OFN1431_n_16779;
wire FE_OFN1432_n_16779;
wire FE_OFN1433_n_16779;
wire FE_OFN1434_n_9372;
wire FE_OFN1435_n_9372;
wire FE_OFN1436_n_9372;
wire FE_OFN1437_n_9372;
wire FE_OFN1438_n_9372;
wire FE_OFN1439_n_9372;
wire FE_OFN1440_n_9372;
wire FE_OFN1441_n_9372;
wire FE_OFN1442_n_11125;
wire FE_OFN1443_n_11125;
wire FE_OFN1444_n_11125;
wire FE_OFN1445_n_11125;
wire FE_OFN1446_n_11125;
wire FE_OFN1447_n_9163;
wire FE_OFN1448_n_9163;
wire FE_OFN1449_n_9163;
wire FE_OFN1450_n_9163;
wire FE_OFN1451_n_10588;
wire FE_OFN1452_n_10588;
wire FE_OFN1453_n_10588;
wire FE_OFN1454_n_11138;
wire FE_OFN1455_n_11138;
wire FE_OFN1456_n_11138;
wire FE_OFN1457_n_11138;
wire FE_OFN1458_n_11138;
wire FE_OFN1459_n_11795;
wire FE_OFN1460_n_11795;
wire FE_OFN1461_n_11795;
wire FE_OFN1462_n_11795;
wire FE_OFN1463_n_10789;
wire FE_OFN1464_n_10789;
wire FE_OFN1465_n_10789;
wire FE_OFN1466_n_10789;
wire FE_OFN1467_n_10789;
wire FE_OFN1468_n_10789;
wire FE_OFN1469_g52675_p;
wire FE_OFN146_g65530_p;
wire FE_OFN1470_g52675_p;
wire FE_OFN1471_g52675_p;
wire FE_OFN1472_g52675_p;
wire FE_OFN1473_n_16637;
wire FE_OFN1474_n_16637;
wire FE_OFN1475_n_16637;
wire FE_OFN1477_n_16637;
wire FE_OFN1478_n_16637;
wire FE_OFN1479_n_16637;
wire FE_OFN147_g65530_p;
wire FE_OFN1480_n_15534;
wire FE_OFN1481_n_15534;
wire FE_OFN1483_n_15534;
wire FE_OFN1484_n_15534;
wire FE_OFN1485_n_15534;
wire FE_OFN1486_n_16992;
wire FE_OFN1487_n_9320;
wire FE_OFN1488_n_9320;
wire FE_OFN1489_n_9320;
wire FE_OFN1490_n_9320;
wire FE_OFN1491_n_9320;
wire FE_OFN1492_n_9320;
wire FE_OFN1493_n_9320;
wire FE_OFN1495_n_15558;
wire FE_OFN1496_n_15558;
wire FE_OFN1497_n_15558;
wire FE_OFN1498_n_15558;
wire FE_OFN1499_n_15558;
wire FE_OFN1500_n_15558;
wire FE_OFN1501_n_15558;
wire FE_OFN1502_n_15558;
wire FE_OFN1503_n_15768;
wire FE_OFN1505_n_15768;
wire FE_OFN1506_n_15768;
wire FE_OFN1507_n_15587;
wire FE_OFN1508_n_15587;
wire FE_OFN1509_n_15587;
wire FE_OFN1510_n_15587;
wire FE_OFN1511_n_15587;
wire FE_OFN1513_n_14987;
wire FE_OFN1514_n_10538;
wire FE_OFN1519_n_10892;
wire FE_OFN1520_n_10892;
wire FE_OFN1521_n_10892;
wire FE_OFN1522_n_10892;
wire FE_OFN1523_n_10892;
wire FE_OFN1524_n_10853;
wire FE_OFN1525_n_10853;
wire FE_OFN1526_n_10853;
wire FE_OFN1527_n_10853;
wire FE_OFN1528_n_10853;
wire FE_OFN1529_n_10853;
wire FE_OFN1530_n_10853;
wire FE_OFN1531_n_10143;
wire FE_OFN1532_n_10143;
wire FE_OFN1533_n_10143;
wire FE_OFN1535_n_10143;
wire FE_OFN1536_n_10143;
wire FE_OFN1537_n_10595;
wire FE_OFN1538_n_10595;
wire FE_OFN1539_n_10595;
wire FE_OFN1540_n_10595;
wire FE_OFN1541_n_10595;
wire FE_OFN1542_n_10566;
wire FE_OFN1543_n_10566;
wire FE_OFN1544_n_10566;
wire FE_OFN1545_n_10566;
wire FE_OFN1546_n_10566;
wire FE_OFN1547_n_10566;
wire FE_OFN1548_n_10566;
wire FE_OFN1549_n_12104;
wire FE_OFN1550_n_12104;
wire FE_OFN1551_n_12104;
wire FE_OFN1552_n_12104;
wire FE_OFN1553_n_12104;
wire FE_OFN1554_n_12104;
wire FE_OFN1556_n_12042;
wire FE_OFN1558_n_12042;
wire FE_OFN1559_n_12042;
wire FE_OFN1560_n_12502;
wire FE_OFN1561_n_12502;
wire FE_OFN1562_n_12502;
wire FE_OFN1563_n_12502;
wire FE_OFN1564_n_12502;
wire FE_OFN1565_n_12502;
wire FE_OFN1566_n_12502;
wire FE_OFN1568_n_11027;
wire FE_OFN1572_n_11027;
wire FE_OFN1573_n_12028;
wire FE_OFN1574_n_12028;
wire FE_OFN1575_n_12028;
wire FE_OFN1576_n_12028;
wire FE_OFN1577_n_12028;
wire FE_OFN1579_n_12306;
wire FE_OFN1581_n_12306;
wire FE_OFN1583_n_12306;
wire FE_OFN1584_n_12306;
wire FE_OFN1585_n_13736;
wire FE_OFN1586_n_13736;
wire FE_OFN1587_n_13736;
wire FE_OFN1588_n_13736;
wire FE_OFN1589_n_13736;
wire FE_OFN1590_n_13741;
wire FE_OFN1591_n_13741;
wire FE_OFN1592_n_13741;
wire FE_OFN1593_n_13741;
wire FE_OFN1596_n_13741;
wire FE_OFN1598_n_13995;
wire FE_OFN1599_n_13995;
wire FE_OFN1600_n_13995;
wire FE_OFN1601_n_13995;
wire FE_OFN1602_n_13995;
wire FE_OFN1603_n_13997;
wire FE_OFN1604_n_13997;
wire FE_OFN1605_n_13997;
wire FE_OFN1606_n_13997;
wire FE_OFN1607_n_2122;
wire FE_OFN1608_n_2122;
wire FE_OFN1609_n_2122;
wire FE_OFN1610_n_2122;
wire FE_OFN1611_n_2122;
wire FE_OFN1612_n_2122;
wire FE_OFN1613_n_1787;
wire FE_OFN1614_n_1787;
wire FE_OFN1615_n_1787;
wire FE_OFN1616_n_1787;
wire FE_OFN1617_n_1787;
wire FE_OFN1618_n_1787;
wire FE_OFN1619_n_1787;
wire FE_OFN1620_n_1787;
wire FE_OFN1621_n_1787;
wire FE_OFN1622_n_4438;
wire FE_OFN1623_n_4438;
wire FE_OFN1624_n_4438;
wire FE_OFN1625_n_4438;
wire FE_OFN1626_n_4438;
wire FE_OFN1627_n_4438;
wire FE_OFN1628_n_4438;
wire FE_OFN1629_n_9531;
wire FE_OFN1630_n_9531;
wire FE_OFN1631_n_9531;
wire FE_OFN1632_n_9531;
wire FE_OFN1633_n_9531;
wire FE_OFN1634_n_9531;
wire FE_OFN1635_n_9531;
wire FE_OFN1636_n_4460;
wire FE_OFN1637_n_4671;
wire FE_OFN1638_n_4671;
wire FE_OFN1639_n_4671;
wire FE_OFN1640_n_4671;
wire FE_OFN1641_n_4671;
wire FE_OFN1642_n_4671;
wire FE_OFN1643_n_4671;
wire FE_OFN1644_n_4671;
wire FE_OFN1645_n_4671;
wire FE_OFN1646_n_9428;
wire FE_OFN1647_n_9428;
wire FE_OFN1648_n_9428;
wire FE_OFN1649_n_9428;
wire FE_OFN1650_n_9428;
wire FE_OFN1651_n_9428;
wire FE_OFN1652_n_9502;
wire FE_OFN1653_n_9502;
wire FE_OFN1654_n_9502;
wire FE_OFN1655_n_9502;
wire FE_OFN1656_n_9502;
wire FE_OFN1657_n_9502;
wire FE_OFN1658_n_4490;
wire FE_OFN1659_n_4490;
wire FE_OFN1660_n_4490;
wire FE_OFN1661_n_4490;
wire FE_OFN1662_n_4490;
wire FE_OFN1663_n_4490;
wire FE_OFN1664_n_9477;
wire FE_OFN1665_n_9477;
wire FE_OFN1666_n_9477;
wire FE_OFN1667_n_9477;
wire FE_OFN1668_n_9477;
wire FE_OFN1669_n_9477;
wire FE_OFN1670_n_9477;
wire FE_OFN1671_n_9477;
wire FE_OFN1672_n_4655;
wire FE_OFN1673_n_4655;
wire FE_OFN1674_n_4655;
wire FE_OFN1675_n_4655;
wire FE_OFN1676_n_4655;
wire FE_OFN1677_n_4655;
wire FE_OFN1678_n_4655;
wire FE_OFN1679_n_4655;
wire FE_OFN1680_n_4655;
wire FE_OFN1681_n_4669;
wire FE_OFN1682_n_4669;
wire FE_OFN1683_n_9528;
wire FE_OFN1684_n_9528;
wire FE_OFN1685_n_9528;
wire FE_OFN1686_n_9528;
wire FE_OFN1687_n_9528;
wire FE_OFN1688_n_9528;
wire FE_OFN1689_n_9528;
wire FE_OFN1690_n_9528;
wire FE_OFN1691_n_9528;
wire FE_OFN1692_n_9528;
wire FE_OFN1693_n_3368;
wire FE_OFN1694_n_3368;
wire FE_OFN1695_n_3368;
wire FE_OFN1696_n_5751;
wire FE_OFN1697_n_5751;
wire FE_OFN1698_n_5751;
wire FE_OFN1699_n_5751;
wire FE_OFN1700_n_5751;
wire FE_OFN1701_n_4868;
wire FE_OFN1702_n_4868;
wire FE_OFN1703_n_4868;
wire FE_OFN1704_n_4868;
wire FE_OFN1705_n_4868;
wire FE_OFN1706_n_4868;
wire FE_OFN1707_n_4868;
wire FE_OFN1708_n_4868;
wire FE_OFN1709_n_4868;
wire FE_OFN1710_n_4868;
wire FE_OFN1711_n_13563;
wire FE_OFN1712_n_13563;
wire FE_OFN1713_n_13650;
wire FE_OFN1714_n_13650;
wire FE_OFN1716_n_16698;
wire FE_OFN1719_n_16891;
wire FE_OFN1720_n_16891;
wire FE_OFN1721_n_16891;
wire FE_OFN1722_n_16891;
wire FE_OFN1723_n_16891;
wire FE_OFN1724_n_16891;
wire FE_OFN1725_n_16891;
wire FE_OFN1726_n_9975;
wire FE_OFN1727_n_9975;
wire FE_OFN1728_n_9975;
wire FE_OFN1729_n_9975;
wire FE_OFN1730_n_9975;
wire FE_OFN1731_n_9975;
wire FE_OFN1732_n_16317;
wire FE_OFN1733_n_16317;
wire FE_OFN1734_n_16317;
wire FE_OFN1735_n_16317;
wire FE_OFN1736_n_16317;
wire FE_OFN1737_n_11019;
wire FE_OFN1738_n_11019;
wire FE_OFN1739_n_11019;
wire FE_OFN1740_n_11019;
wire FE_OFN1741_n_11019;
wire FE_OFN1742_n_11019;
wire FE_OFN1743_n_12004;
wire FE_OFN1744_n_12004;
wire FE_OFN1745_n_12004;
wire FE_OFN1746_n_12004;
wire FE_OFN1747_n_12004;
wire FE_OFN1748_n_12004;
wire FE_OFN1749_n_12004;
wire FE_OFN1751_n_12086;
wire FE_OFN1752_n_12086;
wire FE_OFN1753_n_12086;
wire FE_OFN1754_n_12681;
wire FE_OFN1755_n_12681;
wire FE_OFN1756_n_12681;
wire FE_OFN1757_n_12681;
wire FE_OFN1758_n_10780;
wire FE_OFN1759_n_10780;
wire FE_OFN1760_n_10780;
wire FE_OFN1761_n_10780;
wire FE_OFN1762_n_10780;
wire FE_OFN1767_n_14054;
wire FE_OFN1768_n_14054;
wire FE_OFN1769_n_14054;
wire FE_OFN1770_n_14054;
wire FE_OFN1771_n_14054;
wire FE_OFN1772_n_13800;
wire FE_OFN1773_n_13800;
wire FE_OFN1774_n_13800;
wire FE_OFN1775_n_13800;
wire FE_OFN1776_parchk_pci_ad_reg_in_1222;
wire FE_OFN1777_parchk_pci_ad_reg_in_1222;
wire FE_OFN1778_parchk_pci_ad_reg_in_1222;
wire FE_OFN1779_parchk_pci_ad_reg_in_1221;
wire FE_OFN1780_parchk_pci_ad_reg_in_1221;
wire FE_OFN1781_parchk_pci_ad_reg_in_1221;
wire FE_OFN1782_n_1699;
wire FE_OFN1783_n_1699;
wire FE_OFN1784_n_1699;
wire FE_OFN1785_n_1699;
wire FE_OFN1786_n_1699;
wire FE_OFN1789_n_9823;
wire FE_OFN1790_n_2687;
wire FE_OFN1791_n_9904;
wire FE_OFN1792_n_9904;
wire FE_OFN1793_n_9904;
wire FE_OFN1794_n_9904;
wire FE_OFN1795_n_9904;
wire FE_OFN1796_n_2299;
wire FE_OFN1797_n_2299;
wire FE_OFN1798_n_9690;
wire FE_OFN1799_n_9690;
wire FE_OFN1800_n_9690;
wire FE_OFN1801_n_9690;
wire FE_OFN1802_n_9690;
wire FE_OFN1803_n_9690;
wire FE_OFN1804_n_4501;
wire FE_OFN1805_n_4501;
wire FE_OFN1806_n_4501;
wire FE_OFN1807_n_4501;
wire FE_OFN1808_n_4454;
wire FE_OFN1809_n_4454;
wire FE_OFN1810_n_4454;
wire FE_OFN1811_n_7845;
wire FE_OFN1812_n_7845;
wire FE_OFN1813_n_2919;
wire FE_OFN1814_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid;
wire FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid;
wire FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid;
wire FE_OFN1819_n_2919;
wire FE_OFN186_n_15768;
wire FE_OFN190_n_1193;
wire FE_OFN191_n_1193;
wire FE_OFN1935_n_1781;
wire FE_OFN1936_n_1781;
wire FE_OFN1937_g66085_p;
wire FE_OFN1938_g66085_p;
wire FE_OFN1939_g66095_p;
wire FE_OFN1940_g66095_p;
wire FE_OFN1941_n_3241;
wire FE_OFN1942_n_3241;
wire FE_OFN1943_n_15813;
wire FE_OFN1944_n_15813;
wire FE_OFN1945_n_13784;
wire FE_OFN1946_n_13784;
wire FE_OFN196_n_2683;
wire FE_OFN197_n_2683;
wire FE_OFN198_n_3298;
wire FE_OFN199_n_3298;
wire FE_OFN1_n_4778;
wire FE_OFN200_n_9230;
wire FE_OFN201_n_9230;
wire FE_OFN2020_n_4778;
wire FE_OFN2021_n_4778;
wire FE_OFN2022_n_4778;
wire FE_OFN202_n_9228;
wire FE_OFN203_n_9228;
wire FE_OFN204_n_9140;
wire FE_OFN2051_n_6965;
wire FE_OFN2052_n_6965;
wire FE_OFN2053_n_8831;
wire FE_OFN2054_n_8831;
wire FE_OFN2055_n_8831;
wire FE_OFN2056_n_2117;
wire FE_OFN2057_n_2117;
wire FE_OFN2058_n_13447;
wire FE_OFN2059_n_13447;
wire FE_OFN205_n_9140;
wire FE_OFN2060_g66087_p;
wire FE_OFN2061_g66087_p;
wire FE_OFN2062_n_6391;
wire FE_OFN2063_n_6391;
wire FE_OFN2064_n_6391;
wire FE_OFN2069_n_15978;
wire FE_OFN206_n_9865;
wire FE_OFN2070_n_15978;
wire FE_OFN2071_n_15978;
wire FE_OFN2072_n_15978;
wire FE_OFN2073_n_2723;
wire FE_OFN2074_n_2723;
wire FE_OFN2075_FE_OCPUNCON1952_FE_OFN697_n_16760;
wire FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760;
wire FE_OFN2077_n_8069;
wire FE_OFN2079_n_8069;
wire FE_OFN207_n_9865;
wire FE_OFN2080_n_8176;
wire FE_OFN2081_n_8176;
wire FE_OFN2082_n_8407;
wire FE_OFN2083_n_8407;
wire FE_OFN2084_n_8407;
wire FE_OFN2085_n_8448;
wire FE_OFN2086_n_8448;
wire FE_OFN2088_n_13124;
wire FE_OFN208_n_9126;
wire FE_OFN2092_n_2301;
wire FE_OFN2093_n_2301;
wire FE_OFN2094_n_2520;
wire FE_OFN2095_n_2520;
wire FE_OFN2096_n_2520;
wire FE_OFN2099_n_3281;
wire FE_OFN209_n_9126;
wire FE_OFN2100_n_3281;
wire FE_OFN2101_n_2834;
wire FE_OFN2102_n_2834;
wire FE_OFN2103_g64577_p;
wire FE_OFN2104_g64577_p;
wire FE_OFN2105_g64577_p;
wire FE_OFN2106_g64577_p;
wire FE_OFN2107_n_2047;
wire FE_OFN2108_n_2047;
wire FE_OFN2109_n_2047;
wire FE_OFN210_n_9858;
wire FE_OFN2110_n_2248;
wire FE_OFN2111_n_2248;
wire FE_OFN2112_n_2053;
wire FE_OFN2113_n_2053;
wire FE_OFN2114_wishbone_slave_unit_pci_initiator_if_data_source;
wire FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source;
wire FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source;
wire FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source;
wire FE_OFN2119_wishbone_slave_unit_pci_initiator_if_data_source;
wire FE_OFN211_n_9858;
wire FE_OFN2121_n_2687;
wire FE_OFN2123_n_16497;
wire FE_OFN2124_n_16497;
wire FE_OFN2125_n_16497;
wire FE_OFN2126_n_16497;
wire FE_OFN2127_n_16497;
wire FE_OFN2128_n_16497;
wire FE_OFN2129_n_16720;
wire FE_OFN212_n_9124;
wire FE_OFN2130_n_10588;
wire FE_OFN2131_n_10588;
wire FE_OFN2132_n_13124;
wire FE_OFN2133_n_13124;
wire FE_OFN2134_n_13124;
wire FE_OFN2135_n_13124;
wire FE_OFN2136_n_13124;
wire FE_OFN2137_n_15534;
wire FE_OFN2139_n_16992;
wire FE_OFN213_n_9124;
wire FE_OFN2140_n_16992;
wire FE_OFN2141_n_16992;
wire FE_OFN2142_n_16992;
wire FE_OFN2143_n_16992;
wire FE_OFN2144_n_16992;
wire FE_OFN2145_n_16992;
wire FE_OFN2146_n_9320;
wire FE_OFN2147_n_10595;
wire FE_OFN2148_n_10595;
wire FE_OFN2149_n_10595;
wire FE_OFN214_n_9856;
wire FE_OFN2150_n_10595;
wire FE_OFN2151_n_16439;
wire FE_OFN2152_n_16439;
wire FE_OFN2153_n_16439;
wire FE_OFN2154_n_16439;
wire FE_OFN2155_n_16439;
wire FE_OFN2156_n_16439;
wire FE_OFN2157_n_16439;
wire FE_OFN2158_n_16439;
wire FE_OFN2159_n_16301;
wire FE_OFN215_n_9856;
wire FE_OFN2160_n_16301;
wire FE_OFN2161_n_16301;
wire FE_OFN2162_n_16301;
wire FE_OFN2163_n_16301;
wire FE_OFN2164_n_16301;
wire FE_OFN2165_n_16301;
wire FE_OFN2166_n_8567;
wire FE_OFN2167_n_8567;
wire FE_OFN2168_n_8567;
wire FE_OFN2169_n_8567;
wire FE_OFN216_n_9889;
wire FE_OFN2170_n_8567;
wire FE_OFN2171_n_8567;
wire FE_OFN2172_n_8567;
wire FE_OFN2173_n_8567;
wire FE_OFN2174_n_8567;
wire FE_OFN2175_n_8567;
wire FE_OFN2176_n_8567;
wire FE_OFN2177_n_8567;
wire FE_OFN2178_n_8567;
wire FE_OFN2179_n_8567;
wire FE_OFN217_n_9889;
wire FE_OFN2180_n_8567;
wire FE_OFN2181_n_8567;
wire FE_OFN2182_n_8567;
wire FE_OFN2183_n_8567;
wire FE_OFN2184_n_8567;
wire FE_OFN2185_n_8567;
wire FE_OFN2186_n_8567;
wire FE_OFN2187_n_8567;
wire FE_OFN2188_n_8567;
wire FE_OFN2189_n_8567;
wire FE_OFN218_n_9853;
wire FE_OFN2190_n_8567;
wire FE_OFN2191_n_8567;
wire FE_OFN2192_n_16779;
wire FE_OFN2193_n_9163;
wire FE_OFN2194_n_9163;
wire FE_OFN2195_n_9163;
wire FE_OFN2196_n_9163;
wire FE_OFN2197_n_10256;
wire FE_OFN2198_n_10256;
wire FE_OFN2199_n_10256;
wire FE_OFN219_n_9853;
wire FE_OFN21_n_9372;
wire FE_OFN2200_n_10256;
wire FE_OFN2201_n_12042;
wire FE_OFN2202_n_12042;
wire FE_OFN2203_n_12042;
wire FE_OFN2204_n_12028;
wire FE_OFN2205_n_10538;
wire FE_OFN2206_n_10892;
wire FE_OFN2207_n_10892;
wire FE_OFN2208_n_11795;
wire FE_OFN2209_n_11027;
wire FE_OFN220_n_9846;
wire FE_OFN2210_n_11027;
wire FE_OFN2211_n_8407;
wire FE_OFN2212_n_8407;
wire FE_OFN2213_n_15366;
wire FE_OFN2214_n_15366;
wire FE_OFN2215_n_15366;
wire FE_OFN2216_n_10143;
wire FE_OFN221_n_9846;
wire FE_OFN222_n_9844;
wire FE_OFN223_n_9844;
wire FE_OFN2240_g52675_p;
wire FE_OFN2241_g52675_p;
wire FE_OFN2242_g52675_p;
wire FE_OFN2243_g52675_p;
wire FE_OFN2244_n_4792;
wire FE_OFN2245_n_4792;
wire FE_OFN2246_n_2113;
wire FE_OFN2247_n_2113;
wire FE_OFN2248_n_1790;
wire FE_OFN2249_n_1790;
wire FE_OFN224_n_9122;
wire FE_OFN2250_n_2101;
wire FE_OFN2251_n_2101;
wire FE_OFN2252_n_9687;
wire FE_OFN2253_n_9687;
wire FE_OFN2254_n_9687;
wire FE_OFN2255_n_8060;
wire FE_OFN2256_n_8060;
wire FE_OFN2257_n_8060;
wire FE_OFN2258_n_8060;
wire FE_OFN2259_n_2775;
wire FE_OFN225_n_9122;
wire FE_OFN2260_n_2775;
wire FE_OFN226_n_9841;
wire FE_OFN227_n_9841;
wire FE_OFN228_n_9120;
wire FE_OFN229_n_9120;
wire FE_OFN230_n_9839;
wire FE_OFN231_n_9839;
wire FE_OFN232_n_9876;
wire FE_OFN233_n_9876;
wire FE_OFN234_n_9834;
wire FE_OFN235_n_9834;
wire FE_OFN236_n_9118;
wire FE_OFN237_n_9118;
wire FE_OFN238_n_9832;
wire FE_OFN239_n_9832;
wire FE_OFN240_n_9830;
wire FE_OFN241_n_9830;
wire FE_OFN242_n_9116;
wire FE_OFN243_n_9116;
wire FE_OFN244_n_9114;
wire FE_OFN245_n_9114;
wire FE_OFN246_n_9112;
wire FE_OFN247_n_9112;
wire FE_OFN248_n_9789;
wire FE_OFN250_n_9789;
wire FE_OFN251_n_9868;
wire FE_OFN252_n_9868;
wire FE_OFN253_n_9825;
wire FE_OFN254_n_9825;
wire FE_OFN255_n_8969;
wire FE_OFN256_n_8969;
wire FE_OFN257_n_9862;
wire FE_OFN258_n_9862;
wire FE_OFN259_n_9860;
wire FE_OFN260_n_9860;
wire FE_OFN261_n_9851;
wire FE_OFN262_n_9851;
wire FE_OFN263_n_9849;
wire FE_OFN264_n_9849;
wire FE_OFN265_n_9884;
wire FE_OFN266_n_9884;
wire FE_OFN267_n_9880;
wire FE_OFN268_n_9880;
wire FE_OFN269_n_9836;
wire FE_OFN270_n_9836;
wire FE_OFN271_n_9828;
wire FE_OFN272_n_9828;
wire FE_OFN275_n_9941;
wire FE_OFN276_n_9941;
wire FE_OFN2_n_4778;
wire FE_OFN334_g66081_p;
wire FE_OFN335_g66081_p;
wire FE_OFN336_g66089_p;
wire FE_OFN337_g66089_p;
wire FE_OFN365_n_4093;
wire FE_OFN369_n_4092;
wire FE_OFN3_n_4778;
wire FE_OFN514_n_9697;
wire FE_OFN515_n_9697;
wire FE_OFN516_n_9697;
wire FE_OFN517_n_9697;
wire FE_OFN518_n_9697;
wire FE_OFN519_n_9697;
wire FE_OFN523_n_9428;
wire FE_OFN524_n_9899;
wire FE_OFN525_n_9899;
wire FE_OFN526_n_9899;
wire FE_OFN527_n_9899;
wire FE_OFN528_n_9899;
wire FE_OFN529_n_9899;
wire FE_OFN530_n_9823;
wire FE_OFN531_n_9823;
wire FE_OFN532_n_9823;
wire FE_OFN533_n_9823;
wire FE_OFN534_n_9823;
wire FE_OFN535_n_9823;
wire FE_OFN537_n_9690;
wire FE_OFN539_n_9690;
wire FE_OFN540_n_9690;
wire FE_OFN541_n_9690;
wire FE_OFN542_n_9690;
wire FE_OFN543_n_9690;
wire FE_OFN548_n_9477;
wire FE_OFN549_n_9864;
wire FE_OFN550_n_9864;
wire FE_OFN551_n_9864;
wire FE_OFN552_n_9864;
wire FE_OFN553_n_9864;
wire FE_OFN554_n_9864;
wire FE_OFN555_n_9864;
wire FE_OFN556_n_9864;
wire FE_OFN557_n_9895;
wire FE_OFN558_n_9895;
wire FE_OFN559_n_9895;
wire FE_OFN560_n_9895;
wire FE_OFN561_n_9895;
wire FE_OFN562_n_9895;
wire FE_OFN563_n_9895;
wire FE_OFN564_n_9895;
wire FE_OFN568_n_9528;
wire FE_OFN569_n_9528;
wire FE_OFN572_n_9502;
wire FE_OFN573_n_9902;
wire FE_OFN574_n_9902;
wire FE_OFN575_n_9902;
wire FE_OFN576_n_9902;
wire FE_OFN577_n_9902;
wire FE_OFN579_n_9531;
wire FE_OFN580_n_9531;
wire FE_OFN582_n_9692;
wire FE_OFN583_n_9692;
wire FE_OFN584_n_9692;
wire FE_OFN585_n_9692;
wire FE_OFN587_n_9692;
wire FE_OFN588_n_9692;
wire FE_OFN589_n_9692;
wire FE_OFN590_n_9694;
wire FE_OFN591_n_9694;
wire FE_OFN592_n_9694;
wire FE_OFN593_n_9694;
wire FE_OFN595_n_9694;
wire FE_OFN596_n_9694;
wire FE_OFN597_n_9694;
wire FE_OFN598_n_9687;
wire FE_OFN599_n_9687;
wire FE_OFN600_n_9687;
wire FE_OFN601_n_9687;
wire FE_OFN602_n_9687;
wire FE_OFN603_n_9687;
wire FE_OFN605_n_9904;
wire FE_OFN606_n_9904;
wire FE_OFN607_n_9904;
wire FE_OFN608_n_9904;
wire FE_OFN611_n_4501;
wire FE_OFN612_n_4501;
wire FE_OFN613_n_4501;
wire FE_OFN614_n_4501;
wire FE_OFN615_n_4501;
wire FE_OFN618_n_4490;
wire FE_OFN619_n_4490;
wire FE_OFN620_n_4490;
wire FE_OFN621_n_4409;
wire FE_OFN622_n_4409;
wire FE_OFN623_n_4409;
wire FE_OFN624_n_4409;
wire FE_OFN625_n_4409;
wire FE_OFN627_n_4454;
wire FE_OFN628_n_4454;
wire FE_OFN629_n_4454;
wire FE_OFN630_n_4454;
wire FE_OFN631_n_4454;
wire FE_OFN632_n_4454;
wire FE_OFN633_n_4454;
wire FE_OFN634_n_4454;
wire FE_OFN636_n_4669;
wire FE_OFN638_n_4669;
wire FE_OFN639_n_4669;
wire FE_OFN640_n_4669;
wire FE_OFN641_n_4677;
wire FE_OFN642_n_4677;
wire FE_OFN643_n_4677;
wire FE_OFN644_n_4677;
wire FE_OFN645_n_4497;
wire FE_OFN646_n_4497;
wire FE_OFN647_n_4497;
wire FE_OFN648_n_4497;
wire FE_OFN649_n_4497;
wire FE_OFN650_n_4508;
wire FE_OFN651_n_4508;
wire FE_OFN652_n_4508;
wire FE_OFN653_n_4508;
wire FE_OFN654_n_4508;
wire FE_OFN658_n_4392;
wire FE_OFN659_n_4392;
wire FE_OFN660_n_4392;
wire FE_OFN661_n_4392;
wire FE_OFN662_n_4392;
wire FE_OFN663_n_4495;
wire FE_OFN664_n_4495;
wire FE_OFN665_n_4495;
wire FE_OFN666_n_4495;
wire FE_OFN667_n_4495;
wire FE_OFN668_n_4505;
wire FE_OFN669_n_4505;
wire FE_OFN670_n_4505;
wire FE_OFN671_n_4505;
wire FE_OFN672_n_4505;
wire FE_OFN678_n_4460;
wire FE_OFN679_n_4460;
wire FE_OFN681_n_4460;
wire FE_OFN682_n_4460;
wire FE_OFN683_n_4417;
wire FE_OFN684_n_4417;
wire FE_OFN685_n_4417;
wire FE_OFN686_n_4417;
wire FE_OFN687_n_4417;
wire FE_OFN689_n_4438;
wire FE_OFN697_n_16760;
wire FE_OFN698_n_7845;
wire FE_OFN699_n_7845;
wire FE_OFN700_n_7845;
wire FE_OFN701_n_7845;
wire FE_OFN702_n_7845;
wire FE_OFN703_n_8069;
wire FE_OFN704_n_8069;
wire FE_OFN705_n_8119;
wire FE_OFN706_n_8119;
wire FE_OFN707_n_8119;
wire FE_OFN708_n_8232;
wire FE_OFN709_n_8232;
wire FE_OFN710_n_8232;
wire FE_OFN711_n_8140;
wire FE_OFN712_n_8140;
wire FE_OFN713_n_8140;
wire FE_OFN714_n_8140;
wire FE_OFN715_n_8176;
wire FE_OFN716_n_8176;
wire FE_OFN717_n_8176;
wire FE_OFN718_n_8060;
wire FE_OFN719_n_8060;
wire FE_OFN720_n_8060;
wire FE_OFN732_n_7498;
wire FE_OFN775_n_15366;
wire FE_OFN776_n_15366;
wire FE_OFN777_n_4152;
wire FE_OFN778_n_4152;
wire FE_OFN779_n_2746;
wire FE_OFN780_n_2746;
wire FE_OFN781_n_2746;
wire FE_OFN782_n_2678;
wire FE_OFN783_n_2678;
wire FE_OFN784_n_2678;
wire FE_OFN785_n_2678;
wire FE_OFN786_n_2678;
wire FE_OFN787_n_2678;
wire FE_OFN789_n_2678;
wire FE_OFN792_n_2547;
wire FE_OFN793_n_2547;
wire FE_OFN794_n_2520;
wire FE_OFN795_n_2520;
wire FE_OFN877_g64577_p;
wire FE_OFN881_g64577_p;
wire FE_OFN882_g64577_p;
wire FE_OFN8_n_11877;
wire FE_OFN900_n_4736;
wire FE_OFN901_n_4736;
wire FE_OFN902_n_4736;
wire FE_OFN903_n_4736;
wire FE_OFN904_n_4736;
wire FE_OFN905_n_4736;
wire FE_OFN906_n_4736;
wire FE_OFN908_n_4734;
wire FE_OFN912_n_4727;
wire FE_OFN915_n_4725;
wire FE_OFN916_n_4725;
wire FE_OFN917_n_4725;
wire FE_OFN918_n_4725;
wire FE_OFN923_n_4740;
wire FE_OFN926_n_4730;
wire FE_OFN927_n_4730;
wire FE_OFN928_n_4730;
wire FE_OFN929_n_4730;
wire FE_OFN930_n_4730;
wire FE_OFN934_n_2292;
wire FE_OFN935_n_2292;
wire FE_OFN936_n_2292;
wire FE_OFN937_n_2292;
wire FE_OFN938_n_2292;
wire FE_OFN941_n_2047;
wire FE_OFN944_n_2248;
wire FE_OFN945_n_2248;
wire FE_OFN946_n_2248;
wire FE_OFN947_n_2248;
wire FE_OFN948_n_2248;
wire FE_OFN949_n_2055;
wire FE_OFN950_n_2055;
wire FE_OFN951_n_2055;
wire FE_OFN952_n_2055;
wire FE_OFN953_n_2055;
wire FE_OFN954_n_1699;
wire FE_OFN955_n_1699;
wire FE_OFN956_n_1699;
wire FE_OFN957_n_2299;
wire FE_OFN958_n_2299;
wire FE_OFN959_n_2299;
wire FE_OFN966_n_2233;
wire FE_OFN967_n_2233;
wire FE_OFN968_n_13784;
wire FE_OFN969_n_13784;
wire FE_OFN982_n_2700;
wire FE_OFN983_n_2700;
wire FE_OFN984_n_2697;
wire FE_OFN985_n_2697;
wire FE_OFN986_n_2696;
wire FE_OFN987_n_2696;
wire FE_OFN988_n_574;
wire FE_OFN989_n_574;
wire FE_OFN991_n_2373;
wire FE_OFN992_n_2373;
wire FE_OFN993_n_15366;
wire FE_OFN994_n_15366;
wire FE_OFN995_n_15366;
wire FE_OFN996_n_15366;
wire FE_OFN997_n_15978;
wire FE_OFN999_n_15978;
wire FE_OFN9_n_11877;
wire FE_RN_0_0;
wire FE_RN_100_0;
wire FE_RN_101_0;
wire FE_RN_102_0;
wire FE_RN_103_0;
wire TIMEBOOST_net_12666;
wire FE_RN_105_0;
wire FE_RN_106_0;
wire FE_RN_107_0;
wire FE_RN_108_0;
wire FE_RN_109_0;
wire FE_RN_110_0;
wire FE_RN_111_0;
wire FE_RN_112_0;
wire FE_RN_113_0;
wire FE_RN_114_0;
wire FE_RN_115_0;
wire FE_RN_116_0;
wire TIMEBOOST_net_185;
wire FE_RN_120_0;
wire FE_RN_121_0;
wire FE_RN_122_0;
wire FE_RN_124_0;
wire TIMEBOOST_net_11563;
wire FE_RN_127_0;
wire TIMEBOOST_net_11589;
wire FE_RN_130_0;
wire TIMEBOOST_net_13485;
wire FE_RN_135_0;
wire FE_RN_136_0;
wire FE_RN_137_0;
wire FE_RN_138_0;
wire FE_RN_139_0;
wire FE_RN_140_0;
wire FE_RN_141_0;
wire FE_RN_142_0;
wire FE_RN_143_0;
wire FE_RN_144_0;
wire FE_RN_145_0;
wire FE_RN_146_0;
wire FE_RN_147_0;
wire FE_RN_148_0;
wire FE_RN_149_0;
wire FE_RN_150_0;
wire FE_RN_151_0;
wire TIMEBOOST_net_273;
wire FE_RN_153_0;
wire FE_RN_154_0;
wire TIMEBOOST_net_11662;
wire FE_RN_156_0;
wire FE_RN_158_0;
wire FE_RN_159_0;
wire FE_RN_15_0;
wire FE_RN_160_0;
wire TIMEBOOST_net_221;
wire TIMEBOOST_net_11778;
wire FE_RN_176_0;
wire FE_RN_177_0;
wire FE_RN_178_0;
wire FE_RN_179_0;
wire FE_RN_180_0;
wire FE_RN_181_0;
wire FE_RN_182_0;
wire FE_RN_183_0;
wire FE_RN_184_0;
wire FE_RN_185_0;
wire FE_RN_186_0;
wire FE_RN_187_0;
wire FE_RN_188_0;
wire FE_RN_189_0;
wire FE_RN_18_0;
wire FE_RN_190_0;
wire FE_RN_191_0;
wire FE_RN_192_0;
wire FE_RN_193_0;
wire FE_RN_194_0;
wire FE_RN_195_0;
wire FE_RN_196_0;
wire FE_RN_197_0;
wire FE_RN_198_0;
wire FE_RN_199_0;
wire FE_RN_19_0;
wire FE_RN_200_0;
wire FE_RN_201_0;
wire FE_RN_202_0;
wire FE_RN_203_0;
wire FE_RN_207_0;
wire FE_RN_208_0;
wire FE_RN_209_0;
wire FE_RN_20_0;
wire FE_RN_211_0;
wire TIMEBOOST_net_11564;
wire FE_RN_213_0;
wire FE_RN_214_0;
wire FE_RN_215_0;
wire FE_RN_216_0;
wire FE_RN_217_0;
wire FE_RN_218_0;
wire FE_RN_219_0;
wire FE_RN_220_0;
wire FE_RN_221_0;
wire FE_RN_222_0;
wire FE_RN_223_0;
wire FE_RN_224_0;
wire FE_RN_225_0;
wire FE_RN_226_0;
wire FE_RN_227_0;
wire FE_RN_228_0;
wire FE_RN_229_0;
wire FE_RN_230_0;
wire FE_RN_231_0;
wire FE_RN_232_0;
wire FE_RN_233_0;
wire FE_RN_234_0;
wire FE_RN_235_0;
wire FE_RN_236_0;
wire FE_RN_237_0;
wire FE_RN_238_0;
wire FE_RN_239_0;
wire FE_RN_23_0;
wire FE_RN_240_0;
wire FE_RN_241_0;
wire FE_RN_242_0;
wire FE_RN_243_0;
wire FE_RN_244_0;
wire FE_RN_245_0;
wire FE_RN_246_0;
wire FE_RN_247_0;
wire FE_RN_248_0;
wire FE_RN_249_0;
wire FE_RN_250_0;
wire FE_RN_251_0;
wire FE_RN_259_0;
wire FE_RN_25_0;
wire FE_RN_260_0;
wire FE_RN_261_0;
wire FE_RN_262_0;
wire FE_RN_263_0;
wire FE_RN_264_0;
wire TIMEBOOST_net_9615;
wire TIMEBOOST_net_13786;
wire FE_RN_267_0;
wire FE_RN_268_0;
wire FE_RN_269_0;
wire FE_RN_26_0;
wire FE_RN_270_0;
wire FE_RN_271_0;
wire TIMEBOOST_net_12701;
wire FE_RN_273_0;
wire FE_RN_274_0;
wire FE_RN_275_0;
wire FE_RN_276_0;
wire FE_RN_278_0;
wire FE_RN_279_0;
wire FE_RN_27_0;
wire FE_RN_280_0;
wire FE_RN_281_0;
wire TIMEBOOST_net_13900;
wire FE_RN_283_0;
wire FE_RN_284_0;
wire FE_RN_285_0;
wire TIMEBOOST_net_13966;
wire FE_RN_28_0;
wire FE_RN_294_0;
wire FE_RN_295_0;
wire TIMEBOOST_net_6;
wire FE_RN_299_0;
wire FE_RN_29_0;
wire TIMEBOOST_net_14075;
wire FE_RN_302_0;
wire FE_RN_303_0;
wire FE_RN_304_0;
wire FE_RN_305_0;
wire TIMEBOOST_net_12411;
wire FE_RN_307_0;
wire FE_RN_308_0;
wire FE_RN_309_0;
wire FE_RN_30_0;
wire FE_RN_310_0;
wire FE_RN_311_0;
wire FE_RN_312_0;
wire FE_RN_313_0;
wire FE_RN_314_0;
wire FE_RN_315_0;
wire FE_RN_316_0;
wire FE_RN_317_0;
wire FE_RN_318_0;
wire FE_RN_319_0;
wire FE_RN_31_0;
wire FE_RN_320_0;
wire FE_RN_321_0;
wire FE_RN_322_0;
wire FE_RN_323_0;
wire FE_RN_324_0;
wire FE_RN_325_0;
wire FE_RN_326_0;
wire FE_RN_327_0;
wire FE_RN_328_0;
wire FE_RN_329_0;
wire FE_RN_32_0;
wire FE_RN_330_0;
wire FE_RN_331_0;
wire FE_RN_332_0;
wire FE_RN_333_0;
wire FE_RN_334_0;
wire FE_RN_335_0;
wire FE_RN_336_0;
wire FE_RN_337_0;
wire FE_RN_338_0;
wire FE_RN_339_0;
wire FE_RN_33_0;
wire FE_RN_340_0;
wire FE_RN_341_0;
wire FE_RN_342_0;
wire FE_RN_343_0;
wire FE_RN_344_0;
wire FE_RN_345_0;
wire FE_RN_346_0;
wire FE_RN_347_0;
wire FE_RN_348_0;
wire FE_RN_349_0;
wire FE_RN_34_0;
wire FE_RN_350_0;
wire FE_RN_351_0;
wire FE_RN_352_0;
wire FE_RN_353_0;
wire FE_RN_354_0;
wire FE_RN_355_0;
wire FE_RN_356_0;
wire FE_RN_357_0;
wire FE_RN_358_0;
wire FE_RN_359_0;
wire FE_RN_35_0;
wire FE_RN_360_0;
wire FE_RN_361_0;
wire FE_RN_362_0;
wire TIMEBOOST_net_11813;
wire FE_RN_364_0;
wire FE_RN_365_0;
wire FE_RN_366_0;
wire FE_RN_367_0;
wire FE_RN_368_0;
wire FE_RN_369_0;
wire FE_RN_36_0;
wire FE_RN_370_0;
wire FE_RN_371_0;
wire TIMEBOOST_net_11184;
wire FE_RN_373_0;
wire FE_RN_374_0;
wire TIMEBOOST_net_11185;
wire FE_RN_376_0;
wire FE_RN_377_0;
wire TIMEBOOST_net_5279;
wire TIMEBOOST_net_3736;
wire FE_RN_37_0;
wire TIMEBOOST_net_14915;
wire FE_RN_381_0;
wire FE_RN_382_0;
wire FE_RN_383_0;
wire FE_RN_384_0;
wire FE_RN_385_0;
wire FE_RN_386_0;
wire FE_RN_387_0;
wire FE_RN_388_0;
wire FE_RN_389_0;
wire TIMEBOOST_net_12429;
wire FE_RN_390_0;
wire FE_RN_392_0;
wire FE_RN_393_0;
wire FE_RN_394_0;
wire FE_RN_395_0;
wire FE_RN_396_0;
wire FE_RN_397_0;
wire FE_RN_398_0;
wire FE_RN_399_0;
wire FE_RN_39_0;
wire FE_RN_400_0;
wire FE_RN_401_0;
wire FE_RN_402_0;
wire FE_RN_403_0;
wire FE_RN_404_0;
wire FE_RN_405_0;
wire FE_RN_406_0;
wire FE_RN_407_0;
wire FE_RN_409_0;
wire FE_RN_40_0;
wire FE_RN_410_0;
wire FE_RN_411_0;
wire TIMEBOOST_net_10089;
wire FE_RN_413_0;
wire TIMEBOOST_net_12859;
wire FE_RN_415_0;
wire FE_RN_416_0;
wire FE_RN_417_0;
wire FE_RN_418_0;
wire FE_RN_419_0;
wire FE_RN_41_0;
wire FE_RN_420_0;
wire FE_RN_421_0;
wire FE_RN_422_0;
wire FE_RN_423_0;
wire TIMEBOOST_net_1168;
wire FE_RN_425_0;
wire FE_RN_426_0;
wire FE_RN_427_0;
wire FE_RN_428_0;
wire FE_RN_429_0;
wire FE_RN_42_0;
wire FE_RN_430_0;
wire FE_RN_431_0;
wire FE_RN_432_0;
wire FE_RN_433_0;
wire FE_RN_434_0;
wire FE_RN_435_0;
wire TIMEBOOST_net_10272;
wire FE_RN_437_0;
wire FE_RN_438_0;
wire FE_RN_439_0;
wire FE_RN_43_0;
wire FE_RN_440_0;
wire FE_RN_441_0;
wire FE_RN_442_0;
wire FE_RN_443_0;
wire FE_RN_444_0;
wire FE_RN_445_0;
wire FE_RN_446_0;
wire FE_RN_447_0;
wire FE_RN_448_0;
wire FE_RN_449_0;
wire FE_RN_44_0;
wire FE_RN_450_0;
wire TIMEBOOST_net_1169;
wire FE_RN_452_0;
wire FE_RN_453_0;
wire FE_RN_454_0;
wire FE_RN_455_0;
wire FE_RN_456_0;
wire FE_RN_457_0;
wire FE_RN_458_0;
wire FE_RN_459_0;
wire FE_RN_45_0;
wire FE_RN_460_0;
wire FE_RN_462_0;
wire FE_RN_463_0;
wire FE_RN_464_0;
wire FE_RN_465_0;
wire FE_RN_466_0;
wire FE_RN_467_0;
wire FE_RN_468_0;
wire FE_RN_469_0;
wire FE_RN_46_0;
wire FE_RN_470_0;
wire FE_RN_471_0;
wire FE_RN_472_0;
wire FE_RN_473_0;
wire FE_RN_474_0;
wire FE_RN_475_0;
wire FE_RN_476_0;
wire FE_RN_477_0;
wire FE_RN_478_0;
wire FE_RN_479_0;
wire FE_RN_47_0;
wire FE_RN_480_0;
wire FE_RN_481_0;
wire FE_RN_483_0;
wire FE_RN_484_0;
wire FE_RN_486_0;
wire FE_RN_489_0;
wire FE_RN_48_0;
wire FE_RN_490_0;
wire FE_RN_491_0;
wire FE_RN_493_0;
wire FE_RN_494_0;
wire TIMEBOOST_net_9468;
wire FE_RN_496_0;
wire TIMEBOOST_net_15161;
wire FE_RN_498_0;
wire FE_RN_49_0;
wire FE_RN_500_0;
wire FE_RN_501_0;
wire FE_RN_502_0;
wire FE_RN_503_0;
wire FE_RN_505_0;
wire FE_RN_506_0;
wire FE_RN_507_0;
wire FE_RN_508_0;
wire FE_RN_509_0;
wire TIMEBOOST_net_13278;
wire FE_RN_510_0;
wire FE_RN_511_0;
wire FE_RN_512_0;
wire FE_RN_513_0;
wire FE_RN_514_0;
wire FE_RN_515_0;
wire FE_RN_516_0;
wire FE_RN_517_0;
wire FE_RN_518_0;
wire FE_RN_519_0;
wire FE_RN_51_0;
wire FE_RN_520_0;
wire FE_RN_521_0;
wire FE_RN_522_0;
wire FE_RN_523_0;
wire FE_RN_524_0;
wire FE_RN_525_0;
wire FE_RN_526_0;
wire FE_RN_527_0;
wire FE_RN_528_0;
wire FE_RN_529_0;
wire FE_RN_52_0;
wire FE_RN_530_0;
wire FE_RN_531_0;
wire FE_RN_532_0;
wire FE_RN_533_0;
wire TIMEBOOST_net_174;
wire FE_RN_535_0;
wire TIMEBOOST_net_14498;
wire FE_RN_538_0;
wire FE_RN_539_0;
wire FE_RN_53_0;
wire TIMEBOOST_net_11884;
wire FE_RN_541_0;
wire FE_RN_542_0;
wire TIMEBOOST_net_11186;
wire FE_RN_544_0;
wire FE_RN_545_0;
wire TIMEBOOST_net_11187;
wire FE_RN_547_0;
wire FE_RN_548_0;
wire FE_RN_549_0;
wire TIMEBOOST_net_7;
wire FE_RN_551_0;
wire TIMEBOOST_net_14707;
wire FE_RN_553_0;
wire FE_RN_554_0;
wire FE_RN_555_0;
wire FE_RN_556_0;
wire FE_RN_557_0;
wire FE_RN_558_0;
wire FE_RN_559_0;
wire FE_RN_55_0;
wire FE_RN_560_0;
wire FE_RN_561_0;
wire FE_RN_562_0;
wire TIMEBOOST_net_10866;
wire FE_RN_564_0;
wire FE_RN_565_0;
wire FE_RN_566_0;
wire FE_RN_567_0;
wire FE_RN_568_0;
wire FE_RN_569_0;
wire FE_RN_56_0;
wire FE_RN_570_0;
wire FE_RN_571_0;
wire FE_RN_572_0;
wire FE_RN_573_0;
wire TIMEBOOST_net_12959;
wire TIMEBOOST_net_9376;
wire TIMEBOOST_net_13064;
wire TIMEBOOST_net_12824;
wire FE_RN_578_0;
wire TIMEBOOST_net_12416;
wire FE_RN_57_0;
wire TIMEBOOST_net_9677;
wire FE_RN_581_0;
wire FE_RN_582_0;
wire FE_RN_583_0;
wire FE_RN_584_0;
wire TIMEBOOST_net_14816;
wire TIMEBOOST_net_10944;
wire TIMEBOOST_net_14007;
wire TIMEBOOST_net_12897;
wire FE_RN_589_0;
wire FE_RN_58_0;
wire FE_RN_590_0;
wire FE_RN_591_0;
wire FE_RN_592_0;
wire FE_RN_593_0;
wire FE_RN_594_0;
wire FE_RN_595_0;
wire FE_RN_596_0;
wire FE_RN_597_0;
wire FE_RN_598_0;
wire n_2160;
wire TIMEBOOST_net_12665;
wire FE_RN_600_0;
wire FE_RN_601_0;
wire FE_RN_602_0;
wire FE_RN_603_0;
wire FE_RN_604_0;
wire FE_RN_605_0;
wire FE_RN_606_0;
wire FE_RN_607_0;
wire FE_RN_608_0;
wire FE_RN_609_0;
wire FE_RN_60_0;
wire FE_RN_610_0;
wire FE_RN_611_0;
wire FE_RN_612_0;
wire FE_RN_613_0;
wire FE_RN_614_0;
wire FE_RN_615_0;
wire FE_RN_616_0;
wire FE_RN_617_0;
wire FE_RN_618_0;
wire FE_RN_619_0;
wire FE_RN_61_0;
wire FE_RN_620_0;
wire FE_RN_621_0;
wire FE_RN_622_0;
wire FE_RN_623_0;
wire TIMEBOOST_net_12728;
wire TIMEBOOST_net_14986;
wire FE_RN_626_0;
wire FE_RN_627_0;
wire FE_RN_628_0;
wire TIMEBOOST_net_104;
wire TIMEBOOST_net_14203;
wire TIMEBOOST_net_12690;
wire FE_RN_631_0;
wire FE_RN_632_0;
wire FE_RN_633_0;
wire TIMEBOOST_net_12635;
wire TIMEBOOST_net_14822;
wire FE_RN_636_0;
wire FE_RN_637_0;
wire FE_RN_638_0;
wire TIMEBOOST_net_9385;
wire FE_RN_63_0;
wire TIMEBOOST_net_12680;
wire FE_RN_641_0;
wire FE_RN_642_0;
wire FE_RN_643_0;
wire FE_RN_644_0;
wire FE_RN_645_0;
wire FE_RN_646_0;
wire FE_RN_647_0;
wire FE_RN_648_0;
wire FE_RN_649_0;
wire FE_RN_64_0;
wire FE_RN_650_0;
wire FE_RN_651_0;
wire FE_RN_653_0;
wire FE_RN_654_0;
wire FE_RN_655_0;
wire FE_RN_656_0;
wire FE_RN_657_0;
wire FE_RN_659_0;
wire TIMEBOOST_net_2873;
wire FE_RN_660_0;
wire FE_RN_661_0;
wire FE_RN_662_0;
wire FE_RN_663_0;
wire FE_RN_665_0;
wire FE_RN_666_0;
wire FE_RN_667_0;
wire FE_RN_668_0;
wire FE_RN_669_0;
wire FE_RN_66_0;
wire FE_RN_670_0;
wire FE_RN_671_0;
wire FE_RN_672_0;
wire FE_RN_673_0;
wire FE_RN_674_0;
wire FE_RN_675_0;
wire TIMEBOOST_net_24;
wire FE_RN_677_0;
wire FE_RN_678_0;
wire TIMEBOOST_net_12706;
wire FE_RN_67_0;
wire FE_RN_680_0;
wire FE_RN_681_0;
wire FE_RN_682_0;
wire FE_RN_683_0;
wire FE_RN_684_0;
wire FE_RN_685_0;
wire FE_RN_686_0;
wire TIMEBOOST_net_12729;
wire FE_RN_688_0;
wire FE_RN_689_0;
wire TIMEBOOST_net_13280;
wire TIMEBOOST_net_14981;
wire FE_RN_691_0;
wire FE_RN_693_0;
wire FE_RN_694_0;
wire FE_RN_695_0;
wire FE_RN_697_0;
wire FE_RN_698_0;
wire FE_RN_699_0;
wire FE_RN_69_0;
wire FE_RN_6_0;
wire FE_RN_700_0;
wire FE_RN_701_0;
wire FE_RN_702_0;
wire FE_RN_703_0;
wire FE_RN_704_0;
wire FE_RN_705_0;
wire TIMEBOOST_net_869;
wire FE_RN_707_0;
wire FE_RN_708_0;
wire FE_RN_709_0;
wire FE_RN_70_0;
wire FE_RN_710_0;
wire FE_RN_711_0;
wire TIMEBOOST_net_11183;
wire FE_RN_713_0;
wire FE_RN_714_0;
wire FE_RN_715_0;
wire FE_RN_716_0;
wire FE_RN_717_0;
wire TIMEBOOST_net_12964;
wire FE_RN_71_0;
wire FE_RN_720_0;
wire FE_RN_722_0;
wire FE_RN_723_0;
wire TIMEBOOST_net_13853;
wire FE_RN_725_0;
wire FE_RN_726_0;
wire TIMEBOOST_net_12999;
wire FE_RN_728_0;
wire FE_RN_729_0;
wire FE_RN_72_0;
wire TIMEBOOST_net_13001;
wire FE_RN_731_0;
wire FE_RN_732_0;
wire TIMEBOOST_net_14280;
wire FE_RN_734_0;
wire FE_RN_735_0;
wire FE_RN_736_0;
wire FE_RN_737_0;
wire FE_RN_738_0;
wire FE_RN_739_0;
wire FE_RN_73_0;
wire FE_RN_740_0;
wire FE_RN_741_0;
wire FE_RN_742_0;
wire FE_RN_743_0;
wire FE_RN_744_0;
wire FE_RN_745_0;
wire FE_RN_746_0;
wire FE_RN_747_0;
wire FE_RN_748_0;
wire FE_RN_749_0;
wire TIMEBOOST_net_3515;
wire FE_RN_750_0;
wire FE_RN_751_0;
wire FE_RN_752_0;
wire FE_RN_753_0;
wire FE_RN_754_0;
wire FE_RN_755_0;
wire FE_RN_756_0;
wire FE_RN_758_0;
wire FE_RN_759_0;
wire FE_RN_764_0;
wire FE_RN_767_0;
wire FE_RN_768_0;
wire FE_RN_769_0;
wire TIMEBOOST_net_12952;
wire FE_RN_772_0;
wire FE_RN_773_0;
wire FE_RN_774_0;
wire FE_RN_775_0;
wire FE_RN_776_0;
wire FE_RN_778_0;
wire FE_RN_779_0;
wire FE_RN_780_0;
wire FE_RN_795_0;
wire FE_RN_796_0;
wire FE_RN_797_0;
wire FE_RN_798_0;
wire TIMEBOOST_net_2874;
wire FE_RN_7_0;
wire FE_RN_800_0;
wire FE_RN_801_0;
wire FE_RN_802_0;
wire TIMEBOOST_net_12947;
wire TIMEBOOST_net_12948;
wire FE_RN_805_0;
wire FE_RN_806_0;
wire FE_RN_807_0;
wire TIMEBOOST_net_13181;
wire FE_RN_809_0;
wire FE_RN_810_0;
wire FE_RN_811_0;
wire FE_RN_812_0;
wire TIMEBOOST_net_12951;
wire FE_RN_814_0;
wire FE_RN_815_0;
wire FE_RN_816_0;
wire FE_RN_817_0;
wire FE_RN_818_0;
wire FE_RN_81_0;
wire FE_RN_820_0;
wire FE_RN_821_0;
wire FE_RN_822_0;
wire FE_RN_824_0;
wire TIMEBOOST_net_9408;
wire TIMEBOOST_net_14283;
wire FE_RN_827_0;
wire FE_RN_828_0;
wire FE_RN_829_0;
wire FE_RN_82_0;
wire TIMEBOOST_net_12936;
wire FE_RN_831_0;
wire FE_RN_832_0;
wire FE_RN_833_0;
wire TIMEBOOST_net_12618;
wire FE_RN_835_0;
wire FE_RN_836_0;
wire FE_RN_837_0;
wire FE_RN_838_0;
wire FE_RN_839_0;
wire FE_RN_83_0;
wire FE_RN_840_0;
wire TIMEBOOST_net_709;
wire TIMEBOOST_net_13234;
wire FE_RN_843_0;
wire FE_RN_844_0;
wire FE_RN_845_0;
wire TIMEBOOST_net_12617;
wire FE_RN_847_0;
wire FE_RN_862_0;
wire FE_RN_863_0;
wire FE_RN_87_0;
wire FE_RN_880_0;
wire FE_RN_881_0;
wire FE_RN_882_0;
wire FE_RN_883_0;
wire FE_RN_887_0;
wire FE_RN_888_0;
wire FE_RN_88_0;
wire FE_RN_890_0;
wire FE_RN_893_0;
wire FE_RN_894_0;
wire FE_RN_895_0;
wire FE_RN_896_0;
wire FE_RN_897_0;
wire FE_RN_898_0;
wire FE_RN_899_0;
wire FE_RN_89_0;
wire FE_RN_8_0;
wire FE_RN_900_0;
wire FE_RN_901_0;
wire FE_RN_902_0;
wire FE_RN_904_0;
wire FE_RN_905_0;
wire FE_RN_906_0;
wire FE_RN_907_0;
wire FE_RN_908_0;
wire FE_RN_909_0;
wire FE_RN_90_0;
wire FE_RN_910_0;
wire FE_RN_911_0;
wire FE_RN_912_0;
wire FE_RN_913_0;
wire FE_RN_914_0;
wire FE_RN_915_0;
wire FE_RN_916_0;
wire FE_RN_917_0;
wire FE_RN_91_0;
wire FE_RN_92_0;
wire FE_RN_93_0;
wire FE_RN_94_0;
wire FE_RN_95_0;
wire FE_RN_96_0;
wire FE_RN_97_0;
wire FE_RN_98_0;
wire FE_RN_99_0;
wire FE_RN_9_0;
wire conf_pci_init_complete_out;
wire conf_target_abort_recv_in;
wire conf_w_addr_in;
wire conf_w_addr_in_931;
wire conf_w_addr_in_932;
wire conf_w_addr_in_933;
wire conf_w_addr_in_935;
wire conf_w_addr_in_937;
wire conf_w_addr_in_938;
wire conf_w_addr_in_939;
wire conf_wb_err_addr_in_943;
wire conf_wb_err_addr_in_944;
wire conf_wb_err_addr_in_945;
wire conf_wb_err_addr_in_946;
wire conf_wb_err_addr_in_947;
wire conf_wb_err_addr_in_948;
wire conf_wb_err_addr_in_949;
wire conf_wb_err_addr_in_950;
wire conf_wb_err_addr_in_951;
wire conf_wb_err_addr_in_952;
wire conf_wb_err_addr_in_953;
wire conf_wb_err_addr_in_954;
wire conf_wb_err_addr_in_955;
wire conf_wb_err_addr_in_956;
wire conf_wb_err_addr_in_957;
wire conf_wb_err_addr_in_958;
wire conf_wb_err_addr_in_959;
wire conf_wb_err_addr_in_960;
wire conf_wb_err_addr_in_961;
wire conf_wb_err_addr_in_962;
wire conf_wb_err_addr_in_963;
wire conf_wb_err_addr_in_964;
wire conf_wb_err_addr_in_965;
wire conf_wb_err_addr_in_966;
wire conf_wb_err_addr_in_967;
wire conf_wb_err_addr_in_968;
wire conf_wb_err_addr_in_969;
wire conf_wb_err_addr_in_970;
wire conf_wb_err_addr_in_971;
wire conf_wb_err_bc_in;
wire conf_wb_err_bc_in_846;
wire conf_wb_err_bc_in_847;
wire conf_wb_err_bc_in_848;
wire configuration_cache_line_size_reg;
wire configuration_cache_line_size_reg_2996;
wire configuration_command_bit;
wire configuration_icr_bit2_0;
wire configuration_icr_bit_2961;
wire configuration_icr_bit_2967;
wire configuration_int_meta;
wire configuration_interrupt_line;
wire configuration_interrupt_line_37;
wire configuration_interrupt_line_38;
wire configuration_interrupt_line_39;
wire configuration_interrupt_line_40;
wire configuration_interrupt_line_41;
wire configuration_interrupt_line_42;
wire configuration_interrupt_line_43;
wire configuration_interrupt_out_reg_Q;
wire configuration_isr_bit_1457;
wire configuration_isr_bit_1461;
wire configuration_isr_bit_2975;
wire configuration_isr_bit_618;
wire configuration_isr_bit_631;
wire configuration_meta_cache_lsize_to_wb_bits;
wire configuration_meta_cache_lsize_to_wb_bits_926;
wire configuration_meta_cache_lsize_to_wb_bits_927;
wire configuration_meta_cache_lsize_to_wb_bits_928;
wire configuration_meta_cache_lsize_to_wb_bits_929;
wire configuration_meta_cache_lsize_to_wb_bits_930;
wire configuration_meta_cache_lsize_to_wb_bits_931;
wire configuration_meta_command_bit;
wire configuration_meta_pci_err_cs_bits;
wire configuration_pci_err_addr;
wire configuration_pci_err_addr_471;
wire configuration_pci_err_addr_472;
wire configuration_pci_err_addr_473;
wire configuration_pci_err_addr_474;
wire configuration_pci_err_addr_475;
wire configuration_pci_err_addr_476;
wire configuration_pci_err_addr_477;
wire configuration_pci_err_addr_478;
wire configuration_pci_err_addr_479;
wire configuration_pci_err_addr_480;
wire configuration_pci_err_addr_481;
wire configuration_pci_err_addr_482;
wire configuration_pci_err_addr_483;
wire configuration_pci_err_addr_484;
wire configuration_pci_err_addr_485;
wire configuration_pci_err_addr_486;
wire configuration_pci_err_addr_487;
wire configuration_pci_err_addr_488;
wire configuration_pci_err_addr_489;
wire configuration_pci_err_addr_490;
wire configuration_pci_err_addr_491;
wire configuration_pci_err_addr_492;
wire configuration_pci_err_addr_493;
wire configuration_pci_err_addr_494;
wire configuration_pci_err_addr_495;
wire configuration_pci_err_addr_496;
wire configuration_pci_err_addr_497;
wire configuration_pci_err_addr_498;
wire configuration_pci_err_addr_499;
wire configuration_pci_err_addr_500;
wire configuration_pci_err_addr_501;
wire configuration_pci_err_cs_bit0;
wire configuration_pci_err_cs_bit10;
wire configuration_pci_err_cs_bit31_24;
wire configuration_pci_err_cs_bit8;
wire configuration_pci_err_cs_bit9;
wire configuration_pci_err_cs_bit_464;
wire configuration_pci_err_cs_bit_465;
wire configuration_pci_err_cs_bit_466;
wire configuration_pci_err_cs_bit_467;
wire configuration_pci_err_cs_bit_468;
wire configuration_pci_err_cs_bit_469;
wire configuration_pci_err_cs_bit_470;
wire configuration_pci_err_data;
wire configuration_pci_err_data_502;
wire configuration_pci_err_data_503;
wire configuration_pci_err_data_504;
wire configuration_pci_err_data_505;
wire configuration_pci_err_data_506;
wire configuration_pci_err_data_507;
wire configuration_pci_err_data_508;
wire configuration_pci_err_data_509;
wire configuration_pci_err_data_510;
wire configuration_pci_err_data_511;
wire configuration_pci_err_data_512;
wire configuration_pci_err_data_513;
wire configuration_pci_err_data_514;
wire configuration_pci_err_data_515;
wire configuration_pci_err_data_516;
wire configuration_pci_err_data_517;
wire configuration_pci_err_data_518;
wire configuration_pci_err_data_519;
wire configuration_pci_err_data_520;
wire configuration_pci_err_data_521;
wire configuration_pci_err_data_522;
wire configuration_pci_err_data_523;
wire configuration_pci_err_data_524;
wire configuration_pci_err_data_525;
wire configuration_pci_err_data_526;
wire configuration_pci_err_data_527;
wire configuration_pci_err_data_528;
wire configuration_pci_err_data_529;
wire configuration_pci_err_data_530;
wire configuration_pci_err_data_531;
wire configuration_pci_err_data_532;
wire configuration_rst_inactive;
wire configuration_rst_inactive_sync;
wire configuration_set_isr_bit2;
wire configuration_set_isr_bit2_reg_Q;
wire configuration_set_pci_err_cs_bit8;
wire configuration_set_pci_err_cs_bit8_reg_Q;
wire configuration_status_bit8;
wire configuration_status_bit_322;
wire configuration_status_bit_351;
wire configuration_status_bit_379;
wire configuration_status_bit_407;
wire configuration_status_bit_435;
wire configuration_sync_cache_lsize_to_wb_bits_reg_2__Q;
wire configuration_sync_cache_lsize_to_wb_bits_reg_3__Q;
wire configuration_sync_cache_lsize_to_wb_bits_reg_4__Q;
wire configuration_sync_command_bit0;
wire configuration_sync_command_bit1;
wire configuration_sync_command_bit2;
wire configuration_sync_command_bit6;
wire configuration_sync_command_bit8;
wire configuration_sync_init_complete;
wire configuration_sync_isr_2_del_bit_reg_Q;
wire configuration_sync_isr_2_delayed_bckp_bit;
wire configuration_sync_isr_2_delayed_bckp_bit_reg_Q;
wire configuration_sync_isr_2_delayed_del_bit;
wire configuration_sync_isr_2_delayed_del_bit_reg_Q;
wire configuration_sync_isr_2_meta_bckp_bit;
wire configuration_sync_isr_2_meta_del_bit;
wire configuration_sync_isr_2_sync_bckp_bit;
wire configuration_sync_isr_2_sync_del_bit;
wire configuration_sync_pci_err_cs_8_del_bit_reg_Q;
wire configuration_sync_pci_err_cs_8_delayed_bckp_bit;
wire configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg_Q;
wire configuration_sync_pci_err_cs_8_delayed_del_bit;
wire configuration_sync_pci_err_cs_8_delayed_del_bit_reg_Q;
wire configuration_sync_pci_err_cs_8_meta_bckp_bit;
wire configuration_sync_pci_err_cs_8_meta_del_bit;
wire configuration_sync_pci_err_cs_8_sync_bckp_bit;
wire configuration_sync_pci_err_cs_8_sync_del_bit;
wire configuration_wb_err_addr;
wire configuration_wb_err_addr_533;
wire configuration_wb_err_addr_534;
wire configuration_wb_err_addr_535;
wire configuration_wb_err_addr_536;
wire configuration_wb_err_addr_537;
wire configuration_wb_err_addr_538;
wire configuration_wb_err_addr_539;
wire configuration_wb_err_addr_540;
wire configuration_wb_err_addr_541;
wire configuration_wb_err_addr_542;
wire configuration_wb_err_addr_543;
wire configuration_wb_err_addr_544;
wire configuration_wb_err_addr_545;
wire configuration_wb_err_addr_546;
wire configuration_wb_err_addr_547;
wire configuration_wb_err_addr_548;
wire configuration_wb_err_addr_549;
wire configuration_wb_err_addr_550;
wire configuration_wb_err_addr_551;
wire configuration_wb_err_addr_552;
wire configuration_wb_err_addr_553;
wire configuration_wb_err_addr_554;
wire configuration_wb_err_addr_555;
wire configuration_wb_err_addr_556;
wire configuration_wb_err_addr_557;
wire configuration_wb_err_addr_558;
wire configuration_wb_err_addr_559;
wire configuration_wb_err_addr_560;
wire configuration_wb_err_addr_561;
wire configuration_wb_err_addr_562;
wire configuration_wb_err_addr_563;
wire configuration_wb_err_cs_bit0;
wire configuration_wb_err_cs_bit31_24;
wire configuration_wb_err_cs_bit8;
wire configuration_wb_err_cs_bit9;
wire configuration_wb_err_cs_bit_564;
wire configuration_wb_err_cs_bit_565;
wire configuration_wb_err_cs_bit_566;
wire configuration_wb_err_cs_bit_567;
wire configuration_wb_err_cs_bit_568;
wire configuration_wb_err_cs_bit_569;
wire configuration_wb_err_cs_bit_570;
wire configuration_wb_err_data;
wire configuration_wb_err_data_571;
wire configuration_wb_err_data_572;
wire configuration_wb_err_data_573;
wire configuration_wb_err_data_574;
wire configuration_wb_err_data_575;
wire configuration_wb_err_data_576;
wire configuration_wb_err_data_577;
wire configuration_wb_err_data_578;
wire configuration_wb_err_data_579;
wire configuration_wb_err_data_580;
wire configuration_wb_err_data_581;
wire configuration_wb_err_data_582;
wire configuration_wb_err_data_583;
wire configuration_wb_err_data_584;
wire configuration_wb_err_data_585;
wire configuration_wb_err_data_586;
wire configuration_wb_err_data_587;
wire configuration_wb_err_data_588;
wire configuration_wb_err_data_589;
wire configuration_wb_err_data_590;
wire configuration_wb_err_data_591;
wire configuration_wb_err_data_592;
wire configuration_wb_err_data_593;
wire configuration_wb_err_data_594;
wire configuration_wb_err_data_595;
wire configuration_wb_err_data_596;
wire configuration_wb_err_data_597;
wire configuration_wb_err_data_598;
wire configuration_wb_err_data_599;
wire configuration_wb_err_data_600;
wire configuration_wb_err_data_601;
wire g15_p;
wire g17_p;
wire g22_p;
wire g52252_p;
wire g52253_p;
wire TIMEBOOST_net_13944;
wire TIMEBOOST_net_11145;
wire g52393_sb;
wire TIMEBOOST_net_13941;
wire TIMEBOOST_net_11146;
wire g52394_sb;
wire TIMEBOOST_net_14022;
wire TIMEBOOST_net_10731;
wire g52395_sb;
wire TIMEBOOST_net_14041;
wire g52396_db;
wire g52396_sb;
wire TIMEBOOST_net_14078;
wire g52397_db;
wire g52397_sb;
wire TIMEBOOST_net_14299;
wire g52398_db;
wire g52398_sb;
wire TIMEBOOST_net_14258;
wire g52399_db;
wire g52399_sb;
wire TIMEBOOST_net_14240;
wire g52400_db;
wire g52400_sb;
wire TIMEBOOST_net_14374;
wire g52401_db;
wire g52401_sb;
wire TIMEBOOST_net_14013;
wire TIMEBOOST_net_10811;
wire g52402_sb;
wire TIMEBOOST_net_13947;
wire g52403_db;
wire g52403_sb;
wire TIMEBOOST_net_14296;
wire g52404_db;
wire g52404_sb;
wire TIMEBOOST_net_14259;
wire TIMEBOOST_net_13757;
wire g52405_sb;
wire TIMEBOOST_net_14304;
wire TIMEBOOST_net_10600;
wire TIMEBOOST_net_13939;
wire g52440_db;
wire g52440_sb;
wire TIMEBOOST_net_14021;
wire TIMEBOOST_net_10737;
wire g52441_sb;
wire TIMEBOOST_net_14291;
wire TIMEBOOST_net_13791;
wire g52442_sb;
wire TIMEBOOST_net_14018;
wire g52443_db;
wire g52443_sb;
wire TIMEBOOST_net_14019;
wire TIMEBOOST_net_10781;
wire g52444_sb;
wire TIMEBOOST_net_14322;
wire g52445_db;
wire TIMEBOOST_net_14086;
wire TIMEBOOST_net_11162;
wire g52446_sb;
wire TIMEBOOST_net_14564;
wire g52447_db;
wire g52447_sb;
wire TIMEBOOST_net_14617;
wire g52448_db;
wire g52448_sb;
wire TIMEBOOST_net_13940;
wire g52449_db;
wire g52449_sb;
wire TIMEBOOST_net_13952;
wire g52450_db;
wire g52450_sb;
wire TIMEBOOST_net_14330;
wire g52451_db;
wire g52451_sb;
wire TIMEBOOST_net_14083;
wire TIMEBOOST_net_13761;
wire g52452_sb;
wire TIMEBOOST_net_14288;
wire TIMEBOOST_net_10812;
wire TIMEBOOST_net_13985;
wire g52454_db;
wire g52454_sb;
wire TIMEBOOST_net_13984;
wire g52455_db;
wire g52455_sb;
wire g52456_da;
wire TIMEBOOST_net_12847;
wire g52456_sb;
wire g52457_da;
wire g65240_da;
wire g52457_sb;
wire g52458_da;
wire g65236_da;
wire g52458_sb;
wire TIMEBOOST_net_14343;
wire TIMEBOOST_net_12895;
wire g52459_sb;
wire g52460_da;
wire TIMEBOOST_net_1441;
wire g52460_sb;
wire g52461_da;
wire TIMEBOOST_net_12850;
wire g52461_sb;
wire TIMEBOOST_net_14650;
wire TIMEBOOST_net_12890;
wire g52462_sb;
wire g52463_da;
wire TIMEBOOST_net_12851;
wire g52463_sb;
wire g52464_da;
wire TIMEBOOST_net_12852;
wire g52464_sb;
wire g52465_da;
wire TIMEBOOST_net_13169;
wire g52466_da;
wire TIMEBOOST_net_13135;
wire g52466_sb;
wire g52467_da;
wire TIMEBOOST_net_12891;
wire TIMEBOOST_net_14647;
wire TIMEBOOST_net_12949;
wire g52469_da;
wire TIMEBOOST_net_13170;
wire g52470_da;
wire TIMEBOOST_net_13123;
wire g52470_sb;
wire g52471_da;
wire TIMEBOOST_net_12885;
wire g52472_da;
wire TIMEBOOST_net_12881;
wire g52473_da;
wire g65235_da;
wire g52474_da;
wire TIMEBOOST_net_12860;
wire TIMEBOOST_net_12961;
wire TIMEBOOST_net_12965;
wire g52476_da;
wire TIMEBOOST_net_12861;
wire g52476_sb;
wire g52477_da;
wire TIMEBOOST_net_1439;
wire g52477_sb;
wire g52478_da;
wire TIMEBOOST_net_12869;
wire g52478_sb;
wire g52479_da;
wire TIMEBOOST_net_12967;
wire g52479_sb;
wire g52480_da;
wire TIMEBOOST_net_12957;
wire g52481_da;
wire TIMEBOOST_net_13139;
wire g52482_da;
wire TIMEBOOST_net_2805;
wire g52482_sb;
wire g52483_da;
wire TIMEBOOST_net_13175;
wire g52484_da;
wire TIMEBOOST_net_13136;
wire g52485_da;
wire TIMEBOOST_net_12889;
wire g52495_p;
wire g52496_p;
wire g52497_p;
wire g52498_p;
wire TIMEBOOST_net_15156;
wire TIMEBOOST_net_14795;
wire g52503_sb;
wire TIMEBOOST_net_6210;
wire TIMEBOOST_net_13230;
wire g52504_sb;
wire TIMEBOOST_net_15160;
wire TIMEBOOST_net_12925;
wire g52505_sb;
wire TIMEBOOST_net_15175;
wire TIMEBOOST_net_13231;
wire g52506_sb;
wire TIMEBOOST_net_15085;
wire TIMEBOOST_net_12929;
wire g52507_sb;
wire TIMEBOOST_net_15138;
wire TIMEBOOST_net_12926;
wire g52508_sb;
wire TIMEBOOST_net_12950;
wire g52509_sb;
wire TIMEBOOST_net_15153;
wire TIMEBOOST_net_12928;
wire g52510_sb;
wire TIMEBOOST_net_15164;
wire TIMEBOOST_net_12916;
wire g52511_sb;
wire TIMEBOOST_net_15165;
wire TIMEBOOST_net_12921;
wire g52512_sb;
wire TIMEBOOST_net_15204;
wire TIMEBOOST_net_12919;
wire g52513_sb;
wire TIMEBOOST_net_15166;
wire TIMEBOOST_net_12917;
wire g52514_sb;
wire TIMEBOOST_net_13156;
wire g52515_sb;
wire g65216_da;
wire g52516_sb;
wire TIMEBOOST_net_12934;
wire g52517_sb;
wire TIMEBOOST_net_15167;
wire n_1598;
wire g52518_sb;
wire TIMEBOOST_net_15148;
wire TIMEBOOST_net_13244;
wire g52519_sb;
wire TIMEBOOST_net_15168;
wire TIMEBOOST_net_12898;
wire g52520_sb;
wire TIMEBOOST_net_15169;
wire TIMEBOOST_net_12901;
wire g52521_sb;
wire TIMEBOOST_net_15170;
wire TIMEBOOST_net_12900;
wire g52522_sb;
wire TIMEBOOST_net_15171;
wire TIMEBOOST_net_12906;
wire g52523_sb;
wire TIMEBOOST_net_15172;
wire TIMEBOOST_net_12892;
wire g52524_sb;
wire TIMEBOOST_net_13162;
wire g52525_sb;
wire TIMEBOOST_net_15140;
wire TIMEBOOST_net_12899;
wire g52526_sb;
wire g64827_db;
wire g52527_sb;
wire TIMEBOOST_net_13167;
wire g52528_sb;
wire TIMEBOOST_net_15149;
wire TIMEBOOST_net_13245;
wire g52529_sb;
wire TIMEBOOST_net_13168;
wire g52530_sb;
wire TIMEBOOST_net_15150;
wire TIMEBOOST_net_13246;
wire g52531_sb;
wire TIMEBOOST_net_15151;
wire TIMEBOOST_net_13243;
wire g52532_sb;
wire TIMEBOOST_net_15152;
wire TIMEBOOST_net_13236;
wire g52533_sb;
wire TIMEBOOST_net_15162;
wire TIMEBOOST_net_13226;
wire g52534_sb;
wire TIMEBOOST_net_10951;
wire TIMEBOOST_net_12694;
wire g52590_sb;
wire TIMEBOOST_net_10952;
wire TIMEBOOST_net_12688;
wire g52591_sb;
wire TIMEBOOST_net_10953;
wire TIMEBOOST_net_12647;
wire g52592_sb;
wire TIMEBOOST_net_10954;
wire TIMEBOOST_net_12669;
wire g52593_sb;
wire TIMEBOOST_net_13041;
wire TIMEBOOST_net_15216;
wire g52594_sb;
wire TIMEBOOST_net_12990;
wire TIMEBOOST_net_15261;
wire g52595_sb;
wire TIMEBOOST_net_12997;
wire TIMEBOOST_net_15262;
wire g52596_sb;
wire TIMEBOOST_net_13013;
wire g52597_db;
wire g52597_sb;
wire TIMEBOOST_net_12987;
wire TIMEBOOST_net_15263;
wire g52598_sb;
wire TIMEBOOST_net_12992;
wire TIMEBOOST_net_15264;
wire g52599_sb;
wire TIMEBOOST_net_13015;
wire g52600_db;
wire g52600_sb;
wire TIMEBOOST_net_12993;
wire TIMEBOOST_net_15265;
wire g52601_sb;
wire TIMEBOOST_net_12989;
wire g52602_db;
wire g52602_sb;
wire TIMEBOOST_net_12979;
wire TIMEBOOST_net_15266;
wire g52603_sb;
wire TIMEBOOST_net_13030;
wire TIMEBOOST_net_15217;
wire g52604_sb;
wire TIMEBOOST_net_1540;
wire TIMEBOOST_net_15267;
wire g52605_sb;
wire TIMEBOOST_net_13009;
wire g52606_db;
wire g52606_sb;
wire TIMEBOOST_net_12991;
wire TIMEBOOST_net_15268;
wire g52607_sb;
wire TIMEBOOST_net_1542;
wire TIMEBOOST_net_15269;
wire g52608_sb;
wire TIMEBOOST_net_13019;
wire g52609_sb;
wire TIMEBOOST_net_1555;
wire g52610_sb;
wire TIMEBOOST_net_12962;
wire g52611_sb;
wire TIMEBOOST_net_12963;
wire g52612_sb;
wire TIMEBOOST_net_13004;
wire g52614_db;
wire g52614_sb;
wire TIMEBOOST_net_13020;
wire g52616_sb;
wire TIMEBOOST_net_14184;
wire TIMEBOOST_net_15218;
wire g52617_sb;
wire TIMEBOOST_net_13036;
wire g52618_db;
wire g52618_sb;
wire TIMEBOOST_net_13033;
wire g52619_db;
wire g52619_sb;
wire TIMEBOOST_net_13850;
wire g52620_sb;
wire TIMEBOOST_net_13018;
wire g52621_db;
wire g52621_sb;
wire TIMEBOOST_net_13031;
wire g52622_sb;
wire g52623_p;
wire g52624_da;
wire g52624_db;
wire g52624_sb;
wire TIMEBOOST_net_4495;
wire g52625_db;
wire g52625_sb;
wire g52626_da;
wire TIMEBOOST_net_9938;
wire g52626_sb;
wire TIMEBOOST_net_13279;
wire TIMEBOOST_net_10766;
wire g52627_sb;
wire TIMEBOOST_net_4496;
wire g52628_db;
wire g52628_sb;
wire TIMEBOOST_net_10679;
wire TIMEBOOST_net_15178;
wire g52629_sb;
wire TIMEBOOST_net_4876;
wire TIMEBOOST_net_12392;
wire g52630_sb;
wire g52631_da;
wire TIMEBOOST_net_14428;
wire g52631_sb;
wire g52632_da;
wire g52632_db;
wire g52632_sb;
wire TIMEBOOST_net_10680;
wire g52633_db;
wire g52633_sb;
wire g52634_da;
wire TIMEBOOST_net_9955;
wire g52634_sb;
wire g52635_da;
wire g52635_db;
wire g52635_sb;
wire TIMEBOOST_net_4497;
wire g52636_db;
wire g52636_sb;
wire g52637_da;
wire TIMEBOOST_net_14129;
wire g52637_sb;
wire TIMEBOOST_net_4498;
wire g52638_db;
wire g52638_sb;
wire TIMEBOOST_net_4499;
wire g52639_db;
wire g52639_sb;
wire TIMEBOOST_net_4500;
wire TIMEBOOST_net_14344;
wire TIMEBOOST_net_10655;
wire g52641_db;
wire g52641_sb;
wire TIMEBOOST_net_4633;
wire g52642_db;
wire g52642_sb;
wire g52643_da;
wire g52643_db;
wire g52643_sb;
wire TIMEBOOST_net_10681;
wire g52644_db;
wire g52644_sb;
wire TIMEBOOST_net_13735;
wire g52645_db;
wire g52645_sb;
wire TIMEBOOST_net_10682;
wire g52646_db;
wire g52646_sb;
wire TIMEBOOST_net_3355;
wire TIMEBOOST_net_260;
wire g52647_sb;
wire TIMEBOOST_net_4637;
wire g52648_db;
wire g52648_sb;
wire TIMEBOOST_net_3356;
wire TIMEBOOST_net_12294;
wire g52650_da;
wire TIMEBOOST_net_15177;
wire g52650_sb;
wire TIMEBOOST_net_13736;
wire g52651_db;
wire g52651_sb;
wire TIMEBOOST_net_4502;
wire g52652_db;
wire g52652_sb;
wire TIMEBOOST_net_10492;
wire g52653_db;
wire g52653_sb;
wire g52675_p;
wire g52714_p;
wire g52865_p;
wire TIMEBOOST_net_13933;
wire TIMEBOOST_net_13935;
wire g52876_sb;
wire TIMEBOOST_net_14447;
wire g53897_db;
wire g52877_sb;
wire TIMEBOOST_net_14030;
wire TIMEBOOST_net_13956;
wire g52878_sb;
wire TIMEBOOST_net_10995;
wire TIMEBOOST_net_14087;
wire g52879_sb;
wire TIMEBOOST_net_10997;
wire TIMEBOOST_net_14088;
wire g52880_sb;
wire TIMEBOOST_net_10998;
wire TIMEBOOST_net_14031;
wire g52881_sb;
wire g52_p;
wire g53011_p;
wire g53012_p;
wire g53014_p;
wire g53015_p;
wire g53016_p;
wire g53017_p;
wire g53018_p;
wire g53022_p;
wire g53026_p;
wire g53031_p;
wire g53035_p;
wire g53039_p;
wire g53069_p;
wire g53071_p;
wire g53072_p;
wire g53073_p;
wire g53074_p;
wire g53075_p;
wire g53076_p;
wire g53077_p;
wire g53078_p;
wire g53079_p;
wire g53080_p;
wire g53082_p;
wire g53083_p;
wire g53084_p;
wire g53087_p;
wire g53098_p;
wire TIMEBOOST_net_13040;
wire TIMEBOOST_net_11898;
wire g53141_p;
wire g53142_p;
wire g53154_p;
wire g53155_p;
wire g53158_p;
wire g53159_p;
wire g53163_p;
wire g53167_p;
wire g53170_p;
wire g53171_p;
wire g53174_p;
wire g53175_p;
wire g53182_p;
wire g53183_p;
wire g53187_p;
wire g53199_p;
wire g53203_p;
wire g53206_p;
wire g53207_p;
wire g53210_p;
wire g53211_p;
wire g53214_p;
wire g53222_p;
wire g53223_p;
wire g53226_p;
wire g53230_p;
wire g53231_p;
wire g53234_p;
wire g53235_p;
wire g53238_p;
wire g53239_p;
wire g53242_p;
wire g53243_p;
wire g53250_p;
wire g53251_p;
wire g53254_p;
wire g53255_p;
wire g53258_p;
wire g53259_p;
wire g53262_p;
wire g53263_p;
wire g53267_p;
wire g53268_p;
wire g53275_p;
wire g53276_p;
wire g53288_p;
wire g53289_p;
wire g53298_p;
wire g53301_p;
wire g53302_p;
wire g53310_p;
wire g53314_p;
wire g53709_p;
wire g53726_p;
wire g53729_p;
wire g53752_p;
wire TIMEBOOST_net_648;
wire TIMEBOOST_net_13988;
wire TIMEBOOST_net_10594;
wire g53891_db;
wire TIMEBOOST_net_14349;
wire g53892_db;
wire g53892_sb;
wire TIMEBOOST_net_14119;
wire g53893_db;
wire TIMEBOOST_net_14043;
wire TIMEBOOST_net_10839;
wire g53897_sb;
wire TIMEBOOST_net_11654;
wire TIMEBOOST_net_14054;
wire g53898_sb;
wire TIMEBOOST_net_11656;
wire TIMEBOOST_net_14274;
wire g53899_sb;
wire TIMEBOOST_net_11600;
wire TIMEBOOST_net_14364;
wire g53900_sb;
wire TIMEBOOST_net_11605;
wire TIMEBOOST_net_13961;
wire g53901_sb;
wire TIMEBOOST_net_11608;
wire TIMEBOOST_net_14061;
wire g53902_sb;
wire TIMEBOOST_net_11609;
wire TIMEBOOST_net_14062;
wire g53903_sb;
wire TIMEBOOST_net_11611;
wire TIMEBOOST_net_14460;
wire g53904_sb;
wire TIMEBOOST_net_11620;
wire TIMEBOOST_net_14128;
wire g53905_sb;
wire TIMEBOOST_net_11623;
wire TIMEBOOST_net_14016;
wire g53906_sb;
wire TIMEBOOST_net_11627;
wire TIMEBOOST_net_14555;
wire g53907_sb;
wire TIMEBOOST_net_11599;
wire TIMEBOOST_net_14025;
wire g53908_sb;
wire TIMEBOOST_net_11602;
wire TIMEBOOST_net_14026;
wire g53909_sb;
wire TIMEBOOST_net_11615;
wire TIMEBOOST_net_14032;
wire g53910_sb;
wire TIMEBOOST_net_11625;
wire TIMEBOOST_net_14435;
wire g53911_sb;
wire TIMEBOOST_net_11626;
wire TIMEBOOST_net_13998;
wire g53912_sb;
wire TIMEBOOST_net_11699;
wire TIMEBOOST_net_13999;
wire g53913_sb;
wire TIMEBOOST_net_11700;
wire TIMEBOOST_net_14530;
wire g53914_sb;
wire TIMEBOOST_net_11904;
wire TIMEBOOST_net_14001;
wire g53915_sb;
wire TIMEBOOST_net_11883;
wire TIMEBOOST_net_14438;
wire g53916_sb;
wire TIMEBOOST_net_11494;
wire TIMEBOOST_net_14000;
wire g53917_sb;
wire TIMEBOOST_net_11901;
wire TIMEBOOST_net_14077;
wire g53918_sb;
wire TIMEBOOST_net_11902;
wire TIMEBOOST_net_13993;
wire g53919_sb;
wire TIMEBOOST_net_11903;
wire TIMEBOOST_net_14572;
wire g53920_sb;
wire TIMEBOOST_net_11880;
wire TIMEBOOST_net_14260;
wire g53921_sb;
wire TIMEBOOST_net_11881;
wire TIMEBOOST_net_14355;
wire g53922_sb;
wire TIMEBOOST_net_11882;
wire TIMEBOOST_net_14542;
wire g53923_sb;
wire TIMEBOOST_net_11484;
wire TIMEBOOST_net_14003;
wire g53924_sb;
wire TIMEBOOST_net_11772;
wire TIMEBOOST_net_11193;
wire g53925_sb;
wire TIMEBOOST_net_11483;
wire TIMEBOOST_net_14379;
wire g53926_sb;
wire TIMEBOOST_net_11702;
wire TIMEBOOST_net_14531;
wire g53927_sb;
wire TIMEBOOST_net_11705;
wire TIMEBOOST_net_14005;
wire g53928_sb;
wire TIMEBOOST_net_11900;
wire TIMEBOOST_net_14127;
wire g53929_sb;
wire TIMEBOOST_net_11706;
wire TIMEBOOST_net_14036;
wire g53930_sb;
wire TIMEBOOST_net_11879;
wire TIMEBOOST_net_13967;
wire g53931_sb;
wire TIMEBOOST_net_11877;
wire TIMEBOOST_net_14527;
wire g53932_sb;
wire TIMEBOOST_net_9348;
wire TIMEBOOST_net_13831;
wire TIMEBOOST_net_4895;
wire TIMEBOOST_net_11322;
wire TIMEBOOST_net_14546;
wire TIMEBOOST_net_11359;
wire g53937_sb;
wire TIMEBOOST_net_10405;
wire TIMEBOOST_net_13795;
wire TIMEBOOST_net_4896;
wire TIMEBOOST_net_14321;
wire g53939_sb;
wire TIMEBOOST_net_11361;
wire TIMEBOOST_net_15213;
wire g53940_sb;
wire TIMEBOOST_net_13224;
wire TIMEBOOST_net_11255;
wire TIMEBOOST_net_11587;
wire g53942_db;
wire g53943_da;
wire TIMEBOOST_net_11324;
wire g53944_da;
wire TIMEBOOST_net_11254;
wire g53945_da;
wire TIMEBOOST_net_11323;
wire TIMEBOOST_net_10148;
wire TIMEBOOST_net_14800;
wire g53946_sb;
wire g53947_da;
wire TIMEBOOST_net_11325;
wire g53990_p;
wire TIMEBOOST_net_9643;
wire TIMEBOOST_net_10949;
wire g54030_sb;
wire TIMEBOOST_net_9380;
wire g54038_db;
wire g54038_sb;
wire g54039_da;
wire g54039_db;
wire g54039_sb;
wire TIMEBOOST_net_14825;
wire TIMEBOOST_net_4877;
wire g54040_sb;
wire g54131_da;
wire TIMEBOOST_net_10723;
wire g54131_sb;
wire TIMEBOOST_net_10764;
wire TIMEBOOST_net_4577;
wire g54132_sb;
wire TIMEBOOST_net_10765;
wire TIMEBOOST_net_4578;
wire g54133_sb;
wire TIMEBOOST_net_10746;
wire TIMEBOOST_net_10493;
wire g54134_sb;
wire TIMEBOOST_net_10747;
wire TIMEBOOST_net_13737;
wire g54135_sb;
wire g54137_da;
wire g54137_db;
wire g54137_sb;
wire TIMEBOOST_net_10176;
wire TIMEBOOST_net_10683;
wire g54138_sb;
wire g54139_da;
wire TIMEBOOST_net_10684;
wire TIMEBOOST_net_13789;
wire TIMEBOOST_net_4579;
wire g54140_sb;
wire TIMEBOOST_net_10177;
wire TIMEBOOST_net_10685;
wire g54141_sb;
wire TIMEBOOST_net_5234;
wire TIMEBOOST_net_10902;
wire g54143_sb;
wire TIMEBOOST_net_10506;
wire TIMEBOOST_net_10686;
wire g54144_sb;
wire TIMEBOOST_net_4795;
wire TIMEBOOST_net_4646;
wire g54145_sb;
wire TIMEBOOST_net_13788;
wire TIMEBOOST_net_4580;
wire g54146_sb;
wire TIMEBOOST_net_4796;
wire g54147_db;
wire g54147_sb;
wire TIMEBOOST_net_11028;
wire TIMEBOOST_net_10905;
wire g54148_sb;
wire TIMEBOOST_net_4797;
wire TIMEBOOST_net_10687;
wire g54149_sb;
wire g54150_da;
wire TIMEBOOST_net_10372;
wire g54150_sb;
wire TIMEBOOST_net_10885;
wire TIMEBOOST_net_10907;
wire g54151_sb;
wire g54152_da;
wire TIMEBOOST_net_10688;
wire g54152_sb;
wire TIMEBOOST_net_10184;
wire TIMEBOOST_net_10689;
wire g54153_sb;
wire TIMEBOOST_net_10185;
wire TIMEBOOST_net_10690;
wire g54154_sb;
wire g54155_da;
wire TIMEBOOST_net_2305;
wire g54155_sb;
wire g54157_da;
wire TIMEBOOST_net_4651;
wire g54157_sb;
wire TIMEBOOST_net_10186;
wire TIMEBOOST_net_10691;
wire g54158_sb;
wire TIMEBOOST_net_14885;
wire TIMEBOOST_net_12797;
wire g54160_sb;
wire TIMEBOOST_net_4801;
wire TIMEBOOST_net_4653;
wire g54161_sb;
wire TIMEBOOST_net_14886;
wire TIMEBOOST_net_14142;
wire TIMEBOOST_net_10187;
wire TIMEBOOST_net_4654;
wire g54164_sb;
wire TIMEBOOST_net_14890;
wire TIMEBOOST_net_14141;
wire TIMEBOOST_net_51;
wire TIMEBOOST_net_9383;
wire g54167_sb;
wire TIMEBOOST_net_14294;
wire TIMEBOOST_net_10911;
wire g54168_sb;
wire TIMEBOOST_net_14037;
wire TIMEBOOST_net_10913;
wire g54169_sb;
wire TIMEBOOST_net_14354;
wire TIMEBOOST_net_10914;
wire g54170_sb;
wire TIMEBOOST_net_12394;
wire g54171_sb;
wire TIMEBOOST_net_14289;
wire TIMEBOOST_net_13779;
wire g54172_sb;
wire TIMEBOOST_net_14366;
wire TIMEBOOST_net_10915;
wire g54173_sb;
wire g54174_da;
wire TIMEBOOST_net_14199;
wire g54174_sb;
wire TIMEBOOST_net_10802;
wire g54175_db;
wire g54175_sb;
wire g54176_da;
wire TIMEBOOST_net_10916;
wire g54176_sb;
wire TIMEBOOST_net_10886;
wire TIMEBOOST_net_10918;
wire g54177_sb;
wire TIMEBOOST_net_10887;
wire g54178_db;
wire g54178_sb;
wire TIMEBOOST_net_10888;
wire TIMEBOOST_net_10937;
wire g54179_sb;
wire g54180_da;
wire TIMEBOOST_net_10726;
wire g54180_sb;
wire g54181_da;
wire TIMEBOOST_net_10940;
wire g54181_sb;
wire TIMEBOOST_net_13946;
wire g54182_db;
wire g54182_sb;
wire TIMEBOOST_net_10889;
wire TIMEBOOST_net_10941;
wire g54183_sb;
wire TIMEBOOST_net_14327;
wire g54184_db;
wire g54184_sb;
wire g54185_da;
wire TIMEBOOST_net_14177;
wire g54185_sb;
wire TIMEBOOST_net_10890;
wire TIMEBOOST_net_10942;
wire g54186_sb;
wire TIMEBOOST_net_10891;
wire TIMEBOOST_net_10950;
wire g54187_sb;
wire TIMEBOOST_net_14376;
wire g54188_db;
wire g54188_sb;
wire TIMEBOOST_net_14104;
wire g54189_db;
wire g54189_sb;
wire TIMEBOOST_net_10892;
wire TIMEBOOST_net_10957;
wire g54190_sb;
wire TIMEBOOST_net_10893;
wire TIMEBOOST_net_10978;
wire g54191_sb;
wire TIMEBOOST_net_10894;
wire TIMEBOOST_net_10980;
wire g54192_sb;
wire TIMEBOOST_net_10895;
wire TIMEBOOST_net_10981;
wire g54193_sb;
wire TIMEBOOST_net_10803;
wire TIMEBOOST_net_870;
wire g54194_sb;
wire TIMEBOOST_net_10900;
wire TIMEBOOST_net_10983;
wire g54195_sb;
wire TIMEBOOST_net_14105;
wire g54196_db;
wire g54196_sb;
wire TIMEBOOST_net_10938;
wire TIMEBOOST_net_10987;
wire g54197_sb;
wire TIMEBOOST_net_9345;
wire g54198_db;
wire g54198_sb;
wire TIMEBOOST_net_14282;
wire g54199_db;
wire g54199_sb;
wire TIMEBOOST_net_10939;
wire g54200_db;
wire g54200_sb;
wire TIMEBOOST_net_9346;
wire g54201_db;
wire g54201_sb;
wire g54202_da;
wire TIMEBOOST_net_10988;
wire g54202_sb;
wire TIMEBOOST_net_14130;
wire TIMEBOOST_net_4552;
wire g54203_sb;
wire TIMEBOOST_net_19;
wire TIMEBOOST_net_12227;
wire TIMEBOOST_net_53;
wire TIMEBOOST_net_14153;
wire g54205_sb;
wire TIMEBOOST_net_14900;
wire TIMEBOOST_net_14457;
wire TIMEBOOST_net_12674;
wire g54207_sb;
wire TIMEBOOST_net_12642;
wire TIMEBOOST_net_12165;
wire TIMEBOOST_net_12695;
wire TIMEBOOST_net_11446;
wire g54209_sb;
wire TIMEBOOST_net_58;
wire TIMEBOOST_net_2900;
wire TIMEBOOST_net_59;
wire TIMEBOOST_net_12800;
wire TIMEBOOST_net_60;
wire TIMEBOOST_net_12753;
wire TIMEBOOST_net_61;
wire TIMEBOOST_net_12801;
wire TIMEBOOST_net_20;
wire TIMEBOOST_net_12228;
wire TIMEBOOST_net_62;
wire TIMEBOOST_net_12754;
wire TIMEBOOST_net_63;
wire TIMEBOOST_net_12802;
wire g54216_sb;
wire TIMEBOOST_net_64;
wire TIMEBOOST_net_2906;
wire TIMEBOOST_net_65;
wire TIMEBOOST_net_12755;
wire TIMEBOOST_net_66;
wire TIMEBOOST_net_12758;
wire g54219_sb;
wire TIMEBOOST_net_21;
wire TIMEBOOST_net_12229;
wire TIMEBOOST_net_67;
wire TIMEBOOST_net_3650;
wire TIMEBOOST_net_68;
wire TIMEBOOST_net_12759;
wire TIMEBOOST_net_69;
wire TIMEBOOST_net_12814;
wire TIMEBOOST_net_70;
wire TIMEBOOST_net_12815;
wire TIMEBOOST_net_71;
wire TIMEBOOST_net_12816;
wire TIMEBOOST_net_72;
wire TIMEBOOST_net_12817;
wire TIMEBOOST_net_73;
wire TIMEBOOST_net_12818;
wire TIMEBOOST_net_74;
wire TIMEBOOST_net_12819;
wire TIMEBOOST_net_22;
wire g54229_db;
wire TIMEBOOST_net_75;
wire TIMEBOOST_net_12820;
wire TIMEBOOST_net_76;
wire TIMEBOOST_net_12821;
wire TIMEBOOST_net_77;
wire TIMEBOOST_net_12822;
wire TIMEBOOST_net_78;
wire TIMEBOOST_net_12823;
wire TIMEBOOST_net_14057;
wire TIMEBOOST_net_10693;
wire g54234_sb;
wire TIMEBOOST_net_10763;
wire TIMEBOOST_net_4581;
wire g54235_sb;
wire TIMEBOOST_net_10188;
wire TIMEBOOST_net_10694;
wire g54236_sb;
wire TIMEBOOST_net_14917;
wire TIMEBOOST_net_10695;
wire g54237_sb;
wire TIMEBOOST_net_10189;
wire TIMEBOOST_net_4658;
wire g54238_sb;
wire TIMEBOOST_net_13774;
wire TIMEBOOST_net_10636;
wire g54239_sb;
wire TIMEBOOST_net_14543;
wire TIMEBOOST_net_11899;
wire g54244_sb;
wire TIMEBOOST_net_13992;
wire TIMEBOOST_net_4553;
wire g54304_sb;
wire g54305_da;
wire g54305_db;
wire g54305_sb;
wire g54306_da;
wire g54306_db;
wire g54306_sb;
wire g54309_da;
wire g54309_db;
wire g54309_sb;
wire g54310_da;
wire g54310_db;
wire g54310_sb;
wire g54311_da;
wire g54311_db;
wire g54311_sb;
wire g54312_da;
wire g54312_db;
wire g54312_sb;
wire g54314_da;
wire g54314_db;
wire g54314_sb;
wire g54315_da;
wire g54315_db;
wire g54315_sb;
wire TIMEBOOST_net_910;
wire TIMEBOOST_net_4414;
wire g54316_sb;
wire g54317_da;
wire g54317_db;
wire g54317_sb;
wire TIMEBOOST_net_10392;
wire g54318_db;
wire g54318_sb;
wire g54319_da;
wire TIMEBOOST_net_4879;
wire g54319_sb;
wire g54320_da;
wire TIMEBOOST_net_14072;
wire g54320_sb;
wire TIMEBOOST_net_10833;
wire g54321_db;
wire g54321_sb;
wire g54322_da;
wire g54322_db;
wire g54322_sb;
wire g54323_da;
wire TIMEBOOST_net_14297;
wire g54323_sb;
wire g54324_da;
wire g54324_db;
wire g54324_sb;
wire g54325_da;
wire g54325_db;
wire g54325_sb;
wire TIMEBOOST_net_14467;
wire TIMEBOOST_net_14646;
wire g54326_sb;
wire TIMEBOOST_net_12396;
wire TIMEBOOST_net_10727;
wire g54328_sb;
wire g54329_p;
wire TIMEBOOST_net_10842;
wire g54330_db;
wire g54330_sb;
wire g54331_da;
wire g54331_db;
wire g54331_sb;
wire TIMEBOOST_net_4752;
wire TIMEBOOST_net_14175;
wire g54332_sb;
wire TIMEBOOST_net_14298;
wire TIMEBOOST_net_10500;
wire g54333_sb;
wire TIMEBOOST_net_9333;
wire TIMEBOOST_net_4556;
wire g54334_sb;
wire TIMEBOOST_net_9334;
wire TIMEBOOST_net_10728;
wire g54335_sb;
wire g54336_da;
wire g54336_db;
wire g54336_sb;
wire TIMEBOOST_net_13032;
wire g54337_sb;
wire TIMEBOOST_net_9358;
wire TIMEBOOST_net_11790;
wire g54338_sb;
wire TIMEBOOST_net_11886;
wire TIMEBOOST_net_14937;
wire g54339_sb;
wire TIMEBOOST_net_11887;
wire TIMEBOOST_net_2042;
wire g54340_sb;
wire TIMEBOOST_net_11888;
wire TIMEBOOST_net_14938;
wire g54341_sb;
wire TIMEBOOST_net_11889;
wire n_14087;
wire g54342_sb;
wire TIMEBOOST_net_11890;
wire TIMEBOOST_net_14039;
wire g54343_sb;
wire TIMEBOOST_net_11891;
wire TIMEBOOST_net_14333;
wire g54344_sb;
wire TIMEBOOST_net_11769;
wire TIMEBOOST_net_14607;
wire g54345_sb;
wire TIMEBOOST_net_11824;
wire TIMEBOOST_net_10778;
wire g54346_sb;
wire TIMEBOOST_net_11715;
wire TIMEBOOST_net_2048;
wire g54347_sb;
wire TIMEBOOST_net_11716;
wire TIMEBOOST_net_13980;
wire g54348_sb;
wire TIMEBOOST_net_13929;
wire TIMEBOOST_net_11568;
wire g54349_sb;
wire TIMEBOOST_net_11717;
wire TIMEBOOST_net_14218;
wire g54350_sb;
wire TIMEBOOST_net_11718;
wire TIMEBOOST_net_14196;
wire g54351_sb;
wire TIMEBOOST_net_11770;
wire TIMEBOOST_net_14206;
wire g54352_sb;
wire TIMEBOOST_net_2018;
wire TIMEBOOST_net_11710;
wire g54353_sb;
wire TIMEBOOST_net_9359;
wire TIMEBOOST_net_11825;
wire g54354_sb;
wire TIMEBOOST_net_11773;
wire TIMEBOOST_net_14188;
wire g54355_sb;
wire TIMEBOOST_net_11775;
wire TIMEBOOST_net_14192;
wire g54356_sb;
wire TIMEBOOST_net_14074;
wire TIMEBOOST_net_11873;
wire g54357_sb;
wire TIMEBOOST_net_9360;
wire TIMEBOOST_net_11875;
wire g54358_sb;
wire TIMEBOOST_net_14347;
wire TIMEBOOST_net_11876;
wire g54359_sb;
wire TIMEBOOST_net_14338;
wire TIMEBOOST_net_11711;
wire g54360_sb;
wire TIMEBOOST_net_2024;
wire TIMEBOOST_net_11712;
wire g54361_sb;
wire TIMEBOOST_net_2025;
wire TIMEBOOST_net_11713;
wire g54362_sb;
wire TIMEBOOST_net_14253;
wire TIMEBOOST_net_11714;
wire g54363_sb;
wire TIMEBOOST_net_14547;
wire TIMEBOOST_net_11707;
wire g54364_sb;
wire TIMEBOOST_net_2028;
wire TIMEBOOST_net_11721;
wire g54365_sb;
wire TIMEBOOST_net_14009;
wire TIMEBOOST_net_11722;
wire g54366_sb;
wire TIMEBOOST_net_14540;
wire TIMEBOOST_net_11730;
wire g54367_sb;
wire TIMEBOOST_net_11776;
wire TIMEBOOST_net_13844;
wire g54368_sb;
wire TIMEBOOST_net_11777;
wire TIMEBOOST_net_10777;
wire g54369_sb;
wire g54453_p;
wire g54456_p;
wire g54458_p;
wire g54465_p;
wire TIMEBOOST_net_13021;
wire g54471_sb;
wire TIMEBOOST_net_13854;
wire g54472_sb;
wire TIMEBOOST_net_13856;
wire g54484_sb;
wire TIMEBOOST_net_14181;
wire g54485_sb;
wire TIMEBOOST_net_13039;
wire g54486_sb;
wire TIMEBOOST_net_6487;
wire TIMEBOOST_net_13005;
wire g54487_sb;
wire n_12062;
wire g62000_db;
wire g54488_sb;
wire TIMEBOOST_net_695;
wire TIMEBOOST_net_13034;
wire g54489_sb;
wire n_12410;
wire TIMEBOOST_net_13017;
wire g54490_sb;
wire n_12183;
wire TIMEBOOST_net_13023;
wire g54491_sb;
wire TIMEBOOST_net_14183;
wire g54492_sb;
wire TIMEBOOST_net_13043;
wire g54493_sb;
wire TIMEBOOST_net_6438;
wire TIMEBOOST_net_13011;
wire g54494_sb;
wire TIMEBOOST_net_13029;
wire g54495_sb;
wire g54568_p;
wire g54569_p;
wire g54572_p;
wire g54573_p;
wire g54574_p;
wire g54579_p;
wire g54580_p;
wire g54581_p;
wire g54586_p;
wire g54587_p;
wire g54591_p;
wire g54593_p;
wire g54594_p;
wire g54595_p;
wire g54596_p;
wire g54597_p;
wire g54601_p;
wire g54603_p;
wire g54606_p;
wire TIMEBOOST_net_13287;
wire g55851_sb;
wire TIMEBOOST_net_13288;
wire g55852_sb;
wire TIMEBOOST_net_13289;
wire g55853_sb;
wire TIMEBOOST_net_12645;
wire TIMEBOOST_net_2057;
wire g56933_sb;
wire TIMEBOOST_net_9608;
wire TIMEBOOST_net_6439;
wire g56934_sb;
wire g57030_p;
wire g57033_p;
wire TIMEBOOST_net_11784;
wire TIMEBOOST_net_13804;
wire g57034_sb;
wire TIMEBOOST_net_13803;
wire g57035_sb;
wire TIMEBOOST_net_11786;
wire TIMEBOOST_net_13801;
wire g57036_sb;
wire TIMEBOOST_net_6032;
wire TIMEBOOST_net_13802;
wire g57037_sb;
wire TIMEBOOST_net_11965;
wire TIMEBOOST_net_13797;
wire g57038_sb;
wire TIMEBOOST_net_13142;
wire g57039_sb;
wire TIMEBOOST_net_13143;
wire g57040_sb;
wire TIMEBOOST_net_11966;
wire TIMEBOOST_net_13796;
wire g57041_sb;
wire TIMEBOOST_net_11917;
wire TIMEBOOST_net_13798;
wire g57042_sb;
wire TIMEBOOST_net_11918;
wire TIMEBOOST_net_13799;
wire g57043_sb;
wire TIMEBOOST_net_13895;
wire TIMEBOOST_net_11893;
wire g57044_sb;
wire TIMEBOOST_net_11919;
wire TIMEBOOST_net_13792;
wire g57045_sb;
wire TIMEBOOST_net_13144;
wire g57046_sb;
wire TIMEBOOST_net_13322;
wire TIMEBOOST_net_11878;
wire g57047_sb;
wire TIMEBOOST_net_11920;
wire TIMEBOOST_net_10828;
wire g57048_sb;
wire TIMEBOOST_net_13145;
wire g57049_sb;
wire TIMEBOOST_net_13146;
wire g57050_sb;
wire TIMEBOOST_net_11928;
wire TIMEBOOST_net_13689;
wire g57051_sb;
wire TIMEBOOST_net_11906;
wire TIMEBOOST_net_13690;
wire g57052_sb;
wire TIMEBOOST_net_11907;
wire TIMEBOOST_net_13691;
wire g57053_sb;
wire TIMEBOOST_net_11908;
wire TIMEBOOST_net_13163;
wire TIMEBOOST_net_13147;
wire g57055_sb;
wire TIMEBOOST_net_11909;
wire TIMEBOOST_net_13692;
wire g57056_sb;
wire TIMEBOOST_net_11910;
wire TIMEBOOST_net_13693;
wire g57057_sb;
wire TIMEBOOST_net_13148;
wire g57058_sb;
wire TIMEBOOST_net_13149;
wire g57059_sb;
wire TIMEBOOST_net_13150;
wire g57060_sb;
wire TIMEBOOST_net_11911;
wire TIMEBOOST_net_13694;
wire g57061_sb;
wire TIMEBOOST_net_11912;
wire TIMEBOOST_net_4373;
wire g57062_sb;
wire TIMEBOOST_net_13321;
wire TIMEBOOST_net_11747;
wire g57063_sb;
wire TIMEBOOST_net_13151;
wire g57064_sb;
wire TIMEBOOST_net_11943;
wire TIMEBOOST_net_13695;
wire g57065_sb;
wire TIMEBOOST_net_11913;
wire TIMEBOOST_net_13696;
wire g57066_sb;
wire TIMEBOOST_net_13128;
wire g57067_sb;
wire TIMEBOOST_net_11914;
wire TIMEBOOST_net_13697;
wire g57068_sb;
wire TIMEBOOST_net_15207;
wire TIMEBOOST_net_13698;
wire g57069_sb;
wire TIMEBOOST_net_11739;
wire TIMEBOOST_net_13699;
wire g57070_sb;
wire TIMEBOOST_net_11944;
wire TIMEBOOST_net_4371;
wire g57071_sb;
wire TIMEBOOST_net_14664;
wire TIMEBOOST_net_13665;
wire g57072_sb;
wire TIMEBOOST_net_11750;
wire TIMEBOOST_net_13664;
wire g57073_sb;
wire TIMEBOOST_net_13152;
wire g57074_sb;
wire TIMEBOOST_net_11785;
wire TIMEBOOST_net_13667;
wire g57075_sb;
wire TIMEBOOST_net_13126;
wire g57076_sb;
wire TIMEBOOST_net_14663;
wire TIMEBOOST_net_13669;
wire g57077_sb;
wire TIMEBOOST_net_13313;
wire g57078_db;
wire g57078_sb;
wire TIMEBOOST_net_926;
wire TIMEBOOST_net_11569;
wire g57079_sb;
wire TIMEBOOST_net_11787;
wire TIMEBOOST_net_13670;
wire g57080_sb;
wire TIMEBOOST_net_6058;
wire TIMEBOOST_net_13589;
wire g57081_sb;
wire TIMEBOOST_net_11788;
wire TIMEBOOST_net_10934;
wire g57082_sb;
wire TIMEBOOST_net_11789;
wire n_13436;
wire g57083_sb;
wire TIMEBOOST_net_11986;
wire n_4768;
wire g57084_sb;
wire TIMEBOOST_net_11987;
wire n_4770;
wire g57085_sb;
wire TIMEBOOST_net_11988;
wire n_4772;
wire g57086_sb;
wire TIMEBOOST_net_11989;
wire n_4773;
wire g57087_sb;
wire TIMEBOOST_net_11921;
wire n_4774;
wire g57088_sb;
wire TIMEBOOST_net_11926;
wire n_4775;
wire g57089_sb;
wire TIMEBOOST_net_11927;
wire TIMEBOOST_net_13659;
wire g57090_sb;
wire TIMEBOOST_net_11929;
wire n_4779;
wire g57091_sb;
wire TIMEBOOST_net_11930;
wire n_4760;
wire g57092_sb;
wire TIMEBOOST_net_6463;
wire TIMEBOOST_net_13108;
wire g57093_sb;
wire TIMEBOOST_net_6464;
wire TIMEBOOST_net_13109;
wire g57094_sb;
wire TIMEBOOST_net_14692;
wire n_4748;
wire g57095_sb;
wire TIMEBOOST_net_14691;
wire TIMEBOOST_net_13633;
wire g57096_sb;
wire TIMEBOOST_net_11947;
wire TIMEBOOST_net_13623;
wire g57097_sb;
wire TIMEBOOST_net_11948;
wire TIMEBOOST_net_13632;
wire g57098_sb;
wire TIMEBOOST_net_11949;
wire TIMEBOOST_net_13622;
wire g57099_sb;
wire TIMEBOOST_net_11950;
wire TIMEBOOST_net_13621;
wire g57100_sb;
wire TIMEBOOST_net_11951;
wire TIMEBOOST_net_13620;
wire g57101_sb;
wire TIMEBOOST_net_11952;
wire TIMEBOOST_net_13619;
wire g57102_sb;
wire TIMEBOOST_net_11953;
wire TIMEBOOST_net_13618;
wire g57103_sb;
wire TIMEBOOST_net_11954;
wire TIMEBOOST_net_13617;
wire g57104_sb;
wire TIMEBOOST_net_11955;
wire TIMEBOOST_net_13634;
wire g57105_sb;
wire TIMEBOOST_net_11974;
wire TIMEBOOST_net_13616;
wire g57106_sb;
wire TIMEBOOST_net_11975;
wire TIMEBOOST_net_13635;
wire g57107_sb;
wire TIMEBOOST_net_11767;
wire TIMEBOOST_net_13615;
wire g57108_sb;
wire TIMEBOOST_net_6465;
wire TIMEBOOST_net_3887;
wire g57109_sb;
wire TIMEBOOST_net_12000;
wire TIMEBOOST_net_13614;
wire g57110_sb;
wire TIMEBOOST_net_12160;
wire TIMEBOOST_net_13153;
wire g57111_sb;
wire TIMEBOOST_net_11458;
wire TIMEBOOST_net_6430;
wire g57112_sb;
wire TIMEBOOST_net_12001;
wire TIMEBOOST_net_4611;
wire g57113_sb;
wire TIMEBOOST_net_11971;
wire TIMEBOOST_net_4609;
wire g57114_sb;
wire TIMEBOOST_net_10815;
wire g57115_db;
wire g57115_sb;
wire TIMEBOOST_net_12006;
wire TIMEBOOST_net_4541;
wire g57116_sb;
wire TIMEBOOST_net_14579;
wire g57117_db;
wire g57117_sb;
wire TIMEBOOST_net_11946;
wire TIMEBOOST_net_4606;
wire g57118_sb;
wire TIMEBOOST_net_12190;
wire TIMEBOOST_net_13154;
wire g57119_sb;
wire TIMEBOOST_net_12007;
wire TIMEBOOST_net_4605;
wire g57120_sb;
wire TIMEBOOST_net_12018;
wire TIMEBOOST_net_14506;
wire g57121_sb;
wire TIMEBOOST_net_11967;
wire TIMEBOOST_net_13712;
wire g57122_sb;
wire TIMEBOOST_net_13894;
wire TIMEBOOST_net_11748;
wire g57123_sb;
wire TIMEBOOST_net_11962;
wire TIMEBOOST_net_14507;
wire g57124_sb;
wire TIMEBOOST_net_11963;
wire TIMEBOOST_net_13713;
wire g57125_sb;
wire TIMEBOOST_net_11964;
wire TIMEBOOST_net_14581;
wire g57126_sb;
wire TIMEBOOST_net_11969;
wire TIMEBOOST_net_14419;
wire g57127_sb;
wire TIMEBOOST_net_11991;
wire TIMEBOOST_net_13714;
wire g57128_sb;
wire TIMEBOOST_net_11992;
wire TIMEBOOST_net_13715;
wire g57129_sb;
wire TIMEBOOST_net_11993;
wire TIMEBOOST_net_13716;
wire g57130_sb;
wire TIMEBOOST_net_12008;
wire TIMEBOOST_net_13717;
wire g57131_sb;
wire TIMEBOOST_net_12009;
wire TIMEBOOST_net_14421;
wire g57132_sb;
wire TIMEBOOST_net_12010;
wire TIMEBOOST_net_4533;
wire g57133_sb;
wire TIMEBOOST_net_12011;
wire TIMEBOOST_net_13748;
wire g57134_sb;
wire TIMEBOOST_net_12012;
wire TIMEBOOST_net_13613;
wire g57135_sb;
wire TIMEBOOST_net_12013;
wire TIMEBOOST_net_4629;
wire g57136_sb;
wire TIMEBOOST_net_12184;
wire TIMEBOOST_net_13155;
wire g57137_sb;
wire TIMEBOOST_net_12014;
wire TIMEBOOST_net_4623;
wire g57138_sb;
wire TIMEBOOST_net_12015;
wire TIMEBOOST_net_13721;
wire g57139_sb;
wire TIMEBOOST_net_13290;
wire g57140_db;
wire g57140_sb;
wire TIMEBOOST_net_12016;
wire TIMEBOOST_net_4545;
wire g57141_sb;
wire TIMEBOOST_net_12017;
wire TIMEBOOST_net_4544;
wire g57142_sb;
wire TIMEBOOST_net_13864;
wire TIMEBOOST_net_11758;
wire g57143_sb;
wire TIMEBOOST_net_6469;
wire TIMEBOOST_net_13157;
wire g57144_sb;
wire TIMEBOOST_net_12022;
wire TIMEBOOST_net_13722;
wire g57145_sb;
wire TIMEBOOST_net_6470;
wire TIMEBOOST_net_13158;
wire g57146_sb;
wire TIMEBOOST_net_11940;
wire TIMEBOOST_net_14599;
wire g57147_sb;
wire TIMEBOOST_net_13865;
wire g57148_db;
wire g57148_sb;
wire TIMEBOOST_net_11973;
wire TIMEBOOST_net_13723;
wire g57149_sb;
wire TIMEBOOST_net_12005;
wire TIMEBOOST_net_13724;
wire g57150_sb;
wire TIMEBOOST_net_12004;
wire TIMEBOOST_net_4572;
wire g57151_sb;
wire TIMEBOOST_net_11972;
wire TIMEBOOST_net_4532;
wire g57152_sb;
wire TIMEBOOST_net_13292;
wire g57153_db;
wire g57153_sb;
wire TIMEBOOST_net_12181;
wire TIMEBOOST_net_13159;
wire g57154_sb;
wire TIMEBOOST_net_11922;
wire TIMEBOOST_net_13756;
wire g57155_sb;
wire TIMEBOOST_net_11924;
wire TIMEBOOST_net_13707;
wire g57156_sb;
wire TIMEBOOST_net_12195;
wire TIMEBOOST_net_13706;
wire g57157_sb;
wire TIMEBOOST_net_13866;
wire TIMEBOOST_net_11759;
wire g57158_sb;
wire TIMEBOOST_net_11925;
wire TIMEBOOST_net_13677;
wire g57159_sb;
wire TIMEBOOST_net_13868;
wire g57160_db;
wire g57160_sb;
wire TIMEBOOST_net_12003;
wire TIMEBOOST_net_13728;
wire g57161_sb;
wire TIMEBOOST_net_12020;
wire TIMEBOOST_net_13709;
wire g57162_sb;
wire TIMEBOOST_net_6473;
wire TIMEBOOST_net_13726;
wire g57163_sb;
wire TIMEBOOST_net_12021;
wire TIMEBOOST_net_14583;
wire g57164_sb;
wire TIMEBOOST_net_11979;
wire TIMEBOOST_net_14582;
wire g57165_sb;
wire TIMEBOOST_net_11998;
wire TIMEBOOST_net_10869;
wire g57166_sb;
wire TIMEBOOST_net_11978;
wire TIMEBOOST_net_14584;
wire g57167_sb;
wire TIMEBOOST_net_11980;
wire TIMEBOOST_net_14585;
wire g57168_sb;
wire TIMEBOOST_net_11981;
wire TIMEBOOST_net_14594;
wire g57169_sb;
wire TIMEBOOST_net_11771;
wire TIMEBOOST_net_10870;
wire g57170_sb;
wire TIMEBOOST_net_11982;
wire TIMEBOOST_net_14593;
wire g57171_sb;
wire TIMEBOOST_net_6474;
wire TIMEBOOST_net_13160;
wire g57172_sb;
wire TIMEBOOST_net_11983;
wire TIMEBOOST_net_13731;
wire g57173_sb;
wire TIMEBOOST_net_13161;
wire g57174_sb;
wire TIMEBOOST_net_13165;
wire g57175_sb;
wire TIMEBOOST_net_12019;
wire TIMEBOOST_net_14431;
wire g57176_sb;
wire TIMEBOOST_net_12002;
wire TIMEBOOST_net_14432;
wire g57177_sb;
wire TIMEBOOST_net_10816;
wire g57178_db;
wire g57178_sb;
wire TIMEBOOST_net_6477;
wire TIMEBOOST_net_13166;
wire g57179_sb;
wire TIMEBOOST_net_11936;
wire TIMEBOOST_net_13732;
wire g57180_sb;
wire TIMEBOOST_net_13291;
wire TIMEBOOST_net_13264;
wire g57181_sb;
wire TIMEBOOST_net_11937;
wire TIMEBOOST_net_10871;
wire g57182_sb;
wire TIMEBOOST_net_11941;
wire TIMEBOOST_net_14588;
wire g57183_sb;
wire TIMEBOOST_net_13869;
wire TIMEBOOST_net_11723;
wire g57184_sb;
wire TIMEBOOST_net_11942;
wire TIMEBOOST_net_14410;
wire g57185_sb;
wire TIMEBOOST_net_13293;
wire TIMEBOOST_net_6431;
wire g57186_sb;
wire TIMEBOOST_net_13294;
wire TIMEBOOST_net_11724;
wire g57187_sb;
wire TIMEBOOST_net_11945;
wire TIMEBOOST_net_13746;
wire g57188_sb;
wire TIMEBOOST_net_11976;
wire TIMEBOOST_net_13794;
wire g57189_sb;
wire TIMEBOOST_net_11977;
wire g52441_db;
wire g57190_sb;
wire TIMEBOOST_net_11985;
wire TIMEBOOST_net_13790;
wire g57191_sb;
wire TIMEBOOST_net_11994;
wire TIMEBOOST_net_14590;
wire g57192_sb;
wire TIMEBOOST_net_11995;
wire TIMEBOOST_net_13729;
wire g57193_sb;
wire TIMEBOOST_net_6478;
wire TIMEBOOST_net_13130;
wire g57194_sb;
wire TIMEBOOST_net_11996;
wire TIMEBOOST_net_13730;
wire g57195_sb;
wire TIMEBOOST_net_11997;
wire TIMEBOOST_net_13751;
wire g57196_sb;
wire TIMEBOOST_net_11923;
wire TIMEBOOST_net_4688;
wire g57197_sb;
wire TIMEBOOST_net_13295;
wire TIMEBOOST_net_6432;
wire g57198_sb;
wire TIMEBOOST_net_6479;
wire TIMEBOOST_net_13171;
wire g57199_sb;
wire TIMEBOOST_net_13296;
wire g57200_sb;
wire TIMEBOOST_net_11933;
wire TIMEBOOST_net_4687;
wire g57201_sb;
wire TIMEBOOST_net_11934;
wire TIMEBOOST_net_13745;
wire g57202_sb;
wire TIMEBOOST_net_13297;
wire n_1566;
wire g57203_sb;
wire TIMEBOOST_net_11935;
wire TIMEBOOST_net_14306;
wire g57204_sb;
wire TIMEBOOST_net_11956;
wire TIMEBOOST_net_14512;
wire g57205_sb;
wire TIMEBOOST_net_11957;
wire TIMEBOOST_net_14598;
wire g57206_sb;
wire TIMEBOOST_net_13172;
wire g57207_sb;
wire TIMEBOOST_net_11958;
wire TIMEBOOST_net_10872;
wire g57208_sb;
wire TIMEBOOST_net_11959;
wire TIMEBOOST_net_13720;
wire g57209_sb;
wire TIMEBOOST_net_13298;
wire TIMEBOOST_net_6434;
wire g57210_sb;
wire TIMEBOOST_net_11968;
wire TIMEBOOST_net_4631;
wire g57211_sb;
wire TIMEBOOST_net_11970;
wire n_4758;
wire g57212_sb;
wire TIMEBOOST_net_11999;
wire TIMEBOOST_net_4678;
wire g57213_sb;
wire TIMEBOOST_net_6481;
wire TIMEBOOST_net_13173;
wire g57214_sb;
wire TIMEBOOST_net_13718;
wire g57215_sb;
wire TIMEBOOST_net_11938;
wire TIMEBOOST_net_13719;
wire g57216_sb;
wire TIMEBOOST_net_12025;
wire TIMEBOOST_net_13749;
wire g57217_sb;
wire TIMEBOOST_net_11939;
wire TIMEBOOST_net_13778;
wire g57218_sb;
wire TIMEBOOST_net_10788;
wire TIMEBOOST_net_11760;
wire g57219_sb;
wire TIMEBOOST_net_11931;
wire TIMEBOOST_net_14589;
wire g57220_sb;
wire TIMEBOOST_net_6483;
wire TIMEBOOST_net_13174;
wire g57221_sb;
wire TIMEBOOST_net_13299;
wire TIMEBOOST_net_11725;
wire g57222_sb;
wire TIMEBOOST_net_11932;
wire TIMEBOOST_net_14587;
wire g57223_sb;
wire TIMEBOOST_net_13131;
wire g57224_sb;
wire TIMEBOOST_net_13176;
wire g57225_sb;
wire TIMEBOOST_net_11960;
wire TIMEBOOST_net_14314;
wire g57226_sb;
wire TIMEBOOST_net_11961;
wire TIMEBOOST_net_4673;
wire g57227_sb;
wire TIMEBOOST_net_6161;
wire TIMEBOOST_net_13752;
wire g57228_sb;
wire TIMEBOOST_net_6486;
wire TIMEBOOST_net_13164;
wire g57229_sb;
wire TIMEBOOST_net_12194;
wire TIMEBOOST_net_13134;
wire g57230_sb;
wire TIMEBOOST_net_12023;
wire TIMEBOOST_net_13753;
wire g57231_sb;
wire TIMEBOOST_net_13112;
wire g57232_sb;
wire TIMEBOOST_net_11984;
wire TIMEBOOST_net_13754;
wire g57233_sb;
wire TIMEBOOST_net_13177;
wire g57234_sb;
wire TIMEBOOST_net_6490;
wire TIMEBOOST_net_13138;
wire g57235_sb;
wire TIMEBOOST_net_11990;
wire TIMEBOOST_net_4663;
wire g57236_sb;
wire TIMEBOOST_net_6165;
wire TIMEBOOST_net_4657;
wire g57237_sb;
wire TIMEBOOST_net_13300;
wire TIMEBOOST_net_11761;
wire g57238_sb;
wire TIMEBOOST_net_6491;
wire TIMEBOOST_net_13178;
wire g57239_sb;
wire TIMEBOOST_net_6166;
wire TIMEBOOST_net_13733;
wire g57240_sb;
wire TIMEBOOST_net_6167;
wire TIMEBOOST_net_14600;
wire g57241_sb;
wire TIMEBOOST_net_6492;
wire TIMEBOOST_net_13179;
wire g57242_sb;
wire TIMEBOOST_net_6168;
wire TIMEBOOST_net_13734;
wire g57243_sb;
wire TIMEBOOST_net_6169;
wire TIMEBOOST_net_13711;
wire g57244_sb;
wire TIMEBOOST_net_6493;
wire TIMEBOOST_net_13180;
wire g57245_sb;
wire TIMEBOOST_net_12064;
wire TIMEBOOST_net_4650;
wire g57246_sb;
wire TIMEBOOST_net_6171;
wire TIMEBOOST_net_13755;
wire g57247_sb;
wire TIMEBOOST_net_12057;
wire TIMEBOOST_net_4648;
wire g57248_sb;
wire TIMEBOOST_net_6494;
wire TIMEBOOST_net_13124;
wire g57249_sb;
wire TIMEBOOST_net_12063;
wire TIMEBOOST_net_13750;
wire g57250_sb;
wire TIMEBOOST_net_12048;
wire TIMEBOOST_net_14601;
wire g57251_sb;
wire TIMEBOOST_net_12049;
wire TIMEBOOST_net_4566;
wire g57252_sb;
wire TIMEBOOST_net_12050;
wire TIMEBOOST_net_13738;
wire g57253_sb;
wire TIMEBOOST_net_12051;
wire TIMEBOOST_net_13739;
wire g57254_sb;
wire TIMEBOOST_net_12061;
wire TIMEBOOST_net_13725;
wire g57255_sb;
wire TIMEBOOST_net_6495;
wire TIMEBOOST_net_13740;
wire g57256_sb;
wire TIMEBOOST_net_12060;
wire TIMEBOOST_net_13741;
wire g57257_sb;
wire TIMEBOOST_net_13060;
wire g57258_sb;
wire TIMEBOOST_net_13096;
wire g57259_sb;
wire TIMEBOOST_net_13301;
wire g57260_sb;
wire TIMEBOOST_net_12042;
wire TIMEBOOST_net_13742;
wire g57261_sb;
wire TIMEBOOST_net_12027;
wire TIMEBOOST_net_13743;
wire g57262_sb;
wire TIMEBOOST_net_12043;
wire TIMEBOOST_net_4583;
wire g57263_sb;
wire TIMEBOOST_net_12046;
wire TIMEBOOST_net_10931;
wire g57264_sb;
wire TIMEBOOST_net_12038;
wire TIMEBOOST_net_14511;
wire g57265_sb;
wire TIMEBOOST_net_12039;
wire TIMEBOOST_net_13744;
wire g57266_sb;
wire TIMEBOOST_net_12040;
wire TIMEBOOST_net_13704;
wire g57267_sb;
wire TIMEBOOST_net_6498;
wire TIMEBOOST_net_13097;
wire g57268_sb;
wire TIMEBOOST_net_12041;
wire TIMEBOOST_net_14559;
wire g57269_sb;
wire TIMEBOOST_net_13302;
wire TIMEBOOST_net_11762;
wire g57270_sb;
wire TIMEBOOST_net_6499;
wire TIMEBOOST_net_13058;
wire g57271_sb;
wire TIMEBOOST_net_12045;
wire TIMEBOOST_net_13658;
wire g57272_sb;
wire TIMEBOOST_net_12029;
wire TIMEBOOST_net_13702;
wire g57273_sb;
wire TIMEBOOST_net_12037;
wire TIMEBOOST_net_13703;
wire g57274_sb;
wire TIMEBOOST_net_12044;
wire TIMEBOOST_net_13674;
wire g57275_sb;
wire TIMEBOOST_net_12047;
wire TIMEBOOST_net_13675;
wire g57276_sb;
wire TIMEBOOST_net_12052;
wire TIMEBOOST_net_10932;
wire g57277_sb;
wire TIMEBOOST_net_12053;
wire TIMEBOOST_net_13676;
wire g57278_sb;
wire TIMEBOOST_net_12054;
wire TIMEBOOST_net_13678;
wire g57279_sb;
wire TIMEBOOST_net_12055;
wire TIMEBOOST_net_13679;
wire g57280_sb;
wire TIMEBOOST_net_6500;
wire TIMEBOOST_net_13129;
wire g57281_sb;
wire TIMEBOOST_net_12056;
wire TIMEBOOST_net_13680;
wire g57282_sb;
wire TIMEBOOST_net_6501;
wire TIMEBOOST_net_13065;
wire g57283_sb;
wire TIMEBOOST_net_13066;
wire g57284_sb;
wire TIMEBOOST_net_10817;
wire TIMEBOOST_net_11763;
wire g57285_sb;
wire TIMEBOOST_net_12058;
wire TIMEBOOST_net_13681;
wire g57286_sb;
wire TIMEBOOST_net_12059;
wire TIMEBOOST_net_13682;
wire g57287_sb;
wire TIMEBOOST_net_12062;
wire TIMEBOOST_net_13683;
wire g57288_sb;
wire TIMEBOOST_net_12028;
wire TIMEBOOST_net_13684;
wire g57289_sb;
wire TIMEBOOST_net_13867;
wire TIMEBOOST_net_11764;
wire g57290_sb;
wire TIMEBOOST_net_13303;
wire TIMEBOOST_net_6436;
wire g57291_sb;
wire TIMEBOOST_net_12035;
wire TIMEBOOST_net_13685;
wire g57292_sb;
wire TIMEBOOST_net_12036;
wire TIMEBOOST_net_10933;
wire g57293_sb;
wire TIMEBOOST_net_12030;
wire TIMEBOOST_net_13686;
wire g57294_sb;
wire TIMEBOOST_net_12031;
wire TIMEBOOST_net_13687;
wire g57295_sb;
wire TIMEBOOST_net_12032;
wire TIMEBOOST_net_13688;
wire g57296_sb;
wire TIMEBOOST_net_12033;
wire TIMEBOOST_net_4374;
wire g57297_sb;
wire TIMEBOOST_net_12034;
wire TIMEBOOST_net_13663;
wire g57298_sb;
wire TIMEBOOST_net_6209;
wire TIMEBOOST_net_13668;
wire g57299_sb;
wire TIMEBOOST_net_13884;
wire g57300_db;
wire g57300_sb;
wire TIMEBOOST_net_12024;
wire n_4753;
wire g57301_sb;
wire TIMEBOOST_net_12138;
wire TIMEBOOST_net_13777;
wire g57302_sb;
wire TIMEBOOST_net_12139;
wire TIMEBOOST_net_10929;
wire g57303_sb;
wire TIMEBOOST_net_12140;
wire TIMEBOOST_net_13771;
wire g57304_sb;
wire TIMEBOOST_net_12141;
wire TIMEBOOST_net_13762;
wire g57305_sb;
wire TIMEBOOST_net_12142;
wire g52395_db;
wire g57306_sb;
wire TIMEBOOST_net_12143;
wire TIMEBOOST_net_13758;
wire g57307_sb;
wire TIMEBOOST_net_12144;
wire TIMEBOOST_net_13727;
wire g57308_sb;
wire TIMEBOOST_net_12145;
wire TIMEBOOST_net_13644;
wire g57309_sb;
wire TIMEBOOST_net_12137;
wire TIMEBOOST_net_13647;
wire g57310_sb;
wire TIMEBOOST_net_12136;
wire TIMEBOOST_net_13652;
wire g57311_sb;
wire TIMEBOOST_net_12146;
wire TIMEBOOST_net_13639;
wire g57312_sb;
wire TIMEBOOST_net_13067;
wire g57313_sb;
wire TIMEBOOST_net_12147;
wire TIMEBOOST_net_13638;
wire g57314_sb;
wire TIMEBOOST_net_12206;
wire TIMEBOOST_net_13641;
wire g57315_sb;
wire TIMEBOOST_net_13068;
wire g57316_sb;
wire TIMEBOOST_net_12148;
wire TIMEBOOST_net_13653;
wire g57317_sb;
wire TIMEBOOST_net_12149;
wire TIMEBOOST_net_13637;
wire g57318_sb;
wire TIMEBOOST_net_6225;
wire TIMEBOOST_net_13651;
wire g57319_sb;
wire TIMEBOOST_net_6226;
wire TIMEBOOST_net_14557;
wire g57320_sb;
wire TIMEBOOST_net_10641;
wire TIMEBOOST_net_14558;
wire g57321_sb;
wire TIMEBOOST_net_10786;
wire TIMEBOOST_net_11779;
wire g57322_sb;
wire TIMEBOOST_net_13305;
wire TIMEBOOST_net_12187;
wire g57323_sb;
wire TIMEBOOST_net_6228;
wire TIMEBOOST_net_14515;
wire g57324_sb;
wire TIMEBOOST_net_11472;
wire TIMEBOOST_net_13648;
wire g57325_sb;
wire TIMEBOOST_net_12072;
wire TIMEBOOST_net_13642;
wire g57326_sb;
wire TIMEBOOST_net_12150;
wire TIMEBOOST_net_13611;
wire g57327_sb;
wire TIMEBOOST_net_6232;
wire TIMEBOOST_net_14176;
wire g57328_sb;
wire TIMEBOOST_net_12156;
wire TIMEBOOST_net_13608;
wire g57329_sb;
wire TIMEBOOST_net_12157;
wire TIMEBOOST_net_2300;
wire g57330_sb;
wire TIMEBOOST_net_10787;
wire g57331_db;
wire g57331_sb;
wire TIMEBOOST_net_12151;
wire TIMEBOOST_net_2301;
wire g57332_sb;
wire TIMEBOOST_net_12070;
wire TIMEBOOST_net_11192;
wire g57333_sb;
wire TIMEBOOST_net_12071;
wire TIMEBOOST_net_13955;
wire g57334_sb;
wire TIMEBOOST_net_12073;
wire TIMEBOOST_net_14027;
wire g57335_sb;
wire TIMEBOOST_net_12074;
wire TIMEBOOST_net_11168;
wire g57336_sb;
wire TIMEBOOST_net_6240;
wire TIMEBOOST_net_14066;
wire g57337_sb;
wire TIMEBOOST_net_6241;
wire TIMEBOOST_net_2307;
wire g57338_sb;
wire TIMEBOOST_net_6242;
wire TIMEBOOST_net_14160;
wire g57339_sb;
wire TIMEBOOST_net_13069;
wire g57340_sb;
wire TIMEBOOST_net_13070;
wire g57341_sb;
wire TIMEBOOST_net_6243;
wire TIMEBOOST_net_2309;
wire g57342_sb;
wire TIMEBOOST_net_6244;
wire TIMEBOOST_net_2310;
wire g57343_sb;
wire TIMEBOOST_net_6245;
wire TIMEBOOST_net_13957;
wire g57344_sb;
wire TIMEBOOST_net_13071;
wire g57345_sb;
wire TIMEBOOST_net_6246;
wire TIMEBOOST_net_13551;
wire g57346_sb;
wire TIMEBOOST_net_2529;
wire TIMEBOOST_net_11780;
wire g57347_sb;
wire TIMEBOOST_net_6247;
wire TIMEBOOST_net_13626;
wire g57348_sb;
wire TIMEBOOST_net_6248;
wire TIMEBOOST_net_13559;
wire g57349_sb;
wire TIMEBOOST_net_6249;
wire TIMEBOOST_net_13473;
wire g57350_sb;
wire TIMEBOOST_net_13474;
wire g57351_sb;
wire TIMEBOOST_net_14549;
wire g57352_sb;
wire TIMEBOOST_net_10814;
wire TIMEBOOST_net_11726;
wire g57353_sb;
wire TIMEBOOST_net_4341;
wire g57354_sb;
wire TIMEBOOST_net_13609;
wire g57355_sb;
wire TIMEBOOST_net_6510;
wire TIMEBOOST_net_13072;
wire g57356_sb;
wire TIMEBOOST_net_6253;
wire TIMEBOOST_net_13584;
wire g57357_sb;
wire TIMEBOOST_net_14550;
wire g57358_sb;
wire TIMEBOOST_net_13568;
wire g57359_sb;
wire TIMEBOOST_net_13645;
wire g57360_sb;
wire TIMEBOOST_net_13631;
wire g57361_sb;
wire TIMEBOOST_net_13628;
wire g57362_sb;
wire TIMEBOOST_net_13565;
wire g57363_sb;
wire TIMEBOOST_net_6511;
wire TIMEBOOST_net_13073;
wire g57364_sb;
wire TIMEBOOST_net_13566;
wire g57365_sb;
wire TIMEBOOST_net_13627;
wire g57366_sb;
wire TIMEBOOST_net_13074;
wire g57367_sb;
wire TIMEBOOST_net_6262;
wire TIMEBOOST_net_13486;
wire g57368_sb;
wire TIMEBOOST_net_12084;
wire TIMEBOOST_net_13552;
wire g57369_sb;
wire TIMEBOOST_net_13484;
wire TIMEBOOST_net_12188;
wire g57370_sb;
wire TIMEBOOST_net_6264;
wire TIMEBOOST_net_13570;
wire g57371_sb;
wire TIMEBOOST_net_6265;
wire TIMEBOOST_net_13636;
wire g57372_sb;
wire TIMEBOOST_net_6266;
wire TIMEBOOST_net_13556;
wire g57373_sb;
wire TIMEBOOST_net_13640;
wire g57374_sb;
wire n_13466;
wire g57375_sb;
wire TIMEBOOST_net_13603;
wire g57376_sb;
wire TIMEBOOST_net_6513;
wire TIMEBOOST_net_13075;
wire g57377_sb;
wire n_13460;
wire g57378_sb;
wire TIMEBOOST_net_13076;
wire g57379_sb;
wire TIMEBOOST_net_6271;
wire TIMEBOOST_net_13604;
wire g57380_sb;
wire TIMEBOOST_net_14182;
wire g57381_sb;
wire TIMEBOOST_net_13488;
wire g57382_sb;
wire TIMEBOOST_net_13482;
wire g57383_sb;
wire TIMEBOOST_net_13492;
wire g57384_sb;
wire TIMEBOOST_net_13493;
wire g57385_sb;
wire TIMEBOOST_net_13606;
wire g57386_sb;
wire TIMEBOOST_net_6515;
wire TIMEBOOST_net_13077;
wire g57387_sb;
wire TIMEBOOST_net_14418;
wire g57388_sb;
wire TIMEBOOST_net_13646;
wire g57389_sb;
wire TIMEBOOST_net_13851;
wire g57390_sb;
wire TIMEBOOST_net_13852;
wire g57391_sb;
wire TIMEBOOST_net_13625;
wire g57392_sb;
wire TIMEBOOST_net_13624;
wire g57393_sb;
wire TIMEBOOST_net_9310;
wire g57394_db;
wire g57394_sb;
wire TIMEBOOST_net_10789;
wire g57395_db;
wire g57395_sb;
wire TIMEBOOST_net_13567;
wire g57396_sb;
wire TIMEBOOST_net_13569;
wire g57397_sb;
wire TIMEBOOST_net_13649;
wire g57398_sb;
wire TIMEBOOST_net_6287;
wire TIMEBOOST_net_13553;
wire g57399_sb;
wire TIMEBOOST_net_6288;
wire TIMEBOOST_net_13555;
wire g57400_sb;
wire TIMEBOOST_net_12164;
wire TIMEBOOST_net_13605;
wire g57401_sb;
wire TIMEBOOST_net_6516;
wire TIMEBOOST_net_13078;
wire g57402_sb;
wire TIMEBOOST_net_11327;
wire g57403_sb;
wire TIMEBOOST_net_13010;
wire TIMEBOOST_net_11781;
wire g57404_sb;
wire TIMEBOOST_net_13079;
wire g57405_sb;
wire TIMEBOOST_net_6518;
wire TIMEBOOST_net_13082;
wire g57406_sb;
wire TIMEBOOST_net_6291;
wire TIMEBOOST_net_13607;
wire g57407_sb;
wire TIMEBOOST_net_12162;
wire TIMEBOOST_net_13472;
wire g57408_sb;
wire TIMEBOOST_net_6293;
wire TIMEBOOST_net_14551;
wire g57409_sb;
wire TIMEBOOST_net_12163;
wire TIMEBOOST_net_14552;
wire g57410_sb;
wire TIMEBOOST_net_12101;
wire TIMEBOOST_net_13592;
wire g57411_sb;
wire TIMEBOOST_net_12103;
wire TIMEBOOST_net_14553;
wire g57412_sb;
wire TIMEBOOST_net_6519;
wire TIMEBOOST_net_13083;
wire g57413_sb;
wire TIMEBOOST_net_12104;
wire TIMEBOOST_net_13475;
wire g57414_sb;
wire TIMEBOOST_net_6520;
wire TIMEBOOST_net_4798;
wire g57415_sb;
wire TIMEBOOST_net_12105;
wire TIMEBOOST_net_13593;
wire g57416_sb;
wire TIMEBOOST_net_12127;
wire TIMEBOOST_net_14554;
wire g57417_sb;
wire TIMEBOOST_net_12128;
wire TIMEBOOST_net_13594;
wire g57418_sb;
wire TIMEBOOST_net_12129;
wire TIMEBOOST_net_13610;
wire g57419_sb;
wire TIMEBOOST_net_12119;
wire TIMEBOOST_net_13595;
wire g57420_sb;
wire TIMEBOOST_net_14096;
wire TIMEBOOST_net_11727;
wire g57421_sb;
wire TIMEBOOST_net_12122;
wire TIMEBOOST_net_13476;
wire g57422_sb;
wire TIMEBOOST_net_13477;
wire g57423_sb;
wire TIMEBOOST_net_12108;
wire TIMEBOOST_net_13596;
wire g57424_sb;
wire TIMEBOOST_net_13597;
wire g57425_sb;
wire TIMEBOOST_net_13598;
wire g57426_sb;
wire TIMEBOOST_net_12112;
wire TIMEBOOST_net_13599;
wire g57427_sb;
wire TIMEBOOST_net_12115;
wire TIMEBOOST_net_13478;
wire g57428_sb;
wire TIMEBOOST_net_12117;
wire TIMEBOOST_net_13601;
wire g57429_sb;
wire TIMEBOOST_net_12124;
wire TIMEBOOST_net_13479;
wire g57430_sb;
wire TIMEBOOST_net_1724;
wire g57431_sb;
wire TIMEBOOST_net_12126;
wire TIMEBOOST_net_13480;
wire g57432_sb;
wire TIMEBOOST_net_12102;
wire TIMEBOOST_net_13495;
wire g57433_sb;
wire TIMEBOOST_net_13600;
wire g57434_sb;
wire TIMEBOOST_net_12111;
wire TIMEBOOST_net_13494;
wire g57435_sb;
wire TIMEBOOST_net_12120;
wire TIMEBOOST_net_4355;
wire g57436_sb;
wire TIMEBOOST_net_12121;
wire TIMEBOOST_net_14178;
wire g57437_sb;
wire TIMEBOOST_net_13489;
wire g57438_sb;
wire TIMEBOOST_net_13585;
wire g57439_sb;
wire TIMEBOOST_net_12107;
wire TIMEBOOST_net_14539;
wire g57440_sb;
wire TIMEBOOST_net_12110;
wire TIMEBOOST_net_1751;
wire g57441_sb;
wire TIMEBOOST_net_13044;
wire g57442_sb;
wire TIMEBOOST_net_12113;
wire TIMEBOOST_net_13586;
wire g57443_sb;
wire TIMEBOOST_net_13269;
wire TIMEBOOST_net_11445;
wire g57444_sb;
wire TIMEBOOST_net_13270;
wire TIMEBOOST_net_6440;
wire g57445_sb;
wire TIMEBOOST_net_13046;
wire g57446_sb;
wire TIMEBOOST_net_12114;
wire TIMEBOOST_net_14538;
wire g57447_sb;
wire TIMEBOOST_net_13271;
wire TIMEBOOST_net_11782;
wire g57448_sb;
wire TIMEBOOST_net_6525;
wire TIMEBOOST_net_13045;
wire g57449_sb;
wire TIMEBOOST_net_13057;
wire g57450_sb;
wire TIMEBOOST_net_13229;
wire TIMEBOOST_net_13272;
wire g57451_sb;
wire TIMEBOOST_net_12116;
wire TIMEBOOST_net_1846;
wire g57452_sb;
wire TIMEBOOST_net_12118;
wire TIMEBOOST_net_1844;
wire g57453_sb;
wire TIMEBOOST_net_12123;
wire TIMEBOOST_net_13588;
wire g57454_sb;
wire TIMEBOOST_net_12125;
wire TIMEBOOST_net_13487;
wire g57455_sb;
wire TIMEBOOST_net_12106;
wire TIMEBOOST_net_14517;
wire g57456_sb;
wire TIMEBOOST_net_13954;
wire TIMEBOOST_net_11728;
wire g57457_sb;
wire TIMEBOOST_net_12109;
wire TIMEBOOST_net_13468;
wire g57458_sb;
wire TIMEBOOST_net_6329;
wire TIMEBOOST_net_13554;
wire g57459_sb;
wire TIMEBOOST_net_6330;
wire TIMEBOOST_net_13548;
wire g57460_sb;
wire TIMEBOOST_net_6527;
wire TIMEBOOST_net_13088;
wire g57461_sb;
wire TIMEBOOST_net_13549;
wire g57462_sb;
wire TIMEBOOST_net_14221;
wire g57463_sb;
wire TIMEBOOST_net_6528;
wire TIMEBOOST_net_13084;
wire g57464_sb;
wire TIMEBOOST_net_13550;
wire g57465_sb;
wire TIMEBOOST_net_13562;
wire g57466_sb;
wire TIMEBOOST_net_13490;
wire g57467_sb;
wire TIMEBOOST_net_13085;
wire g57468_sb;
wire TIMEBOOST_net_6530;
wire TIMEBOOST_net_13049;
wire g57469_sb;
wire TIMEBOOST_net_13276;
wire n_1582;
wire g57470_sb;
wire TIMEBOOST_net_6531;
wire TIMEBOOST_net_13491;
wire g57471_sb;
wire TIMEBOOST_net_6532;
wire TIMEBOOST_net_13267;
wire g57472_sb;
wire TIMEBOOST_net_13469;
wire g57473_sb;
wire TIMEBOOST_net_6337;
wire TIMEBOOST_net_14510;
wire g57474_sb;
wire TIMEBOOST_net_13056;
wire g57475_sb;
wire TIMEBOOST_net_2408;
wire g57476_sb;
wire TIMEBOOST_net_2409;
wire g57477_sb;
wire TIMEBOOST_net_13266;
wire TIMEBOOST_net_13274;
wire g57478_sb;
wire TIMEBOOST_net_10432;
wire g57479_sb;
wire TIMEBOOST_net_6341;
wire TIMEBOOST_net_14219;
wire g57480_sb;
wire TIMEBOOST_net_2412;
wire g57481_sb;
wire TIMEBOOST_net_13360;
wire g57482_sb;
wire TIMEBOOST_net_13454;
wire g57483_sb;
wire TIMEBOOST_net_13463;
wire g57484_sb;
wire TIMEBOOST_net_6534;
wire TIMEBOOST_net_13051;
wire g57485_sb;
wire TIMEBOOST_net_13464;
wire g57486_sb;
wire TIMEBOOST_net_13086;
wire g57487_sb;
wire TIMEBOOST_net_13447;
wire g57488_sb;
wire TIMEBOOST_net_14067;
wire g57489_db;
wire g57489_sb;
wire TIMEBOOST_net_13452;
wire g57490_sb;
wire TIMEBOOST_net_13453;
wire g57491_sb;
wire TIMEBOOST_net_579;
wire g57492_sb;
wire TIMEBOOST_net_13446;
wire g57493_sb;
wire TIMEBOOST_net_11338;
wire g57494_sb;
wire TIMEBOOST_net_1726;
wire g57495_sb;
wire TIMEBOOST_net_337;
wire g57496_sb;
wire TIMEBOOST_net_13425;
wire g57497_sb;
wire TIMEBOOST_net_13429;
wire g57498_sb;
wire TIMEBOOST_net_12170;
wire TIMEBOOST_net_13427;
wire g57499_sb;
wire TIMEBOOST_net_13430;
wire g57500_sb;
wire TIMEBOOST_net_6359;
wire TIMEBOOST_net_11339;
wire g57501_sb;
wire TIMEBOOST_net_13440;
wire g57502_sb;
wire TIMEBOOST_net_6361;
wire TIMEBOOST_net_2431;
wire g57503_sb;
wire TIMEBOOST_net_12098;
wire TIMEBOOST_net_11340;
wire g57504_sb;
wire TIMEBOOST_net_6536;
wire TIMEBOOST_net_13052;
wire g57505_sb;
wire TIMEBOOST_net_12099;
wire TIMEBOOST_net_13439;
wire g57506_sb;
wire TIMEBOOST_net_12088;
wire TIMEBOOST_net_13438;
wire g57507_sb;
wire TIMEBOOST_net_12089;
wire TIMEBOOST_net_13437;
wire g57508_sb;
wire TIMEBOOST_net_12095;
wire TIMEBOOST_net_13436;
wire g57509_sb;
wire TIMEBOOST_net_13275;
wire TIMEBOOST_net_6441;
wire g57510_sb;
wire TIMEBOOST_net_12093;
wire TIMEBOOST_net_13433;
wire g57511_sb;
wire TIMEBOOST_net_12094;
wire TIMEBOOST_net_13434;
wire g57512_sb;
wire TIMEBOOST_net_12097;
wire TIMEBOOST_net_13428;
wire g57513_sb;
wire TIMEBOOST_net_12085;
wire TIMEBOOST_net_13435;
wire g57514_sb;
wire TIMEBOOST_net_12091;
wire TIMEBOOST_net_13426;
wire g57515_sb;
wire TIMEBOOST_net_12100;
wire g57516_db;
wire TIMEBOOST_net_12096;
wire TIMEBOOST_net_13431;
wire g57517_sb;
wire TIMEBOOST_net_12201;
wire TIMEBOOST_net_13061;
wire g57518_sb;
wire TIMEBOOST_net_6374;
wire n_3914;
wire g57519_sb;
wire TIMEBOOST_net_12086;
wire TIMEBOOST_net_13408;
wire g57520_sb;
wire TIMEBOOST_net_12202;
wire TIMEBOOST_net_13063;
wire g57521_sb;
wire TIMEBOOST_net_12203;
wire TIMEBOOST_net_13053;
wire g57522_sb;
wire TIMEBOOST_net_12092;
wire TIMEBOOST_net_13409;
wire g57523_sb;
wire TIMEBOOST_net_6377;
wire TIMEBOOST_net_2446;
wire g57524_sb;
wire TIMEBOOST_net_12197;
wire g53938_da;
wire g57525_sb;
wire TIMEBOOST_net_12068;
wire TIMEBOOST_net_13411;
wire g57526_sb;
wire TIMEBOOST_net_6380;
wire TIMEBOOST_net_13403;
wire g57527_sb;
wire TIMEBOOST_net_12204;
wire TIMEBOOST_net_13054;
wire g57528_sb;
wire TIMEBOOST_net_9367;
wire TIMEBOOST_net_11729;
wire g57529_sb;
wire TIMEBOOST_net_6381;
wire TIMEBOOST_net_13404;
wire g57530_sb;
wire TIMEBOOST_net_6382;
wire TIMEBOOST_net_13405;
wire g57531_sb;
wire TIMEBOOST_net_12205;
wire TIMEBOOST_net_13081;
wire g57532_sb;
wire TIMEBOOST_net_6383;
wire TIMEBOOST_net_4245;
wire g57533_sb;
wire TIMEBOOST_net_6384;
wire TIMEBOOST_net_13407;
wire g57534_sb;
wire TIMEBOOST_net_6385;
wire TIMEBOOST_net_13406;
wire g57535_sb;
wire TIMEBOOST_net_6542;
wire TIMEBOOST_net_13062;
wire g57536_sb;
wire TIMEBOOST_net_13237;
wire TIMEBOOST_net_6442;
wire g57537_sb;
wire TIMEBOOST_net_12172;
wire TIMEBOOST_net_13393;
wire g57538_sb;
wire TIMEBOOST_net_6387;
wire TIMEBOOST_net_13394;
wire g57539_sb;
wire TIMEBOOST_net_12180;
wire TIMEBOOST_net_13087;
wire g57540_sb;
wire TIMEBOOST_net_12182;
wire TIMEBOOST_net_13089;
wire g57541_sb;
wire TIMEBOOST_net_12183;
wire TIMEBOOST_net_13090;
wire g57542_sb;
wire TIMEBOOST_net_2540;
wire g57543_db;
wire g57543_sb;
wire TIMEBOOST_net_12185;
wire TIMEBOOST_net_13050;
wire g57544_sb;
wire TIMEBOOST_net_6388;
wire TIMEBOOST_net_13396;
wire g57545_sb;
wire TIMEBOOST_net_12026;
wire TIMEBOOST_net_13395;
wire g57546_sb;
wire TIMEBOOST_net_6547;
wire TIMEBOOST_net_13091;
wire g57547_sb;
wire TIMEBOOST_net_6390;
wire TIMEBOOST_net_13397;
wire g57548_sb;
wire TIMEBOOST_net_6391;
wire TIMEBOOST_net_13415;
wire g57549_sb;
wire TIMEBOOST_net_13241;
wire TIMEBOOST_net_4129;
wire g57550_sb;
wire TIMEBOOST_net_6392;
wire TIMEBOOST_net_13390;
wire g57551_sb;
wire TIMEBOOST_net_6393;
wire TIMEBOOST_net_13392;
wire g57552_sb;
wire TIMEBOOST_net_6394;
wire TIMEBOOST_net_13388;
wire g57553_sb;
wire TIMEBOOST_net_6395;
wire TIMEBOOST_net_13380;
wire g57554_sb;
wire TIMEBOOST_net_6396;
wire TIMEBOOST_net_13381;
wire g57555_sb;
wire TIMEBOOST_net_6397;
wire TIMEBOOST_net_13382;
wire g57556_sb;
wire TIMEBOOST_net_12087;
wire TIMEBOOST_net_13383;
wire g57557_sb;
wire TIMEBOOST_net_12189;
wire TIMEBOOST_net_13092;
wire g57558_sb;
wire TIMEBOOST_net_13094;
wire g57559_sb;
wire TIMEBOOST_net_12090;
wire TIMEBOOST_net_13455;
wire g57560_sb;
wire TIMEBOOST_net_6550;
wire TIMEBOOST_net_13048;
wire g57561_sb;
wire TIMEBOOST_net_12218;
wire TIMEBOOST_net_13080;
wire g57562_sb;
wire TIMEBOOST_net_12219;
wire TIMEBOOST_net_13095;
wire g57563_sb;
wire TIMEBOOST_net_6400;
wire TIMEBOOST_net_13456;
wire g57564_sb;
wire TIMEBOOST_net_13932;
wire g57565_db;
wire g57565_sb;
wire TIMEBOOST_net_12217;
wire TIMEBOOST_net_13055;
wire g57566_sb;
wire TIMEBOOST_net_13216;
wire g57567_sb;
wire TIMEBOOST_net_6401;
wire TIMEBOOST_net_11337;
wire g57568_sb;
wire TIMEBOOST_net_11406;
wire TIMEBOOST_net_13457;
wire g57569_sb;
wire TIMEBOOST_net_6403;
wire TIMEBOOST_net_13458;
wire g57570_sb;
wire TIMEBOOST_net_14548;
wire TIMEBOOST_net_11816;
wire g57571_sb;
wire TIMEBOOST_net_6404;
wire TIMEBOOST_net_13459;
wire g57572_sb;
wire TIMEBOOST_net_12216;
wire TIMEBOOST_net_13022;
wire g57573_sb;
wire TIMEBOOST_net_6405;
wire TIMEBOOST_net_13460;
wire g57574_sb;
wire TIMEBOOST_net_12069;
wire TIMEBOOST_net_13467;
wire g57575_sb;
wire TIMEBOOST_net_10743;
wire TIMEBOOST_net_13384;
wire g57576_sb;
wire TIMEBOOST_net_6408;
wire TIMEBOOST_net_2477;
wire g57577_sb;
wire TIMEBOOST_net_13218;
wire TIMEBOOST_net_11817;
wire g57578_sb;
wire TIMEBOOST_net_6409;
wire TIMEBOOST_net_13461;
wire g57579_sb;
wire TIMEBOOST_net_6410;
wire TIMEBOOST_net_13462;
wire g57580_sb;
wire TIMEBOOST_net_12220;
wire TIMEBOOST_net_13849;
wire g57581_sb;
wire TIMEBOOST_net_6556;
wire TIMEBOOST_net_13361;
wire g57582_sb;
wire TIMEBOOST_net_6411;
wire TIMEBOOST_net_13352;
wire g57583_sb;
wire TIMEBOOST_net_13347;
wire g57584_sb;
wire TIMEBOOST_net_6413;
wire g57585_db;
wire TIMEBOOST_net_6557;
wire TIMEBOOST_net_13024;
wire g57586_sb;
wire TIMEBOOST_net_6414;
wire TIMEBOOST_net_13353;
wire g57587_sb;
wire TIMEBOOST_net_6558;
wire TIMEBOOST_net_14179;
wire g57588_sb;
wire TIMEBOOST_net_13354;
wire g57589_sb;
wire TIMEBOOST_net_6416;
wire TIMEBOOST_net_13355;
wire g57590_sb;
wire TIMEBOOST_net_6559;
wire TIMEBOOST_net_13356;
wire g57591_sb;
wire TIMEBOOST_net_6417;
wire TIMEBOOST_net_13357;
wire g57592_sb;
wire TIMEBOOST_net_6418;
wire TIMEBOOST_net_13345;
wire g57593_sb;
wire TIMEBOOST_net_6560;
wire TIMEBOOST_net_13014;
wire g57594_sb;
wire TIMEBOOST_net_6419;
wire TIMEBOOST_net_13385;
wire g57595_sb;
wire TIMEBOOST_net_6420;
wire TIMEBOOST_net_13348;
wire g57596_sb;
wire TIMEBOOST_net_6421;
wire TIMEBOOST_net_4106;
wire g57597_sb;
wire TIMEBOOST_net_6422;
wire TIMEBOOST_net_13317;
wire g57598_sb;
wire g57779_da;
wire TIMEBOOST_net_15221;
wire g57780_da;
wire TIMEBOOST_net_11885;
wire g57780_sb;
wire g57781_da;
wire TIMEBOOST_net_11874;
wire TIMEBOOST_net_12646;
wire TIMEBOOST_net_14633;
wire TIMEBOOST_net_12681;
wire TIMEBOOST_net_10779;
wire TIMEBOOST_net_12697;
wire TIMEBOOST_net_14337;
wire TIMEBOOST_net_12699;
wire TIMEBOOST_net_2037;
wire TIMEBOOST_net_12641;
wire TIMEBOOST_net_14792;
wire g57787_da;
wire TIMEBOOST_net_2039;
wire g57788_da;
wire TIMEBOOST_net_10827;
wire g57789_da;
wire TIMEBOOST_net_14936;
wire TIMEBOOST_net_13991;
wire g57790_sb;
wire TIMEBOOST_net_14053;
wire TIMEBOOST_net_1997;
wire g57794_da;
wire g57794_db;
wire g57794_sb;
wire g57795_da;
wire TIMEBOOST_net_15223;
wire g57795_sb;
wire TIMEBOOST_net_14669;
wire TIMEBOOST_net_14563;
wire TIMEBOOST_net_9609;
wire TIMEBOOST_net_13963;
wire g57797_sb;
wire TIMEBOOST_net_3025;
wire TIMEBOOST_net_14099;
wire TIMEBOOST_net_14993;
wire TIMEBOOST_net_14360;
wire TIMEBOOST_net_3027;
wire TIMEBOOST_net_14038;
wire TIMEBOOST_net_3028;
wire TIMEBOOST_net_14011;
wire TIMEBOOST_net_14094;
wire TIMEBOOST_net_14014;
wire g57856_p;
wire g57863_p;
wire g57864_p;
wire TIMEBOOST_net_13318;
wire TIMEBOOST_net_13268;
wire g57875_sb;
wire g57876_p;
wire g57878_p;
wire g57890_da;
wire g57890_db;
wire g57890_sb;
wire TIMEBOOST_net_10862;
wire g57891_db;
wire g57891_sb;
wire g57892_da;
wire g57892_db;
wire g57892_sb;
wire TIMEBOOST_net_12311;
wire g57893_db;
wire g57893_sb;
wire TIMEBOOST_net_10863;
wire g57894_db;
wire g57894_sb;
wire TIMEBOOST_net_10864;
wire g57895_db;
wire g57895_sb;
wire TIMEBOOST_net_13542;
wire g57896_db;
wire g57896_sb;
wire TIMEBOOST_net_10865;
wire g57897_db;
wire g57897_sb;
wire TIMEBOOST_net_10876;
wire g57898_db;
wire g57898_sb;
wire TIMEBOOST_net_3335;
wire g57899_db;
wire g57899_sb;
wire TIMEBOOST_net_10883;
wire g57900_db;
wire g57900_sb;
wire g57901_da;
wire g57901_db;
wire g57901_sb;
wire TIMEBOOST_net_9557;
wire g57902_db;
wire g57902_sb;
wire TIMEBOOST_net_10884;
wire g57903_db;
wire g57903_sb;
wire TIMEBOOST_net_10903;
wire g57904_db;
wire g57904_sb;
wire g57905_da;
wire g57905_db;
wire g57905_sb;
wire TIMEBOOST_net_11029;
wire g57906_db;
wire g57906_sb;
wire g57907_da;
wire g57907_db;
wire g57907_sb;
wire TIMEBOOST_net_13319;
wire TIMEBOOST_net_13265;
wire g57908_sb;
wire TIMEBOOST_net_13113;
wire TIMEBOOST_net_14729;
wire g57909_sb;
wire TIMEBOOST_net_509;
wire TIMEBOOST_net_12581;
wire g57910_sb;
wire TIMEBOOST_net_510;
wire TIMEBOOST_net_12444;
wire g57911_sb;
wire g57912_da;
wire g57912_db;
wire g57912_sb;
wire TIMEBOOST_net_13526;
wire g57913_db;
wire g57913_sb;
wire TIMEBOOST_net_13527;
wire g57914_db;
wire g57914_sb;
wire TIMEBOOST_net_511;
wire TIMEBOOST_net_3193;
wire g57915_sb;
wire TIMEBOOST_net_512;
wire TIMEBOOST_net_9543;
wire g57916_sb;
wire g57917_da;
wire g57917_db;
wire g57917_sb;
wire g57918_da;
wire g57918_db;
wire g57918_sb;
wire TIMEBOOST_net_4309;
wire g57919_db;
wire g57919_sb;
wire TIMEBOOST_net_10488;
wire g57920_db;
wire g57920_sb;
wire g57921_da;
wire g57921_db;
wire g57921_sb;
wire TIMEBOOST_net_12784;
wire g57922_db;
wire g57922_sb;
wire TIMEBOOST_net_4855;
wire TIMEBOOST_net_3195;
wire g57923_sb;
wire TIMEBOOST_net_10805;
wire TIMEBOOST_net_3196;
wire g57924_sb;
wire TIMEBOOST_net_515;
wire TIMEBOOST_net_9548;
wire g57925_sb;
wire TIMEBOOST_net_4311;
wire g57926_db;
wire g57926_sb;
wire TIMEBOOST_net_12783;
wire g57927_db;
wire g57927_sb;
wire TIMEBOOST_net_9792;
wire g57928_db;
wire g57928_sb;
wire TIMEBOOST_net_10806;
wire TIMEBOOST_net_3198;
wire g57929_sb;
wire TIMEBOOST_net_9800;
wire g57930_db;
wire g57930_sb;
wire g57931_da;
wire g57931_db;
wire g57931_sb;
wire TIMEBOOST_net_10491;
wire g57932_db;
wire g57932_sb;
wire TIMEBOOST_net_13557;
wire g57933_db;
wire g57933_sb;
wire TIMEBOOST_net_10807;
wire g57934_db;
wire g57934_sb;
wire TIMEBOOST_net_4314;
wire g57935_db;
wire g57935_sb;
wire TIMEBOOST_net_9801;
wire g57936_db;
wire g57936_sb;
wire TIMEBOOST_net_4315;
wire g57937_db;
wire g57937_sb;
wire TIMEBOOST_net_4316;
wire g57938_db;
wire g57938_sb;
wire TIMEBOOST_net_10808;
wire TIMEBOOST_net_3199;
wire g57939_sb;
wire TIMEBOOST_net_3432;
wire g57940_db;
wire g57940_sb;
wire TIMEBOOST_net_3433;
wire g57941_db;
wire g57941_sb;
wire TIMEBOOST_net_321;
wire g57942_db;
wire g57942_sb;
wire TIMEBOOST_net_3434;
wire g57943_db;
wire TIMEBOOST_net_4317;
wire g57944_db;
wire g57944_sb;
wire TIMEBOOST_net_13558;
wire g57945_db;
wire g57945_sb;
wire TIMEBOOST_net_13560;
wire g57946_db;
wire g57946_sb;
wire TIMEBOOST_net_14514;
wire g57947_db;
wire g57947_sb;
wire TIMEBOOST_net_10809;
wire TIMEBOOST_net_3200;
wire g57948_sb;
wire g57949_da;
wire g57949_db;
wire g57949_sb;
wire g57950_da;
wire g57950_db;
wire TIMEBOOST_net_13561;
wire g57951_db;
wire g57951_sb;
wire TIMEBOOST_net_4321;
wire g57952_db;
wire g57952_sb;
wire g57953_da;
wire g57953_db;
wire g57953_sb;
wire g57954_da;
wire g57954_db;
wire g57954_sb;
wire TIMEBOOST_net_10810;
wire TIMEBOOST_net_3201;
wire TIMEBOOST_net_10804;
wire TIMEBOOST_net_3202;
wire g57956_sb;
wire TIMEBOOST_net_522;
wire TIMEBOOST_net_3203;
wire g57957_sb;
wire TIMEBOOST_net_13571;
wire g57958_db;
wire g57958_sb;
wire g57959_da;
wire g57959_db;
wire g57959_sb;
wire g57960_da;
wire g57960_db;
wire TIMEBOOST_net_5193;
wire TIMEBOOST_net_3204;
wire g57961_sb;
wire g57962_da;
wire g57962_db;
wire g57963_da;
wire g57963_db;
wire g57964_da;
wire g57964_db;
wire g57964_sb;
wire g57965_da;
wire g57965_db;
wire g57965_sb;
wire TIMEBOOST_net_10769;
wire TIMEBOOST_net_12259;
wire g57967_da;
wire g57967_db;
wire g57968_da;
wire g57968_db;
wire g57968_sb;
wire TIMEBOOST_net_4323;
wire g57969_db;
wire g57969_sb;
wire g57970_da;
wire g57970_db;
wire g57970_sb;
wire TIMEBOOST_net_525;
wire TIMEBOOST_net_3206;
wire g57971_sb;
wire g57972_da;
wire g57972_db;
wire g57972_sb;
wire TIMEBOOST_net_3435;
wire g57973_db;
wire g57973_sb;
wire TIMEBOOST_net_322;
wire TIMEBOOST_net_14969;
wire g57975_da;
wire g57975_db;
wire g57975_sb;
wire TIMEBOOST_net_10495;
wire g57976_db;
wire TIMEBOOST_net_10498;
wire g57977_db;
wire g57977_sb;
wire n_3426;
wire TIMEBOOST_net_3147;
wire g57978_sb;
wire TIMEBOOST_net_14790;
wire TIMEBOOST_net_3148;
wire g57979_sb;
wire TIMEBOOST_net_12888;
wire g57980_db;
wire g57980_sb;
wire TIMEBOOST_net_10499;
wire g57981_db;
wire g57981_sb;
wire TIMEBOOST_net_10501;
wire g57982_db;
wire g57982_sb;
wire TIMEBOOST_net_13577;
wire g57983_db;
wire g57983_sb;
wire TIMEBOOST_net_9541;
wire g57984_db;
wire g57984_sb;
wire TIMEBOOST_net_528;
wire TIMEBOOST_net_3149;
wire g57985_sb;
wire TIMEBOOST_net_12785;
wire g57986_db;
wire g57986_sb;
wire TIMEBOOST_net_10102;
wire TIMEBOOST_net_3150;
wire g57987_sb;
wire TIMEBOOST_net_530;
wire TIMEBOOST_net_3151;
wire g57988_sb;
wire TIMEBOOST_net_13578;
wire g57989_db;
wire g57989_sb;
wire g57990_da;
wire g57990_db;
wire g57990_sb;
wire TIMEBOOST_net_9793;
wire TIMEBOOST_net_15010;
wire g57991_sb;
wire TIMEBOOST_net_531;
wire TIMEBOOST_net_3152;
wire g57992_sb;
wire TIMEBOOST_net_12781;
wire g57993_db;
wire g57993_sb;
wire TIMEBOOST_net_13002;
wire g57994_db;
wire g57994_sb;
wire TIMEBOOST_net_4330;
wire g57995_db;
wire g57995_sb;
wire TIMEBOOST_net_532;
wire TIMEBOOST_net_3153;
wire g57996_sb;
wire g57997_da;
wire g57997_db;
wire g57997_sb;
wire TIMEBOOST_net_12872;
wire g57998_db;
wire TIMEBOOST_net_10502;
wire g57999_db;
wire g57999_sb;
wire g58000_da;
wire g58000_db;
wire g58000_sb;
wire TIMEBOOST_net_533;
wire TIMEBOOST_net_3154;
wire g58001_sb;
wire g58002_da;
wire g58002_db;
wire g58002_sb;
wire TIMEBOOST_net_12427;
wire g58003_db;
wire g58003_sb;
wire TIMEBOOST_net_4332;
wire g58004_db;
wire g58004_sb;
wire TIMEBOOST_net_12871;
wire g58005_db;
wire g58005_sb;
wire TIMEBOOST_net_4333;
wire g58006_db;
wire g58006_sb;
wire g58007_da;
wire g58007_db;
wire g58008_da;
wire g58008_db;
wire g58008_sb;
wire TIMEBOOST_net_10729;
wire TIMEBOOST_net_12430;
wire g58009_sb;
wire TIMEBOOST_net_535;
wire TIMEBOOST_net_3099;
wire g58010_sb;
wire g58011_da;
wire g58011_db;
wire g58011_sb;
wire TIMEBOOST_net_10503;
wire g58012_db;
wire g58012_sb;
wire TIMEBOOST_net_4335;
wire g58013_db;
wire g58013_sb;
wire TIMEBOOST_net_13336;
wire g58014_db;
wire g58014_sb;
wire g58015_da;
wire g58015_db;
wire g58015_sb;
wire g58016_da;
wire g58016_db;
wire g58016_sb;
wire TIMEBOOST_net_14609;
wire TIMEBOOST_net_12560;
wire g58017_sb;
wire TIMEBOOST_net_10385;
wire TIMEBOOST_net_12561;
wire g58018_sb;
wire TIMEBOOST_net_13760;
wire TIMEBOOST_net_12562;
wire g58019_sb;
wire g58020_da;
wire g58020_db;
wire g58020_sb;
wire g58021_da;
wire g58021_db;
wire g58021_sb;
wire TIMEBOOST_net_12419;
wire TIMEBOOST_net_14751;
wire g58022_sb;
wire g58023_da;
wire g58023_db;
wire g58023_sb;
wire g58024_da;
wire g58024_db;
wire g58024_sb;
wire TIMEBOOST_net_13377;
wire g58025_db;
wire g58025_sb;
wire TIMEBOOST_net_4338;
wire g58026_db;
wire g58026_sb;
wire TIMEBOOST_net_539;
wire g64856_db;
wire g58027_sb;
wire TIMEBOOST_net_4339;
wire TIMEBOOST_net_14696;
wire g58028_sb;
wire g58029_da;
wire g58029_db;
wire g58029_sb;
wire g58030_da;
wire g58030_db;
wire g58030_sb;
wire g58031_da;
wire g58031_db;
wire g58031_sb;
wire TIMEBOOST_net_540;
wire TIMEBOOST_net_12517;
wire g58032_sb;
wire g58033_da;
wire g58033_db;
wire g58033_sb;
wire TIMEBOOST_net_13536;
wire g58034_db;
wire g58034_sb;
wire TIMEBOOST_net_10524;
wire g58035_db;
wire g58035_sb;
wire g58036_da;
wire g58036_db;
wire g58036_sb;
wire g58037_da;
wire g58037_db;
wire g58037_sb;
wire TIMEBOOST_net_10526;
wire g58038_db;
wire g58039_da;
wire g58039_db;
wire g58039_sb;
wire TIMEBOOST_net_541;
wire g58040_db;
wire g58040_sb;
wire TIMEBOOST_net_542;
wire TIMEBOOST_net_3053;
wire g58041_sb;
wire TIMEBOOST_net_188;
wire g58042_db;
wire g58042_sb;
wire TIMEBOOST_net_4342;
wire TIMEBOOST_net_14742;
wire g58043_sb;
wire g58044_da;
wire g58044_db;
wire g58044_sb;
wire TIMEBOOST_net_13375;
wire g58045_db;
wire g58045_sb;
wire TIMEBOOST_net_9710;
wire g58046_db;
wire g58046_sb;
wire TIMEBOOST_net_4769;
wire g58047_db;
wire g58047_sb;
wire TIMEBOOST_net_4770;
wire g58048_db;
wire g58048_sb;
wire TIMEBOOST_net_543;
wire g58049_db;
wire g58049_sb;
wire TIMEBOOST_net_4344;
wire g58050_db;
wire g58050_sb;
wire TIMEBOOST_net_3342;
wire TIMEBOOST_net_12350;
wire g58051_sb;
wire TIMEBOOST_net_12976;
wire g58052_db;
wire g58052_sb;
wire TIMEBOOST_net_13114;
wire TIMEBOOST_net_12289;
wire g58053_sb;
wire TIMEBOOST_net_181;
wire g58054_db;
wire TIMEBOOST_net_4345;
wire TIMEBOOST_net_1091;
wire g58055_sb;
wire TIMEBOOST_net_544;
wire g58056_db;
wire g58056_sb;
wire TIMEBOOST_net_10368;
wire g58057_db;
wire g58057_sb;
wire g58058_da;
wire g58058_db;
wire g58058_sb;
wire TIMEBOOST_net_4347;
wire g58059_db;
wire g58059_sb;
wire TIMEBOOST_net_4348;
wire TIMEBOOST_net_12371;
wire g58060_sb;
wire TIMEBOOST_net_545;
wire g64939_db;
wire TIMEBOOST_net_4056;
wire TIMEBOOST_net_14689;
wire g58062_sb;
wire TIMEBOOST_net_13535;
wire g58063_db;
wire g58063_sb;
wire TIMEBOOST_net_323;
wire g58064_db;
wire TIMEBOOST_net_182;
wire g58065_db;
wire g58066_da;
wire g58066_db;
wire g58066_sb;
wire TIMEBOOST_net_13337;
wire g58067_db;
wire TIMEBOOST_net_4771;
wire TIMEBOOST_net_9853;
wire g58068_sb;
wire g58069_da;
wire g58069_db;
wire g58069_sb;
wire TIMEBOOST_net_546;
wire TIMEBOOST_net_12520;
wire g58070_sb;
wire TIMEBOOST_net_14144;
wire TIMEBOOST_net_12839;
wire g58071_sb;
wire g58072_da;
wire g58072_db;
wire g58072_sb;
wire g58073_da;
wire g58073_db;
wire g58073_sb;
wire TIMEBOOST_net_4350;
wire g58074_db;
wire g58074_sb;
wire TIMEBOOST_net_324;
wire g58075_db;
wire g58075_sb;
wire g58076_da;
wire g58076_db;
wire g58076_sb;
wire g58077_da;
wire g58077_db;
wire g58077_sb;
wire TIMEBOOST_net_548;
wire TIMEBOOST_net_12750;
wire g58078_sb;
wire TIMEBOOST_net_549;
wire TIMEBOOST_net_12837;
wire g58079_sb;
wire g58080_da;
wire g58080_db;
wire g58080_sb;
wire TIMEBOOST_net_13534;
wire g58081_db;
wire g58081_sb;
wire g58082_da;
wire g58082_db;
wire g58082_sb;
wire TIMEBOOST_net_550;
wire TIMEBOOST_net_12794;
wire g58083_sb;
wire g58084_da;
wire g58084_db;
wire g58084_sb;
wire g58085_da;
wire g58085_db;
wire TIMEBOOST_net_13378;
wire g58086_db;
wire g58086_sb;
wire g58087_da;
wire g58087_db;
wire g58087_sb;
wire TIMEBOOST_net_551;
wire g65679_da;
wire g58088_sb;
wire g58089_da;
wire g58089_db;
wire g58089_sb;
wire g58090_da;
wire g58090_db;
wire g58090_sb;
wire g58091_da;
wire g58091_db;
wire g58091_sb;
wire g58092_da;
wire g58092_db;
wire g58092_sb;
wire TIMEBOOST_net_10635;
wire TIMEBOOST_net_12721;
wire g58093_sb;
wire TIMEBOOST_net_9713;
wire g58094_db;
wire g58094_sb;
wire TIMEBOOST_net_13402;
wire g58095_db;
wire g58095_sb;
wire TIMEBOOST_net_4352;
wire g58096_db;
wire g58096_sb;
wire g58097_da;
wire g58097_db;
wire g58097_sb;
wire TIMEBOOST_net_4271;
wire TIMEBOOST_net_12500;
wire g58099_da;
wire g58099_db;
wire g58099_sb;
wire TIMEBOOST_net_10510;
wire g58100_db;
wire g58100_sb;
wire g58101_da;
wire g58101_db;
wire g58101_sb;
wire TIMEBOOST_net_12445;
wire g58102_db;
wire g58102_sb;
wire TIMEBOOST_net_3436;
wire g58103_db;
wire g58103_sb;
wire g58104_da;
wire g58104_db;
wire g58104_sb;
wire TIMEBOOST_net_4503;
wire TIMEBOOST_net_14336;
wire g58105_sb;
wire TIMEBOOST_net_326;
wire g58106_db;
wire g58106_sb;
wire TIMEBOOST_net_10733;
wire TIMEBOOST_net_14162;
wire g58107_sb;
wire TIMEBOOST_net_14429;
wire TIMEBOOST_net_12307;
wire g58108_sb;
wire g58109_da;
wire g58109_db;
wire TIMEBOOST_net_327;
wire g58110_db;
wire g58110_sb;
wire TIMEBOOST_net_328;
wire g58111_db;
wire g58111_sb;
wire TIMEBOOST_net_329;
wire g58112_db;
wire g58112_sb;
wire g58113_da;
wire g58113_db;
wire g58113_sb;
wire g58114_da;
wire g58114_db;
wire g58114_sb;
wire TIMEBOOST_net_13930;
wire g58115_db;
wire g58115_sb;
wire TIMEBOOST_net_556;
wire TIMEBOOST_net_14164;
wire g58116_sb;
wire TIMEBOOST_net_557;
wire TIMEBOOST_net_12667;
wire g58117_sb;
wire TIMEBOOST_net_330;
wire g58118_db;
wire g58118_sb;
wire g58119_da;
wire g58119_db;
wire g58119_sb;
wire TIMEBOOST_net_9951;
wire TIMEBOOST_net_14873;
wire g58120_sb;
wire TIMEBOOST_net_558;
wire g58121_db;
wire TIMEBOOST_net_12611;
wire TIMEBOOST_net_12308;
wire g58123_da;
wire g58123_db;
wire g58123_sb;
wire TIMEBOOST_net_331;
wire g58124_db;
wire g58124_sb;
wire TIMEBOOST_net_332;
wire g58125_db;
wire g58125_sb;
wire TIMEBOOST_net_14055;
wire TIMEBOOST_net_12644;
wire g58126_sb;
wire TIMEBOOST_net_4354;
wire g58127_db;
wire g58127_sb;
wire g58128_da;
wire g58128_db;
wire g58128_sb;
wire TIMEBOOST_net_333;
wire g58129_db;
wire g58129_sb;
wire TIMEBOOST_net_334;
wire g58130_db;
wire g58130_sb;
wire TIMEBOOST_net_13785;
wire TIMEBOOST_net_14357;
wire TIMEBOOST_net_9708;
wire g58132_db;
wire g58132_sb;
wire g58133_da;
wire g58133_db;
wire g58133_sb;
wire TIMEBOOST_net_335;
wire g58134_db;
wire g58135_da;
wire g58135_db;
wire TIMEBOOST_net_336;
wire g58136_db;
wire g58136_sb;
wire TIMEBOOST_net_10424;
wire TIMEBOOST_net_12309;
wire g58138_da;
wire g58138_db;
wire g58138_sb;
wire TIMEBOOST_net_13970;
wire TIMEBOOST_net_12518;
wire g58139_sb;
wire TIMEBOOST_net_562;
wire TIMEBOOST_net_12497;
wire g58140_sb;
wire g58141_da;
wire g58141_db;
wire g58141_sb;
wire g58142_da;
wire g58142_db;
wire g58142_sb;
wire TIMEBOOST_net_10511;
wire g58143_db;
wire g58143_sb;
wire TIMEBOOST_net_13587;
wire g58144_db;
wire g58144_sb;
wire g58145_da;
wire g58145_db;
wire g58145_sb;
wire g58146_da;
wire g58146_db;
wire g58146_sb;
wire TIMEBOOST_net_563;
wire TIMEBOOST_net_12466;
wire g58147_sb;
wire TIMEBOOST_net_14323;
wire TIMEBOOST_net_3108;
wire g58148_sb;
wire TIMEBOOST_net_13996;
wire TIMEBOOST_net_12902;
wire g58149_sb;
wire g58150_da;
wire g58150_db;
wire g58150_sb;
wire g58151_da;
wire g58151_db;
wire TIMEBOOST_net_13282;
wire g58152_db;
wire g58152_sb;
wire TIMEBOOST_net_14521;
wire TIMEBOOST_net_3110;
wire g58153_sb;
wire g58154_da;
wire g58154_db;
wire g58154_sb;
wire g58155_da;
wire g58155_db;
wire TIMEBOOST_net_10528;
wire g58156_db;
wire g58156_sb;
wire g58157_da;
wire g58157_db;
wire TIMEBOOST_net_14076;
wire TIMEBOOST_net_12479;
wire g58158_sb;
wire g58159_da;
wire g58159_db;
wire g58159_sb;
wire g58160_da;
wire g58160_db;
wire g58160_sb;
wire TIMEBOOST_net_338;
wire TIMEBOOST_net_12481;
wire g58161_sb;
wire g58162_da;
wire g58162_db;
wire g58162_sb;
wire TIMEBOOST_net_568;
wire TIMEBOOST_net_12482;
wire g58163_sb;
wire g58164_da;
wire g58164_db;
wire g58164_sb;
wire TIMEBOOST_net_12365;
wire g58165_db;
wire g58165_sb;
wire TIMEBOOST_net_10529;
wire g58166_db;
wire g58167_da;
wire g58167_db;
wire g58167_sb;
wire TIMEBOOST_net_4740;
wire g58168_db;
wire TIMEBOOST_net_10530;
wire g58169_db;
wire g58169_sb;
wire TIMEBOOST_net_569;
wire TIMEBOOST_net_12234;
wire g58170_sb;
wire TIMEBOOST_net_570;
wire TIMEBOOST_net_12235;
wire g58171_sb;
wire TIMEBOOST_net_3437;
wire g58172_db;
wire g58172_sb;
wire g58173_da;
wire g58173_db;
wire g58173_sb;
wire TIMEBOOST_net_4360;
wire g58174_db;
wire g58174_sb;
wire TIMEBOOST_net_10402;
wire g58175_db;
wire g58175_sb;
wire TIMEBOOST_net_3438;
wire g58176_db;
wire g58176_sb;
wire TIMEBOOST_net_571;
wire TIMEBOOST_net_12236;
wire g58177_sb;
wire TIMEBOOST_net_10880;
wire TIMEBOOST_net_12276;
wire g58178_sb;
wire TIMEBOOST_net_573;
wire TIMEBOOST_net_3211;
wire g58179_sb;
wire TIMEBOOST_net_13666;
wire g58180_db;
wire g58180_sb;
wire g58181_da;
wire g58181_db;
wire g58181_sb;
wire TIMEBOOST_net_9958;
wire g58182_db;
wire g58182_sb;
wire TIMEBOOST_net_9802;
wire g58183_db;
wire g58183_sb;
wire TIMEBOOST_net_9803;
wire g58184_db;
wire g58184_sb;
wire TIMEBOOST_net_4363;
wire g58185_db;
wire g58185_sb;
wire TIMEBOOST_net_4364;
wire g58186_db;
wire g58186_sb;
wire TIMEBOOST_net_574;
wire TIMEBOOST_net_9538;
wire g58187_sb;
wire TIMEBOOST_net_14525;
wire g58188_db;
wire g58188_sb;
wire TIMEBOOST_net_3441;
wire g58189_db;
wire g58189_sb;
wire TIMEBOOST_net_13661;
wire TIMEBOOST_net_14970;
wire g58190_sb;
wire TIMEBOOST_net_13660;
wire g58191_db;
wire g58191_sb;
wire TIMEBOOST_net_575;
wire TIMEBOOST_net_3213;
wire g58192_sb;
wire TIMEBOOST_net_3442;
wire g58193_db;
wire g58193_sb;
wire TIMEBOOST_net_10601;
wire g58194_db;
wire g58194_sb;
wire TIMEBOOST_net_13544;
wire g58195_db;
wire g58195_sb;
wire g58196_da;
wire g58196_db;
wire g58196_sb;
wire TIMEBOOST_net_4368;
wire g58197_db;
wire g58197_sb;
wire g58198_da;
wire g58198_db;
wire g58198_sb;
wire TIMEBOOST_net_10767;
wire TIMEBOOST_net_12474;
wire g58199_sb;
wire TIMEBOOST_net_577;
wire TIMEBOOST_net_12460;
wire g58200_sb;
wire g58201_da;
wire g58201_db;
wire g58201_sb;
wire g58202_da;
wire g58202_db;
wire g58202_sb;
wire TIMEBOOST_net_4369;
wire g58203_db;
wire g58203_sb;
wire TIMEBOOST_net_4370;
wire g58204_db;
wire g58204_sb;
wire g58205_da;
wire g58205_db;
wire g58205_sb;
wire TIMEBOOST_net_14796;
wire g58206_sb;
wire TIMEBOOST_net_10427;
wire g58207_db;
wire g58207_sb;
wire TIMEBOOST_net_580;
wire g58208_db;
wire g58208_sb;
wire g58209_da;
wire g58209_db;
wire g58209_sb;
wire TIMEBOOST_net_3351;
wire g58210_db;
wire g58210_sb;
wire g58211_da;
wire g58211_db;
wire g58211_sb;
wire TIMEBOOST_net_581;
wire TIMEBOOST_net_12461;
wire g58212_sb;
wire g58213_da;
wire g58213_db;
wire g58213_sb;
wire g58214_da;
wire g58214_db;
wire g58214_sb;
wire TIMEBOOST_net_10602;
wire g58215_db;
wire g58215_sb;
wire g58216_da;
wire g58216_db;
wire g58216_sb;
wire TIMEBOOST_net_582;
wire TIMEBOOST_net_3118;
wire g58217_sb;
wire g58218_da;
wire g58218_db;
wire g58218_sb;
wire g58219_da;
wire g58219_db;
wire g58219_sb;
wire g58220_da;
wire g58220_db;
wire g58220_sb;
wire g58221_da;
wire g58221_db;
wire g58221_sb;
wire TIMEBOOST_net_583;
wire TIMEBOOST_net_12462;
wire g58222_sb;
wire g58223_da;
wire g58223_db;
wire g58223_sb;
wire TIMEBOOST_net_3352;
wire g58224_db;
wire g58224_sb;
wire TIMEBOOST_net_340;
wire g58225_db;
wire g58225_sb;
wire g58226_da;
wire g58226_db;
wire TIMEBOOST_net_9586;
wire g58227_db;
wire g58227_sb;
wire TIMEBOOST_net_10608;
wire g58228_db;
wire g58228_sb;
wire TIMEBOOST_net_584;
wire TIMEBOOST_net_13101;
wire g58229_sb;
wire TIMEBOOST_net_9805;
wire g58230_db;
wire g58230_sb;
wire TIMEBOOST_net_10748;
wire TIMEBOOST_net_14350;
wire g58231_sb;
wire g58232_da;
wire g58232_db;
wire g58232_sb;
wire TIMEBOOST_net_10611;
wire g58233_db;
wire g58233_sb;
wire TIMEBOOST_net_4375;
wire g58234_db;
wire g58234_sb;
wire TIMEBOOST_net_4505;
wire TIMEBOOST_net_14372;
wire g58235_sb;
wire TIMEBOOST_net_3445;
wire g58236_db;
wire g58236_sb;
wire TIMEBOOST_net_585;
wire TIMEBOOST_net_12286;
wire g58237_sb;
wire TIMEBOOST_net_586;
wire TIMEBOOST_net_9578;
wire g58238_sb;
wire TIMEBOOST_net_587;
wire TIMEBOOST_net_9579;
wire g58239_sb;
wire TIMEBOOST_net_4772;
wire TIMEBOOST_net_12224;
wire g58240_sb;
wire g58241_da;
wire g58241_db;
wire TIMEBOOST_net_4506;
wire TIMEBOOST_net_14461;
wire g58242_sb;
wire g58243_da;
wire g58243_db;
wire g58243_sb;
wire TIMEBOOST_net_588;
wire TIMEBOOST_net_9575;
wire g58244_sb;
wire TIMEBOOST_net_3446;
wire g58245_db;
wire TIMEBOOST_net_9807;
wire g58246_db;
wire TIMEBOOST_net_10489;
wire g58247_db;
wire g58248_da;
wire g58248_db;
wire TIMEBOOST_net_589;
wire TIMEBOOST_net_9535;
wire g58250_da;
wire g58250_db;
wire TIMEBOOST_net_3353;
wire TIMEBOOST_net_15011;
wire g58251_sb;
wire g58252_da;
wire g58252_db;
wire g58252_sb;
wire TIMEBOOST_net_590;
wire TIMEBOOST_net_3220;
wire TIMEBOOST_net_10496;
wire TIMEBOOST_net_14389;
wire g58254_sb;
wire TIMEBOOST_net_9808;
wire g58255_db;
wire g58255_sb;
wire TIMEBOOST_net_13443;
wire g58256_db;
wire g58256_sb;
wire TIMEBOOST_net_9809;
wire g58257_db;
wire g58257_sb;
wire TIMEBOOST_net_4508;
wire TIMEBOOST_net_14392;
wire g58258_sb;
wire TIMEBOOST_net_4378;
wire g58259_db;
wire TIMEBOOST_net_11176;
wire TIMEBOOST_net_9539;
wire g58260_sb;
wire TIMEBOOST_net_5299;
wire TIMEBOOST_net_13987;
wire g58261_sb;
wire TIMEBOOST_net_3222;
wire g58262_db;
wire g58262_sb;
wire TIMEBOOST_net_4509;
wire TIMEBOOST_net_14409;
wire g58263_sb;
wire TIMEBOOST_net_3651;
wire g58264_db;
wire g58264_sb;
wire g58265_da;
wire g58265_db;
wire g58265_sb;
wire TIMEBOOST_net_3652;
wire g58266_db;
wire g58266_sb;
wire TIMEBOOST_net_12836;
wire g58267_db;
wire g58267_sb;
wire TIMEBOOST_net_183;
wire g58268_db;
wire g58268_sb;
wire TIMEBOOST_net_184;
wire g58269_db;
wire g58269_sb;
wire TIMEBOOST_net_14257;
wire g58270_db;
wire g58270_sb;
wire TIMEBOOST_net_10045;
wire g58271_db;
wire g58271_sb;
wire TIMEBOOST_net_14310;
wire TIMEBOOST_net_4773;
wire g58272_sb;
wire TIMEBOOST_net_14241;
wire TIMEBOOST_net_4774;
wire g58273_sb;
wire TIMEBOOST_net_10046;
wire g58274_db;
wire g58274_sb;
wire TIMEBOOST_net_10047;
wire g58275_db;
wire g58275_sb;
wire TIMEBOOST_net_10048;
wire g58276_db;
wire g58276_sb;
wire TIMEBOOST_net_4219;
wire g58277_db;
wire g58277_sb;
wire TIMEBOOST_net_4220;
wire g58278_db;
wire g58278_sb;
wire TIMEBOOST_net_4221;
wire g58279_db;
wire g58279_sb;
wire TIMEBOOST_net_14242;
wire TIMEBOOST_net_10818;
wire g58280_sb;
wire TIMEBOOST_net_14456;
wire TIMEBOOST_net_9339;
wire g58281_sb;
wire TIMEBOOST_net_14243;
wire TIMEBOOST_net_4776;
wire g58282_sb;
wire TIMEBOOST_net_4222;
wire g58283_db;
wire g58283_sb;
wire TIMEBOOST_net_4223;
wire g58284_db;
wire g58284_sb;
wire TIMEBOOST_net_4224;
wire g58285_db;
wire g58285_sb;
wire TIMEBOOST_net_14244;
wire TIMEBOOST_net_4777;
wire g58286_sb;
wire TIMEBOOST_net_4225;
wire g58287_db;
wire g58287_sb;
wire TIMEBOOST_net_4226;
wire g58288_db;
wire g58288_sb;
wire TIMEBOOST_net_4227;
wire g58289_db;
wire g58289_sb;
wire TIMEBOOST_net_10389;
wire g58290_db;
wire g58290_sb;
wire TIMEBOOST_net_14245;
wire TIMEBOOST_net_4778;
wire g58291_sb;
wire TIMEBOOST_net_13445;
wire g58292_db;
wire g58292_sb;
wire TIMEBOOST_net_10390;
wire g58293_db;
wire g58293_sb;
wire TIMEBOOST_net_13444;
wire g58294_db;
wire g58294_sb;
wire TIMEBOOST_net_10391;
wire g58295_db;
wire g58295_sb;
wire TIMEBOOST_net_4233;
wire TIMEBOOST_net_14415;
wire g58296_sb;
wire TIMEBOOST_net_4234;
wire g58297_db;
wire g58297_sb;
wire TIMEBOOST_net_4235;
wire g58298_db;
wire g58298_sb;
wire TIMEBOOST_net_9283;
wire TIMEBOOST_net_10140;
wire g58299_sb;
wire TIMEBOOST_net_14311;
wire TIMEBOOST_net_9340;
wire g58300_sb;
wire TIMEBOOST_net_4236;
wire g58301_db;
wire g58301_sb;
wire TIMEBOOST_net_4237;
wire g58302_db;
wire g58302_sb;
wire TIMEBOOST_net_4238;
wire g58303_db;
wire g58303_sb;
wire TIMEBOOST_net_4239;
wire g58304_db;
wire g58304_sb;
wire TIMEBOOST_net_4240;
wire g58305_db;
wire g58305_sb;
wire TIMEBOOST_net_4241;
wire TIMEBOOST_net_14452;
wire g58306_sb;
wire g58307_da;
wire g58307_db;
wire g58307_sb;
wire TIMEBOOST_net_12734;
wire TIMEBOOST_net_592;
wire g58308_sb;
wire TIMEBOOST_net_3655;
wire TIMEBOOST_net_593;
wire g58309_sb;
wire TIMEBOOST_net_3656;
wire g58310_db;
wire g58310_sb;
wire g58311_da;
wire TIMEBOOST_net_10480;
wire g58311_sb;
wire g58312_da;
wire g58312_db;
wire g58312_sb;
wire TIMEBOOST_net_3657;
wire TIMEBOOST_net_14824;
wire g58313_sb;
wire TIMEBOOST_net_3658;
wire g58314_db;
wire g58314_sb;
wire TIMEBOOST_net_3659;
wire TIMEBOOST_net_594;
wire g58315_sb;
wire TIMEBOOST_net_9957;
wire TIMEBOOST_net_595;
wire g58316_sb;
wire TIMEBOOST_net_3661;
wire TIMEBOOST_net_596;
wire g58317_sb;
wire g58318_da;
wire g58318_db;
wire g58318_sb;
wire TIMEBOOST_net_3662;
wire g58319_db;
wire g58319_sb;
wire g58320_da;
wire g58320_db;
wire g58320_sb;
wire TIMEBOOST_net_3663;
wire TIMEBOOST_net_597;
wire g58321_sb;
wire TIMEBOOST_net_9954;
wire g58322_db;
wire g58322_sb;
wire TIMEBOOST_net_3665;
wire g58323_db;
wire g58323_sb;
wire g58324_da;
wire g58324_db;
wire g58324_sb;
wire g58325_da;
wire g58325_db;
wire g58325_sb;
wire TIMEBOOST_net_9937;
wire TIMEBOOST_net_10985;
wire g58326_sb;
wire g58327_da;
wire g58327_db;
wire g58327_sb;
wire g58328_da;
wire g58328_db;
wire g58328_sb;
wire g58329_da;
wire g58329_db;
wire g58329_sb;
wire TIMEBOOST_net_3667;
wire g58330_db;
wire g58330_sb;
wire TIMEBOOST_net_9950;
wire g58331_db;
wire g58331_sb;
wire TIMEBOOST_net_3669;
wire g58332_db;
wire g58332_sb;
wire TIMEBOOST_net_15051;
wire TIMEBOOST_net_10141;
wire g58333_sb;
wire TIMEBOOST_net_3670;
wire TIMEBOOST_net_599;
wire g58334_sb;
wire g58335_da;
wire g58335_db;
wire g58335_sb;
wire TIMEBOOST_net_3671;
wire g58336_db;
wire g58336_sb;
wire g58337_da;
wire g58337_db;
wire g58337_sb;
wire TIMEBOOST_net_3672;
wire g58338_db;
wire g58338_sb;
wire TIMEBOOST_net_3673;
wire g58339_db;
wire g58339_sb;
wire TIMEBOOST_net_9933;
wire g58340_db;
wire g58340_sb;
wire TIMEBOOST_net_4779;
wire TIMEBOOST_net_14137;
wire g58341_sb;
wire TIMEBOOST_net_4242;
wire TIMEBOOST_net_600;
wire g58342_sb;
wire TIMEBOOST_net_4243;
wire TIMEBOOST_net_601;
wire g58343_sb;
wire TIMEBOOST_net_4244;
wire g58344_db;
wire g58344_sb;
wire TIMEBOOST_net_10400;
wire g58345_db;
wire g58345_sb;
wire TIMEBOOST_net_10401;
wire g58346_db;
wire g58346_sb;
wire TIMEBOOST_net_4247;
wire g58347_db;
wire g58347_sb;
wire TIMEBOOST_net_4780;
wire TIMEBOOST_net_14133;
wire g58348_sb;
wire TIMEBOOST_net_4248;
wire g58349_db;
wire g58349_sb;
wire TIMEBOOST_net_13254;
wire TIMEBOOST_net_602;
wire g58350_sb;
wire TIMEBOOST_net_11331;
wire TIMEBOOST_net_14070;
wire g58351_sb;
wire TIMEBOOST_net_10200;
wire g58352_db;
wire g58352_sb;
wire TIMEBOOST_net_4251;
wire g58353_db;
wire g58353_sb;
wire TIMEBOOST_net_4252;
wire g58354_db;
wire g58354_sb;
wire TIMEBOOST_net_4253;
wire TIMEBOOST_net_603;
wire g58355_sb;
wire TIMEBOOST_net_4254;
wire g58356_db;
wire g58356_sb;
wire TIMEBOOST_net_4255;
wire g58357_db;
wire g58357_sb;
wire TIMEBOOST_net_4256;
wire g58358_db;
wire g58358_sb;
wire TIMEBOOST_net_4257;
wire g58359_db;
wire g58359_sb;
wire TIMEBOOST_net_4258;
wire TIMEBOOST_net_604;
wire g58360_sb;
wire TIMEBOOST_net_4259;
wire g58361_db;
wire g58361_sb;
wire TIMEBOOST_net_4260;
wire g58362_db;
wire g58362_sb;
wire TIMEBOOST_net_10403;
wire g58363_db;
wire g58363_sb;
wire TIMEBOOST_net_4262;
wire g58364_db;
wire g58364_sb;
wire TIMEBOOST_net_9983;
wire TIMEBOOST_net_14528;
wire g58365_sb;
wire TIMEBOOST_net_11334;
wire TIMEBOOST_net_14134;
wire g58366_sb;
wire g58367_da;
wire TIMEBOOST_net_4614;
wire TIMEBOOST_net_4263;
wire TIMEBOOST_net_605;
wire g58368_sb;
wire TIMEBOOST_net_4264;
wire g58369_db;
wire g58369_sb;
wire TIMEBOOST_net_4265;
wire g58370_db;
wire g58370_sb;
wire TIMEBOOST_net_4266;
wire g58371_db;
wire g58371_sb;
wire TIMEBOOST_net_4267;
wire g58372_db;
wire g58372_sb;
wire TIMEBOOST_net_10744;
wire TIMEBOOST_net_14136;
wire g58373_sb;
wire TIMEBOOST_net_4268;
wire g58374_db;
wire g58374_sb;
wire TIMEBOOST_net_12257;
wire TIMEBOOST_net_4380;
wire g58375_sb;
wire TIMEBOOST_net_3675;
wire TIMEBOOST_net_606;
wire g58376_sb;
wire TIMEBOOST_net_3676;
wire TIMEBOOST_net_607;
wire g58377_sb;
wire TIMEBOOST_net_9932;
wire g58378_db;
wire g58378_sb;
wire g58379_da;
wire g58379_db;
wire g58379_sb;
wire TIMEBOOST_net_4510;
wire TIMEBOOST_net_14445;
wire g58380_sb;
wire TIMEBOOST_net_4511;
wire TIMEBOOST_net_14194;
wire g58381_sb;
wire g58382_da;
wire g58382_db;
wire g58382_sb;
wire TIMEBOOST_net_9985;
wire g58383_db;
wire g58383_sb;
wire TIMEBOOST_net_9984;
wire TIMEBOOST_net_608;
wire g58384_sb;
wire TIMEBOOST_net_12914;
wire TIMEBOOST_net_609;
wire g58385_sb;
wire TIMEBOOST_net_4512;
wire TIMEBOOST_net_14073;
wire g58386_sb;
wire TIMEBOOST_net_4513;
wire g58387_db;
wire g58387_sb;
wire TIMEBOOST_net_12842;
wire g58388_db;
wire g58388_sb;
wire g58389_da;
wire g58389_db;
wire g58389_sb;
wire TIMEBOOST_net_3682;
wire TIMEBOOST_net_610;
wire g58390_sb;
wire TIMEBOOST_net_12912;
wire g58391_db;
wire g58391_sb;
wire TIMEBOOST_net_3684;
wire g58392_db;
wire g58392_sb;
wire g58393_da;
wire g58393_db;
wire g58393_sb;
wire TIMEBOOST_net_10670;
wire TIMEBOOST_net_13942;
wire g58394_sb;
wire TIMEBOOST_net_9945;
wire TIMEBOOST_net_10481;
wire g58395_sb;
wire TIMEBOOST_net_3685;
wire g58396_db;
wire g58396_sb;
wire g58397_da;
wire g58397_db;
wire g58397_sb;
wire TIMEBOOST_net_10671;
wire g58398_db;
wire g58398_sb;
wire g58399_da;
wire g58399_db;
wire g58399_sb;
wire TIMEBOOST_net_4516;
wire TIMEBOOST_net_13978;
wire g58400_sb;
wire TIMEBOOST_net_14576;
wire TIMEBOOST_net_13122;
wire g58401_sb;
wire TIMEBOOST_net_13035;
wire TIMEBOOST_net_13506;
wire g58402_sb;
wire TIMEBOOST_net_13326;
wire TIMEBOOST_net_611;
wire g58403_sb;
wire g58404_da;
wire g58404_db;
wire g58404_sb;
wire TIMEBOOST_net_4517;
wire TIMEBOOST_net_14317;
wire g58405_sb;
wire TIMEBOOST_net_3688;
wire g58406_db;
wire g58406_sb;
wire TIMEBOOST_net_4518;
wire TIMEBOOST_net_14303;
wire g58407_sb;
wire TIMEBOOST_net_15053;
wire TIMEBOOST_net_10482;
wire g58408_sb;
wire TIMEBOOST_net_15054;
wire g58409_db;
wire g58409_sb;
wire TIMEBOOST_net_11030;
wire g58410_db;
wire g58410_sb;
wire g58411_da;
wire g58411_db;
wire g58411_sb;
wire TIMEBOOST_net_11031;
wire g58412_db;
wire g58412_sb;
wire TIMEBOOST_net_11032;
wire g58413_db;
wire g58413_sb;
wire TIMEBOOST_net_9810;
wire g58414_db;
wire g58414_sb;
wire TIMEBOOST_net_11035;
wire g58415_db;
wire g58415_sb;
wire g58416_da;
wire g58416_db;
wire g58416_sb;
wire TIMEBOOST_net_9582;
wire g58417_db;
wire g58417_sb;
wire TIMEBOOST_net_3689;
wire g58418_db;
wire g58418_sb;
wire TIMEBOOST_net_13343;
wire g58419_db;
wire g58419_sb;
wire TIMEBOOST_net_13342;
wire TIMEBOOST_net_612;
wire g58420_sb;
wire TIMEBOOST_net_9993;
wire TIMEBOOST_net_613;
wire g58421_sb;
wire TIMEBOOST_net_13572;
wire TIMEBOOST_net_9299;
wire g58422_sb;
wire g58423_da;
wire g58423_db;
wire g58423_sb;
wire g58424_da;
wire TIMEBOOST_net_10483;
wire g58424_sb;
wire TIMEBOOST_net_3694;
wire g58425_db;
wire g58425_sb;
wire TIMEBOOST_net_3695;
wire TIMEBOOST_net_614;
wire g58426_sb;
wire TIMEBOOST_net_13222;
wire TIMEBOOST_net_10740;
wire g58427_sb;
wire g58428_da;
wire g58428_db;
wire g58428_sb;
wire TIMEBOOST_net_10004;
wire g58429_db;
wire g58429_sb;
wire TIMEBOOST_net_3698;
wire g58430_db;
wire g58430_sb;
wire TIMEBOOST_net_14091;
wire g58431_db;
wire g58431_sb;
wire TIMEBOOST_net_12910;
wire g58432_db;
wire g58432_sb;
wire g58433_da;
wire g58433_db;
wire g58433_sb;
wire TIMEBOOST_net_3701;
wire TIMEBOOST_net_14541;
wire g58434_sb;
wire g58435_da;
wire g58435_db;
wire g58435_sb;
wire g58436_da;
wire g58436_db;
wire g58436_sb;
wire g58437_da;
wire g58437_db;
wire g58437_sb;
wire TIMEBOOST_net_3702;
wire TIMEBOOST_net_13979;
wire g58438_sb;
wire TIMEBOOST_net_14265;
wire g58439_db;
wire g58439_sb;
wire TIMEBOOST_net_14565;
wire TIMEBOOST_net_10142;
wire g58440_sb;
wire TIMEBOOST_net_3704;
wire TIMEBOOST_net_617;
wire g58441_sb;
wire TIMEBOOST_net_13327;
wire g58442_db;
wire g58442_sb;
wire g58443_da;
wire g58443_db;
wire g58443_sb;
wire TIMEBOOST_net_3706;
wire g58444_db;
wire g58444_sb;
wire g58445_da;
wire g58445_db;
wire g58445_sb;
wire TIMEBOOST_net_11037;
wire TIMEBOOST_net_14414;
wire g58446_sb;
wire g58447_da;
wire g58447_db;
wire g58447_sb;
wire TIMEBOOST_net_4269;
wire g58448_db;
wire g58448_sb;
wire g58449_da;
wire g58449_db;
wire g58449_sb;
wire TIMEBOOST_net_12862;
wire TIMEBOOST_net_618;
wire g58450_sb;
wire TIMEBOOST_net_3708;
wire g58451_db;
wire g58451_sb;
wire TIMEBOOST_net_3709;
wire g58452_db;
wire g58452_sb;
wire TIMEBOOST_net_3710;
wire g58453_db;
wire g58453_sb;
wire TIMEBOOST_net_3711;
wire g58454_db;
wire g58454_sb;
wire TIMEBOOST_net_12177;
wire TIMEBOOST_net_14080;
wire g58455_sb;
wire TIMEBOOST_net_12207;
wire TIMEBOOST_net_14451;
wire g58456_sb;
wire TIMEBOOST_net_6570;
wire TIMEBOOST_net_1820;
wire g58457_sb;
wire TIMEBOOST_net_12215;
wire TIMEBOOST_net_12339;
wire g58458_sb;
wire TIMEBOOST_net_12198;
wire TIMEBOOST_net_1822;
wire g58459_sb;
wire TIMEBOOST_net_12222;
wire TIMEBOOST_net_1823;
wire g58460_sb;
wire TIMEBOOST_net_12221;
wire TIMEBOOST_net_1824;
wire g58461_sb;
wire TIMEBOOST_net_12223;
wire TIMEBOOST_net_1825;
wire g58462_sb;
wire TIMEBOOST_net_6576;
wire TIMEBOOST_net_1826;
wire g58463_sb;
wire TIMEBOOST_net_6577;
wire TIMEBOOST_net_14765;
wire g58464_sb;
wire TIMEBOOST_net_6578;
wire TIMEBOOST_net_1828;
wire g58465_sb;
wire TIMEBOOST_net_6579;
wire TIMEBOOST_net_12278;
wire g58466_sb;
wire TIMEBOOST_net_6580;
wire TIMEBOOST_net_12790;
wire g58467_sb;
wire TIMEBOOST_net_6581;
wire TIMEBOOST_net_1831;
wire g58468_sb;
wire TIMEBOOST_net_1832;
wire g58469_sb;
wire TIMEBOOST_net_9354;
wire g58470_sb;
wire TIMEBOOST_net_1834;
wire g58471_sb;
wire TIMEBOOST_net_1835;
wire g58472_sb;
wire TIMEBOOST_net_1836;
wire g58473_sb;
wire TIMEBOOST_net_1837;
wire g58474_sb;
wire TIMEBOOST_net_12744;
wire g58475_sb;
wire TIMEBOOST_net_1839;
wire g58476_sb;
wire TIMEBOOST_net_6571;
wire TIMEBOOST_net_1840;
wire g58477_sb;
wire TIMEBOOST_net_12275;
wire g58478_sb;
wire TIMEBOOST_net_1842;
wire g58479_sb;
wire TIMEBOOST_net_1843;
wire g58480_sb;
wire n_12023;
wire TIMEBOOST_net_10507;
wire g58481_sb;
wire TIMEBOOST_net_1845;
wire g58482_sb;
wire n_12328;
wire TIMEBOOST_net_10508;
wire g58483_sb;
wire n_12312;
wire TIMEBOOST_net_14578;
wire g58484_sb;
wire TIMEBOOST_net_1848;
wire g58485_sb;
wire TIMEBOOST_net_14545;
wire g58486_sb;
wire TIMEBOOST_net_4270;
wire TIMEBOOST_net_11892;
wire g58487_sb;
wire TIMEBOOST_net_13221;
wire TIMEBOOST_net_620;
wire g58488_sb;
wire TIMEBOOST_net_13328;
wire TIMEBOOST_net_13273;
wire g58489_sb;
wire g58490_p;
wire g58569_p;
wire TIMEBOOST_net_6423;
wire TIMEBOOST_net_13311;
wire g58574_sb;
wire TIMEBOOST_net_14307;
wire TIMEBOOST_net_11765;
wire g58576_sb;
wire g58582_p;
wire TIMEBOOST_net_13219;
wire TIMEBOOST_net_13253;
wire g58586_sb;
wire TIMEBOOST_net_13026;
wire g58587_sb;
wire TIMEBOOST_net_6562;
wire TIMEBOOST_net_13338;
wire g58588_sb;
wire TIMEBOOST_net_6424;
wire TIMEBOOST_net_13331;
wire g58589_sb;
wire TIMEBOOST_net_6425;
wire TIMEBOOST_net_13333;
wire g58590_sb;
wire TIMEBOOST_net_6426;
wire TIMEBOOST_net_13316;
wire g58591_sb;
wire TIMEBOOST_net_13217;
wire TIMEBOOST_net_13257;
wire g58592_sb;
wire TIMEBOOST_net_6427;
wire TIMEBOOST_net_13308;
wire g58593_sb;
wire TIMEBOOST_net_13027;
wire TIMEBOOST_net_13255;
wire g58594_sb;
wire TIMEBOOST_net_13037;
wire g58595_sb;
wire TIMEBOOST_net_6564;
wire TIMEBOOST_net_13025;
wire g58596_sb;
wire TIMEBOOST_net_6428;
wire TIMEBOOST_net_13309;
wire g58597_sb;
wire g58598_da;
wire g58598_db;
wire g58598_sb;
wire g58599_p;
wire TIMEBOOST_net_13951;
wire g58600_db;
wire g58600_sb;
wire TIMEBOOST_net_12825;
wire TIMEBOOST_net_12709;
wire g58601_sb;
wire TIMEBOOST_net_466;
wire TIMEBOOST_net_4489;
wire g58605_sb;
wire TIMEBOOST_net_6565;
wire TIMEBOOST_net_13038;
wire g58606_sb;
wire TIMEBOOST_net_14284;
wire TIMEBOOST_net_13256;
wire g58607_sb;
wire TIMEBOOST_net_6429;
wire TIMEBOOST_net_14509;
wire g58608_sb;
wire TIMEBOOST_net_6566;
wire TIMEBOOST_net_13012;
wire g58609_sb;
wire TIMEBOOST_net_14285;
wire g58610_sb;
wire TIMEBOOST_net_3988;
wire TIMEBOOST_net_14033;
wire g58611_sb;
wire TIMEBOOST_net_14302;
wire TIMEBOOST_net_11493;
wire g58616_sb;
wire TIMEBOOST_net_13110;
wire TIMEBOOST_net_11536;
wire g58617_sb;
wire TIMEBOOST_net_13127;
wire TIMEBOOST_net_11734;
wire g58618_sb;
wire TIMEBOOST_net_13140;
wire TIMEBOOST_net_11735;
wire g58619_sb;
wire TIMEBOOST_net_13141;
wire TIMEBOOST_net_11736;
wire g58620_sb;
wire TIMEBOOST_net_3926;
wire TIMEBOOST_net_11783;
wire g58621_sb;
wire g58622_da;
wire g58622_db;
wire g58622_sb;
wire TIMEBOOST_net_13960;
wire g58630_db;
wire g58630_sb;
wire TIMEBOOST_net_14093;
wire g58631_db;
wire g58631_sb;
wire TIMEBOOST_net_14368;
wire g58632_db;
wire g58632_sb;
wire TIMEBOOST_net_2007;
wire g58633_db;
wire g58633_sb;
wire TIMEBOOST_net_14568;
wire g58634_db;
wire g58634_sb;
wire TIMEBOOST_net_9357;
wire g58635_db;
wire g58635_sb;
wire TIMEBOOST_net_10453;
wire TIMEBOOST_net_14373;
wire g58636_sb;
wire TIMEBOOST_net_12826;
wire TIMEBOOST_net_12793;
wire g58640_sb;
wire TIMEBOOST_net_14024;
wire TIMEBOOST_net_12076;
wire g58652_sb;
wire TIMEBOOST_net_14278;
wire TIMEBOOST_net_12077;
wire g58653_sb;
wire TIMEBOOST_net_14002;
wire TIMEBOOST_net_12078;
wire g58654_sb;
wire TIMEBOOST_net_14468;
wire TIMEBOOST_net_12079;
wire g58655_sb;
wire g58656_p;
wire g58692_p;
wire g58695_p;
wire g58742_p;
wire g58744_p;
wire g58759_p;
wire g58760_p;
wire g58761_p;
wire g58763_p;
wire g58764_p;
wire TIMEBOOST_net_106;
wire g58767_db;
wire g58767_sb;
wire TIMEBOOST_net_3226;
wire TIMEBOOST_net_133;
wire g58768_sb;
wire TIMEBOOST_net_12316;
wire TIMEBOOST_net_134;
wire g58769_sb;
wire TIMEBOOST_net_31;
wire g58770_db;
wire g58770_sb;
wire TIMEBOOST_net_107;
wire TIMEBOOST_net_12730;
wire g58771_sb;
wire TIMEBOOST_net_12636;
wire TIMEBOOST_net_14667;
wire g58772_sb;
wire TIMEBOOST_net_109;
wire TIMEBOOST_net_12731;
wire g58773_sb;
wire TIMEBOOST_net_32;
wire g58774_db;
wire g58774_sb;
wire TIMEBOOST_net_33;
wire g58775_db;
wire g58775_sb;
wire TIMEBOOST_net_3227;
wire TIMEBOOST_net_135;
wire g58776_sb;
wire TIMEBOOST_net_3228;
wire TIMEBOOST_net_136;
wire g58777_sb;
wire TIMEBOOST_net_12315;
wire TIMEBOOST_net_137;
wire g58778_sb;
wire TIMEBOOST_net_3732;
wire g58779_db;
wire g58779_sb;
wire TIMEBOOST_net_29;
wire g58780_db;
wire TIMEBOOST_net_14758;
wire TIMEBOOST_net_80;
wire TIMEBOOST_net_12318;
wire TIMEBOOST_net_138;
wire g58782_sb;
wire TIMEBOOST_net_34;
wire TIMEBOOST_net_14985;
wire g58783_sb;
wire TIMEBOOST_net_35;
wire TIMEBOOST_net_14960;
wire TIMEBOOST_net_111;
wire TIMEBOOST_net_15007;
wire g58785_sb;
wire TIMEBOOST_net_112;
wire g58786_db;
wire g58786_sb;
wire TIMEBOOST_net_12516;
wire TIMEBOOST_net_139;
wire g58787_sb;
wire TIMEBOOST_net_113;
wire TIMEBOOST_net_12795;
wire g58788_sb;
wire TIMEBOOST_net_14884;
wire TIMEBOOST_net_12752;
wire g58789_sb;
wire TIMEBOOST_net_114;
wire g58790_db;
wire g58790_sb;
wire TIMEBOOST_net_14846;
wire g58791_db;
wire g58791_sb;
wire TIMEBOOST_net_12313;
wire TIMEBOOST_net_140;
wire g58792_sb;
wire TIMEBOOST_net_36;
wire g58793_db;
wire g58793_sb;
wire TIMEBOOST_net_37;
wire g58794_db;
wire g58794_sb;
wire TIMEBOOST_net_116;
wire g58795_db;
wire g58795_sb;
wire TIMEBOOST_net_38;
wire g58796_db;
wire TIMEBOOST_net_117;
wire g58797_db;
wire g58797_sb;
wire TIMEBOOST_net_118;
wire TIMEBOOST_net_12796;
wire g58798_sb;
wire TIMEBOOST_net_10460;
wire TIMEBOOST_net_12366;
wire g58799_sb;
wire TIMEBOOST_net_14920;
wire g58800_sb;
wire TIMEBOOST_net_12956;
wire g58801_sb;
wire TIMEBOOST_net_12955;
wire g58802_sb;
wire TIMEBOOST_net_12954;
wire g58803_sb;
wire TIMEBOOST_net_14596;
wire TIMEBOOST_net_12953;
wire g58804_sb;
wire TIMEBOOST_net_14597;
wire TIMEBOOST_net_12940;
wire g58805_sb;
wire TIMEBOOST_net_15260;
wire TIMEBOOST_net_12941;
wire g58806_sb;
wire TIMEBOOST_net_15258;
wire TIMEBOOST_net_12942;
wire g58807_sb;
wire TIMEBOOST_net_15237;
wire TIMEBOOST_net_12943;
wire g58808_sb;
wire TIMEBOOST_net_15238;
wire TIMEBOOST_net_12944;
wire g58809_sb;
wire TIMEBOOST_net_15226;
wire TIMEBOOST_net_12935;
wire g58810_sb;
wire TIMEBOOST_net_15240;
wire TIMEBOOST_net_12938;
wire g58811_sb;
wire TIMEBOOST_net_15241;
wire TIMEBOOST_net_12945;
wire g58812_sb;
wire TIMEBOOST_net_15242;
wire TIMEBOOST_net_12933;
wire g58813_sb;
wire TIMEBOOST_net_15243;
wire TIMEBOOST_net_13258;
wire g58814_sb;
wire TIMEBOOST_net_15246;
wire TIMEBOOST_net_13259;
wire g58815_sb;
wire TIMEBOOST_net_15247;
wire TIMEBOOST_net_13233;
wire g58816_sb;
wire TIMEBOOST_net_15248;
wire TIMEBOOST_net_13047;
wire g58817_sb;
wire TIMEBOOST_net_15249;
wire TIMEBOOST_net_13261;
wire g58818_sb;
wire TIMEBOOST_net_15250;
wire TIMEBOOST_net_13006;
wire g58819_sb;
wire TIMEBOOST_net_15251;
wire TIMEBOOST_net_13111;
wire g58820_sb;
wire TIMEBOOST_net_15235;
wire TIMEBOOST_net_13260;
wire g58821_sb;
wire TIMEBOOST_net_15225;
wire TIMEBOOST_net_13232;
wire g58822_sb;
wire TIMEBOOST_net_15232;
wire TIMEBOOST_net_13242;
wire g58823_sb;
wire TIMEBOOST_net_15233;
wire TIMEBOOST_net_12978;
wire g58824_sb;
wire TIMEBOOST_net_15234;
wire TIMEBOOST_net_13235;
wire g58825_sb;
wire TIMEBOOST_net_15239;
wire TIMEBOOST_net_13228;
wire g58826_sb;
wire TIMEBOOST_net_15253;
wire TIMEBOOST_net_13238;
wire g58827_sb;
wire TIMEBOOST_net_15236;
wire TIMEBOOST_net_13247;
wire g58828_sb;
wire TIMEBOOST_net_15231;
wire TIMEBOOST_net_13059;
wire g58829_sb;
wire TIMEBOOST_net_15254;
wire TIMEBOOST_net_13028;
wire g58830_sb;
wire TIMEBOOST_net_15255;
wire TIMEBOOST_net_13016;
wire g58831_sb;
wire TIMEBOOST_net_15230;
wire TIMEBOOST_net_13042;
wire g58832_sb;
wire TIMEBOOST_net_15244;
wire TIMEBOOST_net_1554;
wire g58833_sb;
wire TIMEBOOST_net_15228;
wire TIMEBOOST_net_1539;
wire g58834_sb;
wire TIMEBOOST_net_15229;
wire TIMEBOOST_net_13250;
wire g58835_sb;
wire TIMEBOOST_net_15222;
wire TIMEBOOST_net_13227;
wire g58836_sb;
wire TIMEBOOST_net_6541;
wire TIMEBOOST_net_9347;
wire g58837_sb;
wire TIMEBOOST_net_6540;
wire TIMEBOOST_net_10595;
wire g58838_sb;
wire TIMEBOOST_net_6539;
wire TIMEBOOST_net_14571;
wire g58839_sb;
wire TIMEBOOST_net_10597;
wire g58840_sb;
wire TIMEBOOST_net_6537;
wire TIMEBOOST_net_10599;
wire g58841_sb;
wire TIMEBOOST_net_14446;
wire TIMEBOOST_net_6567;
wire g58842_sb;
wire TIMEBOOST_net_10109;
wire TIMEBOOST_net_14443;
wire g58843_sb;
wire TIMEBOOST_net_14674;
wire TIMEBOOST_net_10858;
wire g59082_sb;
wire g59086_p;
wire TIMEBOOST_net_14836;
wire TIMEBOOST_net_10859;
wire g59089_sb;
wire TIMEBOOST_net_14798;
wire TIMEBOOST_net_5430;
wire g59090_sb;
wire TIMEBOOST_net_14776;
wire TIMEBOOST_net_13612;
wire TIMEBOOST_net_738;
wire TIMEBOOST_net_10709;
wire g59092_sb;
wire TIMEBOOST_net_10598;
wire TIMEBOOST_net_14523;
wire g59093_sb;
wire g59095_p;
wire TIMEBOOST_net_10110;
wire TIMEBOOST_net_14058;
wire g59096_sb;
wire TIMEBOOST_net_11012;
wire TIMEBOOST_net_10596;
wire g59097_sb;
wire TIMEBOOST_net_1662;
wire TIMEBOOST_net_5431;
wire g59098_sb;
wire TIMEBOOST_net_12254;
wire TIMEBOOST_net_5432;
wire g59109_sb;
wire TIMEBOOST_net_15044;
wire TIMEBOOST_net_5433;
wire g59110_sb;
wire TIMEBOOST_net_14401;
wire TIMEBOOST_net_5434;
wire g59111_sb;
wire TIMEBOOST_net_14402;
wire TIMEBOOST_net_10179;
wire g59112_sb;
wire TIMEBOOST_net_14403;
wire TIMEBOOST_net_5436;
wire g59113_sb;
wire TIMEBOOST_net_14404;
wire TIMEBOOST_net_5437;
wire TIMEBOOST_net_14405;
wire TIMEBOOST_net_5438;
wire TIMEBOOST_net_14406;
wire TIMEBOOST_net_5439;
wire TIMEBOOST_net_14444;
wire TIMEBOOST_net_5440;
wire TIMEBOOST_net_14574;
wire TIMEBOOST_net_10180;
wire g59118_sb;
wire TIMEBOOST_net_14340;
wire TIMEBOOST_net_5442;
wire TIMEBOOST_net_14341;
wire TIMEBOOST_net_10632;
wire TIMEBOOST_net_467;
wire TIMEBOOST_net_10725;
wire g59121_sb;
wire TIMEBOOST_net_11189;
wire TIMEBOOST_net_904;
wire g59122_sb;
wire TIMEBOOST_net_9362;
wire TIMEBOOST_net_11182;
wire g59123_sb;
wire g59124_p;
wire g59125_p;
wire TIMEBOOST_net_14422;
wire g59126_db;
wire g59126_sb;
wire g59127_p;
wire g59128_p;
wire g59129_p;
wire g59196_p;
wire g59198_p;
wire g59199_p;
wire g59201_p;
wire g59206_p;
wire TIMEBOOST_net_3989;
wire TIMEBOOST_net_12649;
wire g59226_sb;
wire g59227_p;
wire g59228_p;
wire g59229_p;
wire TIMEBOOST_net_10125;
wire TIMEBOOST_net_14921;
wire g59230_sb;
wire TIMEBOOST_net_10126;
wire TIMEBOOST_net_14922;
wire g59231_sb;
wire TIMEBOOST_net_350;
wire TIMEBOOST_net_13190;
wire g59232_p;
wire TIMEBOOST_net_10711;
wire TIMEBOOST_net_10749;
wire g59234_sb;
wire g59239_da;
wire TIMEBOOST_net_11326;
wire g59239_sb;
wire g59240_da;
wire g59240_db;
wire g59240_sb;
wire g59296_p;
wire g59300_p;
wire g59331_p;
wire g59344_p;
wire g59345_p;
wire g59346_p;
wire g59347_p;
wire TIMEBOOST_net_12358;
wire g59350_db;
wire g59350_sb;
wire g59364_p;
wire g59367_p;
wire TIMEBOOST_net_899;
wire g59368_db;
wire g59368_sb;
wire TIMEBOOST_net_900;
wire g59369_db;
wire g59369_sb;
wire TIMEBOOST_net_4565;
wire TIMEBOOST_net_4897;
wire g59370_sb;
wire TIMEBOOST_net_4659;
wire TIMEBOOST_net_4898;
wire g59371_sb;
wire TIMEBOOST_net_10646;
wire TIMEBOOST_net_4899;
wire g59372_sb;
wire TIMEBOOST_net_915;
wire TIMEBOOST_net_4900;
wire g59373_sb;
wire g59374_p;
wire g59377_p;
wire TIMEBOOST_net_4567;
wire TIMEBOOST_net_4901;
wire g59378_sb;
wire TIMEBOOST_net_12566;
wire TIMEBOOST_net_4902;
wire g59379_sb;
wire TIMEBOOST_net_11814;
wire TIMEBOOST_net_4903;
wire g59380_sb;
wire TIMEBOOST_net_4660;
wire g59381_db;
wire g59381_sb;
wire TIMEBOOST_net_9363;
wire TIMEBOOST_net_11840;
wire g59382_sb;
wire TIMEBOOST_net_468;
wire g59383_db;
wire g59383_sb;
wire TIMEBOOST_net_12671;
wire TIMEBOOST_net_10780;
wire g59384_sb;
wire g59385_p;
wire g59386_p;
wire TIMEBOOST_net_13806;
wire TIMEBOOST_net_5444;
wire g59387_sb;
wire g59388_p;
wire g59389_p;
wire g59622_p;
wire g59623_p;
wire g59627_p;
wire g59659_p;
wire g59665_p;
wire g59666_p;
wire g59670_p;
wire g59674_p;
wire g59721_p;
wire g59761_p;
wire TIMEBOOST_net_11791;
wire TIMEBOOST_net_14301;
wire g59763_sb;
wire TIMEBOOST_net_3229;
wire TIMEBOOST_net_12519;
wire TIMEBOOST_net_14365;
wire g59783_p;
wire g59785_p;
wire g59790_p;
wire g59791_p;
wire g59793_p;
wire g59794_p;
wire g59795_p;
wire TIMEBOOST_net_1857;
wire g59796_db;
wire g59796_sb;
wire TIMEBOOST_net_5307;
wire TIMEBOOST_net_1184;
wire g59797_sb;
wire TIMEBOOST_net_10820;
wire TIMEBOOST_net_14287;
wire g59798_sb;
wire g59799_da;
wire TIMEBOOST_net_10993;
wire g59799_sb;
wire TIMEBOOST_net_9364;
wire TIMEBOOST_net_10979;
wire g59800_sb;
wire TIMEBOOST_net_11256;
wire TIMEBOOST_net_14008;
wire g59801_sb;
wire g59802_p;
wire g59803_p;
wire g59804_da;
wire TIMEBOOST_net_11014;
wire g59804_sb;
wire g59805_da;
wire TIMEBOOST_net_11015;
wire g59805_sb;
wire TIMEBOOST_net_13882;
wire TIMEBOOST_net_11019;
wire g59806_sb;
wire g59807_da;
wire TIMEBOOST_net_11022;
wire g59807_sb;
wire TIMEBOOST_net_14668;
wire TIMEBOOST_net_11023;
wire g59808_sb;
wire TIMEBOOST_net_15015;
wire TIMEBOOST_net_11024;
wire g59809_sb;
wire g60298_p;
wire g60304_p;
wire g60307_p;
wire g60310_p;
wire g60319_p;
wire g60321_p;
wire g60330_p;
wire g60339_p;
wire g60345_p;
wire TIMEBOOST_net_3219;
wire TIMEBOOST_net_4090;
wire g60407_sb;
wire TIMEBOOST_net_12242;
wire TIMEBOOST_net_10469;
wire TIMEBOOST_net_10703;
wire TIMEBOOST_net_14342;
wire g60409_sb;
wire g60414_p;
wire g60415_p;
wire g60557_p;
wire g60591_p;
wire TIMEBOOST_net_3990;
wire TIMEBOOST_net_14167;
wire g60603_sb;
wire TIMEBOOST_net_14709;
wire TIMEBOOST_net_13883;
wire g60604_sb;
wire TIMEBOOST_net_14716;
wire TIMEBOOST_net_13880;
wire g60605_sb;
wire TIMEBOOST_net_14717;
wire TIMEBOOST_net_13871;
wire g60606_sb;
wire TIMEBOOST_net_14719;
wire TIMEBOOST_net_13889;
wire g60607_sb;
wire TIMEBOOST_net_14675;
wire TIMEBOOST_net_13873;
wire g60608_sb;
wire TIMEBOOST_net_14820;
wire TIMEBOOST_net_13890;
wire g60609_sb;
wire TIMEBOOST_net_14805;
wire TIMEBOOST_net_13888;
wire g60610_sb;
wire TIMEBOOST_net_14817;
wire TIMEBOOST_net_13862;
wire g60611_sb;
wire TIMEBOOST_net_14806;
wire TIMEBOOST_net_13879;
wire g60612_sb;
wire TIMEBOOST_net_14725;
wire TIMEBOOST_net_13887;
wire g60613_sb;
wire TIMEBOOST_net_14857;
wire TIMEBOOST_net_13885;
wire g60614_sb;
wire TIMEBOOST_net_14858;
wire TIMEBOOST_net_13886;
wire g60615_sb;
wire TIMEBOOST_net_15022;
wire TIMEBOOST_net_13891;
wire g60616_sb;
wire TIMEBOOST_net_14681;
wire TIMEBOOST_net_13863;
wire g60617_sb;
wire TIMEBOOST_net_14682;
wire TIMEBOOST_net_13893;
wire g60618_sb;
wire TIMEBOOST_net_14799;
wire TIMEBOOST_net_13877;
wire g60619_sb;
wire TIMEBOOST_net_14390;
wire TIMEBOOST_net_13870;
wire g60620_sb;
wire TIMEBOOST_net_14391;
wire TIMEBOOST_net_13878;
wire g60621_sb;
wire TIMEBOOST_net_14335;
wire TIMEBOOST_net_11190;
wire g60622_sb;
wire TIMEBOOST_net_14513;
wire TIMEBOOST_net_13874;
wire g60623_sb;
wire TIMEBOOST_net_14320;
wire TIMEBOOST_net_13872;
wire g60624_sb;
wire TIMEBOOST_net_14383;
wire TIMEBOOST_net_11178;
wire g60625_sb;
wire TIMEBOOST_net_14481;
wire TIMEBOOST_net_13876;
wire g60626_sb;
wire TIMEBOOST_net_14535;
wire TIMEBOOST_net_11179;
wire g60627_sb;
wire TIMEBOOST_net_14384;
wire TIMEBOOST_net_13875;
wire g60628_sb;
wire TIMEBOOST_net_14387;
wire TIMEBOOST_net_13892;
wire g60629_sb;
wire TIMEBOOST_net_14459;
wire TIMEBOOST_net_13861;
wire g60630_sb;
wire TIMEBOOST_net_14482;
wire TIMEBOOST_net_13857;
wire g60631_sb;
wire TIMEBOOST_net_1524;
wire TIMEBOOST_net_13858;
wire g60632_sb;
wire TIMEBOOST_net_14462;
wire TIMEBOOST_net_14518;
wire g60633_sb;
wire TIMEBOOST_net_14829;
wire g52444_db;
wire g60634_sb;
wire TIMEBOOST_net_1484;
wire TIMEBOOST_net_13841;
wire g60635_sb;
wire TIMEBOOST_net_14695;
wire TIMEBOOST_net_13836;
wire g60636_sb;
wire TIMEBOOST_net_14813;
wire TIMEBOOST_net_11191;
wire g60637_sb;
wire TIMEBOOST_net_14827;
wire TIMEBOOST_net_5288;
wire g60638_sb;
wire TIMEBOOST_net_14666;
wire TIMEBOOST_net_10692;
wire g60639_sb;
wire TIMEBOOST_net_14848;
wire TIMEBOOST_net_10461;
wire g60640_sb;
wire TIMEBOOST_net_14888;
wire TIMEBOOST_net_13842;
wire g60641_sb;
wire TIMEBOOST_net_14832;
wire TIMEBOOST_net_13835;
wire g60642_sb;
wire TIMEBOOST_net_1492;
wire TIMEBOOST_net_13843;
wire g60643_sb;
wire TIMEBOOST_net_14362;
wire TIMEBOOST_net_4821;
wire g60644_sb;
wire TIMEBOOST_net_14363;
wire TIMEBOOST_net_4820;
wire g60645_sb;
wire TIMEBOOST_net_9912;
wire TIMEBOOST_net_5291;
wire g60646_sb;
wire TIMEBOOST_net_15083;
wire TIMEBOOST_net_4819;
wire g60647_sb;
wire TIMEBOOST_net_14524;
wire TIMEBOOST_net_13848;
wire g60648_sb;
wire TIMEBOOST_net_14483;
wire TIMEBOOST_net_13834;
wire g60649_sb;
wire TIMEBOOST_net_14686;
wire TIMEBOOST_net_13833;
wire g60650_sb;
wire TIMEBOOST_net_14687;
wire TIMEBOOST_net_524;
wire g60651_sb;
wire TIMEBOOST_net_14685;
wire n_13452;
wire g60652_sb;
wire TIMEBOOST_net_14812;
wire TIMEBOOST_net_13832;
wire g60653_sb;
wire TIMEBOOST_net_1503;
wire TIMEBOOST_net_13830;
wire g60654_sb;
wire TIMEBOOST_net_14847;
wire TIMEBOOST_net_13827;
wire g60655_sb;
wire TIMEBOOST_net_14190;
wire TIMEBOOST_net_13826;
wire g60656_sb;
wire TIMEBOOST_net_9995;
wire TIMEBOOST_net_13825;
wire g60657_sb;
wire TIMEBOOST_net_14193;
wire TIMEBOOST_net_10124;
wire g60658_sb;
wire TIMEBOOST_net_14394;
wire TIMEBOOST_net_13810;
wire g60659_sb;
wire TIMEBOOST_net_1509;
wire TIMEBOOST_net_13811;
wire g60660_sb;
wire TIMEBOOST_net_14395;
wire TIMEBOOST_net_13815;
wire g60661_sb;
wire TIMEBOOST_net_14380;
wire TIMEBOOST_net_13822;
wire g60662_sb;
wire TIMEBOOST_net_1512;
wire TIMEBOOST_net_13814;
wire g60663_sb;
wire TIMEBOOST_net_14381;
wire TIMEBOOST_net_5293;
wire g60664_sb;
wire TIMEBOOST_net_14385;
wire TIMEBOOST_net_13817;
wire g60665_sb;
wire TIMEBOOST_net_14386;
wire TIMEBOOST_net_10129;
wire g60666_sb;
wire TIMEBOOST_net_13220;
wire TIMEBOOST_net_13809;
wire g60667_sb;
wire TIMEBOOST_net_9992;
wire TIMEBOOST_net_13808;
wire g60668_sb;
wire TIMEBOOST_net_1518;
wire TIMEBOOST_net_10130;
wire g60669_sb;
wire TIMEBOOST_net_14967;
wire TIMEBOOST_net_13807;
wire g60670_sb;
wire TIMEBOOST_net_10304;
wire TIMEBOOST_net_13304;
wire g60671_sb;
wire TIMEBOOST_net_3992;
wire TIMEBOOST_net_905;
wire g60672_sb;
wire TIMEBOOST_net_1520;
wire TIMEBOOST_net_13816;
wire g60673_sb;
wire TIMEBOOST_net_12937;
wire TIMEBOOST_net_10475;
wire g60674_sb;
wire TIMEBOOST_net_4700;
wire g60675_db;
wire g60675_sb;
wire g60676_da;
wire g60676_db;
wire g60676_sb;
wire g60677_da;
wire g60677_db;
wire g60677_sb;
wire g60678_da;
wire g60678_db;
wire g60678_sb;
wire g60679_da;
wire TIMEBOOST_net_10956;
wire g60679_sb;
wire TIMEBOOST_net_10782;
wire TIMEBOOST_net_14923;
wire g60681_sb;
wire g60682_da;
wire TIMEBOOST_net_11565;
wire g60682_sb;
wire g60686_da;
wire g60686_db;
wire g60686_sb;
wire TIMEBOOST_net_10546;
wire g60687_db;
wire g60687_sb;
wire TIMEBOOST_net_166;
wire TIMEBOOST_net_12676;
wire g60688_sb;
wire TIMEBOOST_net_154;
wire TIMEBOOST_net_3001;
wire g60689_sb;
wire TIMEBOOST_net_3994;
wire TIMEBOOST_net_9449;
wire g60690_sb;
wire TIMEBOOST_net_13821;
wire TIMEBOOST_net_11360;
wire g60691_sb;
wire TIMEBOOST_net_12648;
wire g60692_db;
wire g60692_sb;
wire g60693_p;
wire g60694_p;
wire g60695_p;
wire g60696_p;
wire TIMEBOOST_net_86;
wire g61569_p;
wire g61570_p;
wire g61572_p;
wire g61575_p;
wire g61581_p;
wire g61582_p;
wire g61597_p;
wire g61606_p;
wire g61617_p;
wire TIMEBOOST_net_172;
wire g61618_BP;
wire g61618_p;
wire g61622_p;
wire g61636_p;
wire g61637_p;
wire g61654_p;
wire TIMEBOOST_net_14868;
wire TIMEBOOST_net_10170;
wire g61676_sb;
wire g61689_p;
wire g61693_p;
wire TIMEBOOST_net_10799;
wire g61697_db;
wire g61697_sb;
wire TIMEBOOST_net_10800;
wire g61698_db;
wire g61698_sb;
wire TIMEBOOST_net_9388;
wire TIMEBOOST_net_10539;
wire g61699_sb;
wire TIMEBOOST_net_10638;
wire TIMEBOOST_net_11143;
wire g61700_sb;
wire TIMEBOOST_net_12632;
wire TIMEBOOST_net_10131;
wire g61701_sb;
wire TIMEBOOST_net_10212;
wire TIMEBOOST_net_12472;
wire g61702_sb;
wire TIMEBOOST_net_10213;
wire TIMEBOOST_net_13533;
wire g61703_sb;
wire TIMEBOOST_net_13708;
wire TIMEBOOST_net_277;
wire g61704_sb;
wire TIMEBOOST_net_9917;
wire g61705_db;
wire g61705_sb;
wire TIMEBOOST_net_4585;
wire TIMEBOOST_net_278;
wire g61706_sb;
wire g61707_db;
wire g61707_sb;
wire TIMEBOOST_net_3873;
wire TIMEBOOST_net_13532;
wire g61708_sb;
wire TIMEBOOST_net_10236;
wire TIMEBOOST_net_12776;
wire g61709_sb;
wire TIMEBOOST_net_10237;
wire TIMEBOOST_net_12775;
wire g61710_sb;
wire TIMEBOOST_net_12582;
wire TIMEBOOST_net_10147;
wire g61711_sb;
wire TIMEBOOST_net_12363;
wire TIMEBOOST_net_13199;
wire g61712_sb;
wire TIMEBOOST_net_3517;
wire g61713_db;
wire TIMEBOOST_net_5118;
wire TIMEBOOST_net_699;
wire g61714_sb;
wire TIMEBOOST_net_10238;
wire TIMEBOOST_net_13531;
wire g61715_sb;
wire TIMEBOOST_net_12711;
wire TIMEBOOST_net_10132;
wire g61716_sb;
wire TIMEBOOST_net_3877;
wire TIMEBOOST_net_13529;
wire g61717_sb;
wire TIMEBOOST_net_4586;
wire TIMEBOOST_net_279;
wire g61718_sb;
wire TIMEBOOST_net_12370;
wire g61719_sb;
wire TIMEBOOST_net_12322;
wire TIMEBOOST_net_13200;
wire g61720_sb;
wire TIMEBOOST_net_12314;
wire TIMEBOOST_net_13201;
wire g61721_sb;
wire TIMEBOOST_net_4587;
wire TIMEBOOST_net_280;
wire g61722_sb;
wire TIMEBOOST_net_370;
wire g61723_sb;
wire TIMEBOOST_net_12310;
wire TIMEBOOST_net_13334;
wire g61724_sb;
wire TIMEBOOST_net_10867;
wire g65076_db;
wire g61725_sb;
wire TIMEBOOST_net_10239;
wire TIMEBOOST_net_12514;
wire g61726_sb;
wire TIMEBOOST_net_3189;
wire TIMEBOOST_net_10112;
wire g61727_sb;
wire TIMEBOOST_net_12305;
wire TIMEBOOST_net_10113;
wire g61728_sb;
wire TIMEBOOST_net_12319;
wire TIMEBOOST_net_10114;
wire g61729_sb;
wire TIMEBOOST_net_375;
wire TIMEBOOST_net_10115;
wire g61730_sb;
wire TIMEBOOST_net_12293;
wire TIMEBOOST_net_10116;
wire g61731_sb;
wire TIMEBOOST_net_12981;
wire g61732_db;
wire g61732_sb;
wire TIMEBOOST_net_4880;
wire TIMEBOOST_net_495;
wire g61733_sb;
wire TIMEBOOST_net_13324;
wire g61734_db;
wire g61734_sb;
wire TIMEBOOST_net_4082;
wire g61735_db;
wire g61735_sb;
wire TIMEBOOST_net_4083;
wire g61736_db;
wire g61736_sb;
wire TIMEBOOST_net_4881;
wire TIMEBOOST_net_496;
wire g61737_sb;
wire TIMEBOOST_net_4084;
wire g61738_db;
wire g61738_sb;
wire TIMEBOOST_net_10650;
wire TIMEBOOST_net_281;
wire g61739_sb;
wire TIMEBOOST_net_4085;
wire g61740_db;
wire g61740_sb;
wire TIMEBOOST_net_4086;
wire TIMEBOOST_net_12513;
wire g61741_sb;
wire TIMEBOOST_net_4087;
wire g61742_db;
wire g61742_sb;
wire TIMEBOOST_net_4088;
wire g61743_db;
wire g61743_sb;
wire TIMEBOOST_net_14916;
wire TIMEBOOST_net_10783;
wire g61744_sb;
wire TIMEBOOST_net_4589;
wire TIMEBOOST_net_12246;
wire g61745_sb;
wire TIMEBOOST_net_3995;
wire g61746_db;
wire g61746_sb;
wire TIMEBOOST_net_469;
wire TIMEBOOST_net_10117;
wire g61747_sb;
wire TIMEBOOST_net_4089;
wire g61748_db;
wire g61748_sb;
wire TIMEBOOST_net_3996;
wire g61749_db;
wire g61749_sb;
wire TIMEBOOST_net_3191;
wire TIMEBOOST_net_10273;
wire g61750_sb;
wire TIMEBOOST_net_9324;
wire TIMEBOOST_net_283;
wire g61751_sb;
wire TIMEBOOST_net_470;
wire g61752_db;
wire g61752_sb;
wire TIMEBOOST_net_471;
wire TIMEBOOST_net_4149;
wire g61753_sb;
wire TIMEBOOST_net_472;
wire TIMEBOOST_net_4150;
wire g61754_sb;
wire TIMEBOOST_net_473;
wire TIMEBOOST_net_10274;
wire g61755_sb;
wire TIMEBOOST_net_4882;
wire TIMEBOOST_net_14065;
wire g61756_sb;
wire TIMEBOOST_net_10352;
wire TIMEBOOST_net_10118;
wire g61757_sb;
wire TIMEBOOST_net_14145;
wire TIMEBOOST_net_10119;
wire g61758_sb;
wire TIMEBOOST_net_12312;
wire TIMEBOOST_net_10275;
wire g61759_sb;
wire TIMEBOOST_net_14146;
wire TIMEBOOST_net_10120;
wire g61760_sb;
wire TIMEBOOST_net_9325;
wire TIMEBOOST_net_284;
wire g61761_sb;
wire TIMEBOOST_net_4883;
wire TIMEBOOST_net_498;
wire g61762_sb;
wire TIMEBOOST_net_12298;
wire TIMEBOOST_net_10121;
wire g61763_sb;
wire g61764_db;
wire g61764_sb;
wire TIMEBOOST_net_10666;
wire g61765_db;
wire g61765_sb;
wire TIMEBOOST_net_12333;
wire g61766_db;
wire g61766_sb;
wire TIMEBOOST_net_10673;
wire g61767_db;
wire g61767_sb;
wire TIMEBOOST_net_10548;
wire g61768_db;
wire g61768_sb;
wire TIMEBOOST_net_10656;
wire TIMEBOOST_net_10443;
wire g61769_sb;
wire TIMEBOOST_net_14861;
wire TIMEBOOST_net_10276;
wire g61770_sb;
wire TIMEBOOST_net_4607;
wire g61771_db;
wire g61771_sb;
wire TIMEBOOST_net_351;
wire g61772_db;
wire g61772_sb;
wire TIMEBOOST_net_12320;
wire TIMEBOOST_net_10122;
wire g61773_sb;
wire TIMEBOOST_net_12317;
wire TIMEBOOST_net_10123;
wire g61774_sb;
wire TIMEBOOST_net_10665;
wire g61775_db;
wire g61775_sb;
wire TIMEBOOST_net_10111;
wire g61776_db;
wire TIMEBOOST_net_4610;
wire g61777_db;
wire g61777_sb;
wire TIMEBOOST_net_4884;
wire TIMEBOOST_net_5231;
wire g61778_sb;
wire TIMEBOOST_net_10669;
wire g61779_db;
wire g61779_sb;
wire TIMEBOOST_net_3188;
wire TIMEBOOST_net_10277;
wire g61780_sb;
wire TIMEBOOST_net_10550;
wire g61781_db;
wire g61781_sb;
wire TIMEBOOST_net_750;
wire TIMEBOOST_net_10784;
wire g61782_sb;
wire TIMEBOOST_net_10672;
wire g61783_db;
wire g61783_sb;
wire TIMEBOOST_net_12273;
wire TIMEBOOST_net_4161;
wire g61784_sb;
wire TIMEBOOST_net_4591;
wire TIMEBOOST_net_15003;
wire g61785_sb;
wire TIMEBOOST_net_4592;
wire TIMEBOOST_net_9639;
wire g61786_sb;
wire TIMEBOOST_net_4593;
wire TIMEBOOST_net_288;
wire g61787_sb;
wire TIMEBOOST_net_3170;
wire TIMEBOOST_net_4162;
wire g61788_sb;
wire TIMEBOOST_net_12283;
wire TIMEBOOST_net_4163;
wire g61789_sb;
wire TIMEBOOST_net_10657;
wire TIMEBOOST_net_289;
wire g61790_sb;
wire TIMEBOOST_net_12263;
wire TIMEBOOST_net_4164;
wire g61791_sb;
wire TIMEBOOST_net_3218;
wire TIMEBOOST_net_10367;
wire g61792_sb;
wire TIMEBOOST_net_12280;
wire TIMEBOOST_net_4166;
wire g61793_sb;
wire TIMEBOOST_net_9309;
wire TIMEBOOST_net_290;
wire g61794_sb;
wire TIMEBOOST_net_12326;
wire TIMEBOOST_net_13329;
wire g61795_sb;
wire TIMEBOOST_net_10668;
wire g61796_db;
wire g61796_sb;
wire TIMEBOOST_net_4608;
wire g61797_db;
wire g61797_sb;
wire TIMEBOOST_net_12269;
wire g61798_db;
wire g61798_sb;
wire TIMEBOOST_net_12297;
wire TIMEBOOST_net_4168;
wire g61799_sb;
wire TIMEBOOST_net_12292;
wire TIMEBOOST_net_4169;
wire g61800_sb;
wire TIMEBOOST_net_10310;
wire TIMEBOOST_net_12512;
wire g61801_sb;
wire TIMEBOOST_net_9312;
wire TIMEBOOST_net_291;
wire g61802_sb;
wire TIMEBOOST_net_12284;
wire TIMEBOOST_net_14185;
wire g61803_sb;
wire TIMEBOOST_net_10311;
wire TIMEBOOST_net_9724;
wire g61804_sb;
wire TIMEBOOST_net_12327;
wire TIMEBOOST_net_293;
wire g61805_sb;
wire TIMEBOOST_net_9315;
wire TIMEBOOST_net_294;
wire g61806_sb;
wire TIMEBOOST_net_1097;
wire g61807_db;
wire g61807_sb;
wire TIMEBOOST_net_4016;
wire TIMEBOOST_net_12643;
wire g61808_sb;
wire TIMEBOOST_net_14879;
wire g61809_db;
wire g61809_sb;
wire TIMEBOOST_net_12296;
wire g61810_db;
wire g61810_sb;
wire TIMEBOOST_net_12402;
wire TIMEBOOST_net_295;
wire g61811_sb;
wire TIMEBOOST_net_4017;
wire TIMEBOOST_net_13524;
wire g61812_sb;
wire TIMEBOOST_net_12295;
wire TIMEBOOST_net_4170;
wire g61813_sb;
wire TIMEBOOST_net_4595;
wire TIMEBOOST_net_296;
wire g61814_sb;
wire TIMEBOOST_net_751;
wire TIMEBOOST_net_4764;
wire g61815_sb;
wire TIMEBOOST_net_3237;
wire TIMEBOOST_net_13523;
wire g61816_sb;
wire TIMEBOOST_net_10836;
wire TIMEBOOST_net_15163;
wire g61817_sb;
wire TIMEBOOST_net_12303;
wire TIMEBOOST_net_4171;
wire g61818_sb;
wire TIMEBOOST_net_3265;
wire TIMEBOOST_net_10354;
wire g61819_sb;
wire TIMEBOOST_net_12930;
wire TIMEBOOST_net_12607;
wire g61820_sb;
wire TIMEBOOST_net_4596;
wire TIMEBOOST_net_297;
wire g61821_sb;
wire TIMEBOOST_net_4885;
wire TIMEBOOST_net_10388;
wire g61822_sb;
wire TIMEBOOST_net_9530;
wire TIMEBOOST_net_10369;
wire g61823_sb;
wire TIMEBOOST_net_12332;
wire TIMEBOOST_net_4174;
wire g61824_sb;
wire TIMEBOOST_net_10824;
wire TIMEBOOST_net_501;
wire g61825_sb;
wire TIMEBOOST_net_3225;
wire TIMEBOOST_net_13100;
wire g61826_sb;
wire TIMEBOOST_net_4887;
wire TIMEBOOST_net_9317;
wire g61827_sb;
wire TIMEBOOST_net_10837;
wire TIMEBOOST_net_3765;
wire g61828_sb;
wire TIMEBOOST_net_12651;
wire TIMEBOOST_net_14426;
wire g61829_sb;
wire TIMEBOOST_net_12302;
wire TIMEBOOST_net_4176;
wire g61830_sb;
wire TIMEBOOST_net_14089;
wire g61831_db;
wire g61832_p;
wire g61833_p;
wire g61834_p;
wire TIMEBOOST_net_4568;
wire TIMEBOOST_net_4904;
wire g61835_sb;
wire TIMEBOOST_net_621;
wire g61836_db;
wire g61836_sb;
wire TIMEBOOST_net_13969;
wire g61837_db;
wire g61837_sb;
wire g61838_p;
wire g61839_p;
wire TIMEBOOST_net_13003;
wire g61840_db;
wire g61840_sb;
wire TIMEBOOST_net_13008;
wire g61841_db;
wire g61841_sb;
wire TIMEBOOST_net_723;
wire g61842_db;
wire g61842_sb;
wire TIMEBOOST_net_11355;
wire TIMEBOOST_net_703;
wire g61843_sb;
wire g61846_p;
wire g61850_p;
wire g61851_p;
wire TIMEBOOST_net_14255;
wire TIMEBOOST_net_14924;
wire g61855_sb;
wire TIMEBOOST_net_11330;
wire TIMEBOOST_net_14930;
wire g61856_sb;
wire g61857_p;
wire TIMEBOOST_net_4675;
wire g61858_db;
wire g61858_sb;
wire TIMEBOOST_net_4676;
wire g61859_db;
wire g61859_sb;
wire TIMEBOOST_net_4888;
wire TIMEBOOST_net_503;
wire g61860_sb;
wire TIMEBOOST_net_3176;
wire TIMEBOOST_net_4177;
wire g61861_sb;
wire TIMEBOOST_net_12247;
wire TIMEBOOST_net_4178;
wire g61862_sb;
wire TIMEBOOST_net_4677;
wire g61863_db;
wire g61863_sb;
wire TIMEBOOST_net_10702;
wire g61864_db;
wire g61864_sb;
wire TIMEBOOST_net_4679;
wire g61865_db;
wire g61865_sb;
wire TIMEBOOST_net_9285;
wire g61866_db;
wire g61866_sb;
wire TIMEBOOST_net_14169;
wire TIMEBOOST_net_14449;
wire g61867_sb;
wire TIMEBOOST_net_4680;
wire TIMEBOOST_net_3174;
wire g61868_sb;
wire TIMEBOOST_net_4615;
wire TIMEBOOST_net_1236;
wire g61869_sb;
wire TIMEBOOST_net_4681;
wire g61870_db;
wire g61870_sb;
wire TIMEBOOST_net_9284;
wire TIMEBOOST_net_10376;
wire g61871_sb;
wire TIMEBOOST_net_4682;
wire TIMEBOOST_net_300;
wire g61872_sb;
wire TIMEBOOST_net_13943;
wire TIMEBOOST_net_10127;
wire g61873_sb;
wire TIMEBOOST_net_14586;
wire TIMEBOOST_net_10377;
wire g61874_sb;
wire TIMEBOOST_net_9350;
wire TIMEBOOST_net_9298;
wire g61875_sb;
wire TIMEBOOST_net_9280;
wire TIMEBOOST_net_10378;
wire g61876_sb;
wire TIMEBOOST_net_10704;
wire g61877_db;
wire g61877_sb;
wire TIMEBOOST_net_10840;
wire TIMEBOOST_net_11259;
wire g61878_sb;
wire TIMEBOOST_net_4683;
wire g61879_db;
wire g61879_sb;
wire TIMEBOOST_net_12382;
wire g61880_db;
wire g61880_sb;
wire TIMEBOOST_net_9351;
wire TIMEBOOST_net_302;
wire g61881_sb;
wire TIMEBOOST_net_9281;
wire TIMEBOOST_net_10379;
wire g61882_sb;
wire TIMEBOOST_net_9286;
wire TIMEBOOST_net_4183;
wire g61883_sb;
wire TIMEBOOST_net_12255;
wire TIMEBOOST_net_4184;
wire g61884_sb;
wire TIMEBOOST_net_9323;
wire g61885_db;
wire g61885_sb;
wire TIMEBOOST_net_3194;
wire TIMEBOOST_net_4185;
wire g61886_sb;
wire TIMEBOOST_net_14079;
wire g61887_db;
wire g61887_sb;
wire TIMEBOOST_net_649;
wire TIMEBOOST_net_10380;
wire g61888_sb;
wire TIMEBOOST_net_4873;
wire g61889_db;
wire g61889_sb;
wire TIMEBOOST_net_650;
wire TIMEBOOST_net_13323;
wire g61890_sb;
wire TIMEBOOST_net_10813;
wire g61891_db;
wire g61891_sb;
wire TIMEBOOST_net_12065;
wire TIMEBOOST_net_10205;
wire g61892_sb;
wire TIMEBOOST_net_10190;
wire g61893_db;
wire g61893_sb;
wire TIMEBOOST_net_10736;
wire g61894_db;
wire g61894_sb;
wire TIMEBOOST_net_11197;
wire g61895_db;
wire g61895_sb;
wire TIMEBOOST_net_4867;
wire g61896_db;
wire TIMEBOOST_net_4868;
wire g61897_db;
wire g61897_sb;
wire TIMEBOOST_net_4869;
wire g61898_db;
wire TIMEBOOST_net_4870;
wire g61899_db;
wire g61899_sb;
wire TIMEBOOST_net_652;
wire TIMEBOOST_net_4189;
wire g61900_sb;
wire TIMEBOOST_net_653;
wire TIMEBOOST_net_10371;
wire g61901_sb;
wire TIMEBOOST_net_10844;
wire TIMEBOOST_net_705;
wire g61902_sb;
wire TIMEBOOST_net_10191;
wire g61903_db;
wire g61903_sb;
wire TIMEBOOST_net_4871;
wire g61904_db;
wire g61904_sb;
wire TIMEBOOST_net_10175;
wire TIMEBOOST_net_12306;
wire g61905_sb;
wire TIMEBOOST_net_654;
wire TIMEBOOST_net_4191;
wire g61906_sb;
wire TIMEBOOST_net_12634;
wire g61907_db;
wire g61907_sb;
wire TIMEBOOST_net_10166;
wire TIMEBOOST_net_12272;
wire g61908_sb;
wire TIMEBOOST_net_10167;
wire g61909_db;
wire g61909_sb;
wire TIMEBOOST_net_4810;
wire TIMEBOOST_net_305;
wire g61910_sb;
wire TIMEBOOST_net_655;
wire TIMEBOOST_net_4192;
wire g61911_sb;
wire TIMEBOOST_net_685;
wire g61912_db;
wire g61912_sb;
wire TIMEBOOST_net_4811;
wire TIMEBOOST_net_306;
wire g61913_sb;
wire TIMEBOOST_net_4812;
wire TIMEBOOST_net_307;
wire g61914_sb;
wire TIMEBOOST_net_656;
wire TIMEBOOST_net_9934;
wire g61915_sb;
wire TIMEBOOST_net_9935;
wire g61916_sb;
wire TIMEBOOST_net_10882;
wire TIMEBOOST_net_706;
wire g61917_sb;
wire TIMEBOOST_net_4872;
wire g61918_db;
wire g61918_sb;
wire TIMEBOOST_net_4813;
wire TIMEBOOST_net_308;
wire g61919_sb;
wire TIMEBOOST_net_3879;
wire TIMEBOOST_net_13522;
wire TIMEBOOST_net_12650;
wire TIMEBOOST_net_14281;
wire g61921_sb;
wire TIMEBOOST_net_3880;
wire g61922_db;
wire TIMEBOOST_net_1128;
wire g61923_db;
wire g61923_sb;
wire TIMEBOOST_net_10240;
wire TIMEBOOST_net_13521;
wire g61924_sb;
wire TIMEBOOST_net_13520;
wire g61925_sb;
wire TIMEBOOST_net_12328;
wire TIMEBOOST_net_4195;
wire g61926_sb;
wire TIMEBOOST_net_12304;
wire TIMEBOOST_net_13341;
wire g61927_sb;
wire TIMEBOOST_net_3883;
wire TIMEBOOST_net_13519;
wire TIMEBOOST_net_3884;
wire g61929_db;
wire g61929_sb;
wire TIMEBOOST_net_10243;
wire TIMEBOOST_net_12353;
wire g61930_sb;
wire TIMEBOOST_net_10244;
wire TIMEBOOST_net_13518;
wire g61931_sb;
wire TIMEBOOST_net_10245;
wire TIMEBOOST_net_13517;
wire g61932_sb;
wire TIMEBOOST_net_10215;
wire TIMEBOOST_net_12748;
wire g61933_sb;
wire TIMEBOOST_net_13118;
wire TIMEBOOST_net_12361;
wire g61934_sb;
wire TIMEBOOST_net_13119;
wire TIMEBOOST_net_13516;
wire TIMEBOOST_net_10896;
wire TIMEBOOST_net_707;
wire g61936_sb;
wire TIMEBOOST_net_10658;
wire TIMEBOOST_net_309;
wire g61937_sb;
wire TIMEBOOST_net_13386;
wire TIMEBOOST_net_13515;
wire TIMEBOOST_net_3892;
wire g61939_db;
wire g61939_sb;
wire TIMEBOOST_net_12855;
wire TIMEBOOST_net_9936;
wire g61940_sb;
wire TIMEBOOST_net_13901;
wire TIMEBOOST_net_14325;
wire g61941_sb;
wire TIMEBOOST_net_9381;
wire TIMEBOOST_net_14305;
wire g61942_sb;
wire TIMEBOOST_net_12386;
wire g61943_db;
wire g61943_sb;
wire TIMEBOOST_net_4598;
wire TIMEBOOST_net_3121;
wire g61944_sb;
wire TIMEBOOST_net_734;
wire TIMEBOOST_net_14232;
wire g61945_sb;
wire TIMEBOOST_net_12271;
wire TIMEBOOST_net_10155;
wire g61946_sb;
wire TIMEBOOST_net_12282;
wire TIMEBOOST_net_10156;
wire g61947_sb;
wire TIMEBOOST_net_735;
wire TIMEBOOST_net_14448;
wire g61948_sb;
wire TIMEBOOST_net_3893;
wire g61949_db;
wire g61949_sb;
wire TIMEBOOST_net_736;
wire TIMEBOOST_net_14560;
wire g61950_sb;
wire TIMEBOOST_net_12265;
wire TIMEBOOST_net_10160;
wire g61951_sb;
wire TIMEBOOST_net_737;
wire TIMEBOOST_net_10381;
wire g61952_sb;
wire TIMEBOOST_net_3518;
wire g61953_db;
wire TIMEBOOST_net_10659;
wire TIMEBOOST_net_311;
wire g61954_sb;
wire TIMEBOOST_net_12983;
wire TIMEBOOST_net_12066;
wire g61955_sb;
wire TIMEBOOST_net_12751;
wire g61956_db;
wire g61956_sb;
wire TIMEBOOST_net_623;
wire g61957_db;
wire g61957_sb;
wire TIMEBOOST_net_12984;
wire TIMEBOOST_net_12844;
wire g61958_sb;
wire TIMEBOOST_net_624;
wire g61959_db;
wire g61959_sb;
wire TIMEBOOST_net_12393;
wire g61960_db;
wire TIMEBOOST_net_12985;
wire g61961_db;
wire g61961_sb;
wire TIMEBOOST_net_1130;
wire g61962_db;
wire g61962_sb;
wire TIMEBOOST_net_739;
wire g61963_db;
wire g61963_sb;
wire TIMEBOOST_net_14131;
wire g61964_db;
wire TIMEBOOST_net_625;
wire g61965_db;
wire g61965_sb;
wire TIMEBOOST_net_9321;
wire g61966_db;
wire TIMEBOOST_net_12299;
wire g61967_db;
wire TIMEBOOST_net_12373;
wire g61968_db;
wire TIMEBOOST_net_13922;
wire g61969_db;
wire TIMEBOOST_net_9319;
wire g61970_db;
wire TIMEBOOST_net_14871;
wire g61971_db;
wire TIMEBOOST_net_11000;
wire g61972_db;
wire TIMEBOOST_net_14789;
wire g61973_db;
wire TIMEBOOST_net_11008;
wire g61974_db;
wire TIMEBOOST_net_1134;
wire g61975_db;
wire TIMEBOOST_net_11002;
wire g61976_db;
wire TIMEBOOST_net_9320;
wire g61977_db;
wire TIMEBOOST_net_11003;
wire g61978_db;
wire TIMEBOOST_net_1135;
wire g61979_db;
wire TIMEBOOST_net_1136;
wire g61980_db;
wire TIMEBOOST_net_11006;
wire g61981_db;
wire TIMEBOOST_net_11005;
wire g61982_db;
wire TIMEBOOST_net_1137;
wire g61983_db;
wire TIMEBOOST_net_9328;
wire g61984_db;
wire TIMEBOOST_net_1138;
wire g61985_db;
wire TIMEBOOST_net_9322;
wire g61986_db;
wire TIMEBOOST_net_1139;
wire g61987_db;
wire TIMEBOOST_net_12400;
wire g61988_db;
wire TIMEBOOST_net_1140;
wire g61989_db;
wire TIMEBOOST_net_3894;
wire TIMEBOOST_net_13514;
wire g61990_sb;
wire TIMEBOOST_net_4890;
wire TIMEBOOST_net_505;
wire g61991_sb;
wire TIMEBOOST_net_3895;
wire TIMEBOOST_net_13513;
wire g61992_sb;
wire TIMEBOOST_net_12261;
wire TIMEBOOST_net_10193;
wire g61993_sb;
wire TIMEBOOST_net_3896;
wire g61994_db;
wire g61994_sb;
wire TIMEBOOST_net_12267;
wire TIMEBOOST_net_4203;
wire g61995_sb;
wire TIMEBOOST_net_3897;
wire g61996_db;
wire TIMEBOOST_net_3898;
wire TIMEBOOST_net_12509;
wire g61997_sb;
wire TIMEBOOST_net_12260;
wire TIMEBOOST_net_4204;
wire g61998_sb;
wire TIMEBOOST_net_3899;
wire TIMEBOOST_net_12508;
wire g61999_sb;
wire TIMEBOOST_net_12270;
wire TIMEBOOST_net_10128;
wire g62000_sb;
wire TIMEBOOST_net_408;
wire TIMEBOOST_net_4205;
wire g62001_sb;
wire TIMEBOOST_net_409;
wire TIMEBOOST_net_4206;
wire g62002_sb;
wire TIMEBOOST_net_10227;
wire TIMEBOOST_net_12507;
wire g62003_sb;
wire TIMEBOOST_net_10228;
wire TIMEBOOST_net_9744;
wire TIMEBOOST_net_477;
wire TIMEBOOST_net_14171;
wire g62005_sb;
wire TIMEBOOST_net_10660;
wire TIMEBOOST_net_3400;
wire g62006_sb;
wire TIMEBOOST_net_10229;
wire TIMEBOOST_net_13507;
wire g62007_sb;
wire TIMEBOOST_net_10280;
wire g62008_db;
wire TIMEBOOST_net_10353;
wire TIMEBOOST_net_14656;
wire g62009_sb;
wire TIMEBOOST_net_9326;
wire TIMEBOOST_net_313;
wire g62010_sb;
wire TIMEBOOST_net_591;
wire TIMEBOOST_net_14248;
wire g62011_sb;
wire TIMEBOOST_net_12237;
wire TIMEBOOST_net_12475;
wire g62012_sb;
wire TIMEBOOST_net_480;
wire TIMEBOOST_net_14655;
wire g62013_sb;
wire TIMEBOOST_net_481;
wire TIMEBOOST_net_4765;
wire g62014_sb;
wire TIMEBOOST_net_4601;
wire TIMEBOOST_net_10091;
wire g62015_sb;
wire TIMEBOOST_net_482;
wire TIMEBOOST_net_14654;
wire g62016_sb;
wire TIMEBOOST_net_4891;
wire TIMEBOOST_net_506;
wire g62017_sb;
wire TIMEBOOST_net_12238;
wire TIMEBOOST_net_4766;
wire g62018_sb;
wire TIMEBOOST_net_4892;
wire TIMEBOOST_net_507;
wire g62019_sb;
wire TIMEBOOST_net_10897;
wire TIMEBOOST_net_15112;
wire g62020_sb;
wire TIMEBOOST_net_14819;
wire g62021_db;
wire TIMEBOOST_net_12243;
wire TIMEBOOST_net_14653;
wire g62022_sb;
wire TIMEBOOST_net_4893;
wire TIMEBOOST_net_13950;
wire g62023_sb;
wire TIMEBOOST_net_12661;
wire TIMEBOOST_net_4767;
wire g62024_sb;
wire TIMEBOOST_net_12244;
wire g62025_db;
wire g62025_sb;
wire TIMEBOOST_net_12662;
wire TIMEBOOST_net_4768;
wire g62026_sb;
wire TIMEBOOST_net_3178;
wire TIMEBOOST_net_14652;
wire g62027_sb;
wire TIMEBOOST_net_3175;
wire TIMEBOOST_net_14651;
wire g62028_sb;
wire TIMEBOOST_net_3197;
wire TIMEBOOST_net_10043;
wire g62029_sb;
wire TIMEBOOST_net_11332;
wire TIMEBOOST_net_14791;
wire g62030_sb;
wire TIMEBOOST_net_14892;
wire TIMEBOOST_net_4492;
wire g62031_sb;
wire TIMEBOOST_net_11407;
wire TIMEBOOST_net_14756;
wire g62032_sb;
wire TIMEBOOST_net_13909;
wire TIMEBOOST_net_10497;
wire g62033_sb;
wire TIMEBOOST_net_12232;
wire TIMEBOOST_net_11033;
wire g62034_sb;
wire TIMEBOOST_net_1427;
wire TIMEBOOST_net_14433;
wire g62035_sb;
wire TIMEBOOST_net_5448;
wire TIMEBOOST_net_12377;
wire g62036_sb;
wire TIMEBOOST_net_1428;
wire TIMEBOOST_net_14295;
wire g62037_sb;
wire TIMEBOOST_net_1429;
wire TIMEBOOST_net_11034;
wire g62038_sb;
wire TIMEBOOST_net_14505;
wire TIMEBOOST_net_11036;
wire g62039_sb;
wire TIMEBOOST_net_1431;
wire TIMEBOOST_net_11333;
wire g62040_sb;
wire TIMEBOOST_net_14492;
wire TIMEBOOST_net_14434;
wire g62041_sb;
wire TIMEBOOST_net_1433;
wire TIMEBOOST_net_11177;
wire g62042_sb;
wire TIMEBOOST_net_12996;
wire TIMEBOOST_net_12376;
wire g62043_sb;
wire TIMEBOOST_net_11342;
wire TIMEBOOST_net_12383;
wire g62044_sb;
wire TIMEBOOST_net_14318;
wire TIMEBOOST_net_11208;
wire g62045_sb;
wire TIMEBOOST_net_11343;
wire TIMEBOOST_net_12362;
wire g62046_sb;
wire TIMEBOOST_net_14495;
wire TIMEBOOST_net_11180;
wire g62047_sb;
wire TIMEBOOST_net_1436;
wire TIMEBOOST_net_5593;
wire g62048_sb;
wire TIMEBOOST_net_1437;
wire TIMEBOOST_net_5592;
wire g62049_sb;
wire TIMEBOOST_net_14476;
wire TIMEBOOST_net_13995;
wire g62050_sb;
wire TIMEBOOST_net_11344;
wire TIMEBOOST_net_14759;
wire g62051_sb;
wire TIMEBOOST_net_10001;
wire TIMEBOOST_net_13902;
wire g62052_sb;
wire TIMEBOOST_net_10002;
wire TIMEBOOST_net_11181;
wire g62053_sb;
wire TIMEBOOST_net_11345;
wire TIMEBOOST_net_14951;
wire g62054_sb;
wire TIMEBOOST_net_11346;
wire TIMEBOOST_net_13214;
wire g62055_sb;
wire TIMEBOOST_net_10003;
wire TIMEBOOST_net_13903;
wire g62056_sb;
wire TIMEBOOST_net_11347;
wire TIMEBOOST_net_1164;
wire g62057_sb;
wire TIMEBOOST_net_3177;
wire TIMEBOOST_net_14234;
wire g62058_sb;
wire TIMEBOOST_net_1442;
wire TIMEBOOST_net_13904;
wire g62059_sb;
wire TIMEBOOST_net_1443;
wire TIMEBOOST_net_13905;
wire g62060_sb;
wire TIMEBOOST_net_11348;
wire TIMEBOOST_net_1165;
wire g62061_sb;
wire TIMEBOOST_net_11349;
wire TIMEBOOST_net_1166;
wire g62062_sb;
wire TIMEBOOST_net_1444;
wire TIMEBOOST_net_13906;
wire g62063_sb;
wire TIMEBOOST_net_11350;
wire TIMEBOOST_net_13401;
wire g62064_sb;
wire TIMEBOOST_net_1445;
wire n_13214;
wire g62065_sb;
wire TIMEBOOST_net_10661;
wire TIMEBOOST_net_315;
wire g62066_sb;
wire TIMEBOOST_net_5313;
wire TIMEBOOST_net_12367;
wire g62067_sb;
wire TIMEBOOST_net_9365;
wire TIMEBOOST_net_11041;
wire g62068_sb;
wire TIMEBOOST_net_4603;
wire TIMEBOOST_net_316;
wire g62069_sb;
wire TIMEBOOST_net_10663;
wire TIMEBOOST_net_317;
wire g62070_sb;
wire TIMEBOOST_net_3179;
wire TIMEBOOST_net_14453;
wire g62071_sb;
wire TIMEBOOST_net_3187;
wire TIMEBOOST_net_10471;
wire g62072_sb;
wire TIMEBOOST_net_4562;
wire TIMEBOOST_net_10773;
wire g62073_sb;
wire TIMEBOOST_net_808;
wire TIMEBOOST_net_10774;
wire g62074_sb;
wire TIMEBOOST_net_809;
wire TIMEBOOST_net_10775;
wire g62075_sb;
wire TIMEBOOST_net_810;
wire TIMEBOOST_net_4822;
wire g62076_sb;
wire TIMEBOOST_net_432;
wire TIMEBOOST_net_10472;
wire g62077_sb;
wire TIMEBOOST_net_3168;
wire TIMEBOOST_net_10473;
wire g62078_sb;
wire TIMEBOOST_net_811;
wire TIMEBOOST_net_4823;
wire g62079_sb;
wire TIMEBOOST_net_9678;
wire TIMEBOOST_net_4824;
wire g62080_sb;
wire TIMEBOOST_net_4398;
wire TIMEBOOST_net_4825;
wire g62081_sb;
wire TIMEBOOST_net_10989;
wire n_10257;
wire g62082_sb;
wire TIMEBOOST_net_10990;
wire g62083_sb;
wire TIMEBOOST_net_10991;
wire TIMEBOOST_net_11013;
wire g62084_sb;
wire TIMEBOOST_net_10992;
wire TIMEBOOST_net_662;
wire g62085_sb;
wire TIMEBOOST_net_10994;
wire TIMEBOOST_net_663;
wire g62086_sb;
wire TIMEBOOST_net_10996;
wire TIMEBOOST_net_664;
wire g62087_sb;
wire TIMEBOOST_net_10999;
wire TIMEBOOST_net_10785;
wire g62088_sb;
wire TIMEBOOST_net_11001;
wire TIMEBOOST_net_666;
wire g62089_sb;
wire TIMEBOOST_net_12245;
wire TIMEBOOST_net_10474;
wire g62090_sb;
wire TIMEBOOST_net_4399;
wire TIMEBOOST_net_4826;
wire g62091_sb;
wire TIMEBOOST_net_11004;
wire TIMEBOOST_net_12803;
wire g62092_sb;
wire TIMEBOOST_net_4400;
wire TIMEBOOST_net_4827;
wire g62093_sb;
wire TIMEBOOST_net_3212;
wire TIMEBOOST_net_4096;
wire g62094_sb;
wire TIMEBOOST_net_9282;
wire TIMEBOOST_net_4097;
wire g62095_sb;
wire TIMEBOOST_net_4401;
wire TIMEBOOST_net_4828;
wire g62096_sb;
wire TIMEBOOST_net_4402;
wire TIMEBOOST_net_4829;
wire g62097_sb;
wire TIMEBOOST_net_4403;
wire TIMEBOOST_net_4830;
wire g62098_sb;
wire TIMEBOOST_net_4404;
wire TIMEBOOST_net_10776;
wire g62099_sb;
wire TIMEBOOST_net_4405;
wire TIMEBOOST_net_4832;
wire g62100_sb;
wire TIMEBOOST_net_12240;
wire TIMEBOOST_net_4098;
wire g62101_sb;
wire TIMEBOOST_net_10640;
wire TIMEBOOST_net_4833;
wire g62102_sb;
wire TIMEBOOST_net_822;
wire TIMEBOOST_net_4834;
wire g62103_sb;
wire TIMEBOOST_net_10143;
wire TIMEBOOST_net_14097;
wire g62104_sb;
wire TIMEBOOST_net_10145;
wire TIMEBOOST_net_4835;
wire g62105_sb;
wire TIMEBOOST_net_3192;
wire TIMEBOOST_net_4099;
wire g62106_sb;
wire TIMEBOOST_net_10146;
wire TIMEBOOST_net_4836;
wire g62107_sb;
wire TIMEBOOST_net_13225;
wire TIMEBOOST_net_4837;
wire g62108_sb;
wire TIMEBOOST_net_10153;
wire TIMEBOOST_net_4838;
wire g62109_sb;
wire TIMEBOOST_net_11007;
wire TIMEBOOST_net_668;
wire g62110_sb;
wire TIMEBOOST_net_12291;
wire g62111_db;
wire g62111_sb;
wire TIMEBOOST_net_828;
wire TIMEBOOST_net_10790;
wire g62112_sb;
wire TIMEBOOST_net_829;
wire TIMEBOOST_net_13964;
wire g62113_sb;
wire TIMEBOOST_net_12248;
wire g62114_db;
wire g62114_sb;
wire TIMEBOOST_net_9352;
wire TIMEBOOST_net_3729;
wire g62115_sb;
wire TIMEBOOST_net_12268;
wire g62116_db;
wire g62116_sb;
wire TIMEBOOST_net_11009;
wire TIMEBOOST_net_12605;
wire g62117_sb;
wire TIMEBOOST_net_11010;
wire TIMEBOOST_net_9436;
wire g62118_sb;
wire TIMEBOOST_net_442;
wire g62119_db;
wire g62119_sb;
wire TIMEBOOST_net_11011;
wire TIMEBOOST_net_3742;
wire g62120_sb;
wire TIMEBOOST_net_10791;
wire g62121_sb;
wire TIMEBOOST_net_13202;
wire TIMEBOOST_net_10792;
wire g62122_sb;
wire TIMEBOOST_net_11016;
wire TIMEBOOST_net_673;
wire g62123_sb;
wire TIMEBOOST_net_443;
wire TIMEBOOST_net_10133;
wire g62124_sb;
wire TIMEBOOST_net_11017;
wire TIMEBOOST_net_12599;
wire g62125_sb;
wire TIMEBOOST_net_11018;
wire TIMEBOOST_net_9437;
wire g62126_sb;
wire TIMEBOOST_net_13203;
wire TIMEBOOST_net_10793;
wire g62127_sb;
wire TIMEBOOST_net_13204;
wire TIMEBOOST_net_10794;
wire g62128_sb;
wire TIMEBOOST_net_11020;
wire TIMEBOOST_net_12591;
wire g62129_sb;
wire TIMEBOOST_net_834;
wire TIMEBOOST_net_11194;
wire g62130_sb;
wire TIMEBOOST_net_12689;
wire TIMEBOOST_net_10795;
wire g62131_sb;
wire TIMEBOOST_net_444;
wire TIMEBOOST_net_10134;
wire g62132_sb;
wire TIMEBOOST_net_12266;
wire TIMEBOOST_net_10278;
wire g62133_sb;
wire TIMEBOOST_net_12329;
wire TIMEBOOST_net_10279;
wire g62134_sb;
wire TIMEBOOST_net_10898;
wire TIMEBOOST_net_15155;
wire g62135_sb;
wire TIMEBOOST_net_10901;
wire TIMEBOOST_net_678;
wire g62136_sb;
wire TIMEBOOST_net_12633;
wire TIMEBOOST_net_10796;
wire g62137_sb;
wire TIMEBOOST_net_11021;
wire TIMEBOOST_net_679;
wire g62138_sb;
wire TIMEBOOST_net_2960;
wire TIMEBOOST_net_10797;
wire g62139_sb;
wire TIMEBOOST_net_9353;
wire TIMEBOOST_net_12573;
wire g62140_sb;
wire TIMEBOOST_net_2961;
wire TIMEBOOST_net_10798;
wire g62141_sb;
wire g62219_p;
wire g62220_p;
wire g62221_p;
wire g62223_p;
wire g62254_p;
wire g62264_p;
wire g62285_p;
wire g62312_p;
wire g62318_p;
wire g62319_p;
wire TIMEBOOST_net_1525;
wire g62326_db;
wire g62326_sb;
wire TIMEBOOST_net_11362;
wire TIMEBOOST_net_14880;
wire g62333_sb;
wire TIMEBOOST_net_11363;
wire TIMEBOOST_net_12351;
wire g62334_sb;
wire TIMEBOOST_net_1526;
wire TIMEBOOST_net_11260;
wire g62335_sb;
wire TIMEBOOST_net_11364;
wire TIMEBOOST_net_1206;
wire g62336_sb;
wire TIMEBOOST_net_13915;
wire TIMEBOOST_net_11819;
wire g62337_sb;
wire TIMEBOOST_net_14442;
wire TIMEBOOST_net_11820;
wire g62338_sb;
wire TIMEBOOST_net_11841;
wire TIMEBOOST_net_10513;
wire g62339_sb;
wire TIMEBOOST_net_1527;
wire TIMEBOOST_net_11261;
wire g62340_sb;
wire TIMEBOOST_net_11365;
wire TIMEBOOST_net_1207;
wire g62341_sb;
wire TIMEBOOST_net_11366;
wire TIMEBOOST_net_1208;
wire g62342_sb;
wire TIMEBOOST_net_11367;
wire TIMEBOOST_net_1209;
wire g62343_sb;
wire TIMEBOOST_net_1528;
wire TIMEBOOST_net_5445;
wire g62344_sb;
wire TIMEBOOST_net_11665;
wire TIMEBOOST_net_14028;
wire g62345_sb;
wire TIMEBOOST_net_14370;
wire TIMEBOOST_net_11821;
wire g62346_sb;
wire TIMEBOOST_net_11368;
wire TIMEBOOST_net_1210;
wire g62347_sb;
wire TIMEBOOST_net_11842;
wire TIMEBOOST_net_1675;
wire g62348_sb;
wire TIMEBOOST_net_11369;
wire TIMEBOOST_net_1211;
wire g62349_sb;
wire TIMEBOOST_net_11370;
wire TIMEBOOST_net_1212;
wire g62350_sb;
wire TIMEBOOST_net_11667;
wire TIMEBOOST_net_14095;
wire g62351_sb;
wire TIMEBOOST_net_1529;
wire TIMEBOOST_net_11209;
wire g62352_sb;
wire TIMEBOOST_net_11371;
wire TIMEBOOST_net_3649;
wire g62353_sb;
wire TIMEBOOST_net_11372;
wire TIMEBOOST_net_1214;
wire g62354_sb;
wire TIMEBOOST_net_11843;
wire TIMEBOOST_net_1725;
wire g62355_sb;
wire TIMEBOOST_net_11373;
wire TIMEBOOST_net_1215;
wire g62356_sb;
wire TIMEBOOST_net_1530;
wire TIMEBOOST_net_11210;
wire g62357_sb;
wire TIMEBOOST_net_14345;
wire TIMEBOOST_net_11211;
wire g62358_sb;
wire TIMEBOOST_net_11374;
wire TIMEBOOST_net_1216;
wire g62359_sb;
wire TIMEBOOST_net_11375;
wire TIMEBOOST_net_12338;
wire g62360_sb;
wire TIMEBOOST_net_11376;
wire TIMEBOOST_net_12778;
wire g62361_sb;
wire TIMEBOOST_net_12324;
wire TIMEBOOST_net_11815;
wire g62362_sb;
wire TIMEBOOST_net_11846;
wire TIMEBOOST_net_1676;
wire g62363_sb;
wire TIMEBOOST_net_11377;
wire TIMEBOOST_net_1219;
wire g62364_sb;
wire TIMEBOOST_net_14149;
wire TIMEBOOST_net_11212;
wire g62365_sb;
wire TIMEBOOST_net_12323;
wire g62366_db;
wire g62366_sb;
wire TIMEBOOST_net_11847;
wire TIMEBOOST_net_10425;
wire g62367_sb;
wire TIMEBOOST_net_11848;
wire TIMEBOOST_net_14367;
wire g62368_sb;
wire TIMEBOOST_net_11378;
wire TIMEBOOST_net_13541;
wire g62369_sb;
wire TIMEBOOST_net_11849;
wire TIMEBOOST_net_14436;
wire g62370_sb;
wire TIMEBOOST_net_14143;
wire TIMEBOOST_net_11213;
wire g62371_sb;
wire TIMEBOOST_net_14156;
wire TIMEBOOST_net_11214;
wire g62372_sb;
wire TIMEBOOST_net_11379;
wire TIMEBOOST_net_12656;
wire g62373_sb;
wire TIMEBOOST_net_11380;
wire TIMEBOOST_net_1222;
wire g62374_sb;
wire TIMEBOOST_net_11381;
wire TIMEBOOST_net_13540;
wire g62375_sb;
wire TIMEBOOST_net_11382;
wire TIMEBOOST_net_14831;
wire g62376_sb;
wire TIMEBOOST_net_11383;
wire TIMEBOOST_net_14953;
wire g62377_sb;
wire TIMEBOOST_net_13917;
wire TIMEBOOST_net_11822;
wire g62378_sb;
wire TIMEBOOST_net_11850;
wire TIMEBOOST_net_14532;
wire g62379_sb;
wire TIMEBOOST_net_11384;
wire TIMEBOOST_net_13539;
wire g62380_sb;
wire TIMEBOOST_net_11851;
wire TIMEBOOST_net_14464;
wire g62381_sb;
wire TIMEBOOST_net_11852;
wire TIMEBOOST_net_14499;
wire g62382_sb;
wire TIMEBOOST_net_11385;
wire TIMEBOOST_net_14954;
wire g62383_sb;
wire TIMEBOOST_net_1537;
wire TIMEBOOST_net_10829;
wire g62384_sb;
wire TIMEBOOST_net_11386;
wire TIMEBOOST_net_14956;
wire g62385_sb;
wire TIMEBOOST_net_11387;
wire TIMEBOOST_net_14957;
wire g62386_sb;
wire TIMEBOOST_net_14779;
wire TIMEBOOST_net_11356;
wire g62387_sb;
wire TIMEBOOST_net_11388;
wire TIMEBOOST_net_14958;
wire g62388_sb;
wire TIMEBOOST_net_11389;
wire TIMEBOOST_net_14475;
wire g62389_sb;
wire TIMEBOOST_net_11390;
wire TIMEBOOST_net_14959;
wire g62390_sb;
wire TIMEBOOST_net_11391;
wire TIMEBOOST_net_14881;
wire g62391_sb;
wire TIMEBOOST_net_11392;
wire TIMEBOOST_net_14962;
wire g62392_sb;
wire TIMEBOOST_net_10082;
wire TIMEBOOST_net_13812;
wire g62393_sb;
wire TIMEBOOST_net_11215;
wire g62394_sb;
wire TIMEBOOST_net_11669;
wire TIMEBOOST_net_1860;
wire g62395_sb;
wire TIMEBOOST_net_11859;
wire TIMEBOOST_net_14500;
wire g62396_sb;
wire TIMEBOOST_net_11393;
wire TIMEBOOST_net_14963;
wire g62397_sb;
wire TIMEBOOST_net_11394;
wire TIMEBOOST_net_14964;
wire g62398_sb;
wire TIMEBOOST_net_14138;
wire TIMEBOOST_net_11216;
wire g62399_sb;
wire TIMEBOOST_net_11862;
wire TIMEBOOST_net_14501;
wire g62400_sb;
wire TIMEBOOST_net_11639;
wire TIMEBOOST_net_14081;
wire g62401_sb;
wire TIMEBOOST_net_11865;
wire TIMEBOOST_net_10426;
wire g62402_sb;
wire TIMEBOOST_net_11866;
wire TIMEBOOST_net_12226;
wire g62403_sb;
wire TIMEBOOST_net_11867;
wire TIMEBOOST_net_14348;
wire g62404_sb;
wire TIMEBOOST_net_11395;
wire TIMEBOOST_net_1235;
wire g62405_sb;
wire TIMEBOOST_net_11507;
wire TIMEBOOST_net_14750;
wire g62406_sb;
wire TIMEBOOST_net_11709;
wire TIMEBOOST_net_14430;
wire g62407_sb;
wire TIMEBOOST_net_11719;
wire TIMEBOOST_net_13971;
wire g62408_sb;
wire TIMEBOOST_net_11511;
wire TIMEBOOST_net_14103;
wire g62409_sb;
wire TIMEBOOST_net_11396;
wire TIMEBOOST_net_12777;
wire g62410_sb;
wire TIMEBOOST_net_10084;
wire TIMEBOOST_net_11217;
wire g62411_sb;
wire TIMEBOOST_net_9303;
wire TIMEBOOST_net_11218;
wire g62412_sb;
wire TIMEBOOST_net_11397;
wire TIMEBOOST_net_14875;
wire g62413_sb;
wire TIMEBOOST_net_11398;
wire TIMEBOOST_net_13538;
wire g62414_sb;
wire TIMEBOOST_net_11399;
wire TIMEBOOST_net_13537;
wire g62415_sb;
wire TIMEBOOST_net_11666;
wire TIMEBOOST_net_14071;
wire g62416_sb;
wire TIMEBOOST_net_11400;
wire TIMEBOOST_net_1240;
wire g62417_sb;
wire TIMEBOOST_net_11401;
wire TIMEBOOST_net_1241;
wire g62418_sb;
wire TIMEBOOST_net_11402;
wire TIMEBOOST_net_1242;
wire g62419_sb;
wire TIMEBOOST_net_11403;
wire TIMEBOOST_net_14782;
wire g62420_sb;
wire TIMEBOOST_net_11514;
wire TIMEBOOST_net_1682;
wire g62421_sb;
wire TIMEBOOST_net_11404;
wire TIMEBOOST_net_14785;
wire g62422_sb;
wire TIMEBOOST_net_1544;
wire TIMEBOOST_net_11219;
wire g62423_sb;
wire TIMEBOOST_net_11405;
wire TIMEBOOST_net_14811;
wire g62424_sb;
wire TIMEBOOST_net_11668;
wire TIMEBOOST_net_14423;
wire g62425_sb;
wire TIMEBOOST_net_14591;
wire TIMEBOOST_net_11220;
wire g62426_sb;
wire TIMEBOOST_net_11670;
wire TIMEBOOST_net_13924;
wire g62427_sb;
wire TIMEBOOST_net_9304;
wire TIMEBOOST_net_11221;
wire g62428_sb;
wire TIMEBOOST_net_10355;
wire TIMEBOOST_net_13283;
wire g62429_sb;
wire TIMEBOOST_net_10356;
wire TIMEBOOST_net_14906;
wire g62430_sb;
wire TIMEBOOST_net_11524;
wire TIMEBOOST_net_14328;
wire g62431_sb;
wire TIMEBOOST_net_11526;
wire TIMEBOOST_net_1735;
wire g62432_sb;
wire TIMEBOOST_net_11672;
wire TIMEBOOST_net_13976;
wire g62433_sb;
wire TIMEBOOST_net_11516;
wire TIMEBOOST_net_14502;
wire g62434_sb;
wire TIMEBOOST_net_11518;
wire TIMEBOOST_net_14503;
wire g62435_sb;
wire TIMEBOOST_net_10357;
wire TIMEBOOST_net_14910;
wire g62436_sb;
wire TIMEBOOST_net_10358;
wire TIMEBOOST_net_14907;
wire g62437_sb;
wire TIMEBOOST_net_10359;
wire TIMEBOOST_net_14931;
wire g62438_sb;
wire TIMEBOOST_net_11905;
wire TIMEBOOST_net_14115;
wire g62439_sb;
wire TIMEBOOST_net_14200;
wire TIMEBOOST_net_11257;
wire g62440_sb;
wire TIMEBOOST_net_11523;
wire TIMEBOOST_net_13938;
wire g62441_sb;
wire TIMEBOOST_net_10360;
wire TIMEBOOST_net_14935;
wire g62442_sb;
wire TIMEBOOST_net_10361;
wire TIMEBOOST_net_15038;
wire g62443_sb;
wire TIMEBOOST_net_11651;
wire TIMEBOOST_net_14060;
wire g62444_sb;
wire TIMEBOOST_net_10362;
wire TIMEBOOST_net_14940;
wire g62445_sb;
wire TIMEBOOST_net_11664;
wire TIMEBOOST_net_14286;
wire g62446_sb;
wire TIMEBOOST_net_14371;
wire TIMEBOOST_net_11812;
wire g62447_sb;
wire TIMEBOOST_net_10363;
wire TIMEBOOST_net_14941;
wire g62448_sb;
wire TIMEBOOST_net_10364;
wire TIMEBOOST_net_14961;
wire g62449_sb;
wire TIMEBOOST_net_12251;
wire TIMEBOOST_net_11262;
wire g62450_sb;
wire TIMEBOOST_net_11676;
wire TIMEBOOST_net_14440;
wire g62451_sb;
wire TIMEBOOST_net_10365;
wire TIMEBOOST_net_14965;
wire g62452_sb;
wire TIMEBOOST_net_11528;
wire TIMEBOOST_net_14300;
wire g62453_sb;
wire TIMEBOOST_net_10366;
wire TIMEBOOST_net_14966;
wire g62454_sb;
wire TIMEBOOST_net_11525;
wire TIMEBOOST_net_13916;
wire g62455_sb;
wire TIMEBOOST_net_14191;
wire TIMEBOOST_net_11263;
wire g62456_sb;
wire TIMEBOOST_net_11527;
wire TIMEBOOST_net_1738;
wire g62457_sb;
wire TIMEBOOST_net_11206;
wire TIMEBOOST_net_14987;
wire g62458_sb;
wire TIMEBOOST_net_5527;
wire TIMEBOOST_net_14988;
wire g62459_sb;
wire TIMEBOOST_net_15259;
wire TIMEBOOST_net_11264;
wire g62460_sb;
wire TIMEBOOST_net_11530;
wire TIMEBOOST_net_14195;
wire g62461_sb;
wire TIMEBOOST_net_11409;
wire TIMEBOOST_net_1424;
wire g62462_sb;
wire TIMEBOOST_net_11410;
wire TIMEBOOST_net_14989;
wire g62463_sb;
wire TIMEBOOST_net_11411;
wire TIMEBOOST_net_15202;
wire g62464_sb;
wire TIMEBOOST_net_11531;
wire TIMEBOOST_net_1740;
wire g62465_sb;
wire TIMEBOOST_net_11412;
wire TIMEBOOST_net_13503;
wire g62466_sb;
wire TIMEBOOST_net_11413;
wire TIMEBOOST_net_14971;
wire g62467_sb;
wire TIMEBOOST_net_14672;
wire g62468_db;
wire g62468_sb;
wire TIMEBOOST_net_11537;
wire TIMEBOOST_net_14407;
wire g62469_sb;
wire TIMEBOOST_net_11414;
wire g57797_da;
wire g62470_sb;
wire TIMEBOOST_net_11415;
wire TIMEBOOST_net_13212;
wire g62471_sb;
wire TIMEBOOST_net_11538;
wire TIMEBOOST_net_14491;
wire g62472_sb;
wire TIMEBOOST_net_11539;
wire TIMEBOOST_net_14107;
wire g62473_sb;
wire TIMEBOOST_net_14159;
wire TIMEBOOST_net_11265;
wire g62474_sb;
wire TIMEBOOST_net_11540;
wire TIMEBOOST_net_14490;
wire g62475_sb;
wire n_3287;
wire TIMEBOOST_net_11266;
wire g62476_sb;
wire TIMEBOOST_net_11573;
wire TIMEBOOST_net_14308;
wire g62477_sb;
wire TIMEBOOST_net_11541;
wire TIMEBOOST_net_14472;
wire g62478_sb;
wire TIMEBOOST_net_10083;
wire TIMEBOOST_net_11223;
wire g62479_sb;
wire TIMEBOOST_net_11224;
wire g62480_sb;
wire TIMEBOOST_net_11522;
wire TIMEBOOST_net_13931;
wire g62481_sb;
wire TIMEBOOST_net_11416;
wire TIMEBOOST_net_14972;
wire g62482_sb;
wire TIMEBOOST_net_11417;
wire TIMEBOOST_net_1267;
wire g62483_sb;
wire TIMEBOOST_net_11529;
wire TIMEBOOST_net_13953;
wire g62484_sb;
wire TIMEBOOST_net_14493;
wire TIMEBOOST_net_14735;
wire g62485_sb;
wire TIMEBOOST_net_11733;
wire TIMEBOOST_net_14319;
wire g62486_sb;
wire TIMEBOOST_net_11418;
wire TIMEBOOST_net_14794;
wire g62487_sb;
wire TIMEBOOST_net_11419;
wire TIMEBOOST_net_13211;
wire g62488_sb;
wire TIMEBOOST_net_14155;
wire TIMEBOOST_net_11225;
wire g62489_sb;
wire TIMEBOOST_net_15061;
wire TIMEBOOST_net_11226;
wire g62490_sb;
wire TIMEBOOST_net_11542;
wire TIMEBOOST_net_14473;
wire g62491_sb;
wire TIMEBOOST_net_11420;
wire TIMEBOOST_net_1271;
wire g62492_sb;
wire TIMEBOOST_net_11543;
wire TIMEBOOST_net_1689;
wire g62493_sb;
wire TIMEBOOST_net_1558;
wire TIMEBOOST_net_11227;
wire g62494_sb;
wire TIMEBOOST_net_14382;
wire TIMEBOOST_net_11660;
wire g62495_sb;
wire TIMEBOOST_net_11421;
wire TIMEBOOST_net_12321;
wire g62496_sb;
wire TIMEBOOST_net_11422;
wire TIMEBOOST_net_1273;
wire g62497_sb;
wire TIMEBOOST_net_11737;
wire TIMEBOOST_net_13920;
wire g62498_sb;
wire TIMEBOOST_net_11423;
wire TIMEBOOST_net_9670;
wire g62499_sb;
wire TIMEBOOST_net_9944;
wire TIMEBOOST_net_11228;
wire g62500_sb;
wire TIMEBOOST_net_11740;
wire TIMEBOOST_net_13921;
wire g62501_sb;
wire TIMEBOOST_net_11424;
wire TIMEBOOST_net_15043;
wire g62502_sb;
wire TIMEBOOST_net_14393;
wire TIMEBOOST_net_11229;
wire g62503_sb;
wire TIMEBOOST_net_11741;
wire TIMEBOOST_net_14519;
wire g62504_sb;
wire TIMEBOOST_net_11425;
wire TIMEBOOST_net_14630;
wire g62505_sb;
wire TIMEBOOST_net_11426;
wire TIMEBOOST_net_14648;
wire g62506_sb;
wire TIMEBOOST_net_1561;
wire TIMEBOOST_net_11230;
wire g62507_sb;
wire TIMEBOOST_net_11427;
wire TIMEBOOST_net_14701;
wire g62508_sb;
wire TIMEBOOST_net_11428;
wire TIMEBOOST_net_13208;
wire g62509_sb;
wire TIMEBOOST_net_11429;
wire TIMEBOOST_net_14768;
wire g62510_sb;
wire TIMEBOOST_net_11544;
wire TIMEBOOST_net_14536;
wire g62511_sb;
wire TIMEBOOST_net_12249;
wire TIMEBOOST_net_11231;
wire g62512_sb;
wire TIMEBOOST_net_1563;
wire TIMEBOOST_net_11267;
wire g62513_sb;
wire TIMEBOOST_net_11430;
wire TIMEBOOST_net_14771;
wire g62514_sb;
wire TIMEBOOST_net_1564;
wire TIMEBOOST_net_11575;
wire g62515_sb;
wire TIMEBOOST_net_1565;
wire TIMEBOOST_net_11268;
wire g62516_sb;
wire TIMEBOOST_net_12253;
wire TIMEBOOST_net_11269;
wire g62517_sb;
wire TIMEBOOST_net_11745;
wire TIMEBOOST_net_14413;
wire g62518_sb;
wire TIMEBOOST_net_11749;
wire TIMEBOOST_net_14047;
wire g62519_sb;
wire TIMEBOOST_net_11746;
wire TIMEBOOST_net_14048;
wire g62520_sb;
wire TIMEBOOST_net_11431;
wire TIMEBOOST_net_14700;
wire g62521_sb;
wire TIMEBOOST_net_11432;
wire TIMEBOOST_net_13207;
wire g62522_sb;
wire TIMEBOOST_net_11601;
wire TIMEBOOST_net_14049;
wire g62523_sb;
wire TIMEBOOST_net_11433;
wire TIMEBOOST_net_15040;
wire g62524_sb;
wire TIMEBOOST_net_14388;
wire TIMEBOOST_net_11270;
wire g62525_sb;
wire TIMEBOOST_net_14293;
wire TIMEBOOST_net_11271;
wire g62526_sb;
wire TIMEBOOST_net_11434;
wire TIMEBOOST_net_14787;
wire g62527_sb;
wire TIMEBOOST_net_14147;
wire TIMEBOOST_net_14180;
wire g62528_sb;
wire TIMEBOOST_net_14450;
wire TIMEBOOST_net_11823;
wire g62529_sb;
wire TIMEBOOST_net_14198;
wire TIMEBOOST_net_11272;
wire g62530_sb;
wire TIMEBOOST_net_11435;
wire TIMEBOOST_net_14840;
wire g62531_sb;
wire TIMEBOOST_net_11545;
wire TIMEBOOST_net_10459;
wire g62532_sb;
wire TIMEBOOST_net_11546;
wire TIMEBOOST_net_14441;
wire g62533_sb;
wire TIMEBOOST_net_11547;
wire TIMEBOOST_net_14309;
wire g62534_sb;
wire TIMEBOOST_net_11612;
wire TIMEBOOST_net_14256;
wire g62535_sb;
wire TIMEBOOST_net_11436;
wire TIMEBOOST_net_14777;
wire g62536_sb;
wire TIMEBOOST_net_11437;
wire TIMEBOOST_net_14814;
wire g62537_sb;
wire TIMEBOOST_net_11438;
wire TIMEBOOST_net_14838;
wire g62538_sb;
wire TIMEBOOST_net_14226;
wire TIMEBOOST_net_11273;
wire g62539_sb;
wire TIMEBOOST_net_11548;
wire TIMEBOOST_net_13925;
wire g62540_sb;
wire TIMEBOOST_net_11439;
wire TIMEBOOST_net_14704;
wire g62541_sb;
wire TIMEBOOST_net_11440;
wire TIMEBOOST_net_14708;
wire g62542_sb;
wire TIMEBOOST_net_14227;
wire TIMEBOOST_net_11274;
wire g62543_sb;
wire TIMEBOOST_net_14420;
wire TIMEBOOST_net_11275;
wire g62544_sb;
wire TIMEBOOST_net_14228;
wire TIMEBOOST_net_11276;
wire g62545_sb;
wire TIMEBOOST_net_11441;
wire TIMEBOOST_net_14893;
wire g62546_sb;
wire TIMEBOOST_net_11584;
wire TIMEBOOST_net_14411;
wire g62547_sb;
wire TIMEBOOST_net_11442;
wire TIMEBOOST_net_14769;
wire g62548_sb;
wire TIMEBOOST_net_11443;
wire TIMEBOOST_net_1294;
wire g62549_sb;
wire TIMEBOOST_net_11549;
wire TIMEBOOST_net_10455;
wire g62550_sb;
wire TIMEBOOST_net_14229;
wire TIMEBOOST_net_11277;
wire g62551_sb;
wire TIMEBOOST_net_14230;
wire TIMEBOOST_net_11278;
wire g62552_sb;
wire TIMEBOOST_net_11550;
wire TIMEBOOST_net_13958;
wire g62553_sb;
wire TIMEBOOST_net_11202;
wire TIMEBOOST_net_1295;
wire g62554_sb;
wire TIMEBOOST_net_11447;
wire TIMEBOOST_net_1296;
wire g62555_sb;
wire TIMEBOOST_net_14231;
wire TIMEBOOST_net_11279;
wire g62556_sb;
wire TIMEBOOST_net_14246;
wire TIMEBOOST_net_11280;
wire g62557_sb;
wire TIMEBOOST_net_11595;
wire TIMEBOOST_net_14006;
wire g62558_sb;
wire TIMEBOOST_net_14247;
wire TIMEBOOST_net_13359;
wire g62559_sb;
wire TIMEBOOST_net_11596;
wire TIMEBOOST_net_14051;
wire g62560_sb;
wire TIMEBOOST_net_11674;
wire TIMEBOOST_net_14326;
wire g62561_sb;
wire TIMEBOOST_net_11675;
wire TIMEBOOST_net_13945;
wire g62562_sb;
wire TIMEBOOST_net_11559;
wire TIMEBOOST_net_14602;
wire g62563_sb;
wire TIMEBOOST_net_14312;
wire TIMEBOOST_net_11281;
wire g62564_sb;
wire TIMEBOOST_net_11341;
wire TIMEBOOST_net_1297;
wire g62565_sb;
wire TIMEBOOST_net_11451;
wire TIMEBOOST_net_1298;
wire g62566_sb;
wire TIMEBOOST_net_14562;
wire TIMEBOOST_net_11282;
wire g62567_sb;
wire TIMEBOOST_net_11448;
wire TIMEBOOST_net_14856;
wire g62568_sb;
wire TIMEBOOST_net_11677;
wire TIMEBOOST_net_14520;
wire g62569_sb;
wire TIMEBOOST_net_11566;
wire TIMEBOOST_net_14263;
wire g62570_sb;
wire TIMEBOOST_net_11678;
wire TIMEBOOST_net_14010;
wire g62571_sb;
wire TIMEBOOST_net_11452;
wire TIMEBOOST_net_1300;
wire g62572_sb;
wire TIMEBOOST_net_11453;
wire TIMEBOOST_net_1301;
wire g62573_sb;
wire TIMEBOOST_net_11454;
wire TIMEBOOST_net_1302;
wire g62574_sb;
wire TIMEBOOST_net_14264;
wire g62575_db;
wire g62575_sb;
wire TIMEBOOST_net_11679;
wire TIMEBOOST_net_13959;
wire g62576_sb;
wire TIMEBOOST_net_11455;
wire TIMEBOOST_net_1303;
wire g62577_sb;
wire TIMEBOOST_net_11450;
wire TIMEBOOST_net_14859;
wire g62578_sb;
wire TIMEBOOST_net_5574;
wire TIMEBOOST_net_14826;
wire g62579_sb;
wire TIMEBOOST_net_14466;
wire TIMEBOOST_net_11283;
wire g62580_sb;
wire TIMEBOOST_net_14254;
wire TIMEBOOST_net_11284;
wire g62581_sb;
wire TIMEBOOST_net_14315;
wire TIMEBOOST_net_11285;
wire g62582_sb;
wire TIMEBOOST_net_14262;
wire TIMEBOOST_net_11286;
wire g62583_sb;
wire TIMEBOOST_net_11459;
wire TIMEBOOST_net_14845;
wire g62584_sb;
wire TIMEBOOST_net_11456;
wire TIMEBOOST_net_1307;
wire g62585_sb;
wire TIMEBOOST_net_11457;
wire TIMEBOOST_net_1308;
wire g62586_sb;
wire TIMEBOOST_net_14222;
wire TIMEBOOST_net_11287;
wire g62587_sb;
wire TIMEBOOST_net_11567;
wire TIMEBOOST_net_13948;
wire g62588_sb;
wire TIMEBOOST_net_14223;
wire TIMEBOOST_net_11288;
wire g62589_sb;
wire TIMEBOOST_net_11471;
wire TIMEBOOST_net_1309;
wire g62590_sb;
wire TIMEBOOST_net_11460;
wire TIMEBOOST_net_15009;
wire g62591_sb;
wire TIMEBOOST_net_14235;
wire TIMEBOOST_net_11597;
wire g62592_sb;
wire TIMEBOOST_net_11680;
wire TIMEBOOST_net_14529;
wire g62593_sb;
wire TIMEBOOST_net_11461;
wire TIMEBOOST_net_15005;
wire g62594_sb;
wire g62595_p;
wire TIMEBOOST_net_11462;
wire TIMEBOOST_net_15008;
wire g62596_sb;
wire TIMEBOOST_net_11463;
wire TIMEBOOST_net_1313;
wire g62597_sb;
wire TIMEBOOST_net_11464;
wire TIMEBOOST_net_1314;
wire g62598_sb;
wire TIMEBOOST_net_11681;
wire TIMEBOOST_net_14125;
wire g62599_sb;
wire TIMEBOOST_net_11671;
wire TIMEBOOST_net_14427;
wire g62600_sb;
wire TIMEBOOST_net_11738;
wire TIMEBOOST_net_10470;
wire g62601_sb;
wire TIMEBOOST_net_11465;
wire TIMEBOOST_net_1315;
wire g62602_sb;
wire TIMEBOOST_net_11466;
wire TIMEBOOST_net_1316;
wire g62603_sb;
wire TIMEBOOST_net_11467;
wire TIMEBOOST_net_15046;
wire g62604_sb;
wire TIMEBOOST_net_14217;
wire TIMEBOOST_net_11289;
wire g62605_sb;
wire TIMEBOOST_net_11766;
wire TIMEBOOST_net_14106;
wire g62606_sb;
wire TIMEBOOST_net_14919;
wire g62607_db;
wire g62607_sb;
wire TIMEBOOST_net_11468;
wire TIMEBOOST_net_14870;
wire g62608_sb;
wire TIMEBOOST_net_11469;
wire TIMEBOOST_net_14786;
wire g62609_sb;
wire TIMEBOOST_net_11470;
wire TIMEBOOST_net_14863;
wire g62610_sb;
wire TIMEBOOST_net_14313;
wire TIMEBOOST_net_11290;
wire g62611_sb;
wire TIMEBOOST_net_11686;
wire TIMEBOOST_net_14090;
wire g62612_sb;
wire TIMEBOOST_net_5590;
wire TIMEBOOST_net_14658;
wire g62613_sb;
wire TIMEBOOST_net_11500;
wire TIMEBOOST_net_10458;
wire g62614_sb;
wire TIMEBOOST_net_14209;
wire TIMEBOOST_net_11291;
wire g62615_sb;
wire TIMEBOOST_net_11473;
wire TIMEBOOST_net_14657;
wire g62616_sb;
wire TIMEBOOST_net_10830;
wire TIMEBOOST_net_14877;
wire g62617_sb;
wire TIMEBOOST_net_11604;
wire TIMEBOOST_net_14439;
wire g62618_sb;
wire TIMEBOOST_net_11517;
wire TIMEBOOST_net_12915;
wire g62619_sb;
wire TIMEBOOST_net_14210;
wire TIMEBOOST_net_11292;
wire g62620_sb;
wire TIMEBOOST_net_10831;
wire TIMEBOOST_net_14788;
wire g62621_sb;
wire TIMEBOOST_net_11614;
wire TIMEBOOST_net_14069;
wire g62622_sb;
wire TIMEBOOST_net_11520;
wire TIMEBOOST_net_14110;
wire g62623_sb;
wire TIMEBOOST_net_11474;
wire TIMEBOOST_net_1447;
wire g62624_sb;
wire TIMEBOOST_net_11521;
wire TIMEBOOST_net_14113;
wire g62625_sb;
wire TIMEBOOST_net_11534;
wire TIMEBOOST_net_14116;
wire g62626_sb;
wire TIMEBOOST_net_13962;
wire TIMEBOOST_net_11583;
wire g62627_sb;
wire TIMEBOOST_net_14211;
wire TIMEBOOST_net_11574;
wire g62628_sb;
wire TIMEBOOST_net_11195;
wire TIMEBOOST_net_12911;
wire g62629_sb;
wire TIMEBOOST_net_11535;
wire TIMEBOOST_net_14202;
wire g62630_sb;
wire TIMEBOOST_net_11449;
wire TIMEBOOST_net_14852;
wire g62631_sb;
wire TIMEBOOST_net_11496;
wire TIMEBOOST_net_14205;
wire g62632_sb;
wire TIMEBOOST_net_11618;
wire TIMEBOOST_net_13936;
wire g62633_sb;
wire TIMEBOOST_net_14455;
wire TIMEBOOST_net_11293;
wire g62634_sb;
wire TIMEBOOST_net_11622;
wire TIMEBOOST_net_13926;
wire g62635_sb;
wire TIMEBOOST_net_11630;
wire TIMEBOOST_net_13968;
wire g62636_sb;
wire TIMEBOOST_net_10373;
wire TIMEBOOST_net_14615;
wire g62637_sb;
wire TIMEBOOST_net_14236;
wire TIMEBOOST_net_11351;
wire g62638_sb;
wire TIMEBOOST_net_5598;
wire TIMEBOOST_net_14616;
wire g62639_sb;
wire TIMEBOOST_net_14570;
wire TIMEBOOST_net_11352;
wire g62640_sb;
wire n_3483;
wire TIMEBOOST_net_11294;
wire g62641_sb;
wire TIMEBOOST_net_11476;
wire TIMEBOOST_net_14610;
wire g62642_sb;
wire TIMEBOOST_net_11477;
wire TIMEBOOST_net_14996;
wire g62643_sb;
wire TIMEBOOST_net_11497;
wire TIMEBOOST_net_1755;
wire g62644_sb;
wire TIMEBOOST_net_14273;
wire TIMEBOOST_net_11353;
wire g62645_sb;
wire TIMEBOOST_net_11533;
wire TIMEBOOST_net_14117;
wire g62646_sb;
wire TIMEBOOST_net_11570;
wire TIMEBOOST_net_14316;
wire g62647_sb;
wire TIMEBOOST_net_14271;
wire TIMEBOOST_net_11295;
wire g62648_sb;
wire TIMEBOOST_net_14268;
wire TIMEBOOST_net_14516;
wire g62649_sb;
wire TIMEBOOST_net_14269;
wire TIMEBOOST_net_11296;
wire g62650_sb;
wire TIMEBOOST_net_11478;
wire TIMEBOOST_net_14874;
wire g62651_sb;
wire TIMEBOOST_net_11479;
wire TIMEBOOST_net_13505;
wire g62652_sb;
wire TIMEBOOST_net_14522;
wire TIMEBOOST_net_11297;
wire g62653_sb;
wire TIMEBOOST_net_11571;
wire TIMEBOOST_net_14215;
wire g62654_sb;
wire TIMEBOOST_net_11576;
wire TIMEBOOST_net_14216;
wire g62655_sb;
wire TIMEBOOST_net_11577;
wire TIMEBOOST_net_14764;
wire g62656_sb;
wire TIMEBOOST_net_11480;
wire TIMEBOOST_net_14802;
wire g62657_sb;
wire TIMEBOOST_net_11481;
wire TIMEBOOST_net_14778;
wire g62658_sb;
wire TIMEBOOST_net_11482;
wire TIMEBOOST_net_14867;
wire g62659_sb;
wire TIMEBOOST_net_11682;
wire TIMEBOOST_net_14114;
wire g62660_sb;
wire TIMEBOOST_net_11203;
wire TIMEBOOST_net_14865;
wire g62661_sb;
wire TIMEBOOST_net_14052;
wire TIMEBOOST_net_11826;
wire g62662_sb;
wire TIMEBOOST_net_11683;
wire TIMEBOOST_net_5235;
wire g62663_sb;
wire TIMEBOOST_net_11578;
wire TIMEBOOST_net_14214;
wire g62664_sb;
wire TIMEBOOST_net_11204;
wire TIMEBOOST_net_14746;
wire g62665_sb;
wire TIMEBOOST_net_11684;
wire TIMEBOOST_net_13975;
wire g62666_sb;
wire TIMEBOOST_net_11205;
wire TIMEBOOST_net_14747;
wire g62667_sb;
wire TIMEBOOST_net_14626;
wire TIMEBOOST_net_14803;
wire g62668_sb;
wire TIMEBOOST_net_14213;
wire TIMEBOOST_net_11298;
wire g62669_sb;
wire TIMEBOOST_net_14625;
wire TIMEBOOST_net_14773;
wire g62670_sb;
wire TIMEBOOST_net_14624;
wire TIMEBOOST_net_14869;
wire g62671_sb;
wire TIMEBOOST_net_14623;
wire TIMEBOOST_net_14946;
wire g62672_sb;
wire TIMEBOOST_net_11685;
wire TIMEBOOST_net_13974;
wire g62673_sb;
wire TIMEBOOST_net_11488;
wire TIMEBOOST_net_15016;
wire g62674_sb;
wire TIMEBOOST_net_14174;
wire TIMEBOOST_net_10494;
wire g62675_sb;
wire TIMEBOOST_net_14622;
wire TIMEBOOST_net_14690;
wire g62676_sb;
wire TIMEBOOST_net_11631;
wire TIMEBOOST_net_14266;
wire g62677_sb;
wire TIMEBOOST_net_11844;
wire TIMEBOOST_net_1425;
wire g62678_sb;
wire TIMEBOOST_net_11834;
wire TIMEBOOST_net_9306;
wire g62679_sb;
wire TIMEBOOST_net_11845;
wire TIMEBOOST_net_14761;
wire g62680_sb;
wire TIMEBOOST_net_11485;
wire TIMEBOOST_net_15018;
wire g62681_sb;
wire TIMEBOOST_net_11486;
wire TIMEBOOST_net_15023;
wire g62682_sb;
wire TIMEBOOST_net_14172;
wire TIMEBOOST_net_11299;
wire g62683_sb;
wire TIMEBOOST_net_11487;
wire TIMEBOOST_net_14926;
wire g62684_sb;
wire TIMEBOOST_net_11853;
wire TIMEBOOST_net_14927;
wire g62685_sb;
wire TIMEBOOST_net_14056;
wire TIMEBOOST_net_11827;
wire g62688_sb;
wire TIMEBOOST_net_11854;
wire TIMEBOOST_net_14932;
wire g62689_sb;
wire TIMEBOOST_net_14324;
wire TIMEBOOST_net_11811;
wire g62690_sb;
wire TIMEBOOST_net_11916;
wire TIMEBOOST_net_14608;
wire g62691_sb;
wire TIMEBOOST_net_11855;
wire TIMEBOOST_net_14677;
wire g62693_sb;
wire TIMEBOOST_net_11835;
wire TIMEBOOST_net_14140;
wire g62697_sb;
wire TIMEBOOST_net_11856;
wire TIMEBOOST_net_14944;
wire g62698_sb;
wire g62699_p;
wire TIMEBOOST_net_11836;
wire TIMEBOOST_net_1760;
wire g62701_sb;
wire TIMEBOOST_net_11857;
wire TIMEBOOST_net_15019;
wire g62706_sb;
wire TIMEBOOST_net_14239;
wire TIMEBOOST_net_11300;
wire g62707_sb;
wire TIMEBOOST_net_11858;
wire TIMEBOOST_net_15024;
wire g62710_sb;
wire TIMEBOOST_net_11860;
wire TIMEBOOST_net_14864;
wire g62711_sb;
wire TIMEBOOST_net_14224;
wire TIMEBOOST_net_11301;
wire g62712_sb;
wire TIMEBOOST_net_11861;
wire TIMEBOOST_net_14804;
wire g62713_sb;
wire TIMEBOOST_net_11495;
wire TIMEBOOST_net_14810;
wire g62714_sb;
wire TIMEBOOST_net_11774;
wire TIMEBOOST_net_14743;
wire g62715_sb;
wire TIMEBOOST_net_9349;
wire TIMEBOOST_net_10710;
wire g62716_sb;
wire TIMEBOOST_net_14238;
wire g62719_db;
wire g62719_sb;
wire TIMEBOOST_net_9452;
wire TIMEBOOST_net_13349;
wire g62720_sb;
wire TIMEBOOST_net_12356;
wire TIMEBOOST_net_4905;
wire g62721_sb;
wire TIMEBOOST_net_11040;
wire TIMEBOOST_net_14042;
wire g62722_sb;
wire TIMEBOOST_net_12398;
wire TIMEBOOST_net_4906;
wire g62723_sb;
wire TIMEBOOST_net_10874;
wire g62724_db;
wire TIMEBOOST_net_11042;
wire g64752_db;
wire g62725_sb;
wire TIMEBOOST_net_12337;
wire TIMEBOOST_net_13989;
wire g62726_sb;
wire TIMEBOOST_net_12331;
wire TIMEBOOST_net_4907;
wire g62727_sb;
wire TIMEBOOST_net_11043;
wire TIMEBOOST_net_14017;
wire g62728_sb;
wire TIMEBOOST_net_13780;
wire TIMEBOOST_net_4908;
wire g62729_sb;
wire TIMEBOOST_net_925;
wire TIMEBOOST_net_4909;
wire g62730_sb;
wire TIMEBOOST_net_9355;
wire TIMEBOOST_net_767;
wire g62731_sb;
wire TIMEBOOST_net_10819;
wire TIMEBOOST_net_4910;
wire g62732_sb;
wire TIMEBOOST_net_15245;
wire TIMEBOOST_net_12838;
wire g62733_sb;
wire TIMEBOOST_net_724;
wire g62734_db;
wire g62734_sb;
wire TIMEBOOST_net_4569;
wire TIMEBOOST_net_4911;
wire g62735_sb;
wire TIMEBOOST_net_12720;
wire TIMEBOOST_net_4912;
wire g62736_sb;
wire TIMEBOOST_net_13629;
wire TIMEBOOST_net_4913;
wire g62737_sb;
wire TIMEBOOST_net_13781;
wire g62738_db;
wire g62738_sb;
wire TIMEBOOST_net_5194;
wire TIMEBOOST_net_768;
wire g62739_sb;
wire TIMEBOOST_net_10647;
wire TIMEBOOST_net_13907;
wire g62740_sb;
wire TIMEBOOST_net_14537;
wire TIMEBOOST_net_13913;
wire g62741_sb;
wire TIMEBOOST_net_11064;
wire TIMEBOOST_net_13192;
wire g62742_sb;
wire TIMEBOOST_net_11065;
wire TIMEBOOST_net_13193;
wire g62743_sb;
wire TIMEBOOST_net_933;
wire TIMEBOOST_net_4916;
wire g62744_sb;
wire TIMEBOOST_net_4571;
wire TIMEBOOST_net_4917;
wire g62745_sb;
wire TIMEBOOST_net_12986;
wire TIMEBOOST_net_4918;
wire g62746_sb;
wire TIMEBOOST_net_10652;
wire TIMEBOOST_net_4919;
wire g62747_sb;
wire TIMEBOOST_net_4661;
wire TIMEBOOST_net_14173;
wire g62748_sb;
wire TIMEBOOST_net_937;
wire TIMEBOOST_net_13912;
wire g62749_sb;
wire TIMEBOOST_net_938;
wire TIMEBOOST_net_4922;
wire g62750_sb;
wire TIMEBOOST_net_939;
wire TIMEBOOST_net_10825;
wire g62751_sb;
wire TIMEBOOST_net_11066;
wire TIMEBOOST_net_9592;
wire g62752_sb;
wire TIMEBOOST_net_11068;
wire TIMEBOOST_net_14150;
wire g62753_sb;
wire TIMEBOOST_net_11831;
wire TIMEBOOST_net_14694;
wire g62754_sb;
wire TIMEBOOST_net_11837;
wire TIMEBOOST_net_14905;
wire g62755_sb;
wire TIMEBOOST_net_4924;
wire g62756_sb;
wire TIMEBOOST_net_626;
wire TIMEBOOST_net_10771;
wire g62757_sb;
wire TIMEBOOST_net_11581;
wire TIMEBOOST_net_14044;
wire g62758_sb;
wire TIMEBOOST_net_4662;
wire TIMEBOOST_net_13911;
wire g62759_sb;
wire TIMEBOOST_net_11695;
wire TIMEBOOST_net_14854;
wire g62760_sb;
wire TIMEBOOST_net_11704;
wire TIMEBOOST_net_15197;
wire g62761_sb;
wire TIMEBOOST_net_3891;
wire TIMEBOOST_net_4927;
wire g62762_sb;
wire TIMEBOOST_net_11532;
wire TIMEBOOST_net_14186;
wire g62763_sb;
wire TIMEBOOST_net_13881;
wire TIMEBOOST_net_10826;
wire g62764_sb;
wire TIMEBOOST_net_944;
wire TIMEBOOST_net_14580;
wire g62765_sb;
wire TIMEBOOST_net_10696;
wire TIMEBOOST_net_10772;
wire g62766_sb;
wire TIMEBOOST_net_4664;
wire TIMEBOOST_net_4931;
wire g62767_sb;
wire TIMEBOOST_net_4665;
wire TIMEBOOST_net_13910;
wire g62768_sb;
wire TIMEBOOST_net_10697;
wire TIMEBOOST_net_4933;
wire g62769_sb;
wire TIMEBOOST_net_4573;
wire TIMEBOOST_net_4934;
wire g62770_sb;
wire TIMEBOOST_net_10654;
wire TIMEBOOST_net_4935;
wire g62771_sb;
wire TIMEBOOST_net_10698;
wire TIMEBOOST_net_4936;
wire g62772_sb;
wire TIMEBOOST_net_627;
wire TIMEBOOST_net_13350;
wire g62773_sb;
wire TIMEBOOST_net_9356;
wire TIMEBOOST_net_773;
wire g62774_sb;
wire TIMEBOOST_net_13564;
wire TIMEBOOST_net_4937;
wire g62775_sb;
wire TIMEBOOST_net_4575;
wire TIMEBOOST_net_10904;
wire g62776_sb;
wire TIMEBOOST_net_11335;
wire g62777_db;
wire g62777_sb;
wire TIMEBOOST_net_4668;
wire TIMEBOOST_net_10920;
wire g62778_sb;
wire TIMEBOOST_net_4669;
wire TIMEBOOST_net_10921;
wire g62779_sb;
wire n_14750;
wire g62780_db;
wire g62780_sb;
wire TIMEBOOST_net_10699;
wire TIMEBOOST_net_10922;
wire g62781_sb;
wire TIMEBOOST_net_4576;
wire TIMEBOOST_net_10923;
wire g62782_sb;
wire TIMEBOOST_net_11838;
wire g62783_db;
wire g62783_sb;
wire TIMEBOOST_net_4671;
wire TIMEBOOST_net_10926;
wire g62784_sb;
wire TIMEBOOST_net_11069;
wire TIMEBOOST_net_12702;
wire g62785_sb;
wire TIMEBOOST_net_4672;
wire TIMEBOOST_net_10927;
wire g62786_sb;
wire TIMEBOOST_net_960;
wire TIMEBOOST_net_10928;
wire g62787_sb;
wire TIMEBOOST_net_10700;
wire TIMEBOOST_net_10930;
wire g62788_sb;
wire TIMEBOOST_net_12988;
wire TIMEBOOST_net_10935;
wire g62789_sb;
wire TIMEBOOST_net_10701;
wire TIMEBOOST_net_10958;
wire g62790_sb;
wire TIMEBOOST_net_963;
wire g62791_db;
wire g62791_sb;
wire TIMEBOOST_net_10959;
wire g62792_sb;
wire TIMEBOOST_net_15174;
wire TIMEBOOST_net_10960;
wire g62793_sb;
wire TIMEBOOST_net_15088;
wire TIMEBOOST_net_10961;
wire g62794_sb;
wire TIMEBOOST_net_10962;
wire g62795_sb;
wire TIMEBOOST_net_968;
wire TIMEBOOST_net_10963;
wire g62796_sb;
wire TIMEBOOST_net_15097;
wire TIMEBOOST_net_10964;
wire g62797_sb;
wire TIMEBOOST_net_10734;
wire TIMEBOOST_net_775;
wire TIMEBOOST_net_630;
wire g62799_db;
wire g62799_sb;
wire TIMEBOOST_net_10965;
wire g62800_sb;
wire TIMEBOOST_net_11070;
wire TIMEBOOST_net_776;
wire g62801_sb;
wire TIMEBOOST_net_11071;
wire TIMEBOOST_net_777;
wire g62802_sb;
wire TIMEBOOST_net_971;
wire g62803_db;
wire g62803_sb;
wire TIMEBOOST_net_4894;
wire TIMEBOOST_net_778;
wire TIMEBOOST_net_14329;
wire TIMEBOOST_net_10966;
wire g62805_sb;
wire TIMEBOOST_net_972;
wire TIMEBOOST_net_10967;
wire g62806_sb;
wire TIMEBOOST_net_11408;
wire g62807_db;
wire g62807_sb;
wire TIMEBOOST_net_10735;
wire g62808_db;
wire g62808_sb;
wire TIMEBOOST_net_11072;
wire TIMEBOOST_net_12760;
wire g62809_sb;
wire TIMEBOOST_net_973;
wire TIMEBOOST_net_10968;
wire g62810_sb;
wire TIMEBOOST_net_13783;
wire g62811_db;
wire g62811_sb;
wire TIMEBOOST_net_974;
wire TIMEBOOST_net_10969;
wire g62812_sb;
wire TIMEBOOST_net_975;
wire TIMEBOOST_net_14109;
wire g62813_sb;
wire TIMEBOOST_net_976;
wire TIMEBOOST_net_14533;
wire g62814_sb;
wire TIMEBOOST_net_977;
wire TIMEBOOST_net_10970;
wire g62815_sb;
wire TIMEBOOST_net_978;
wire TIMEBOOST_net_10971;
wire g62816_sb;
wire TIMEBOOST_net_11073;
wire TIMEBOOST_net_780;
wire g62817_sb;
wire TIMEBOOST_net_979;
wire TIMEBOOST_net_10972;
wire g62818_sb;
wire TIMEBOOST_net_980;
wire TIMEBOOST_net_10973;
wire g62819_sb;
wire TIMEBOOST_net_981;
wire TIMEBOOST_net_10974;
wire g62820_sb;
wire TIMEBOOST_net_13312;
wire g62821_db;
wire g62821_sb;
wire TIMEBOOST_net_982;
wire TIMEBOOST_net_10975;
wire g62822_sb;
wire TIMEBOOST_net_983;
wire TIMEBOOST_net_10976;
wire g62823_sb;
wire TIMEBOOST_net_984;
wire TIMEBOOST_net_10977;
wire g62824_sb;
wire TIMEBOOST_net_985;
wire TIMEBOOST_net_11025;
wire g62825_sb;
wire TIMEBOOST_net_11074;
wire TIMEBOOST_net_781;
wire g62826_sb;
wire TIMEBOOST_net_11075;
wire TIMEBOOST_net_12707;
wire g62827_sb;
wire TIMEBOOST_net_11076;
wire n_3427;
wire g62828_sb;
wire TIMEBOOST_net_986;
wire TIMEBOOST_net_11027;
wire g62829_sb;
wire TIMEBOOST_net_11077;
wire TIMEBOOST_net_784;
wire g62830_sb;
wire TIMEBOOST_net_987;
wire TIMEBOOST_net_11044;
wire g62831_sb;
wire TIMEBOOST_net_988;
wire TIMEBOOST_net_11045;
wire g62832_sb;
wire TIMEBOOST_net_989;
wire g62833_db;
wire g62833_sb;
wire TIMEBOOST_net_990;
wire TIMEBOOST_net_11046;
wire g62834_sb;
wire TIMEBOOST_net_10745;
wire g62835_db;
wire g62835_sb;
wire TIMEBOOST_net_11078;
wire TIMEBOOST_net_14866;
wire g62836_sb;
wire TIMEBOOST_net_11079;
wire TIMEBOOST_net_12357;
wire g62837_sb;
wire TIMEBOOST_net_991;
wire TIMEBOOST_net_11047;
wire g62838_sb;
wire TIMEBOOST_net_992;
wire TIMEBOOST_net_11048;
wire g62839_sb;
wire TIMEBOOST_net_993;
wire TIMEBOOST_net_11049;
wire g62840_sb;
wire TIMEBOOST_net_994;
wire TIMEBOOST_net_11050;
wire g62841_sb;
wire TIMEBOOST_net_5210;
wire TIMEBOOST_net_787;
wire g62842_sb;
wire TIMEBOOST_net_6448;
wire g62843_db;
wire g62843_sb;
wire TIMEBOOST_net_634;
wire g62844_db;
wire g62844_sb;
wire TIMEBOOST_net_995;
wire TIMEBOOST_net_11051;
wire g62845_sb;
wire TIMEBOOST_net_996;
wire TIMEBOOST_net_11052;
wire g62846_sb;
wire TIMEBOOST_net_15045;
wire TIMEBOOST_net_11053;
wire g62847_sb;
wire TIMEBOOST_net_725;
wire g62848_db;
wire g62848_sb;
wire TIMEBOOST_net_14850;
wire TIMEBOOST_net_11054;
wire g62849_sb;
wire TIMEBOOST_net_14887;
wire TIMEBOOST_net_11055;
wire g62850_sb;
wire TIMEBOOST_net_635;
wire TIMEBOOST_net_11056;
wire g62851_sb;
wire TIMEBOOST_net_726;
wire g62852_db;
wire g62852_sb;
wire TIMEBOOST_net_11080;
wire TIMEBOOST_net_788;
wire g62853_sb;
wire TIMEBOOST_net_14660;
wire TIMEBOOST_net_11057;
wire g62854_sb;
wire TIMEBOOST_net_14889;
wire TIMEBOOST_net_11058;
wire g62855_sb;
wire TIMEBOOST_net_15012;
wire TIMEBOOST_net_11059;
wire g62856_sb;
wire TIMEBOOST_net_14760;
wire TIMEBOOST_net_11060;
wire g62857_sb;
wire TIMEBOOST_net_636;
wire g62858_db;
wire g62858_sb;
wire TIMEBOOST_net_13782;
wire g62859_db;
wire g62859_sb;
wire TIMEBOOST_net_14882;
wire TIMEBOOST_net_11061;
wire g62860_sb;
wire TIMEBOOST_net_11082;
wire TIMEBOOST_net_14643;
wire g62861_sb;
wire TIMEBOOST_net_1005;
wire TIMEBOOST_net_11062;
wire g62862_sb;
wire TIMEBOOST_net_1006;
wire TIMEBOOST_net_11063;
wire g62863_sb;
wire TIMEBOOST_net_1007;
wire g62864_db;
wire g62864_sb;
wire TIMEBOOST_net_1008;
wire TIMEBOOST_net_11067;
wire g62865_sb;
wire g62873_p;
wire g62874_p;
wire g62875_p;
wire g62876_p;
wire g62877_p;
wire g62879_p;
wire g62880_p;
wire g62881_p;
wire g62882_p;
wire TIMEBOOST_net_14250;
wire TIMEBOOST_net_11232;
wire g62883_sb;
wire TIMEBOOST_net_11864;
wire TIMEBOOST_net_14902;
wire g62884_sb;
wire TIMEBOOST_net_11582;
wire TIMEBOOST_net_14132;
wire g62885_sb;
wire TIMEBOOST_net_11703;
wire TIMEBOOST_net_14918;
wire g62886_sb;
wire TIMEBOOST_net_11708;
wire TIMEBOOST_net_14955;
wire g62887_sb;
wire TIMEBOOST_net_11863;
wire TIMEBOOST_net_14995;
wire g62888_sb;
wire TIMEBOOST_net_11868;
wire TIMEBOOST_net_14872;
wire g62889_sb;
wire TIMEBOOST_net_11869;
wire TIMEBOOST_net_15000;
wire g62890_sb;
wire TIMEBOOST_net_14604;
wire TIMEBOOST_net_11233;
wire g62891_sb;
wire TIMEBOOST_net_11870;
wire TIMEBOOST_net_15001;
wire g62892_sb;
wire TIMEBOOST_net_14577;
wire TIMEBOOST_net_11302;
wire g62893_sb;
wire TIMEBOOST_net_14573;
wire TIMEBOOST_net_11234;
wire g62894_sb;
wire TIMEBOOST_net_11871;
wire TIMEBOOST_net_15002;
wire g62895_sb;
wire TIMEBOOST_net_11752;
wire TIMEBOOST_net_14945;
wire g62896_sb;
wire TIMEBOOST_net_11757;
wire TIMEBOOST_net_15025;
wire g62897_sb;
wire TIMEBOOST_net_11590;
wire TIMEBOOST_net_14092;
wire g62898_sb;
wire TIMEBOOST_net_11519;
wire TIMEBOOST_net_15192;
wire g62899_sb;
wire TIMEBOOST_net_14290;
wire TIMEBOOST_net_11235;
wire g62900_sb;
wire TIMEBOOST_net_11593;
wire TIMEBOOST_net_14004;
wire g62901_sb;
wire TIMEBOOST_net_11598;
wire TIMEBOOST_net_14126;
wire g62902_sb;
wire TIMEBOOST_net_11475;
wire TIMEBOOST_net_14632;
wire g62903_sb;
wire TIMEBOOST_net_14201;
wire TIMEBOOST_net_11303;
wire g62904_sb;
wire TIMEBOOST_net_11490;
wire TIMEBOOST_net_14465;
wire g62905_sb;
wire TIMEBOOST_net_11592;
wire TIMEBOOST_net_14351;
wire g62906_sb;
wire TIMEBOOST_net_14237;
wire TIMEBOOST_net_11304;
wire g62907_sb;
wire TIMEBOOST_net_11792;
wire TIMEBOOST_net_14855;
wire g62908_sb;
wire TIMEBOOST_net_14102;
wire TIMEBOOST_net_11828;
wire g62909_sb;
wire TIMEBOOST_net_14276;
wire TIMEBOOST_net_11305;
wire g62910_sb;
wire TIMEBOOST_net_11489;
wire TIMEBOOST_net_14267;
wire g62911_sb;
wire TIMEBOOST_net_11585;
wire TIMEBOOST_net_14396;
wire g62912_sb;
wire TIMEBOOST_net_11793;
wire TIMEBOOST_net_15050;
wire g62913_sb;
wire TIMEBOOST_net_14575;
wire TIMEBOOST_net_11306;
wire g62914_sb;
wire TIMEBOOST_net_11794;
wire TIMEBOOST_net_13500;
wire g62915_sb;
wire TIMEBOOST_net_14561;
wire TIMEBOOST_net_11307;
wire g62916_sb;
wire TIMEBOOST_net_14225;
wire TIMEBOOST_net_11308;
wire g62917_sb;
wire TIMEBOOST_net_14458;
wire TIMEBOOST_net_11309;
wire g62918_sb;
wire TIMEBOOST_net_11635;
wire TIMEBOOST_net_13949;
wire g62919_sb;
wire TIMEBOOST_net_14534;
wire TIMEBOOST_net_11310;
wire g62920_sb;
wire TIMEBOOST_net_11579;
wire TIMEBOOST_net_10384;
wire g62921_sb;
wire TIMEBOOST_net_11795;
wire TIMEBOOST_net_14952;
wire g62922_sb;
wire TIMEBOOST_net_14339;
wire TIMEBOOST_net_11311;
wire g62923_sb;
wire TIMEBOOST_net_11632;
wire TIMEBOOST_net_10386;
wire g62924_sb;
wire TIMEBOOST_net_14526;
wire g62925_db;
wire g62925_sb;
wire TIMEBOOST_net_11638;
wire TIMEBOOST_net_14361;
wire g62926_sb;
wire TIMEBOOST_net_11796;
wire TIMEBOOST_net_1369;
wire g62927_sb;
wire TIMEBOOST_net_14474;
wire TIMEBOOST_net_11312;
wire g62928_sb;
wire TIMEBOOST_net_14544;
wire TIMEBOOST_net_11313;
wire g62929_sb;
wire TIMEBOOST_net_11797;
wire TIMEBOOST_net_14767;
wire g62930_sb;
wire TIMEBOOST_net_11754;
wire TIMEBOOST_net_14908;
wire g62931_sb;
wire TIMEBOOST_net_11833;
wire TIMEBOOST_net_14611;
wire g62932_sb;
wire TIMEBOOST_net_14272;
wire TIMEBOOST_net_11314;
wire g62933_sb;
wire TIMEBOOST_net_14270;
wire TIMEBOOST_net_11236;
wire g62934_sb;
wire TIMEBOOST_net_10174;
wire TIMEBOOST_net_11237;
wire g62935_sb;
wire TIMEBOOST_net_11720;
wire TIMEBOOST_net_14909;
wire g62936_sb;
wire TIMEBOOST_net_10154;
wire TIMEBOOST_net_11238;
wire g62937_sb;
wire TIMEBOOST_net_11755;
wire TIMEBOOST_net_14912;
wire g62938_sb;
wire TIMEBOOST_net_11634;
wire TIMEBOOST_net_14279;
wire g62939_sb;
wire TIMEBOOST_net_11872;
wire TIMEBOOST_net_14823;
wire g62940_sb;
wire TIMEBOOST_net_11637;
wire TIMEBOOST_net_14662;
wire g62941_sb;
wire TIMEBOOST_net_14375;
wire TIMEBOOST_net_11357;
wire g62942_sb;
wire TIMEBOOST_net_11499;
wire TIMEBOOST_net_1373;
wire g62943_sb;
wire TIMEBOOST_net_11510;
wire TIMEBOOST_net_14821;
wire g62944_sb;
wire TIMEBOOST_net_11659;
wire TIMEBOOST_net_14928;
wire g62945_sb;
wire TIMEBOOST_net_11512;
wire TIMEBOOST_net_15205;
wire g62946_sb;
wire TIMEBOOST_net_11586;
wire TIMEBOOST_net_13982;
wire g62947_sb;
wire TIMEBOOST_net_11591;
wire TIMEBOOST_net_14397;
wire g62948_sb;
wire TIMEBOOST_net_11513;
wire TIMEBOOST_net_5591;
wire g62949_sb;
wire TIMEBOOST_net_11798;
wire TIMEBOOST_net_14730;
wire g62950_sb;
wire TIMEBOOST_net_1633;
wire TIMEBOOST_net_11239;
wire g62951_sb;
wire TIMEBOOST_net_11799;
wire TIMEBOOST_net_14642;
wire g62952_sb;
wire TIMEBOOST_net_11661;
wire TIMEBOOST_net_14929;
wire g62953_sb;
wire TIMEBOOST_net_11800;
wire TIMEBOOST_net_14860;
wire g62954_sb;
wire TIMEBOOST_net_11594;
wire TIMEBOOST_net_14123;
wire g62955_sb;
wire TIMEBOOST_net_11687;
wire TIMEBOOST_net_13983;
wire g62956_sb;
wire TIMEBOOST_net_14111;
wire TIMEBOOST_net_11240;
wire g62957_sb;
wire TIMEBOOST_net_11491;
wire TIMEBOOST_net_14595;
wire g62958_sb;
wire TIMEBOOST_net_11492;
wire TIMEBOOST_net_15062;
wire g62959_sb;
wire TIMEBOOST_net_11701;
wire TIMEBOOST_net_14124;
wire g62960_sb;
wire TIMEBOOST_net_13986;
wire TIMEBOOST_net_11658;
wire g62961_sb;
wire TIMEBOOST_net_11498;
wire TIMEBOOST_net_14862;
wire g62962_sb;
wire TIMEBOOST_net_14112;
wire TIMEBOOST_net_11241;
wire g62963_sb;
wire TIMEBOOST_net_11663;
wire TIMEBOOST_net_14249;
wire g62964_sb;
wire TIMEBOOST_net_11501;
wire TIMEBOOST_net_14752;
wire g62965_sb;
wire TIMEBOOST_net_14567;
wire TIMEBOOST_net_11818;
wire g62966_sb;
wire TIMEBOOST_net_11603;
wire TIMEBOOST_net_14356;
wire g62967_sb;
wire TIMEBOOST_net_11613;
wire TIMEBOOST_net_14353;
wire g62968_sb;
wire TIMEBOOST_net_11572;
wire TIMEBOOST_net_14252;
wire g62969_sb;
wire TIMEBOOST_net_11502;
wire TIMEBOOST_net_1384;
wire g62970_sb;
wire TIMEBOOST_net_11655;
wire TIMEBOOST_net_6059;
wire g62971_sb;
wire TIMEBOOST_net_11503;
wire TIMEBOOST_net_14851;
wire g62972_sb;
wire TIMEBOOST_net_11657;
wire TIMEBOOST_net_14251;
wire g62973_sb;
wire TIMEBOOST_net_11504;
wire TIMEBOOST_net_15060;
wire g62974_sb;
wire TIMEBOOST_net_11673;
wire TIMEBOOST_net_15028;
wire g62975_sb;
wire TIMEBOOST_net_11505;
wire TIMEBOOST_net_15056;
wire g62976_sb;
wire TIMEBOOST_net_11829;
wire TIMEBOOST_net_15029;
wire g62977_sb;
wire TIMEBOOST_net_11641;
wire TIMEBOOST_net_14233;
wire g62978_sb;
wire TIMEBOOST_net_11753;
wire TIMEBOOST_net_14398;
wire g62979_sb;
wire TIMEBOOST_net_13914;
wire TIMEBOOST_net_11830;
wire g62980_sb;
wire TIMEBOOST_net_11636;
wire TIMEBOOST_net_15030;
wire g62981_sb;
wire TIMEBOOST_net_14029;
wire TIMEBOOST_net_11832;
wire g62982_sb;
wire TIMEBOOST_net_11617;
wire TIMEBOOST_net_13997;
wire g62983_sb;
wire TIMEBOOST_net_11506;
wire TIMEBOOST_net_15034;
wire g62984_sb;
wire TIMEBOOST_net_11633;
wire TIMEBOOST_net_15031;
wire g62985_sb;
wire TIMEBOOST_net_11508;
wire TIMEBOOST_net_15041;
wire g62986_sb;
wire TIMEBOOST_net_11640;
wire TIMEBOOST_net_15033;
wire g62987_sb;
wire TIMEBOOST_net_11624;
wire TIMEBOOST_net_14603;
wire g62988_sb;
wire TIMEBOOST_net_11509;
wire TIMEBOOST_net_14762;
wire g62989_sb;
wire TIMEBOOST_net_11606;
wire TIMEBOOST_net_9335;
wire g62990_sb;
wire TIMEBOOST_net_1637;
wire TIMEBOOST_net_11242;
wire g62991_sb;
wire TIMEBOOST_net_11610;
wire TIMEBOOST_net_9336;
wire g62992_sb;
wire TIMEBOOST_net_14035;
wire TIMEBOOST_net_11243;
wire g62993_sb;
wire TIMEBOOST_net_12252;
wire TIMEBOOST_net_11244;
wire g62994_sb;
wire TIMEBOOST_net_1640;
wire TIMEBOOST_net_11245;
wire g62995_sb;
wire TIMEBOOST_net_11616;
wire TIMEBOOST_net_9337;
wire g62996_sb;
wire TIMEBOOST_net_14638;
wire TIMEBOOST_net_11246;
wire g62997_sb;
wire TIMEBOOST_net_11642;
wire TIMEBOOST_net_14463;
wire g62998_sb;
wire TIMEBOOST_net_11515;
wire TIMEBOOST_net_14702;
wire g62999_sb;
wire TIMEBOOST_net_11619;
wire TIMEBOOST_net_15035;
wire g63000_sb;
wire TIMEBOOST_net_11801;
wire TIMEBOOST_net_15058;
wire g63001_sb;
wire TIMEBOOST_net_1642;
wire TIMEBOOST_net_11247;
wire g63002_sb;
wire TIMEBOOST_net_11628;
wire TIMEBOOST_net_9338;
wire g63003_sb;
wire TIMEBOOST_net_11644;
wire TIMEBOOST_net_14606;
wire g63004_sb;
wire TIMEBOOST_net_11742;
wire TIMEBOOST_net_15037;
wire g63005_sb;
wire TIMEBOOST_net_11802;
wire TIMEBOOST_net_14843;
wire g63006_sb;
wire TIMEBOOST_net_11803;
wire TIMEBOOST_net_14837;
wire g63007_sb;
wire TIMEBOOST_net_11646;
wire TIMEBOOST_net_13923;
wire g63008_sb;
wire TIMEBOOST_net_11743;
wire TIMEBOOST_net_14148;
wire g63009_sb;
wire TIMEBOOST_net_1009;
wire TIMEBOOST_net_11090;
wire g63010_sb;
wire TIMEBOOST_net_11804;
wire TIMEBOOST_net_14740;
wire g63011_sb;
wire TIMEBOOST_net_1010;
wire TIMEBOOST_net_11091;
wire g63012_sb;
wire TIMEBOOST_net_4782;
wire g63013_db;
wire g63013_sb;
wire TIMEBOOST_net_11083;
wire TIMEBOOST_net_790;
wire g63014_sb;
wire TIMEBOOST_net_11084;
wire TIMEBOOST_net_14050;
wire g63015_sb;
wire g63016_db;
wire g63016_sb;
wire TIMEBOOST_net_1011;
wire TIMEBOOST_net_11092;
wire g63017_sb;
wire TIMEBOOST_net_11085;
wire TIMEBOOST_net_14454;
wire g63018_sb;
wire TIMEBOOST_net_12407;
wire TIMEBOOST_net_11093;
wire g63019_sb;
wire g63020_db;
wire g63020_sb;
wire TIMEBOOST_net_1013;
wire TIMEBOOST_net_11094;
wire g63021_sb;
wire TIMEBOOST_net_1014;
wire TIMEBOOST_net_11095;
wire g63022_sb;
wire TIMEBOOST_net_1015;
wire TIMEBOOST_net_11096;
wire g63023_sb;
wire TIMEBOOST_net_1016;
wire TIMEBOOST_net_11097;
wire g63024_sb;
wire TIMEBOOST_net_4878;
wire g63025_db;
wire TIMEBOOST_net_11086;
wire TIMEBOOST_net_793;
wire g63026_sb;
wire TIMEBOOST_net_1017;
wire g63027_db;
wire g63027_sb;
wire TIMEBOOST_net_1018;
wire TIMEBOOST_net_11098;
wire g63028_sb;
wire TIMEBOOST_net_11621;
wire TIMEBOOST_net_13919;
wire g63029_sb;
wire TIMEBOOST_net_1019;
wire TIMEBOOST_net_11099;
wire g63030_sb;
wire FE_RN_580_0;
wire g63031_db;
wire g63031_sb;
wire TIMEBOOST_net_1021;
wire TIMEBOOST_net_11100;
wire g63032_sb;
wire TIMEBOOST_net_3443;
wire TIMEBOOST_net_11101;
wire g63033_sb;
wire TIMEBOOST_net_1023;
wire TIMEBOOST_net_11102;
wire g63034_sb;
wire TIMEBOOST_net_1024;
wire TIMEBOOST_net_11103;
wire g63035_sb;
wire TIMEBOOST_net_14661;
wire g63036_db;
wire g63036_sb;
wire TIMEBOOST_net_1026;
wire TIMEBOOST_net_11104;
wire g63037_sb;
wire TIMEBOOST_net_15047;
wire TIMEBOOST_net_11105;
wire g63038_sb;
wire TIMEBOOST_net_9527;
wire g63039_db;
wire g63039_sb;
wire TIMEBOOST_net_12391;
wire TIMEBOOST_net_11106;
wire g63040_sb;
wire TIMEBOOST_net_1029;
wire TIMEBOOST_net_11107;
wire g63041_sb;
wire TIMEBOOST_net_11629;
wire TIMEBOOST_net_14152;
wire g63042_sb;
wire TIMEBOOST_net_11087;
wire TIMEBOOST_net_3985;
wire g63043_sb;
wire TIMEBOOST_net_1030;
wire TIMEBOOST_net_14045;
wire g63044_sb;
wire TIMEBOOST_net_11108;
wire g63045_sb;
wire TIMEBOOST_net_14745;
wire TIMEBOOST_net_11109;
wire g63046_sb;
wire TIMEBOOST_net_718;
wire g63047_db;
wire g63047_sb;
wire TIMEBOOST_net_12995;
wire TIMEBOOST_net_12067;
wire g63048_sb;
wire TIMEBOOST_net_15020;
wire TIMEBOOST_net_11110;
wire g63049_sb;
wire TIMEBOOST_net_15021;
wire TIMEBOOST_net_11111;
wire g63050_sb;
wire TIMEBOOST_net_15203;
wire g63051_db;
wire g63051_sb;
wire TIMEBOOST_net_719;
wire g63052_db;
wire g63052_sb;
wire TIMEBOOST_net_14713;
wire TIMEBOOST_net_11112;
wire g63053_sb;
wire TIMEBOOST_net_14718;
wire TIMEBOOST_net_11113;
wire g63054_sb;
wire TIMEBOOST_net_14720;
wire TIMEBOOST_net_11114;
wire g63055_sb;
wire TIMEBOOST_net_637;
wire g63056_db;
wire g63056_sb;
wire TIMEBOOST_net_638;
wire TIMEBOOST_net_11115;
wire TIMEBOOST_net_12924;
wire TIMEBOOST_net_10374;
wire g63058_sb;
wire TIMEBOOST_net_14722;
wire TIMEBOOST_net_11116;
wire g63059_sb;
wire TIMEBOOST_net_14738;
wire g63060_db;
wire g63060_sb;
wire TIMEBOOST_net_14739;
wire TIMEBOOST_net_11117;
wire g63061_sb;
wire TIMEBOOST_net_14684;
wire TIMEBOOST_net_11118;
wire g63062_sb;
wire TIMEBOOST_net_14774;
wire g63063_db;
wire g63063_sb;
wire TIMEBOOST_net_14775;
wire TIMEBOOST_net_11119;
wire g63064_sb;
wire TIMEBOOST_net_14784;
wire TIMEBOOST_net_11120;
wire g63065_sb;
wire TIMEBOOST_net_14714;
wire TIMEBOOST_net_11121;
wire g63066_sb;
wire TIMEBOOST_net_14715;
wire TIMEBOOST_net_11122;
wire g63067_sb;
wire TIMEBOOST_net_14726;
wire TIMEBOOST_net_11123;
wire g63068_sb;
wire TIMEBOOST_net_14990;
wire TIMEBOOST_net_11126;
wire g63069_sb;
wire TIMEBOOST_net_14992;
wire TIMEBOOST_net_11130;
wire g63070_sb;
wire TIMEBOOST_net_14911;
wire TIMEBOOST_net_11131;
wire g63071_sb;
wire TIMEBOOST_net_14631;
wire TIMEBOOST_net_11133;
wire g63072_sb;
wire TIMEBOOST_net_14736;
wire TIMEBOOST_net_11136;
wire g63073_sb;
wire TIMEBOOST_net_14978;
wire TIMEBOOST_net_11137;
wire g63074_sb;
wire TIMEBOOST_net_14979;
wire TIMEBOOST_net_11139;
wire g63075_sb;
wire TIMEBOOST_net_14741;
wire TIMEBOOST_net_11141;
wire g63076_sb;
wire TIMEBOOST_net_9371;
wire g63077_db;
wire g63077_sb;
wire TIMEBOOST_net_14904;
wire TIMEBOOST_net_11142;
wire g63078_sb;
wire TIMEBOOST_net_15212;
wire TIMEBOOST_net_11144;
wire g63079_sb;
wire TIMEBOOST_net_11088;
wire TIMEBOOST_net_3986;
wire g63080_sb;
wire TIMEBOOST_net_11089;
wire TIMEBOOST_net_3987;
wire g63081_sb;
wire TIMEBOOST_net_14744;
wire TIMEBOOST_net_11147;
wire g63082_sb;
wire TIMEBOOST_net_11124;
wire TIMEBOOST_net_14359;
wire g63083_sb;
wire TIMEBOOST_net_1059;
wire TIMEBOOST_net_11148;
wire g63084_sb;
wire TIMEBOOST_net_9369;
wire TIMEBOOST_net_13351;
wire g63085_sb;
wire TIMEBOOST_net_12998;
wire g63086_db;
wire g63086_sb;
wire TIMEBOOST_net_1060;
wire TIMEBOOST_net_14082;
wire g63087_sb;
wire TIMEBOOST_net_14639;
wire TIMEBOOST_net_11149;
wire g63088_sb;
wire TIMEBOOST_net_12922;
wire TIMEBOOST_net_10375;
wire g63089_sb;
wire TIMEBOOST_net_14706;
wire TIMEBOOST_net_11150;
wire g63090_sb;
wire TIMEBOOST_net_740;
wire g63091_db;
wire g63091_sb;
wire TIMEBOOST_net_11125;
wire g63092_sb;
wire TIMEBOOST_net_11127;
wire TIMEBOOST_net_799;
wire g63093_sb;
wire TIMEBOOST_net_11805;
wire TIMEBOOST_net_15059;
wire g63094_sb;
wire TIMEBOOST_net_14139;
wire g63095_db;
wire g63095_sb;
wire TIMEBOOST_net_742;
wire TIMEBOOST_net_11151;
wire g63096_sb;
wire TIMEBOOST_net_9561;
wire TIMEBOOST_net_11152;
wire g63097_sb;
wire g66424_db;
wire TIMEBOOST_net_11153;
wire g63098_sb;
wire TIMEBOOST_net_11128;
wire TIMEBOOST_net_800;
wire g63099_sb;
wire TIMEBOOST_net_1065;
wire TIMEBOOST_net_11154;
wire g63100_sb;
wire TIMEBOOST_net_14757;
wire g63101_db;
wire g63101_sb;
wire g66422_db;
wire TIMEBOOST_net_11155;
wire g63102_sb;
wire TIMEBOOST_net_1068;
wire TIMEBOOST_net_11156;
wire g63103_sb;
wire TIMEBOOST_net_14727;
wire TIMEBOOST_net_11157;
wire g63104_sb;
wire TIMEBOOST_net_11129;
wire TIMEBOOST_net_801;
wire g63105_sb;
wire TIMEBOOST_net_14734;
wire TIMEBOOST_net_11158;
wire g63106_sb;
wire TIMEBOOST_net_9562;
wire TIMEBOOST_net_11159;
wire g63107_sb;
wire TIMEBOOST_net_11806;
wire TIMEBOOST_net_15057;
wire g63108_sb;
wire TIMEBOOST_net_14925;
wire TIMEBOOST_net_11160;
wire g63109_sb;
wire TIMEBOOST_net_14894;
wire TIMEBOOST_net_11161;
wire g63110_sb;
wire TIMEBOOST_net_14809;
wire TIMEBOOST_net_11163;
wire g63111_sb;
wire TIMEBOOST_net_14896;
wire TIMEBOOST_net_11167;
wire g63112_sb;
wire TIMEBOOST_net_1076;
wire TIMEBOOST_net_10881;
wire g63113_sb;
wire TIMEBOOST_net_1077;
wire TIMEBOOST_net_10841;
wire g63114_sb;
wire TIMEBOOST_net_1078;
wire TIMEBOOST_net_10845;
wire g63115_sb;
wire TIMEBOOST_net_1079;
wire TIMEBOOST_net_10846;
wire g63116_sb;
wire TIMEBOOST_net_12756;
wire g63117_db;
wire g63117_sb;
wire TIMEBOOST_net_14640;
wire TIMEBOOST_net_10847;
wire g63118_sb;
wire TIMEBOOST_net_14659;
wire TIMEBOOST_net_10848;
wire g63119_sb;
wire TIMEBOOST_net_11132;
wire TIMEBOOST_net_4558;
wire g63120_sb;
wire TIMEBOOST_net_1082;
wire TIMEBOOST_net_10849;
wire g63121_sb;
wire TIMEBOOST_net_14984;
wire TIMEBOOST_net_10850;
wire g63122_sb;
wire TIMEBOOST_net_14844;
wire TIMEBOOST_net_10851;
wire g63123_sb;
wire TIMEBOOST_net_13824;
wire g63124_db;
wire g63124_sb;
wire TIMEBOOST_net_14699;
wire TIMEBOOST_net_10852;
wire g63125_sb;
wire TIMEBOOST_net_9370;
wire g63126_db;
wire g63126_sb;
wire TIMEBOOST_net_4789;
wire g63127_db;
wire TIMEBOOST_net_14697;
wire TIMEBOOST_net_10853;
wire g63128_sb;
wire TIMEBOOST_net_15219;
wire TIMEBOOST_net_10854;
wire TIMEBOOST_net_12387;
wire TIMEBOOST_net_10855;
wire g63130_sb;
wire TIMEBOOST_net_9580;
wire TIMEBOOST_net_10856;
wire g63131_sb;
wire TIMEBOOST_net_14897;
wire TIMEBOOST_net_10857;
wire g63132_sb;
wire TIMEBOOST_net_12630;
wire TIMEBOOST_net_11038;
wire g63133_sb;
wire TIMEBOOST_net_13195;
wire TIMEBOOST_net_11164;
wire g63134_sb;
wire TIMEBOOST_net_1092;
wire TIMEBOOST_net_11165;
wire g63135_sb;
wire TIMEBOOST_net_11134;
wire TIMEBOOST_net_4559;
wire g63136_sb;
wire TIMEBOOST_net_11135;
wire TIMEBOOST_net_4560;
wire g63137_sb;
wire TIMEBOOST_net_12923;
wire TIMEBOOST_net_10843;
wire g63138_sb;
wire TIMEBOOST_net_14749;
wire TIMEBOOST_net_11166;
wire g63139_sb;
wire TIMEBOOST_net_1094;
wire TIMEBOOST_net_10832;
wire g63140_sb;
wire TIMEBOOST_net_646;
wire TIMEBOOST_net_4684;
wire g63141_sb;
wire TIMEBOOST_net_1095;
wire TIMEBOOST_net_10834;
wire g63142_sb;
wire TIMEBOOST_net_1096;
wire TIMEBOOST_net_10835;
wire g63143_sb;
wire TIMEBOOST_net_11688;
wire TIMEBOOST_net_12580;
wire g63144_sb;
wire TIMEBOOST_net_1643;
wire TIMEBOOST_net_11248;
wire g63145_sb;
wire TIMEBOOST_net_11807;
wire TIMEBOOST_net_1398;
wire g63146_sb;
wire TIMEBOOST_net_11808;
wire TIMEBOOST_net_14853;
wire g63147_sb;
wire TIMEBOOST_net_11809;
wire TIMEBOOST_net_14710;
wire g63148_sb;
wire TIMEBOOST_net_11810;
wire TIMEBOOST_net_15063;
wire g63149_sb;
wire TIMEBOOST_net_11744;
wire TIMEBOOST_net_15026;
wire g63150_sb;
wire TIMEBOOST_net_1644;
wire TIMEBOOST_net_11249;
wire g63151_sb;
wire TIMEBOOST_net_11138;
wire TIMEBOOST_net_4561;
wire g63152_sb;
wire TIMEBOOST_net_11751;
wire TIMEBOOST_net_15036;
wire g63153_sb;
wire TIMEBOOST_net_1645;
wire g63154_db;
wire g63154_sb;
wire TIMEBOOST_net_11689;
wire TIMEBOOST_net_14416;
wire g63155_sb;
wire TIMEBOOST_net_1646;
wire TIMEBOOST_net_11250;
wire g63156_sb;
wire TIMEBOOST_net_11756;
wire TIMEBOOST_net_15052;
wire g63157_sb;
wire TIMEBOOST_net_11551;
wire TIMEBOOST_net_1405;
wire g63158_sb;
wire TIMEBOOST_net_11648;
wire TIMEBOOST_net_13918;
wire g63159_sb;
wire TIMEBOOST_net_11649;
wire TIMEBOOST_net_13927;
wire g63160_sb;
wire TIMEBOOST_net_11650;
wire TIMEBOOST_net_13990;
wire g63161_sb;
wire TIMEBOOST_net_11552;
wire TIMEBOOST_net_15049;
wire g63162_sb;
wire TIMEBOOST_net_11553;
wire TIMEBOOST_net_15042;
wire g63163_sb;
wire TIMEBOOST_net_1647;
wire TIMEBOOST_net_11251;
wire g63164_sb;
wire TIMEBOOST_net_744;
wire TIMEBOOST_net_4685;
wire g63165_sb;
wire TIMEBOOST_net_11554;
wire TIMEBOOST_net_14634;
wire g63166_sb;
wire TIMEBOOST_net_1648;
wire TIMEBOOST_net_11252;
wire g63167_sb;
wire TIMEBOOST_net_11555;
wire TIMEBOOST_net_15055;
wire g63168_sb;
wire TIMEBOOST_net_9587;
wire TIMEBOOST_net_10838;
wire g63169_sb;
wire TIMEBOOST_net_1098;
wire TIMEBOOST_net_10860;
wire g63170_sb;
wire TIMEBOOST_net_1649;
wire TIMEBOOST_net_11253;
wire g63171_sb;
wire TIMEBOOST_net_12300;
wire TIMEBOOST_net_10873;
wire g63172_sb;
wire TIMEBOOST_net_1650;
wire TIMEBOOST_net_11315;
wire g63173_sb;
wire TIMEBOOST_net_1651;
wire TIMEBOOST_net_11316;
wire g63174_sb;
wire TIMEBOOST_net_1100;
wire TIMEBOOST_net_10875;
wire g63175_sb;
wire TIMEBOOST_net_1101;
wire TIMEBOOST_net_10877;
wire g63176_sb;
wire TIMEBOOST_net_11690;
wire TIMEBOOST_net_14275;
wire g63177_sb;
wire TIMEBOOST_net_11652;
wire TIMEBOOST_net_14063;
wire g63178_sb;
wire TIMEBOOST_net_6447;
wire g63179_db;
wire g63179_sb;
wire TIMEBOOST_net_11556;
wire TIMEBOOST_net_14939;
wire g63180_sb;
wire TIMEBOOST_net_1652;
wire TIMEBOOST_net_11317;
wire g63181_sb;
wire TIMEBOOST_net_1102;
wire TIMEBOOST_net_10878;
wire g63182_sb;
wire TIMEBOOST_net_15201;
wire TIMEBOOST_net_11318;
wire g63183_sb;
wire TIMEBOOST_net_11557;
wire TIMEBOOST_net_14942;
wire g63184_sb;
wire TIMEBOOST_net_11558;
wire TIMEBOOST_net_14943;
wire g63185_sb;
wire TIMEBOOST_net_11691;
wire TIMEBOOST_net_14100;
wire g63186_sb;
wire TIMEBOOST_net_11560;
wire TIMEBOOST_net_14733;
wire g63187_sb;
wire TIMEBOOST_net_1103;
wire TIMEBOOST_net_10879;
wire g63188_sb;
wire TIMEBOOST_net_11561;
wire TIMEBOOST_net_14703;
wire g63189_sb;
wire TIMEBOOST_net_11562;
wire TIMEBOOST_net_14732;
wire g63190_sb;
wire TIMEBOOST_net_1104;
wire TIMEBOOST_net_10899;
wire g63191_sb;
wire TIMEBOOST_net_14399;
wire TIMEBOOST_net_11319;
wire g63192_sb;
wire TIMEBOOST_net_13705;
wire TIMEBOOST_net_4494;
wire g63193_sb;
wire TIMEBOOST_net_12369;
wire TIMEBOOST_net_11081;
wire g63194_sb;
wire TIMEBOOST_net_4701;
wire g63195_db;
wire g63195_sb;
wire TIMEBOOST_net_4702;
wire g63196_db;
wire g63196_sb;
wire TIMEBOOST_net_14400;
wire g63197_db;
wire g63197_sb;
wire TIMEBOOST_net_14913;
wire g63198_db;
wire g63198_sb;
wire TIMEBOOST_net_14914;
wire g63199_db;
wire g63199_sb;
wire g63200_p;
wire g63201_p;
wire TIMEBOOST_net_11320;
wire TIMEBOOST_net_14437;
wire g63202_sb;
wire TIMEBOOST_net_11321;
wire TIMEBOOST_net_14408;
wire g63203_sb;
wire TIMEBOOST_net_13793;
wire TIMEBOOST_net_10868;
wire g63204_sb;
wire g63206_p;
wire g63207_p;
wire g63208_p;
wire g63209_p;
wire g63215_p;
wire g63216_p;
wire g63217_p;
wire g63252_p;
wire g63253_p;
wire g63256_p;
wire g63259_p;
wire g63263_p;
wire g63268_p;
wire g63271_p;
wire g63291_p;
wire g63292_p;
wire g63293_p;
wire g63307_p;
wire g63315_p;
wire g63338_p;
wire g63340_p;
wire g63348_p;
wire g63361_p;
wire g63362_p;
wire g63364_p;
wire TIMEBOOST_net_1105;
wire g63378_db;
wire g63378_sb;
wire TIMEBOOST_net_1106;
wire TIMEBOOST_net_10724;
wire g63392_sb;
wire TIMEBOOST_net_1107;
wire TIMEBOOST_net_13965;
wire g63397_sb;
wire g63409_p;
wire g63422_p;
wire g63423_p;
wire g63424_p;
wire g63426_p;
wire g63428_p;
wire g63429_p;
wire TIMEBOOST_net_12288;
wire TIMEBOOST_net_14665;
wire TIMEBOOST_net_10906;
wire g63431_sb;
wire TIMEBOOST_net_14980;
wire TIMEBOOST_net_10908;
wire g63432_sb;
wire TIMEBOOST_net_14899;
wire TIMEBOOST_net_10910;
wire g63433_sb;
wire TIMEBOOST_net_14901;
wire TIMEBOOST_net_10912;
wire g63434_sb;
wire TIMEBOOST_net_14903;
wire g63435_db;
wire g63435_sb;
wire TIMEBOOST_net_14678;
wire TIMEBOOST_net_10917;
wire g63436_sb;
wire TIMEBOOST_net_14679;
wire TIMEBOOST_net_10919;
wire g63437_sb;
wire TIMEBOOST_net_15027;
wire TIMEBOOST_net_10925;
wire g63438_sb;
wire g63525_p;
wire TIMEBOOST_net_10332;
wire g63530_db;
wire g63530_sb;
wire TIMEBOOST_net_4814;
wire TIMEBOOST_net_4686;
wire g63533_sb;
wire TIMEBOOST_net_15039;
wire g63537_db;
wire g63537_sb;
wire TIMEBOOST_net_10712;
wire g63538_db;
wire g63538_sb;
wire g63539_p;
wire g63542_p;
wire g63543_da;
wire g63543_db;
wire g63543_sb;
wire TIMEBOOST_net_10713;
wire g63544_db;
wire g63544_sb;
wire g63545_da;
wire g63545_db;
wire g63545_sb;
wire g63546_p;
wire TIMEBOOST_net_14189;
wire g63547_db;
wire g63547_sb;
wire TIMEBOOST_net_3155;
wire g63548_db;
wire g63548_sb;
wire TIMEBOOST_net_14556;
wire g63549_db;
wire g63549_sb;
wire TIMEBOOST_net_14728;
wire TIMEBOOST_net_10936;
wire g63550_sb;
wire TIMEBOOST_net_14688;
wire TIMEBOOST_net_10943;
wire g63551_sb;
wire TIMEBOOST_net_14780;
wire TIMEBOOST_net_10946;
wire g63552_sb;
wire TIMEBOOST_net_14781;
wire TIMEBOOST_net_10948;
wire g63553_sb;
wire TIMEBOOST_net_14683;
wire TIMEBOOST_net_11199;
wire g63554_sb;
wire TIMEBOOST_net_12374;
wire TIMEBOOST_net_11200;
wire g63555_sb;
wire TIMEBOOST_net_12378;
wire TIMEBOOST_net_11201;
wire g63556_sb;
wire TIMEBOOST_net_12385;
wire TIMEBOOST_net_10984;
wire g63557_sb;
wire TIMEBOOST_net_12360;
wire g63559_db;
wire g63559_sb;
wire TIMEBOOST_net_14101;
wire g63560_db;
wire g63560_sb;
wire TIMEBOOST_net_14046;
wire g63561_db;
wire g63561_sb;
wire TIMEBOOST_net_13934;
wire g63562_db;
wire g63562_sb;
wire g63563_da;
wire g63563_db;
wire g63563_sb;
wire TIMEBOOST_net_10549;
wire g63564_db;
wire g63564_sb;
wire g63565_da;
wire g63565_db;
wire g63565_sb;
wire g63566_da;
wire g63566_db;
wire g63566_sb;
wire TIMEBOOST_net_10230;
wire g63567_db;
wire g63567_sb;
wire TIMEBOOST_net_10231;
wire g63568_db;
wire g63568_sb;
wire TIMEBOOST_net_4519;
wire g63569_db;
wire g63569_sb;
wire g63570_da;
wire g63570_db;
wire g63570_sb;
wire TIMEBOOST_net_1125;
wire g63571_db;
wire g63571_sb;
wire TIMEBOOST_net_4790;
wire g63572_db;
wire g63572_sb;
wire TIMEBOOST_net_14015;
wire g63573_db;
wire g63573_sb;
wire TIMEBOOST_net_14034;
wire g63574_db;
wire g63574_sb;
wire TIMEBOOST_net_5429;
wire TIMEBOOST_net_14332;
wire g63576_sb;
wire TIMEBOOST_net_9366;
wire TIMEBOOST_net_10955;
wire g63577_sb;
wire g63578_p;
wire g63579_p;
wire g63580_p;
wire g63581_p;
wire TIMEBOOST_net_10370;
wire g63582_db;
wire g63582_sb;
wire TIMEBOOST_net_262;
wire TIMEBOOST_net_14471;
wire TIMEBOOST_net_10135;
wire g63584_db;
wire g63584_sb;
wire TIMEBOOST_net_13344;
wire g63585_db;
wire TIMEBOOST_net_10136;
wire g63586_db;
wire g63586_sb;
wire TIMEBOOST_net_10150;
wire g63587_db;
wire TIMEBOOST_net_10152;
wire g63588_db;
wire g63588_sb;
wire TIMEBOOST_net_12554;
wire TIMEBOOST_net_13362;
wire g63589_sb;
wire TIMEBOOST_net_119;
wire TIMEBOOST_net_12389;
wire g63590_sb;
wire g63591_da;
wire TIMEBOOST_net_4689;
wire g63591_sb;
wire TIMEBOOST_net_12555;
wire g63592_db;
wire g63592_sb;
wire TIMEBOOST_net_683;
wire TIMEBOOST_net_13363;
wire g63593_sb;
wire TIMEBOOST_net_12722;
wire TIMEBOOST_net_13364;
wire g63594_sb;
wire TIMEBOOST_net_12179;
wire TIMEBOOST_net_13365;
wire g63595_sb;
wire TIMEBOOST_net_686;
wire TIMEBOOST_net_13366;
wire g63596_sb;
wire g63597_da;
wire TIMEBOOST_net_10705;
wire g63597_sb;
wire TIMEBOOST_net_9447;
wire TIMEBOOST_net_13367;
wire g63598_sb;
wire g63599_da;
wire g63599_db;
wire g63599_sb;
wire TIMEBOOST_net_3727;
wire TIMEBOOST_net_13368;
wire g63600_sb;
wire TIMEBOOST_net_9448;
wire g63601_db;
wire g63601_sb;
wire g63602_da;
wire g63602_db;
wire g63602_sb;
wire g63603_da;
wire g63603_db;
wire g63603_sb;
wire g63604_da;
wire TIMEBOOST_net_10706;
wire g63604_sb;
wire g63605_da;
wire g63605_db;
wire g63605_sb;
wire g63606_da;
wire TIMEBOOST_net_10707;
wire g63606_sb;
wire g63607_da;
wire g63607_db;
wire g63607_sb;
wire TIMEBOOST_net_12604;
wire TIMEBOOST_net_13369;
wire g63608_sb;
wire g63609_da;
wire TIMEBOOST_net_4693;
wire g63609_sb;
wire TIMEBOOST_net_12606;
wire TIMEBOOST_net_13370;
wire g63610_sb;
wire g63611_da;
wire g63611_db;
wire g63611_sb;
wire g63612_da;
wire TIMEBOOST_net_4694;
wire g63612_sb;
wire g63613_da;
wire g63613_db;
wire g63613_sb;
wire g63614_da;
wire g63614_db;
wire g63614_sb;
wire TIMEBOOST_net_12608;
wire TIMEBOOST_net_13371;
wire g63615_sb;
wire TIMEBOOST_net_12186;
wire g63616_db;
wire g63616_sb;
wire g63617_da;
wire TIMEBOOST_net_10708;
wire g63617_sb;
wire TIMEBOOST_net_12499;
wire g63618_db;
wire g63618_sb;
wire g63619_da;
wire g63619_db;
wire g63619_sb;
wire TIMEBOOST_net_12503;
wire TIMEBOOST_net_13372;
wire g63620_sb;
wire g63621_da;
wire TIMEBOOST_net_4696;
wire g63621_sb;
wire g63891_p;
wire g63892_p;
wire g63895_p;
wire g63902_p;
wire g63916_p;
wire g63922_p;
wire g63925_p;
wire g63935_p;
wire g63939_p;
wire TIMEBOOST_net_3734;
wire TIMEBOOST_net_12388;
wire g63943_p;
wire g63989_p;
wire g64022_p;
wire TIMEBOOST_net_9318;
wire TIMEBOOST_net_10551;
wire g64078_sb;
wire TIMEBOOST_net_10553;
wire g64079_db;
wire g64079_sb;
wire TIMEBOOST_net_4705;
wire g64080_db;
wire g64080_sb;
wire TIMEBOOST_net_10714;
wire g64081_db;
wire g64081_sb;
wire TIMEBOOST_net_4707;
wire g64082_db;
wire g64082_sb;
wire TIMEBOOST_net_10715;
wire g64083_db;
wire g64083_sb;
wire TIMEBOOST_net_10716;
wire g64084_db;
wire g64084_sb;
wire TIMEBOOST_net_3156;
wire g64085_db;
wire g64085_sb;
wire TIMEBOOST_net_10717;
wire g64086_db;
wire g64086_sb;
wire TIMEBOOST_net_9534;
wire g64087_db;
wire g64087_sb;
wire TIMEBOOST_net_4711;
wire g64088_db;
wire g64088_sb;
wire TIMEBOOST_net_4712;
wire g64089_db;
wire g64089_sb;
wire TIMEBOOST_net_10554;
wire g64090_db;
wire g64090_sb;
wire TIMEBOOST_net_10555;
wire g64091_db;
wire g64091_sb;
wire TIMEBOOST_net_10718;
wire g64092_db;
wire g64092_sb;
wire g64093_da;
wire g64093_db;
wire g64093_sb;
wire TIMEBOOST_net_10719;
wire g64094_db;
wire g64094_sb;
wire TIMEBOOST_net_9536;
wire g64095_db;
wire g64095_sb;
wire g64096_da;
wire g64096_db;
wire g64096_sb;
wire TIMEBOOST_net_10631;
wire g64097_db;
wire g64097_sb;
wire TIMEBOOST_net_10171;
wire g64098_db;
wire g64098_sb;
wire TIMEBOOST_net_10172;
wire g64099_db;
wire g64099_sb;
wire TIMEBOOST_net_10720;
wire g64100_db;
wire g64100_sb;
wire g64102_da;
wire g64102_db;
wire g64102_sb;
wire TIMEBOOST_net_10721;
wire g64103_db;
wire g64103_sb;
wire g64105_da;
wire g64105_db;
wire g64105_sb;
wire g64106_da;
wire g64106_db;
wire g64106_sb;
wire TIMEBOOST_net_10173;
wire g64107_db;
wire g64107_sb;
wire g64108_da;
wire g64108_db;
wire g64108_sb;
wire TIMEBOOST_net_4717;
wire g64109_db;
wire g64109_sb;
wire TIMEBOOST_net_10178;
wire g64110_db;
wire g64110_sb;
wire TIMEBOOST_net_4718;
wire g64111_db;
wire g64111_sb;
wire TIMEBOOST_net_4719;
wire g64112_db;
wire g64112_sb;
wire TIMEBOOST_net_13662;
wire g64113_db;
wire g64113_sb;
wire g64114_da;
wire g64114_db;
wire g64114_sb;
wire TIMEBOOST_net_10722;
wire g64115_db;
wire g64115_sb;
wire TIMEBOOST_net_14204;
wire g64116_db;
wire g64116_sb;
wire TIMEBOOST_net_4721;
wire g64117_db;
wire g64117_sb;
wire TIMEBOOST_net_9949;
wire g64118_db;
wire g64118_sb;
wire g64119_da;
wire g64119_db;
wire g64119_sb;
wire g64120_da;
wire g64120_db;
wire g64120_sb;
wire TIMEBOOST_net_12241;
wire g64122_db;
wire g64122_sb;
wire g64123_da;
wire g64123_db;
wire g64123_sb;
wire g64124_p;
wire TIMEBOOST_net_4722;
wire g64125_db;
wire g64125_sb;
wire g64126_da;
wire g64126_db;
wire g64126_sb;
wire TIMEBOOST_net_4468;
wire g64127_db;
wire g64127_sb;
wire TIMEBOOST_net_9532;
wire g64128_db;
wire g64128_sb;
wire g64129_da;
wire g64129_db;
wire g64129_sb;
wire TIMEBOOST_net_9956;
wire g64130_db;
wire g64130_sb;
wire g64131_da;
wire g64131_db;
wire g64131_sb;
wire g64132_da;
wire g64132_db;
wire g64132_sb;
wire TIMEBOOST_net_10490;
wire g64133_db;
wire g64133_sb;
wire TIMEBOOST_net_10504;
wire g64134_db;
wire g64134_sb;
wire TIMEBOOST_net_12920;
wire g64135_db;
wire g64135_sb;
wire TIMEBOOST_net_13897;
wire TIMEBOOST_net_14277;
wire g64136_sb;
wire TIMEBOOST_net_10505;
wire g64137_db;
wire g64137_sb;
wire TIMEBOOST_net_14770;
wire g64138_db;
wire g64138_sb;
wire TIMEBOOST_net_3162;
wire g64139_db;
wire g64139_sb;
wire TIMEBOOST_net_10758;
wire g64140_db;
wire g64140_sb;
wire g64141_da;
wire g64141_db;
wire g64141_sb;
wire TIMEBOOST_net_13499;
wire g64142_db;
wire g64142_sb;
wire g64143_da;
wire g64143_db;
wire g64143_sb;
wire TIMEBOOST_net_3719;
wire g64144_db;
wire g64144_sb;
wire TIMEBOOST_net_10333;
wire g64145_db;
wire g64145_sb;
wire TIMEBOOST_net_14494;
wire g64146_db;
wire g64146_sb;
wire g64147_da;
wire g64147_db;
wire g64147_sb;
wire g64148_da;
wire g64148_db;
wire g64148_sb;
wire TIMEBOOST_net_4725;
wire g64149_db;
wire g64149_sb;
wire TIMEBOOST_net_3720;
wire g64150_db;
wire g64150_sb;
wire TIMEBOOST_net_3721;
wire g64151_db;
wire g64151_sb;
wire g64152_da;
wire g64152_db;
wire g64152_sb;
wire TIMEBOOST_net_3722;
wire g64153_db;
wire g64153_sb;
wire TIMEBOOST_net_14478;
wire g64154_db;
wire g64154_sb;
wire TIMEBOOST_net_3723;
wire g64155_db;
wire g64155_sb;
wire TIMEBOOST_net_3724;
wire g64156_db;
wire g64156_sb;
wire TIMEBOOST_net_13896;
wire g64157_db;
wire g64157_sb;
wire g64158_da;
wire g64158_db;
wire g64158_sb;
wire TIMEBOOST_net_3725;
wire g64159_db;
wire g64159_sb;
wire TIMEBOOST_net_14479;
wire g64160_db;
wire g64160_sb;
wire TIMEBOOST_net_13765;
wire g64161_db;
wire g64161_sb;
wire TIMEBOOST_net_9815;
wire g64162_db;
wire g64162_sb;
wire TIMEBOOST_net_9824;
wire g64163_db;
wire g64163_sb;
wire g64164_da;
wire g64164_db;
wire g64164_sb;
wire TIMEBOOST_net_10759;
wire g64165_db;
wire g64165_sb;
wire TIMEBOOST_net_13508;
wire g64166_db;
wire g64166_sb;
wire g64167_da;
wire g64167_db;
wire g64167_sb;
wire TIMEBOOST_net_9837;
wire g64168_db;
wire g64168_sb;
wire g64169_da;
wire g64169_db;
wire g64169_sb;
wire TIMEBOOST_net_10760;
wire g64170_db;
wire g64170_sb;
wire TIMEBOOST_net_14480;
wire g64171_db;
wire g64171_sb;
wire TIMEBOOST_net_15048;
wire g64172_db;
wire g64172_sb;
wire TIMEBOOST_net_10387;
wire g64173_db;
wire g64173_sb;
wire g64175_da;
wire g64175_db;
wire g64175_sb;
wire g64176_da;
wire g64176_db;
wire g64176_sb;
wire g64177_da;
wire g64177_db;
wire g64177_sb;
wire TIMEBOOST_net_9838;
wire g64178_db;
wire g64178_sb;
wire TIMEBOOST_net_10196;
wire g64179_db;
wire g64179_sb;
wire TIMEBOOST_net_9839;
wire g64180_db;
wire g64180_sb;
wire TIMEBOOST_net_13442;
wire g64181_db;
wire g64181_sb;
wire g64182_da;
wire g64182_db;
wire g64182_sb;
wire TIMEBOOST_net_10739;
wire g64183_db;
wire g64183_sb;
wire TIMEBOOST_net_13441;
wire g64184_db;
wire g64184_sb;
wire g64185_da;
wire g64185_db;
wire g64185_sb;
wire TIMEBOOST_net_13763;
wire g64186_db;
wire g64186_sb;
wire TIMEBOOST_net_9301;
wire TIMEBOOST_net_4060;
wire g64187_sb;
wire g64188_da;
wire g64188_db;
wire g64188_sb;
wire g64189_da;
wire g64189_db;
wire g64189_sb;
wire g64190_da;
wire g64190_db;
wire g64190_sb;
wire g64191_da;
wire g64191_db;
wire g64191_sb;
wire g64192_da;
wire g64192_db;
wire g64192_sb;
wire g64193_da;
wire g64193_db;
wire g64193_sb;
wire g64194_p;
wire TIMEBOOST_net_10738;
wire g64195_db;
wire g64195_sb;
wire g64196_da;
wire g64196_db;
wire g64196_sb;
wire TIMEBOOST_net_3163;
wire g64197_db;
wire g64197_sb;
wire TIMEBOOST_net_13770;
wire g64198_db;
wire g64198_sb;
wire TIMEBOOST_net_3164;
wire g64199_db;
wire g64199_sb;
wire g64200_da;
wire g64200_db;
wire g64200_sb;
wire g64201_da;
wire g64201_db;
wire g64201_sb;
wire TIMEBOOST_net_3165;
wire g64202_db;
wire g64202_sb;
wire g64203_da;
wire g64203_db;
wire g64203_sb;
wire TIMEBOOST_net_4476;
wire g64204_db;
wire g64204_sb;
wire TIMEBOOST_net_10761;
wire g64205_db;
wire g64205_sb;
wire g64206_da;
wire g64206_db;
wire g64206_sb;
wire g64207_da;
wire g64207_db;
wire g64207_sb;
wire TIMEBOOST_net_10157;
wire g64208_db;
wire g64208_sb;
wire TIMEBOOST_net_10762;
wire g64209_db;
wire g64209_sb;
wire g64210_da;
wire g64210_db;
wire g64210_sb;
wire TIMEBOOST_net_10754;
wire g64211_db;
wire g64211_sb;
wire TIMEBOOST_net_10750;
wire g64212_db;
wire g64212_sb;
wire TIMEBOOST_net_10158;
wire g64213_db;
wire g64213_sb;
wire TIMEBOOST_net_10751;
wire g64214_db;
wire g64214_sb;
wire TIMEBOOST_net_10329;
wire g64215_db;
wire g64215_sb;
wire TIMEBOOST_net_9540;
wire g64216_db;
wire g64216_sb;
wire TIMEBOOST_net_10182;
wire g64217_db;
wire g64217_sb;
wire TIMEBOOST_net_10752;
wire g64218_db;
wire g64218_sb;
wire g64219_da;
wire g64219_db;
wire g64219_sb;
wire TIMEBOOST_net_10753;
wire g64220_db;
wire g64220_sb;
wire TIMEBOOST_net_10755;
wire g64221_db;
wire g64221_sb;
wire TIMEBOOST_net_10756;
wire g64222_db;
wire g64222_sb;
wire TIMEBOOST_net_10741;
wire g64223_db;
wire g64223_sb;
wire TIMEBOOST_net_10232;
wire g64224_db;
wire g64224_sb;
wire g64225_da;
wire g64225_db;
wire g64225_sb;
wire g64226_da;
wire g64226_db;
wire g64226_sb;
wire TIMEBOOST_net_9811;
wire g64227_db;
wire g64227_sb;
wire TIMEBOOST_net_10552;
wire g64228_db;
wire g64228_sb;
wire TIMEBOOST_net_10556;
wire g64229_db;
wire g64229_sb;
wire TIMEBOOST_net_10557;
wire g64230_db;
wire g64230_sb;
wire TIMEBOOST_net_4520;
wire g64231_db;
wire g64231_sb;
wire TIMEBOOST_net_10558;
wire g64232_db;
wire g64232_sb;
wire TIMEBOOST_net_10559;
wire g64233_db;
wire g64233_sb;
wire TIMEBOOST_net_10566;
wire g64234_db;
wire g64234_sb;
wire TIMEBOOST_net_4521;
wire g64235_db;
wire g64235_sb;
wire TIMEBOOST_net_10637;
wire g64236_db;
wire g64236_sb;
wire TIMEBOOST_net_10567;
wire g64237_db;
wire g64237_sb;
wire TIMEBOOST_net_10568;
wire g64238_db;
wire g64238_sb;
wire g64239_da;
wire g64239_db;
wire g64239_sb;
wire TIMEBOOST_net_10569;
wire g64240_db;
wire g64240_sb;
wire g64241_da;
wire g64241_db;
wire g64241_sb;
wire TIMEBOOST_net_12287;
wire TIMEBOOST_net_4020;
wire g64242_sb;
wire TIMEBOOST_net_10570;
wire g64243_db;
wire g64243_sb;
wire TIMEBOOST_net_10571;
wire g64244_db;
wire g64244_sb;
wire TIMEBOOST_net_10572;
wire g64245_db;
wire g64245_sb;
wire TIMEBOOST_net_10573;
wire g64246_db;
wire g64246_sb;
wire g64247_da;
wire g64247_db;
wire g64247_sb;
wire TIMEBOOST_net_10575;
wire g64248_db;
wire g64248_sb;
wire TIMEBOOST_net_10576;
wire g64250_db;
wire g64250_sb;
wire TIMEBOOST_net_10577;
wire g64251_db;
wire g64251_sb;
wire TIMEBOOST_net_10578;
wire g64252_db;
wire g64252_sb;
wire g64253_da;
wire g64253_db;
wire g64253_sb;
wire TIMEBOOST_net_3452;
wire g64254_db;
wire g64254_sb;
wire TIMEBOOST_net_12341;
wire TIMEBOOST_net_4021;
wire g64255_sb;
wire TIMEBOOST_net_13376;
wire g64256_db;
wire g64256_sb;
wire TIMEBOOST_net_10579;
wire g64257_db;
wire g64257_sb;
wire TIMEBOOST_net_4523;
wire g64258_db;
wire g64258_sb;
wire TIMEBOOST_net_10580;
wire g64259_db;
wire g64259_sb;
wire TIMEBOOST_net_10535;
wire g64260_db;
wire g64260_sb;
wire g64261_da;
wire g64261_db;
wire g64261_sb;
wire g64262_da;
wire g64262_db;
wire g64262_sb;
wire TIMEBOOST_net_10564;
wire g64263_db;
wire g64263_sb;
wire TIMEBOOST_net_10565;
wire g64264_db;
wire g64264_sb;
wire TIMEBOOST_net_10574;
wire g64265_db;
wire g64265_sb;
wire TIMEBOOST_net_10639;
wire g64266_db;
wire g64266_sb;
wire g64267_da;
wire g64267_db;
wire g64267_sb;
wire TIMEBOOST_net_10233;
wire g64268_db;
wire g64268_sb;
wire g64269_da;
wire g64269_db;
wire g64269_sb;
wire TIMEBOOST_net_10234;
wire g64270_db;
wire g64270_sb;
wire TIMEBOOST_net_10247;
wire g64271_db;
wire g64271_sb;
wire g64272_da;
wire g64272_db;
wire g64272_sb;
wire g64273_da;
wire g64273_db;
wire g64273_sb;
wire g64274_da;
wire g64274_db;
wire g64274_sb;
wire TIMEBOOST_net_10251;
wire g64275_db;
wire g64275_sb;
wire TIMEBOOST_net_10252;
wire g64276_db;
wire g64276_sb;
wire g64277_da;
wire g64277_db;
wire g64277_sb;
wire g64278_da;
wire g64278_db;
wire g64278_sb;
wire TIMEBOOST_net_10253;
wire g64279_db;
wire g64279_sb;
wire TIMEBOOST_net_10254;
wire g64280_db;
wire g64280_sb;
wire g64281_da;
wire g64281_db;
wire g64281_sb;
wire TIMEBOOST_net_10255;
wire g64282_db;
wire g64282_sb;
wire TIMEBOOST_net_10642;
wire g64283_db;
wire g64283_sb;
wire g64284_da;
wire g64284_db;
wire g64284_sb;
wire TIMEBOOST_net_10256;
wire g64285_db;
wire g64285_sb;
wire TIMEBOOST_net_223;
wire TIMEBOOST_net_3331;
wire g64286_sb;
wire g64287_db;
wire g64287_sb;
wire g64288_da;
wire g64288_db;
wire g64288_sb;
wire g64289_db;
wire g64289_sb;
wire g64290_da;
wire g64290_db;
wire g64290_sb;
wire g64291_da;
wire g64291_db;
wire g64291_sb;
wire g64292_db;
wire g64292_sb;
wire g64293_da;
wire g64293_db;
wire g64293_sb;
wire TIMEBOOST_net_167;
wire TIMEBOOST_net_3038;
wire g64295_da;
wire g64295_db;
wire g64295_sb;
wire TIMEBOOST_net_3453;
wire g64296_db;
wire g64296_sb;
wire TIMEBOOST_net_10643;
wire g64297_db;
wire g64297_sb;
wire g64298_db;
wire g64298_sb;
wire TIMEBOOST_net_4527;
wire g64300_db;
wire g64300_sb;
wire TIMEBOOST_net_10222;
wire g64301_db;
wire g64301_sb;
wire g64302_da;
wire g64302_db;
wire g64302_sb;
wire TIMEBOOST_net_168;
wire TIMEBOOST_net_14040;
wire TIMEBOOST_net_10223;
wire g64304_db;
wire g64304_sb;
wire TIMEBOOST_net_224;
wire TIMEBOOST_net_3332;
wire g64306_da;
wire g64306_db;
wire g64306_sb;
wire g64307_da;
wire g64307_db;
wire g64307_sb;
wire TIMEBOOST_net_10644;
wire g64308_db;
wire g64308_sb;
wire g64309_da;
wire g64309_db;
wire g64309_sb;
wire g64310_da;
wire g64310_db;
wire g64310_sb;
wire TIMEBOOST_net_4529;
wire g64311_db;
wire g64311_sb;
wire TIMEBOOST_net_10648;
wire g64312_db;
wire g64312_sb;
wire TIMEBOOST_net_10649;
wire g64313_db;
wire g64313_sb;
wire TIMEBOOST_net_10651;
wire g64314_db;
wire g64314_sb;
wire TIMEBOOST_net_9542;
wire g64315_db;
wire g64315_sb;
wire g64316_da;
wire g64316_db;
wire g64316_sb;
wire TIMEBOOST_net_10224;
wire g64317_db;
wire g64317_sb;
wire TIMEBOOST_net_10653;
wire g64318_db;
wire g64318_sb;
wire TIMEBOOST_net_4534;
wire g64319_db;
wire g64319_sb;
wire g64320_da;
wire g64320_db;
wire g64320_sb;
wire g64321_da;
wire g64321_db;
wire g64321_sb;
wire TIMEBOOST_net_13710;
wire g64322_db;
wire g64322_sb;
wire TIMEBOOST_net_4536;
wire g64323_db;
wire g64323_sb;
wire g64324_da;
wire g64324_db;
wire g64324_sb;
wire TIMEBOOST_net_4537;
wire g64325_db;
wire g64325_sb;
wire TIMEBOOST_net_4538;
wire g64326_db;
wire g64326_sb;
wire TIMEBOOST_net_9798;
wire g64327_db;
wire g64327_sb;
wire TIMEBOOST_net_13654;
wire TIMEBOOST_net_15006;
wire g64328_sb;
wire g64329_da;
wire g64329_db;
wire g64329_sb;
wire g64330_da;
wire g64330_db;
wire g64330_sb;
wire g64331_da;
wire g64331_db;
wire g64331_sb;
wire TIMEBOOST_net_10533;
wire g64332_db;
wire g64332_sb;
wire TIMEBOOST_net_9831;
wire g64333_db;
wire g64333_sb;
wire TIMEBOOST_net_9832;
wire g64334_db;
wire g64334_sb;
wire TIMEBOOST_net_9833;
wire g64335_db;
wire g64335_sb;
wire TIMEBOOST_net_3459;
wire g64336_db;
wire g64336_sb;
wire TIMEBOOST_net_10534;
wire g64337_db;
wire g64337_sb;
wire TIMEBOOST_net_10536;
wire g64339_db;
wire g64339_sb;
wire g64340_da;
wire g64340_db;
wire g64340_sb;
wire TIMEBOOST_net_10537;
wire g64341_db;
wire g64341_sb;
wire TIMEBOOST_net_10541;
wire g64342_db;
wire g64342_sb;
wire g64343_da;
wire g64343_db;
wire g64343_sb;
wire TIMEBOOST_net_13766;
wire g64344_db;
wire g64344_sb;
wire g64345_da;
wire g64345_db;
wire g64345_sb;
wire TIMEBOOST_net_10225;
wire g64346_db;
wire g64346_sb;
wire TIMEBOOST_net_10542;
wire g64347_db;
wire g64347_sb;
wire g64348_da;
wire g64348_db;
wire g64348_sb;
wire g64349_da;
wire g64349_db;
wire g64349_sb;
wire g64350_da;
wire g64350_db;
wire g64350_sb;
wire TIMEBOOST_net_9850;
wire TIMEBOOST_net_14698;
wire g64351_sb;
wire g64352_da;
wire g64352_db;
wire g64352_sb;
wire TIMEBOOST_net_9851;
wire g64353_db;
wire g64353_sb;
wire g64354_da;
wire g64354_db;
wire g64354_sb;
wire TIMEBOOST_net_12601;
wire g64355_sb;
wire g64356_da;
wire g64356_db;
wire g64356_sb;
wire TIMEBOOST_net_3463;
wire g64357_db;
wire g64357_sb;
wire g64358_da;
wire g64358_db;
wire g64358_sb;
wire TIMEBOOST_net_3464;
wire g64359_db;
wire g64359_sb;
wire TIMEBOOST_net_3465;
wire g64360_db;
wire g64360_sb;
wire TIMEBOOST_net_9852;
wire g64361_db;
wire g64361_sb;
wire TIMEBOOST_net_3467;
wire g64362_db;
wire g64362_sb;
wire TIMEBOOST_net_13840;
wire g64363_db;
wire g64363_sb;
wire TIMEBOOST_net_155;
wire TIMEBOOST_net_12622;
wire g64366_da;
wire g64366_db;
wire g64366_sb;
wire g64367_da;
wire g64367_db;
wire g64367_sb;
wire g64368_p;
wire g64369_p;
wire g64370_p;
wire g64371_p;
wire g64375_p;
wire g64376_p;
wire g64377_p;
wire g64378_p;
wire g64379_p;
wire g64380_p;
wire TIMEBOOST_net_14754;
wire g64382_p;
wire g64383_p;
wire g64384_p;
wire g64385_p;
wire g64454_p;
wire g64461_p;
wire g64465_p;
wire g64466_p;
wire g64577_p;
wire g64578_p;
wire g64581_p;
wire g64582_p;
wire g64585_p;
wire g64587_p;
wire g64595_p;
wire g64596_p;
wire g64597_p;
wire g64610_p;
wire g66420_db;
wire g64630_BP;
wire g64630_p;
wire g64631_p;
wire g64632_p;
wire g64633_p;
wire g64639_p;
wire g64643_p;
wire g64646_p;
wire g64671_p;
wire g64678_p;
wire g64687_p;
wire g64694_p;
wire g64697_p;
wire g64700_p;
wire g64701_p;
wire g64702_p;
wire g64704_p;
wire g64705_p;
wire g64707_p;
wire g64712_p;
wire g64727_p;
wire g64736_p;
wire g64740_p;
wire g64746_p;
wire g64747_p;
wire TIMEBOOST_net_3519;
wire g64748_db;
wire g64748_sb;
wire TIMEBOOST_net_3469;
wire TIMEBOOST_net_12528;
wire g64749_sb;
wire TIMEBOOST_net_341;
wire TIMEBOOST_net_12579;
wire g64750_sb;
wire TIMEBOOST_net_13768;
wire g64751_db;
wire g64751_sb;
wire TIMEBOOST_net_3470;
wire TIMEBOOST_net_13509;
wire g64752_sb;
wire TIMEBOOST_net_12868;
wire g64753_db;
wire g64753_sb;
wire TIMEBOOST_net_3231;
wire g64754_db;
wire g64754_sb;
wire TIMEBOOST_net_9918;
wire g64755_db;
wire g64755_sb;
wire TIMEBOOST_net_12867;
wire g64756_db;
wire g64756_sb;
wire TIMEBOOST_net_4022;
wire g64757_db;
wire g64757_sb;
wire TIMEBOOST_net_9919;
wire g64758_db;
wire g64758_sb;
wire TIMEBOOST_net_12597;
wire g64759_db;
wire g64759_sb;
wire TIMEBOOST_net_4616;
wire g64760_db;
wire g64760_sb;
wire TIMEBOOST_net_9920;
wire g64761_db;
wire g64761_sb;
wire TIMEBOOST_net_9817;
wire g64762_db;
wire g64762_sb;
wire TIMEBOOST_net_4617;
wire g64763_db;
wire g64763_sb;
wire TIMEBOOST_net_9818;
wire TIMEBOOST_net_12575;
wire g64764_sb;
wire TIMEBOOST_net_209;
wire TIMEBOOST_net_9640;
wire g64765_sb;
wire TIMEBOOST_net_12448;
wire g64766_sb;
wire TIMEBOOST_net_210;
wire g64767_db;
wire g64767_sb;
wire TIMEBOOST_net_9823;
wire g64768_db;
wire g64768_sb;
wire TIMEBOOST_net_12596;
wire g64769_db;
wire g64769_sb;
wire TIMEBOOST_net_10199;
wire g64770_db;
wire g64770_sb;
wire TIMEBOOST_net_192;
wire g64771_sb;
wire TIMEBOOST_net_9566;
wire g64772_db;
wire g64772_sb;
wire TIMEBOOST_net_4019;
wire TIMEBOOST_net_3131;
wire g64773_sb;
wire TIMEBOOST_net_10201;
wire g64774_db;
wire g64774_sb;
wire TIMEBOOST_net_193;
wire TIMEBOOST_net_12574;
wire g64775_sb;
wire TIMEBOOST_net_9567;
wire g64776_db;
wire g64776_sb;
wire TIMEBOOST_net_10202;
wire g64777_db;
wire g64777_sb;
wire TIMEBOOST_net_194;
wire TIMEBOOST_net_12570;
wire g64778_sb;
wire TIMEBOOST_net_3523;
wire g64779_db;
wire g64779_sb;
wire TIMEBOOST_net_12886;
wire g64780_db;
wire g64780_sb;
wire TIMEBOOST_net_9568;
wire g64781_db;
wire g64781_sb;
wire TIMEBOOST_net_13187;
wire g64782_db;
wire g64782_sb;
wire TIMEBOOST_net_13186;
wire g64783_db;
wire g64783_sb;
wire TIMEBOOST_net_13657;
wire g64784_db;
wire g64784_sb;
wire TIMEBOOST_net_13185;
wire g64785_db;
wire g64785_sb;
wire TIMEBOOST_net_13656;
wire g64786_db;
wire g64786_sb;
wire TIMEBOOST_net_195;
wire TIMEBOOST_net_12569;
wire g64787_sb;
wire TIMEBOOST_net_12435;
wire g64788_db;
wire g64788_sb;
wire TIMEBOOST_net_3524;
wire g64789_db;
wire g64789_sb;
wire TIMEBOOST_net_3525;
wire g64790_db;
wire g64790_sb;
wire TIMEBOOST_net_12436;
wire g64791_db;
wire g64791_sb;
wire TIMEBOOST_net_3526;
wire g64792_db;
wire g64792_sb;
wire TIMEBOOST_net_9921;
wire g64793_db;
wire g64793_sb;
wire TIMEBOOST_net_12364;
wire TIMEBOOST_net_12450;
wire g64794_sb;
wire TIMEBOOST_net_3528;
wire g64795_db;
wire g64795_sb;
wire TIMEBOOST_net_3841;
wire g64796_db;
wire g64796_sb;
wire TIMEBOOST_net_196;
wire TIMEBOOST_net_12571;
wire g64797_sb;
wire TIMEBOOST_net_12780;
wire g64798_db;
wire g64798_sb;
wire TIMEBOOST_net_9650;
wire g64799_db;
wire g64799_sb;
wire TIMEBOOST_net_13764;
wire g64800_db;
wire g64800_sb;
wire TIMEBOOST_net_3529;
wire g64801_db;
wire g64801_sb;
wire TIMEBOOST_net_9922;
wire g64802_db;
wire g64802_sb;
wire TIMEBOOST_net_9923;
wire g64803_db;
wire g64803_sb;
wire TIMEBOOST_net_9924;
wire g64804_db;
wire g64804_sb;
wire TIMEBOOST_net_12927;
wire g64805_db;
wire g64805_sb;
wire TIMEBOOST_net_12932;
wire g64806_db;
wire g64806_sb;
wire TIMEBOOST_net_13769;
wire g64807_db;
wire g64807_sb;
wire TIMEBOOST_net_12779;
wire g64808_db;
wire g64808_sb;
wire TIMEBOOST_net_9569;
wire g64809_db;
wire g64809_sb;
wire TIMEBOOST_net_12485;
wire g64810_db;
wire g64810_sb;
wire TIMEBOOST_net_12876;
wire TIMEBOOST_net_12529;
wire g64811_sb;
wire TIMEBOOST_net_9774;
wire g64812_db;
wire g64812_sb;
wire TIMEBOOST_net_157;
wire g64813_db;
wire g64813_sb;
wire TIMEBOOST_net_187;
wire g64814_db;
wire g64814_sb;
wire TIMEBOOST_net_219;
wire g64815_db;
wire g64815_sb;
wire TIMEBOOST_net_197;
wire TIMEBOOST_net_9593;
wire g64816_sb;
wire TIMEBOOST_net_3471;
wire g64817_db;
wire g64817_sb;
wire TIMEBOOST_net_13575;
wire g64818_db;
wire g64818_sb;
wire TIMEBOOST_net_3306;
wire g64819_db;
wire g64819_sb;
wire TIMEBOOST_net_9856;
wire g64820_db;
wire g64820_sb;
wire TIMEBOOST_net_220;
wire g64821_db;
wire g64821_sb;
wire TIMEBOOST_net_3472;
wire g64822_db;
wire g64822_sb;
wire TIMEBOOST_net_13839;
wire g64823_db;
wire g64823_sb;
wire TIMEBOOST_net_9885;
wire g64824_db;
wire g64824_sb;
wire TIMEBOOST_net_13672;
wire g64825_db;
wire g64825_sb;
wire TIMEBOOST_net_12880;
wire g64826_db;
wire g64826_sb;
wire TIMEBOOST_net_10446;
wire TIMEBOOST_net_13340;
wire g64827_sb;
wire TIMEBOOST_net_13579;
wire g64828_db;
wire g64828_sb;
wire TIMEBOOST_net_9654;
wire g64829_db;
wire g64829_sb;
wire TIMEBOOST_net_9558;
wire TIMEBOOST_net_12406;
wire g64830_sb;
wire TIMEBOOST_net_10447;
wire g64831_db;
wire g64831_sb;
wire TIMEBOOST_net_10448;
wire g64832_db;
wire g64832_sb;
wire TIMEBOOST_net_12375;
wire g64833_db;
wire g64833_sb;
wire TIMEBOOST_net_10634;
wire g64834_db;
wire g64834_sb;
wire TIMEBOOST_net_10449;
wire TIMEBOOST_net_12233;
wire g64835_sb;
wire TIMEBOOST_net_13093;
wire g64836_db;
wire g64836_sb;
wire TIMEBOOST_net_10162;
wire g64837_db;
wire g64837_sb;
wire TIMEBOOST_net_3539;
wire g64838_db;
wire g64838_sb;
wire TIMEBOOST_net_3540;
wire g64839_db;
wire g64839_sb;
wire TIMEBOOST_net_9655;
wire g64840_db;
wire g64840_sb;
wire TIMEBOOST_net_198;
wire g64841_db;
wire g64841_sb;
wire TIMEBOOST_net_12491;
wire g64842_db;
wire g64842_sb;
wire TIMEBOOST_net_9887;
wire TIMEBOOST_net_12531;
wire g64843_sb;
wire TIMEBOOST_net_3844;
wire g64844_db;
wire g64844_sb;
wire TIMEBOOST_net_12492;
wire g64845_db;
wire g64845_sb;
wire TIMEBOOST_net_12493;
wire g64846_db;
wire g64846_sb;
wire TIMEBOOST_net_9888;
wire g64847_db;
wire g64847_sb;
wire TIMEBOOST_net_9889;
wire g64848_db;
wire g64848_sb;
wire TIMEBOOST_net_3479;
wire g64849_db;
wire g64849_sb;
wire TIMEBOOST_net_10543;
wire TIMEBOOST_net_12230;
wire g64850_sb;
wire TIMEBOOST_net_10164;
wire g64851_db;
wire g64851_sb;
wire TIMEBOOST_net_12494;
wire TIMEBOOST_net_258;
wire g64852_sb;
wire TIMEBOOST_net_3545;
wire g64853_db;
wire g64853_sb;
wire TIMEBOOST_net_3546;
wire TIMEBOOST_net_12532;
wire g64854_sb;
wire TIMEBOOST_net_9890;
wire g64855_db;
wire g64855_sb;
wire TIMEBOOST_net_3481;
wire TIMEBOOST_net_13510;
wire g64856_sb;
wire TIMEBOOST_net_3482;
wire g64857_db;
wire g64857_sb;
wire TIMEBOOST_net_9826;
wire g64858_db;
wire g64858_sb;
wire TIMEBOOST_net_10165;
wire g64859_db;
wire g64859_sb;
wire TIMEBOOST_net_10105;
wire g64860_db;
wire g64860_sb;
wire TIMEBOOST_net_12610;
wire g64861_db;
wire g64861_sb;
wire TIMEBOOST_net_13701;
wire g64862_db;
wire g64862_sb;
wire TIMEBOOST_net_10022;
wire g64863_db;
wire g64863_sb;
wire TIMEBOOST_net_4618;
wire g64864_db;
wire g64864_sb;
wire TIMEBOOST_net_10023;
wire g64865_db;
wire g64865_sb;
wire TIMEBOOST_net_15190;
wire g64866_db;
wire g64866_sb;
wire TIMEBOOST_net_4619;
wire g64867_db;
wire g64867_sb;
wire TIMEBOOST_net_14566;
wire TIMEBOOST_net_12576;
wire g64868_sb;
wire TIMEBOOST_net_4620;
wire g64869_db;
wire g64869_sb;
wire TIMEBOOST_net_4621;
wire g64870_db;
wire g64870_sb;
wire TIMEBOOST_net_9820;
wire g64871_db;
wire g64871_sb;
wire TIMEBOOST_net_12878;
wire g64872_db;
wire g64872_sb;
wire TIMEBOOST_net_10676;
wire g64873_db;
wire g64873_sb;
wire TIMEBOOST_net_13374;
wire g64874_db;
wire g64874_sb;
wire TIMEBOOST_net_3547;
wire g64875_db;
wire g64875_sb;
wire TIMEBOOST_net_211;
wire g64876_db;
wire g64876_sb;
wire TIMEBOOST_net_14670;
wire TIMEBOOST_net_3293;
wire g64877_sb;
wire TIMEBOOST_net_3363;
wire TIMEBOOST_net_12452;
wire g64878_sb;
wire TIMEBOOST_net_3483;
wire TIMEBOOST_net_12533;
wire g64879_sb;
wire TIMEBOOST_net_3484;
wire TIMEBOOST_net_12534;
wire g64880_sb;
wire TIMEBOOST_net_12865;
wire TIMEBOOST_net_12535;
wire g64881_sb;
wire TIMEBOOST_net_3548;
wire g64882_db;
wire g64882_sb;
wire TIMEBOOST_net_9891;
wire g64883_db;
wire g64883_sb;
wire TIMEBOOST_net_13838;
wire g64884_db;
wire g64884_sb;
wire TIMEBOOST_net_9914;
wire g64885_db;
wire g64885_sb;
wire TIMEBOOST_net_10192;
wire g64886_db;
wire g64886_sb;
wire TIMEBOOST_net_13837;
wire TIMEBOOST_net_12537;
wire g64887_sb;
wire TIMEBOOST_net_3488;
wire g64888_db;
wire g64888_sb;
wire TIMEBOOST_net_3850;
wire g64889_db;
wire g64889_sb;
wire TIMEBOOST_net_3550;
wire g64890_db;
wire g64890_sb;
wire TIMEBOOST_net_3551;
wire g64891_db;
wire g64891_sb;
wire TIMEBOOST_net_3552;
wire g64892_db;
wire g64892_sb;
wire TIMEBOOST_net_10206;
wire TIMEBOOST_net_12539;
wire g64893_sb;
wire TIMEBOOST_net_12746;
wire TIMEBOOST_net_12540;
wire g64894_sb;
wire TIMEBOOST_net_12745;
wire g64895_db;
wire g64895_sb;
wire TIMEBOOST_net_9589;
wire g64896_db;
wire g64896_sb;
wire TIMEBOOST_net_9896;
wire g64897_db;
wire g64897_sb;
wire TIMEBOOST_net_13860;
wire g64898_db;
wire g64898_sb;
wire TIMEBOOST_net_3310;
wire g64899_db;
wire g64899_sb;
wire TIMEBOOST_net_3311;
wire g64900_db;
wire g64900_sb;
wire TIMEBOOST_net_3553;
wire g64901_db;
wire g64901_sb;
wire TIMEBOOST_net_12536;
wire g64902_db;
wire g64902_sb;
wire TIMEBOOST_net_12401;
wire g64903_db;
wire g64903_sb;
wire TIMEBOOST_net_3277;
wire TIMEBOOST_net_12415;
wire g64904_sb;
wire TIMEBOOST_net_13581;
wire g64905_db;
wire g64905_sb;
wire TIMEBOOST_net_9664;
wire g64906_db;
wire g64906_sb;
wire TIMEBOOST_net_13213;
wire g64907_db;
wire g64907_sb;
wire TIMEBOOST_net_3556;
wire g64908_db;
wire g64908_sb;
wire TIMEBOOST_net_3557;
wire g64909_db;
wire g64909_sb;
wire TIMEBOOST_net_3558;
wire g64910_db;
wire g64910_sb;
wire TIMEBOOST_net_9928;
wire g64911_db;
wire g64911_sb;
wire TIMEBOOST_net_3560;
wire g64912_db;
wire g64912_sb;
wire TIMEBOOST_net_9929;
wire g64913_db;
wire g64913_sb;
wire TIMEBOOST_net_3562;
wire g64914_db;
wire g64914_sb;
wire TIMEBOOST_net_3315;
wire g64915_db;
wire g64915_sb;
wire TIMEBOOST_net_3316;
wire TIMEBOOST_net_12420;
wire g64916_sb;
wire TIMEBOOST_net_13373;
wire g64917_db;
wire g64917_sb;
wire TIMEBOOST_net_9898;
wire TIMEBOOST_net_12541;
wire g64918_sb;
wire TIMEBOOST_net_10450;
wire g64919_db;
wire g64919_sb;
wire TIMEBOOST_net_9559;
wire TIMEBOOST_net_9794;
wire g64920_sb;
wire TIMEBOOST_net_10207;
wire g64921_db;
wire g64921_sb;
wire TIMEBOOST_net_13580;
wire g64922_db;
wire g64922_sb;
wire TIMEBOOST_net_9899;
wire TIMEBOOST_net_12542;
wire g64923_sb;
wire TIMEBOOST_net_12264;
wire TIMEBOOST_net_12845;
wire g64924_sb;
wire TIMEBOOST_net_9825;
wire g64925_db;
wire g64925_sb;
wire TIMEBOOST_net_9746;
wire g64926_db;
wire g64926_sb;
wire TIMEBOOST_net_10208;
wire g64927_db;
wire g64927_sb;
wire TIMEBOOST_net_9900;
wire g64928_db;
wire g64928_sb;
wire TIMEBOOST_net_9901;
wire g64929_db;
wire g64929_sb;
wire TIMEBOOST_net_3497;
wire g64930_db;
wire g64930_sb;
wire TIMEBOOST_net_9769;
wire g64931_db;
wire g64931_sb;
wire TIMEBOOST_net_3566;
wire g64932_db;
wire g64932_sb;
wire TIMEBOOST_net_9969;
wire g64933_db;
wire g64933_sb;
wire TIMEBOOST_net_9970;
wire g64934_db;
wire g64934_sb;
wire TIMEBOOST_net_9971;
wire g64935_db;
wire g64935_sb;
wire TIMEBOOST_net_9902;
wire TIMEBOOST_net_12543;
wire g64936_sb;
wire TIMEBOOST_net_3570;
wire g64937_db;
wire g64937_sb;
wire TIMEBOOST_net_9903;
wire g64938_db;
wire g64938_sb;
wire TIMEBOOST_net_9904;
wire TIMEBOOST_net_13563;
wire g64939_sb;
wire TIMEBOOST_net_3571;
wire g64940_db;
wire g64940_sb;
wire TIMEBOOST_net_15082;
wire g64941_db;
wire g64941_sb;
wire TIMEBOOST_net_10330;
wire g64942_db;
wire g64942_sb;
wire TIMEBOOST_net_4027;
wire TIMEBOOST_net_12714;
wire g64943_sb;
wire TIMEBOOST_net_10347;
wire g64944_db;
wire g64944_sb;
wire TIMEBOOST_net_10348;
wire g64945_db;
wire g64945_sb;
wire TIMEBOOST_net_4030;
wire g64946_db;
wire g64946_sb;
wire TIMEBOOST_net_4031;
wire g64947_db;
wire g64947_sb;
wire g64948_da;
wire g64948_db;
wire g64948_sb;
wire TIMEBOOST_net_4032;
wire g64949_db;
wire g64949_sb;
wire TIMEBOOST_net_4033;
wire g64950_db;
wire g64950_sb;
wire TIMEBOOST_net_4034;
wire g64951_db;
wire g64951_sb;
wire TIMEBOOST_net_10349;
wire g64952_db;
wire g64952_sb;
wire TIMEBOOST_net_199;
wire g64953_db;
wire g64953_sb;
wire TIMEBOOST_net_10350;
wire g64954_db;
wire g64954_sb;
wire TIMEBOOST_net_4037;
wire TIMEBOOST_net_12715;
wire g64955_sb;
wire TIMEBOOST_net_4038;
wire g64956_db;
wire g64956_sb;
wire TIMEBOOST_net_4039;
wire g64957_db;
wire g64957_sb;
wire TIMEBOOST_net_4040;
wire g64958_db;
wire g64958_sb;
wire TIMEBOOST_net_13470;
wire g64959_db;
wire g64959_sb;
wire g64960_da;
wire g64960_db;
wire g64960_sb;
wire TIMEBOOST_net_15189;
wire g64961_db;
wire g64961_sb;
wire TIMEBOOST_net_213;
wire TIMEBOOST_net_9641;
wire g64962_sb;
wire TIMEBOOST_net_3758;
wire g64963_db;
wire g64963_sb;
wire TIMEBOOST_net_3572;
wire g64964_db;
wire TIMEBOOST_net_10677;
wire TIMEBOOST_net_13098;
wire g64965_sb;
wire TIMEBOOST_net_13191;
wire g64966_db;
wire g64966_sb;
wire TIMEBOOST_net_3759;
wire g64967_db;
wire g64967_sb;
wire TIMEBOOST_net_3760;
wire g64968_db;
wire g64968_sb;
wire TIMEBOOST_net_13859;
wire g64969_db;
wire g64969_sb;
wire TIMEBOOST_net_10194;
wire g64970_db;
wire g64970_sb;
wire TIMEBOOST_net_10024;
wire g64971_db;
wire g64971_sb;
wire TIMEBOOST_net_4624;
wire TIMEBOOST_net_10203;
wire g64972_sb;
wire TIMEBOOST_net_4625;
wire TIMEBOOST_net_13099;
wire g64973_sb;
wire TIMEBOOST_net_4041;
wire g64974_db;
wire g64974_sb;
wire TIMEBOOST_net_3573;
wire g64975_db;
wire g64975_sb;
wire TIMEBOOST_net_3763;
wire g64976_db;
wire g64976_sb;
wire TIMEBOOST_net_9905;
wire g64977_db;
wire g64977_sb;
wire TIMEBOOST_net_9953;
wire g64978_db;
wire g64978_sb;
wire TIMEBOOST_net_9812;
wire g64979_db;
wire g64979_sb;
wire TIMEBOOST_net_3575;
wire g64980_db;
wire g64980_sb;
wire TIMEBOOST_net_14772;
wire g64981_db;
wire TIMEBOOST_net_9972;
wire g64982_db;
wire g64982_sb;
wire TIMEBOOST_net_4042;
wire g64983_db;
wire g64983_sb;
wire g64984_da;
wire g64984_db;
wire g64984_sb;
wire TIMEBOOST_net_13249;
wire g64985_db;
wire g64985_sb;
wire TIMEBOOST_net_12359;
wire g64986_db;
wire g64986_sb;
wire TIMEBOOST_net_3577;
wire g64987_db;
wire g64987_sb;
wire TIMEBOOST_net_4043;
wire g64988_db;
wire g64988_sb;
wire TIMEBOOST_net_3578;
wire g64989_db;
wire g64989_sb;
wire TIMEBOOST_net_10195;
wire g64990_db;
wire g64990_sb;
wire TIMEBOOST_net_10544;
wire g64991_db;
wire g64991_sb;
wire TIMEBOOST_net_9906;
wire g64992_db;
wire g64992_sb;
wire TIMEBOOST_net_3579;
wire g64993_db;
wire g64993_sb;
wire TIMEBOOST_net_9907;
wire g64994_db;
wire g64994_sb;
wire TIMEBOOST_net_3580;
wire g64995_db;
wire g64995_sb;
wire TIMEBOOST_net_3581;
wire g64996_db;
wire g64996_sb;
wire TIMEBOOST_net_3582;
wire g64997_db;
wire g64997_sb;
wire TIMEBOOST_net_9908;
wire g64998_db;
wire g64998_sb;
wire TIMEBOOST_net_3856;
wire g64999_db;
wire g64999_sb;
wire TIMEBOOST_net_10545;
wire g65000_db;
wire g65000_sb;
wire TIMEBOOST_net_3857;
wire g65001_db;
wire g65001_sb;
wire TIMEBOOST_net_10343;
wire g65002_db;
wire g65002_sb;
wire TIMEBOOST_net_3583;
wire g65003_db;
wire g65003_sb;
wire TIMEBOOST_net_9714;
wire TIMEBOOST_net_12453;
wire g65004_sb;
wire TIMEBOOST_net_3584;
wire g65005_db;
wire g65005_sb;
wire TIMEBOOST_net_14120;
wire g65006_db;
wire g65006_sb;
wire TIMEBOOST_net_10161;
wire g65007_db;
wire g65007_sb;
wire TIMEBOOST_net_14170;
wire g65008_db;
wire g65008_sb;
wire TIMEBOOST_net_10344;
wire g65009_db;
wire g65009_sb;
wire TIMEBOOST_net_3317;
wire g65010_db;
wire g65010_sb;
wire TIMEBOOST_net_4407;
wire g65011_db;
wire g65011_sb;
wire TIMEBOOST_net_3587;
wire g65012_db;
wire g65012_sb;
wire TIMEBOOST_net_3588;
wire g65013_db;
wire g65013_sb;
wire TIMEBOOST_net_10345;
wire g65014_db;
wire g65014_sb;
wire TIMEBOOST_net_10547;
wire g65015_db;
wire g65015_sb;
wire TIMEBOOST_net_3318;
wire g65016_db;
wire g65016_sb;
wire TIMEBOOST_net_4047;
wire g65017_db;
wire g65017_sb;
wire TIMEBOOST_net_9909;
wire g65018_db;
wire g65018_sb;
wire TIMEBOOST_net_14108;
wire g65019_db;
wire g65019_sb;
wire TIMEBOOST_net_201;
wire g65020_db;
wire g65020_sb;
wire TIMEBOOST_net_3319;
wire g65021_db;
wire g65021_sb;
wire TIMEBOOST_net_9910;
wire g65022_db;
wire g65022_sb;
wire TIMEBOOST_net_4408;
wire g65023_db;
wire g65023_sb;
wire TIMEBOOST_net_3320;
wire g65024_db;
wire g65024_sb;
wire TIMEBOOST_net_12882;
wire g65025_db;
wire g65025_sb;
wire TIMEBOOST_net_3321;
wire TIMEBOOST_net_12421;
wire g65026_sb;
wire TIMEBOOST_net_202;
wire TIMEBOOST_net_12469;
wire g65027_sb;
wire TIMEBOOST_net_9941;
wire g65028_db;
wire g65028_sb;
wire TIMEBOOST_net_3591;
wire g65029_db;
wire g65029_sb;
wire TIMEBOOST_net_3322;
wire g65030_db;
wire g65030_sb;
wire TIMEBOOST_net_13105;
wire g65031_db;
wire g65031_sb;
wire TIMEBOOST_net_12884;
wire g65032_db;
wire g65032_sb;
wire TIMEBOOST_net_3593;
wire TIMEBOOST_net_12422;
wire g65033_sb;
wire TIMEBOOST_net_3594;
wire g65034_db;
wire g65034_sb;
wire TIMEBOOST_net_10451;
wire g65035_db;
wire g65035_sb;
wire TIMEBOOST_net_9813;
wire g65036_db;
wire g65036_sb;
wire TIMEBOOST_net_3595;
wire g65037_db;
wire g65037_sb;
wire TIMEBOOST_net_14161;
wire TIMEBOOST_net_12423;
wire g65038_sb;
wire TIMEBOOST_net_13845;
wire g65039_db;
wire g65039_sb;
wire TIMEBOOST_net_10452;
wire g65040_db;
wire g65040_sb;
wire TIMEBOOST_net_3861;
wire g65041_db;
wire g65041_sb;
wire TIMEBOOST_net_10346;
wire g65042_db;
wire g65042_sb;
wire TIMEBOOST_net_4409;
wire g65043_db;
wire g65043_sb;
wire TIMEBOOST_net_3323;
wire g65044_db;
wire g65044_sb;
wire TIMEBOOST_net_10456;
wire g65045_db;
wire g65045_sb;
wire TIMEBOOST_net_14121;
wire g65046_db;
wire g65046_sb;
wire TIMEBOOST_net_13210;
wire g65047_db;
wire g65047_sb;
wire TIMEBOOST_net_13183;
wire g65048_db;
wire g65048_sb;
wire TIMEBOOST_net_9979;
wire g65049_db;
wire g65049_sb;
wire TIMEBOOST_net_9911;
wire g65050_db;
wire g65050_sb;
wire TIMEBOOST_net_12969;
wire g65051_db;
wire g65051_sb;
wire TIMEBOOST_net_3600;
wire g65052_db;
wire g65052_sb;
wire TIMEBOOST_net_10181;
wire g65053_db;
wire g65053_sb;
wire TIMEBOOST_net_9814;
wire g65054_db;
wire g65054_sb;
wire TIMEBOOST_net_214;
wire TIMEBOOST_net_9649;
wire g65055_sb;
wire TIMEBOOST_net_10183;
wire g65056_db;
wire g65056_sb;
wire TIMEBOOST_net_3172;
wire g65057_db;
wire g65057_sb;
wire TIMEBOOST_net_9816;
wire g65058_db;
wire g65058_sb;
wire TIMEBOOST_net_9819;
wire g65059_db;
wire g65059_sb;
wire TIMEBOOST_net_3367;
wire g65060_db;
wire g65060_sb;
wire TIMEBOOST_net_12619;
wire g65061_db;
wire g65061_sb;
wire TIMEBOOST_net_13773;
wire g65062_db;
wire g65062_sb;
wire TIMEBOOST_net_3601;
wire g65063_db;
wire g65063_sb;
wire TIMEBOOST_net_13747;
wire g65064_db;
wire g65064_sb;
wire TIMEBOOST_net_3602;
wire g65065_db;
wire g65065_sb;
wire TIMEBOOST_net_13772;
wire g65066_db;
wire g65066_sb;
wire TIMEBOOST_net_15191;
wire g65067_db;
wire g65067_sb;
wire TIMEBOOST_net_14064;
wire TIMEBOOST_net_9651;
wire g65068_sb;
wire TIMEBOOST_net_12486;
wire g65069_db;
wire g65069_sb;
wire TIMEBOOST_net_3368;
wire TIMEBOOST_net_12454;
wire g65070_sb;
wire TIMEBOOST_net_9947;
wire g65071_db;
wire g65071_sb;
wire TIMEBOOST_net_3604;
wire g65072_db;
wire g65072_sb;
wire TIMEBOOST_net_12736;
wire g65073_db;
wire g65073_sb;
wire TIMEBOOST_net_10209;
wire TIMEBOOST_net_12545;
wire g65074_sb;
wire TIMEBOOST_net_10163;
wire g65075_db;
wire g65075_sb;
wire TIMEBOOST_net_3508;
wire TIMEBOOST_net_12538;
wire g65076_sb;
wire TIMEBOOST_net_12487;
wire g65077_db;
wire g65077_sb;
wire TIMEBOOST_net_13104;
wire g65078_db;
wire g65078_sb;
wire TIMEBOOST_net_12877;
wire g65079_db;
wire g65079_sb;
wire TIMEBOOST_net_13103;
wire g65080_db;
wire g65080_sb;
wire TIMEBOOST_net_3329;
wire g65081_db;
wire g65081_sb;
wire TIMEBOOST_net_13823;
wire g65082_db;
wire g65082_sb;
wire TIMEBOOST_net_13209;
wire g65083_db;
wire g65083_sb;
wire TIMEBOOST_net_13847;
wire g65084_db;
wire g65084_sb;
wire g65085_da;
wire g65085_db;
wire g65085_sb;
wire TIMEBOOST_net_3509;
wire TIMEBOOST_net_12546;
wire g65086_sb;
wire TIMEBOOST_net_9913;
wire TIMEBOOST_net_12547;
wire g65087_sb;
wire TIMEBOOST_net_3610;
wire g65088_db;
wire g65088_sb;
wire TIMEBOOST_net_3611;
wire g65089_db;
wire g65089_sb;
wire TIMEBOOST_net_12737;
wire g65090_db;
wire g65090_sb;
wire TIMEBOOST_net_3369;
wire g65091_db;
wire g65091_sb;
wire TIMEBOOST_net_216;
wire TIMEBOOST_net_9613;
wire g65092_sb;
wire TIMEBOOST_net_4410;
wire g65093_db;
wire g65093_sb;
wire TIMEBOOST_net_3867;
wire g65094_db;
wire g65094_sb;
wire TIMEBOOST_net_12738;
wire g65095_db;
wire g65095_sb;
wire TIMEBOOST_net_12565;
wire TIMEBOOST_net_12301;
wire g65096_sb;
wire TIMEBOOST_net_13846;
wire g65097_db;
wire g65097_sb;
wire TIMEBOOST_net_13528;
wire g65098_db;
wire g65098_sb;
wire TIMEBOOST_net_9571;
wire g65099_db;
wire g65099_sb;
wire TIMEBOOST_net_10305;
wire TIMEBOOST_net_189;
wire g65210_sb;
wire TIMEBOOST_net_225;
wire g65211_db;
wire g65211_sb;
wire TIMEBOOST_net_171;
wire g65212_db;
wire TIMEBOOST_net_3328;
wire g65213_db;
wire g65213_sb;
wire TIMEBOOST_net_3128;
wire TIMEBOOST_net_13543;
wire g65214_sb;
wire TIMEBOOST_net_3965;
wire TIMEBOOST_net_14711;
wire g65215_sb;
wire TIMEBOOST_net_13339;
wire g65216_db;
wire g65216_sb;
wire TIMEBOOST_net_228;
wire TIMEBOOST_net_12515;
wire g65217_sb;
wire TIMEBOOST_net_3230;
wire TIMEBOOST_net_9688;
wire g65218_sb;
wire TIMEBOOST_net_230;
wire TIMEBOOST_net_12449;
wire g65219_sb;
wire TIMEBOOST_net_231;
wire TIMEBOOST_net_12530;
wire g65220_sb;
wire TIMEBOOST_net_232;
wire TIMEBOOST_net_12511;
wire g65221_sb;
wire TIMEBOOST_net_9931;
wire TIMEBOOST_net_9628;
wire g65222_sb;
wire TIMEBOOST_net_9946;
wire TIMEBOOST_net_9629;
wire g65223_sb;
wire TIMEBOOST_net_235;
wire TIMEBOOST_net_3378;
wire g65224_sb;
wire TIMEBOOST_net_236;
wire g65225_db;
wire g65225_sb;
wire TIMEBOOST_net_237;
wire TIMEBOOST_net_3379;
wire g65226_sb;
wire TIMEBOOST_net_238;
wire TIMEBOOST_net_3380;
wire g65227_sb;
wire TIMEBOOST_net_239;
wire TIMEBOOST_net_3381;
wire g65228_sb;
wire TIMEBOOST_net_3713;
wire TIMEBOOST_net_3382;
wire g65229_sb;
wire TIMEBOOST_net_3714;
wire g65230_db;
wire g65230_sb;
wire TIMEBOOST_net_242;
wire TIMEBOOST_net_3383;
wire g65231_sb;
wire TIMEBOOST_net_243;
wire TIMEBOOST_net_13504;
wire g65232_sb;
wire TIMEBOOST_net_244;
wire TIMEBOOST_net_3385;
wire g65233_sb;
wire TIMEBOOST_net_3966;
wire TIMEBOOST_net_14712;
wire TIMEBOOST_net_13391;
wire g65235_db;
wire g65235_sb;
wire TIMEBOOST_net_13389;
wire g65236_db;
wire g65236_sb;
wire TIMEBOOST_net_245;
wire TIMEBOOST_net_3386;
wire g65237_sb;
wire TIMEBOOST_net_246;
wire TIMEBOOST_net_3387;
wire g65238_sb;
wire TIMEBOOST_net_3967;
wire g65239_db;
wire TIMEBOOST_net_13325;
wire g65240_db;
wire g65240_sb;
wire TIMEBOOST_net_247;
wire TIMEBOOST_net_3388;
wire g65241_sb;
wire TIMEBOOST_net_248;
wire TIMEBOOST_net_9679;
wire g65242_sb;
wire TIMEBOOST_net_249;
wire TIMEBOOST_net_13547;
wire g65243_sb;
wire TIMEBOOST_net_250;
wire TIMEBOOST_net_13546;
wire g65244_sb;
wire TIMEBOOST_net_251;
wire TIMEBOOST_net_12786;
wire g65245_sb;
wire TIMEBOOST_net_252;
wire TIMEBOOST_net_13545;
wire g65246_sb;
wire TIMEBOOST_net_253;
wire TIMEBOOST_net_13502;
wire g65247_sb;
wire TIMEBOOST_net_254;
wire TIMEBOOST_net_12602;
wire g65248_sb;
wire TIMEBOOST_net_255;
wire TIMEBOOST_net_13501;
wire g65249_sb;
wire TIMEBOOST_net_256;
wire TIMEBOOST_net_3397;
wire g65250_sb;
wire TIMEBOOST_net_10757;
wire g65251_db;
wire g65251_sb;
wire g65252_da;
wire g65252_db;
wire g65252_sb;
wire g65254_p;
wire g65255_p;
wire TIMEBOOST_net_3167;
wire TIMEBOOST_net_14968;
wire g65257_p;
wire g65258_p;
wire g65259_p;
wire g65260_p;
wire g65261_p;
wire g65262_da;
wire g65262_db;
wire g65262_sb;
wire g65263_p;
wire g65264_p;
wire g65265_p;
wire g65266_p;
wire g65267_p;
wire g65268_da;
wire TIMEBOOST_net_12408;
wire g65268_sb;
wire TIMEBOOST_net_14973;
wire TIMEBOOST_net_81;
wire g65269_sb;
wire TIMEBOOST_net_23;
wire TIMEBOOST_net_12858;
wire g65270_sb;
wire g65271_da;
wire TIMEBOOST_net_9967;
wire g65271_sb;
wire g65272_da;
wire TIMEBOOST_net_204;
wire g65272_sb;
wire g65273_da;
wire TIMEBOOST_net_9968;
wire g65273_sb;
wire TIMEBOOST_net_14484;
wire TIMEBOOST_net_12833;
wire g65274_sb;
wire g65275_da;
wire TIMEBOOST_net_4411;
wire g65275_sb;
wire TIMEBOOST_net_10287;
wire g65276_db;
wire g65276_sb;
wire TIMEBOOST_net_3969;
wire g65277_db;
wire g65277_sb;
wire TIMEBOOST_net_3970;
wire g65278_db;
wire g65278_sb;
wire g65279_db;
wire g65279_sb;
wire g65280_da;
wire TIMEBOOST_net_3354;
wire g65280_sb;
wire g65281_da;
wire TIMEBOOST_net_3868;
wire g65281_sb;
wire TIMEBOOST_net_10283;
wire g65282_db;
wire g65282_sb;
wire TIMEBOOST_net_3973;
wire g65283_db;
wire g65283_sb;
wire TIMEBOOST_net_10292;
wire g65284_db;
wire g65284_sb;
wire TIMEBOOST_net_10293;
wire g65285_db;
wire g65285_sb;
wire TIMEBOOST_net_9550;
wire TIMEBOOST_net_12467;
wire g65286_sb;
wire g65287_da;
wire TIMEBOOST_net_3869;
wire g65287_sb;
wire TIMEBOOST_net_10288;
wire g65288_db;
wire g65288_sb;
wire TIMEBOOST_net_10302;
wire g65289_db;
wire g65289_sb;
wire g65290_da;
wire TIMEBOOST_net_12568;
wire g65291_da;
wire TIMEBOOST_net_161;
wire g65291_sb;
wire g65292_da;
wire TIMEBOOST_net_12834;
wire g65292_sb;
wire g65293_da;
wire TIMEBOOST_net_9795;
wire g65293_sb;
wire TIMEBOOST_net_12655;
wire g65294_db;
wire g65294_sb;
wire TIMEBOOST_net_13583;
wire TIMEBOOST_net_14649;
wire g65295_sb;
wire TIMEBOOST_net_9784;
wire g65296_db;
wire g65296_sb;
wire TIMEBOOST_net_13582;
wire g65297_db;
wire g65297_sb;
wire TIMEBOOST_net_3778;
wire TIMEBOOST_net_14842;
wire g65298_sb;
wire TIMEBOOST_net_3779;
wire TIMEBOOST_net_14830;
wire g65299_sb;
wire TIMEBOOST_net_15185;
wire TIMEBOOST_net_12841;
wire g65300_sb;
wire TIMEBOOST_net_3781;
wire TIMEBOOST_net_14618;
wire g65301_sb;
wire TIMEBOOST_net_3782;
wire g65302_db;
wire g65302_sb;
wire TIMEBOOST_net_3978;
wire g65303_db;
wire g65303_sb;
wire TIMEBOOST_net_3783;
wire g65304_db;
wire g65304_sb;
wire TIMEBOOST_net_3784;
wire g65305_db;
wire g65305_sb;
wire TIMEBOOST_net_15184;
wire g65306_db;
wire g65306_sb;
wire TIMEBOOST_net_3786;
wire g65307_db;
wire g65307_sb;
wire TIMEBOOST_net_3787;
wire g65308_db;
wire g65308_sb;
wire g65309_da;
wire g65309_db;
wire g65309_sb;
wire g65310_da;
wire g65310_db;
wire g65310_sb;
wire TIMEBOOST_net_3788;
wire g65311_db;
wire g65311_sb;
wire TIMEBOOST_net_14485;
wire TIMEBOOST_net_9653;
wire g65312_sb;
wire TIMEBOOST_net_3789;
wire g65313_db;
wire g65313_sb;
wire TIMEBOOST_net_3790;
wire g65314_db;
wire g65314_sb;
wire TIMEBOOST_net_3791;
wire g65315_db;
wire g65315_sb;
wire g65316_da;
wire TIMEBOOST_net_4412;
wire g65316_sb;
wire TIMEBOOST_net_3792;
wire g65317_db;
wire g65317_sb;
wire TIMEBOOST_net_3793;
wire g65318_db;
wire g65318_sb;
wire TIMEBOOST_net_12654;
wire g65319_db;
wire g65319_sb;
wire g65320_da;
wire TIMEBOOST_net_9796;
wire g65320_sb;
wire TIMEBOOST_net_12653;
wire g65321_db;
wire g65321_sb;
wire g65322_da;
wire TIMEBOOST_net_9790;
wire g65322_sb;
wire TIMEBOOST_net_12640;
wire g65323_db;
wire g65323_sb;
wire TIMEBOOST_net_15183;
wire g65324_db;
wire g65324_sb;
wire g65325_da;
wire TIMEBOOST_net_162;
wire g65325_sb;
wire g65326_da;
wire TIMEBOOST_net_9791;
wire g65326_sb;
wire TIMEBOOST_net_3798;
wire g65327_db;
wire g65327_sb;
wire TIMEBOOST_net_15182;
wire g65328_db;
wire g65328_sb;
wire g65329_da;
wire TIMEBOOST_net_13591;
wire g65329_sb;
wire TIMEBOOST_net_15181;
wire g65330_db;
wire g65330_sb;
wire g65331_da;
wire TIMEBOOST_net_3330;
wire g65331_sb;
wire TIMEBOOST_net_9855;
wire g65332_db;
wire g65332_sb;
wire g65333_da;
wire TIMEBOOST_net_13387;
wire g65333_sb;
wire TIMEBOOST_net_3802;
wire g65334_db;
wire g65334_sb;
wire TIMEBOOST_net_3803;
wire g65335_db;
wire g65335_sb;
wire g65336_da;
wire TIMEBOOST_net_3625;
wire g65336_sb;
wire TIMEBOOST_net_14488;
wire TIMEBOOST_net_3626;
wire g65337_sb;
wire TIMEBOOST_net_3804;
wire g65338_db;
wire g65338_sb;
wire TIMEBOOST_net_10303;
wire g65339_db;
wire g65339_sb;
wire TIMEBOOST_net_12835;
wire TIMEBOOST_net_13121;
wire g65340_sb;
wire g65341_da;
wire TIMEBOOST_net_12856;
wire g65341_sb;
wire TIMEBOOST_net_15180;
wire g65342_db;
wire g65342_sb;
wire TIMEBOOST_net_3806;
wire g65343_db;
wire g65343_sb;
wire TIMEBOOST_net_12349;
wire TIMEBOOST_net_206;
wire TIMEBOOST_net_3807;
wire g65345_db;
wire g65345_sb;
wire TIMEBOOST_net_3808;
wire TIMEBOOST_net_14619;
wire g65346_sb;
wire g65347_da;
wire g65347_sb;
wire TIMEBOOST_net_4272;
wire g65348_db;
wire g65348_sb;
wire TIMEBOOST_net_4273;
wire g65349_db;
wire g65349_sb;
wire g65350_da;
wire TIMEBOOST_net_10730;
wire g65350_sb;
wire TIMEBOOST_net_4274;
wire g65351_db;
wire g65351_sb;
wire TIMEBOOST_net_10399;
wire g65352_db;
wire g65352_sb;
wire TIMEBOOST_net_4276;
wire g65353_db;
wire g65353_sb;
wire TIMEBOOST_net_10398;
wire g65354_db;
wire g65354_sb;
wire TIMEBOOST_net_13262;
wire g65355_db;
wire g65355_sb;
wire TIMEBOOST_net_13412;
wire g65356_db;
wire g65356_sb;
wire TIMEBOOST_net_10159;
wire TIMEBOOST_net_14477;
wire g65357_sb;
wire g65358_da;
wire g65358_sb;
wire TIMEBOOST_net_14197;
wire g65359_sb;
wire TIMEBOOST_net_13263;
wire g65360_db;
wire g65360_sb;
wire g65361_db;
wire g65361_sb;
wire TIMEBOOST_net_10404;
wire g65362_db;
wire g65362_sb;
wire TIMEBOOST_net_4284;
wire g65363_db;
wire g65363_sb;
wire TIMEBOOST_net_10429;
wire g65364_db;
wire g65364_sb;
wire TIMEBOOST_net_13315;
wire g65365_db;
wire g65365_sb;
wire TIMEBOOST_net_15179;
wire g65366_db;
wire g65366_sb;
wire TIMEBOOST_net_15220;
wire g65367_db;
wire g65367_sb;
wire TIMEBOOST_net_10312;
wire g65368_db;
wire g65368_sb;
wire g65369_da;
wire TIMEBOOST_net_9645;
wire g65369_sb;
wire g65370_da;
wire TIMEBOOST_net_12586;
wire g65370_sb;
wire g65371_da;
wire TIMEBOOST_net_12463;
wire g65372_da;
wire TIMEBOOST_net_12733;
wire g65372_sb;
wire g65373_db;
wire g65373_sb;
wire TIMEBOOST_net_10079;
wire TIMEBOOST_net_14705;
wire g65374_sb;
wire g65375_da;
wire TIMEBOOST_net_12740;
wire g65375_sb;
wire g65376_da;
wire g65376_db;
wire g65376_sb;
wire g65377_da;
wire g65377_db;
wire g65377_sb;
wire g65378_da;
wire TIMEBOOST_net_14122;
wire g65378_sb;
wire g65379_da;
wire TIMEBOOST_net_9981;
wire g65379_sb;
wire g65380_da;
wire TIMEBOOST_net_12789;
wire g65380_sb;
wire g65381_da;
wire g65381_sb;
wire TIMEBOOST_net_4287;
wire g65382_db;
wire g65382_sb;
wire TIMEBOOST_net_14207;
wire TIMEBOOST_net_10264;
wire g65383_sb;
wire g65384_da;
wire TIMEBOOST_net_10265;
wire g65384_sb;
wire TIMEBOOST_net_4288;
wire g65385_db;
wire g65385_sb;
wire TIMEBOOST_net_169;
wire TIMEBOOST_net_9368;
wire g65387_da;
wire TIMEBOOST_net_10266;
wire g65387_sb;
wire TIMEBOOST_net_15208;
wire TIMEBOOST_net_14620;
wire g65388_sb;
wire TIMEBOOST_net_13451;
wire g65389_db;
wire g65389_sb;
wire g65390_da;
wire g65390_db;
wire g65390_sb;
wire TIMEBOOST_net_3981;
wire g65391_db;
wire g65391_sb;
wire g65392_da;
wire TIMEBOOST_net_10267;
wire g65392_sb;
wire TIMEBOOST_net_10074;
wire g65393_db;
wire g65393_sb;
wire TIMEBOOST_net_4290;
wire g65394_db;
wire g65394_sb;
wire TIMEBOOST_net_13314;
wire g65395_db;
wire g65395_sb;
wire g65396_da;
wire TIMEBOOST_net_10268;
wire g65396_sb;
wire TIMEBOOST_net_4292;
wire g65397_db;
wire g65397_sb;
wire g65398_db;
wire g65398_sb;
wire TIMEBOOST_net_14489;
wire TIMEBOOST_net_9982;
wire g65399_sb;
wire TIMEBOOST_net_3814;
wire g65400_db;
wire g65400_sb;
wire TIMEBOOST_net_13450;
wire g65401_db;
wire g65401_sb;
wire g65402_da;
wire TIMEBOOST_net_9948;
wire g65402_sb;
wire g65403_da;
wire TIMEBOOST_net_3634;
wire g65403_sb;
wire g65404_db;
wire g65404_sb;
wire TIMEBOOST_net_3816;
wire TIMEBOOST_net_14818;
wire g65405_sb;
wire TIMEBOOST_net_14496;
wire TIMEBOOST_net_12791;
wire g65406_sb;
wire g65407_da;
wire TIMEBOOST_net_12792;
wire g65407_sb;
wire g65408_da;
wire TIMEBOOST_net_13330;
wire g65408_sb;
wire TIMEBOOST_net_14497;
wire TIMEBOOST_net_12830;
wire g65409_sb;
wire TIMEBOOST_net_3983;
wire g65410_db;
wire g65410_sb;
wire g65411_da;
wire TIMEBOOST_net_164;
wire TIMEBOOST_net_3817;
wire g65412_db;
wire g65412_sb;
wire TIMEBOOST_net_3818;
wire g65413_db;
wire g65413_sb;
wire g65414_da;
wire g65414_db;
wire g65414_sb;
wire TIMEBOOST_net_9952;
wire g65415_db;
wire g65415_sb;
wire g65416_da;
wire TIMEBOOST_net_12831;
wire g65416_sb;
wire TIMEBOOST_net_3820;
wire g65417_db;
wire g65417_sb;
wire TIMEBOOST_net_3821;
wire TIMEBOOST_net_14612;
wire g65418_sb;
wire g65419_da;
wire TIMEBOOST_net_12334;
wire g65420_da;
wire g65420_db;
wire g65421_da;
wire TIMEBOOST_net_3639;
wire g65421_sb;
wire TIMEBOOST_net_14504;
wire TIMEBOOST_net_9939;
wire g65422_sb;
wire TIMEBOOST_net_10018;
wire TIMEBOOST_net_3641;
wire g65423_sb;
wire g65424_da;
wire TIMEBOOST_net_3642;
wire g65424_sb;
wire g65425_db;
wire g65425_sb;
wire TIMEBOOST_net_3822;
wire g65426_db;
wire g65426_sb;
wire g65427_da;
wire TIMEBOOST_net_13346;
wire g65427_sb;
wire g65428_da;
wire TIMEBOOST_net_9652;
wire g65428_sb;
wire g65429_da;
wire TIMEBOOST_net_9959;
wire g65429_sb;
wire g65430_da;
wire TIMEBOOST_net_9960;
wire g65430_sb;
wire g65431_da;
wire g65431_db;
wire g65431_sb;
wire TIMEBOOST_net_3823;
wire g65432_db;
wire g65432_sb;
wire TIMEBOOST_net_10103;
wire TIMEBOOST_net_12262;
wire g65433_sb;
wire TIMEBOOST_net_10104;
wire TIMEBOOST_net_14613;
wire g65434_sb;
wire TIMEBOOST_net_10197;
wire TIMEBOOST_net_14614;
wire g65435_sb;
wire g65436_p;
wire g65437_p;
wire g65439_p;
wire g65486_p;
wire g65488_p;
wire g65489_p;
wire g65490_p;
wire g65491_p;
wire g65493_p;
wire g65495_p;
wire g65497_p;
wire g65498_p;
wire g65510_p;
wire g65511_p;
wire g65513_p;
wire g65514_p;
wire g65515_p;
wire g65517_p;
wire g65518_p;
wire g65520_p;
wire g65522_p1;
wire g65522_p2;
wire g65523_p;
wire g65530_p;
wire g65533_p;
wire g65543_p;
wire g65549_p;
wire g65550_p;
wire g65555_p;
wire g65557_p;
wire g65559_p;
wire g65562_p;
wire g65567_p;
wire g65568_p;
wire g65569_p;
wire g65570_p;
wire g65571_p;
wire g65572_p1;
wire g65572_p2;
wire g65573_p;
wire g65583_p;
wire g65588_p;
wire g65590_p;
wire g65595_p;
wire g65614_p;
wire g65617_p;
wire g65626_p;
wire TIMEBOOST_net_13102;
wire g65668_db;
wire g65668_sb;
wire TIMEBOOST_net_9915;
wire TIMEBOOST_net_12548;
wire g65669_sb;
wire TIMEBOOST_net_4051;
wire g65670_db;
wire g65670_sb;
wire TIMEBOOST_net_9755;
wire TIMEBOOST_net_12455;
wire g65671_sb;
wire TIMEBOOST_net_3512;
wire g65672_db;
wire g65672_sb;
wire TIMEBOOST_net_10440;
wire g65673_db;
wire g65673_sb;
wire TIMEBOOST_net_3740;
wire g65674_db;
wire g65674_sb;
wire TIMEBOOST_net_9573;
wire g65675_db;
wire g65675_sb;
wire TIMEBOOST_net_3402;
wire g65676_db;
wire g65676_sb;
wire TIMEBOOST_net_12504;
wire g65677_db;
wire g65677_sb;
wire TIMEBOOST_net_12496;
wire g65678_db;
wire g65678_sb;
wire TIMEBOOST_net_12451;
wire g65679_db;
wire g65679_sb;
wire TIMEBOOST_net_13787;
wire g65680_db;
wire g65680_sb;
wire g65681_da;
wire g65681_db;
wire g65681_sb;
wire TIMEBOOST_net_13498;
wire g65682_db;
wire g65682_sb;
wire TIMEBOOST_net_13116;
wire TIMEBOOST_net_9854;
wire g65683_sb;
wire TIMEBOOST_net_9574;
wire g65684_db;
wire g65684_sb;
wire TIMEBOOST_net_12505;
wire g65685_db;
wire g65685_sb;
wire TIMEBOOST_net_12523;
wire g65686_db;
wire g65686_sb;
wire TIMEBOOST_net_12495;
wire g65687_db;
wire g65687_sb;
wire TIMEBOOST_net_14974;
wire g65688_db;
wire g65688_sb;
wire TIMEBOOST_net_12526;
wire g65689_db;
wire g65689_sb;
wire TIMEBOOST_net_4062;
wire TIMEBOOST_net_14797;
wire g65690_sb;
wire TIMEBOOST_net_9603;
wire g65691_db;
wire g65691_sb;
wire TIMEBOOST_net_12490;
wire g65692_db;
wire g65692_sb;
wire TIMEBOOST_net_12977;
wire g65693_db;
wire g65693_sb;
wire TIMEBOOST_net_9758;
wire g65694_db;
wire g65694_sb;
wire TIMEBOOST_net_12592;
wire g65695_db;
wire g65695_sb;
wire TIMEBOOST_net_3223;
wire TIMEBOOST_net_9604;
wire g65696_sb;
wire TIMEBOOST_net_14975;
wire TIMEBOOST_net_12397;
wire g65697_sb;
wire TIMEBOOST_net_12609;
wire g65698_db;
wire g65698_sb;
wire TIMEBOOST_net_14976;
wire g65699_db;
wire g65699_sb;
wire TIMEBOOST_net_14991;
wire g65700_db;
wire g65700_sb;
wire TIMEBOOST_net_12613;
wire g65701_db;
wire g65701_sb;
wire TIMEBOOST_net_12980;
wire g65702_db;
wire g65702_sb;
wire TIMEBOOST_net_12577;
wire g65703_db;
wire g65703_sb;
wire g65704_db;
wire g65704_sb;
wire TIMEBOOST_net_13530;
wire g65705_db;
wire g65705_sb;
wire TIMEBOOST_net_9489;
wire g65706_db;
wire g65706_sb;
wire TIMEBOOST_net_12200;
wire g65707_db;
wire g65707_sb;
wire TIMEBOOST_net_12433;
wire g65708_db;
wire g65708_sb;
wire TIMEBOOST_net_10334;
wire g65709_db;
wire g65709_sb;
wire TIMEBOOST_net_9605;
wire TIMEBOOST_net_12355;
wire g65710_sb;
wire TIMEBOOST_net_9487;
wire g65711_db;
wire g65711_sb;
wire TIMEBOOST_net_12589;
wire g65712_db;
wire g65712_sb;
wire TIMEBOOST_net_9544;
wire g65713_db;
wire g65713_sb;
wire TIMEBOOST_net_9606;
wire g65714_db;
wire g65714_sb;
wire TIMEBOOST_net_9607;
wire TIMEBOOST_net_287;
wire g65715_sb;
wire TIMEBOOST_net_14636;
wire g65716_db;
wire TIMEBOOST_net_14876;
wire g65717_db;
wire g65717_sb;
wire TIMEBOOST_net_14999;
wire g65718_db;
wire g65718_sb;
wire TIMEBOOST_net_15004;
wire g65719_db;
wire g65719_sb;
wire TIMEBOOST_net_13117;
wire g65720_db;
wire g65720_sb;
wire g65721_da;
wire g65721_db;
wire g65721_sb;
wire TIMEBOOST_net_3407;
wire g65722_db;
wire g65722_sb;
wire TIMEBOOST_net_12747;
wire g65723_db;
wire g65723_sb;
wire TIMEBOOST_net_3999;
wire g65724_db;
wire g65724_sb;
wire TIMEBOOST_net_12343;
wire g65725_db;
wire g65725_sb;
wire TIMEBOOST_net_3263;
wire TIMEBOOST_net_3252;
wire g65726_sb;
wire TIMEBOOST_net_4000;
wire g65727_db;
wire g65727_sb;
wire TIMEBOOST_net_12344;
wire g65728_db;
wire g65728_sb;
wire g65729_p;
wire TIMEBOOST_net_12345;
wire g65730_db;
wire g65730_sb;
wire g65731_da;
wire g65731_db;
wire g65731_sb;
wire TIMEBOOST_net_10335;
wire g65732_db;
wire g65732_sb;
wire g65733_da;
wire g65733_db;
wire g65733_sb;
wire TIMEBOOST_net_12712;
wire TIMEBOOST_net_12354;
wire g65734_sb;
wire TIMEBOOST_net_13251;
wire g65735_db;
wire g65735_sb;
wire TIMEBOOST_net_4002;
wire g65736_db;
wire g65736_sb;
wire TIMEBOOST_net_9611;
wire g65737_db;
wire g65737_sb;
wire g65738_da;
wire g65738_db;
wire g65738_sb;
wire TIMEBOOST_net_12346;
wire g65739_db;
wire g65739_sb;
wire TIMEBOOST_net_12510;
wire g65740_db;
wire g65740_sb;
wire TIMEBOOST_net_13512;
wire g65741_db;
wire g65741_sb;
wire TIMEBOOST_net_13511;
wire g65742_db;
wire g65742_sb;
wire TIMEBOOST_net_12506;
wire g65743_db;
wire g65743_sb;
wire TIMEBOOST_net_3417;
wire g65744_db;
wire g65744_sb;
wire TIMEBOOST_net_15032;
wire g65745_db;
wire g65745_sb;
wire TIMEBOOST_net_12553;
wire g65746_db;
wire g65746_sb;
wire TIMEBOOST_net_10336;
wire g65747_db;
wire g65747_sb;
wire TIMEBOOST_net_4003;
wire g65748_db;
wire g65748_sb;
wire TIMEBOOST_net_12281;
wire TIMEBOOST_net_12887;
wire g65749_sb;
wire TIMEBOOST_net_9545;
wire g65750_db;
wire g65750_sb;
wire TIMEBOOST_net_10337;
wire g65751_db;
wire g65751_sb;
wire g65752_da;
wire g65752_db;
wire g65752_sb;
wire TIMEBOOST_net_14808;
wire g65753_db;
wire g65753_sb;
wire TIMEBOOST_net_12551;
wire g65754_db;
wire g65754_sb;
wire TIMEBOOST_net_9546;
wire g65755_db;
wire g65755_sb;
wire TIMEBOOST_net_9547;
wire g65756_db;
wire g65756_sb;
wire TIMEBOOST_net_3169;
wire g65757_db;
wire TIMEBOOST_net_9779;
wire g65758_db;
wire g65758_sb;
wire TIMEBOOST_net_9595;
wire g65759_db;
wire g65759_sb;
wire TIMEBOOST_net_14807;
wire g65760_db;
wire g65760_sb;
wire TIMEBOOST_net_9553;
wire TIMEBOOST_net_12347;
wire g65761_sb;
wire TIMEBOOST_net_12348;
wire g65762_db;
wire g65762_sb;
wire TIMEBOOST_net_12290;
wire g65763_db;
wire TIMEBOOST_net_3257;
wire g65764_db;
wire g65764_sb;
wire TIMEBOOST_net_3258;
wire TIMEBOOST_net_3289;
wire TIMEBOOST_net_4004;
wire g65766_db;
wire g65766_sb;
wire TIMEBOOST_net_12279;
wire TIMEBOOST_net_3259;
wire g65767_sb;
wire TIMEBOOST_net_13252;
wire TIMEBOOST_net_14721;
wire g65768_sb;
wire TIMEBOOST_net_3260;
wire g65769_db;
wire g65769_sb;
wire TIMEBOOST_net_9560;
wire g65770_db;
wire g65770_sb;
wire TIMEBOOST_net_4006;
wire g65771_db;
wire g65771_sb;
wire TIMEBOOST_net_12621;
wire g65772_db;
wire g65772_sb;
wire TIMEBOOST_net_10338;
wire g65773_db;
wire g65773_sb;
wire TIMEBOOST_net_12590;
wire g65774_db;
wire g65774_sb;
wire TIMEBOOST_net_3752;
wire g65775_db;
wire g65775_sb;
wire TIMEBOOST_net_14841;
wire g65776_db;
wire g65776_sb;
wire TIMEBOOST_net_3180;
wire g65777_db;
wire g65777_sb;
wire TIMEBOOST_net_3181;
wire g65778_db;
wire g65778_sb;
wire TIMEBOOST_net_12552;
wire g65779_db;
wire g65779_sb;
wire g65780_da;
wire g65780_db;
wire g65780_sb;
wire TIMEBOOST_net_14801;
wire TIMEBOOST_net_3262;
wire g65781_sb;
wire TIMEBOOST_net_14637;
wire g65782_db;
wire g65782_sb;
wire TIMEBOOST_net_4007;
wire g65783_db;
wire g65783_sb;
wire TIMEBOOST_net_9581;
wire g65784_db;
wire g65784_sb;
wire TIMEBOOST_net_9616;
wire TIMEBOOST_net_3287;
wire TIMEBOOST_net_4008;
wire TIMEBOOST_net_14723;
wire g65786_sb;
wire TIMEBOOST_net_12931;
wire g65787_db;
wire g65787_sb;
wire TIMEBOOST_net_4009;
wire g65788_db;
wire g65788_sb;
wire TIMEBOOST_net_12498;
wire g65789_db;
wire g65789_sb;
wire TIMEBOOST_net_9549;
wire g65790_db;
wire g65790_sb;
wire TIMEBOOST_net_4010;
wire g65791_db;
wire g65791_sb;
wire TIMEBOOST_net_9552;
wire g65792_db;
wire g65792_sb;
wire TIMEBOOST_net_4011;
wire g65793_db;
wire g65793_sb;
wire TIMEBOOST_net_9537;
wire g65794_db;
wire g65794_sb;
wire TIMEBOOST_net_14680;
wire g65795_db;
wire g65795_sb;
wire TIMEBOOST_net_12909;
wire TIMEBOOST_net_12352;
wire TIMEBOOST_net_257;
wire TIMEBOOST_net_12593;
wire g65797_sb;
wire g65798_db;
wire g65798_sb;
wire TIMEBOOST_net_4013;
wire g65799_db;
wire g65799_sb;
wire TIMEBOOST_net_12563;
wire g65800_db;
wire g65800_sb;
wire g65801_p;
wire TIMEBOOST_net_14753;
wire g65802_db;
wire g65802_sb;
wire TIMEBOOST_net_3084;
wire g65803_db;
wire g65803_sb;
wire TIMEBOOST_net_9797;
wire g65804_db;
wire g65804_sb;
wire TIMEBOOST_net_3185;
wire g65805_db;
wire g65805_sb;
wire TIMEBOOST_net_3186;
wire g65806_db;
wire g65806_sb;
wire TIMEBOOST_net_4071;
wire g65807_db;
wire g65807_sb;
wire TIMEBOOST_net_83;
wire TIMEBOOST_net_9528;
wire g65808_p;
wire TIMEBOOST_net_10269;
wire g65809_db;
wire g65809_sb;
wire TIMEBOOST_net_87;
wire TIMEBOOST_net_12691;
wire g65810_sb;
wire TIMEBOOST_net_10270;
wire g65811_db;
wire g65811_sb;
wire TIMEBOOST_net_10271;
wire g65812_db;
wire g65812_sb;
wire TIMEBOOST_net_352;
wire g65813_db;
wire g65813_sb;
wire TIMEBOOST_net_10214;
wire g65814_db;
wire g65814_sb;
wire TIMEBOOST_net_4626;
wire g65815_db;
wire g65815_sb;
wire TIMEBOOST_net_13115;
wire g65816_db;
wire g65816_sb;
wire TIMEBOOST_net_218;
wire TIMEBOOST_net_3333;
wire TIMEBOOST_net_3937;
wire g65818_db;
wire g65818_sb;
wire TIMEBOOST_net_3938;
wire g65819_db;
wire g65819_sb;
wire TIMEBOOST_net_4627;
wire TIMEBOOST_net_14208;
wire g65820_sb;
wire TIMEBOOST_net_10216;
wire g65821_db;
wire g65821_sb;
wire TIMEBOOST_net_14470;
wire g65822_db;
wire g65822_sb;
wire g65823_db;
wire g65823_sb;
wire TIMEBOOST_net_9287;
wire TIMEBOOST_net_14486;
wire g65824_sb;
wire g65825_da;
wire g65825_db;
wire g65825_sb;
wire TIMEBOOST_net_9288;
wire TIMEBOOST_net_10218;
wire g65826_sb;
wire g65827_da;
wire g65827_db;
wire g65827_sb;
wire TIMEBOOST_net_13449;
wire TIMEBOOST_net_14487;
wire g65828_sb;
wire TIMEBOOST_net_12231;
wire g65829_sb;
wire TIMEBOOST_net_12239;
wire TIMEBOOST_net_3943;
wire g65830_sb;
wire TIMEBOOST_net_9291;
wire TIMEBOOST_net_9942;
wire g65831_sb;
wire TIMEBOOST_net_12225;
wire TIMEBOOST_net_3945;
wire g65832_sb;
wire TIMEBOOST_net_12250;
wire TIMEBOOST_net_9943;
wire g65833_sb;
wire TIMEBOOST_net_12258;
wire TIMEBOOST_net_10284;
wire g65834_sb;
wire TIMEBOOST_net_12672;
wire TIMEBOOST_net_12677;
wire g65835_sb;
wire TIMEBOOST_net_13448;
wire g65836_db;
wire g65836_sb;
wire TIMEBOOST_net_12256;
wire TIMEBOOST_net_10285;
wire g65837_sb;
wire TIMEBOOST_net_10454;
wire g65838_db;
wire g65838_sb;
wire g65839_da;
wire g65839_db;
wire g65839_sb;
wire TIMEBOOST_net_10430;
wire g65840_db;
wire g65840_sb;
wire TIMEBOOST_net_4298;
wire TIMEBOOST_net_632;
wire g65841_sb;
wire g65842_da;
wire g65842_db;
wire g65842_sb;
wire TIMEBOOST_net_10457;
wire g65843_db;
wire g65843_sb;
wire g65844_da;
wire g65844_db;
wire g65844_sb;
wire TIMEBOOST_net_4300;
wire g65845_db;
wire g65845_sb;
wire TIMEBOOST_net_12274;
wire TIMEBOOST_net_3949;
wire g65846_sb;
wire TIMEBOOST_net_3085;
wire g65847_db;
wire g65847_sb;
wire TIMEBOOST_net_10742;
wire TIMEBOOST_net_14331;
wire g65848_sb;
wire TIMEBOOST_net_141;
wire TIMEBOOST_net_14949;
wire g65849_sb;
wire TIMEBOOST_net_3086;
wire TIMEBOOST_net_12399;
wire g65850_sb;
wire TIMEBOOST_net_9551;
wire g65851_db;
wire g65851_sb;
wire TIMEBOOST_net_12442;
wire g65852_db;
wire g65852_sb;
wire TIMEBOOST_net_15210;
wire g65853_db;
wire g65853_sb;
wire g65854_da;
wire g65854_db;
wire g65854_sb;
wire TIMEBOOST_net_10286;
wire g65855_db;
wire g65855_sb;
wire TIMEBOOST_net_10540;
wire TIMEBOOST_net_14412;
wire g65856_sb;
wire TIMEBOOST_net_9588;
wire TIMEBOOST_net_12657;
wire g65857_sb;
wire TIMEBOOST_net_3173;
wire TIMEBOOST_net_720;
wire g65858_sb;
wire TIMEBOOST_net_4484;
wire TIMEBOOST_net_14377;
wire g65859_sb;
wire TIMEBOOST_net_14947;
wire g65860_db;
wire g65860_sb;
wire TIMEBOOST_net_12612;
wire g65861_db;
wire g65861_sb;
wire g65862_da;
wire g65862_db;
wire g65862_sb;
wire TIMEBOOST_net_143;
wire g58068_db;
wire g65863_sb;
wire TIMEBOOST_net_12342;
wire TIMEBOOST_net_14424;
wire TIMEBOOST_net_14165;
wire g65865_db;
wire g65865_sb;
wire TIMEBOOST_net_12432;
wire g65866_db;
wire g65866_sb;
wire TIMEBOOST_net_14948;
wire g65867_db;
wire g65867_sb;
wire TIMEBOOST_net_12918;
wire g65868_db;
wire g65868_sb;
wire g65869_da;
wire g65869_db;
wire g65869_sb;
wire TIMEBOOST_net_3016;
wire g65870_db;
wire g65870_sb;
wire TIMEBOOST_net_3984;
wire g65871_db;
wire g65871_sb;
wire g65872_da;
wire g65872_db;
wire g65872_sb;
wire g65873_db;
wire g65873_sb;
wire TIMEBOOST_net_13277;
wire g65874_db;
wire g65874_sb;
wire TIMEBOOST_net_3017;
wire g65875_db;
wire g65875_sb;
wire TIMEBOOST_net_208;
wire TIMEBOOST_net_3334;
wire g65876_sb;
wire TIMEBOOST_net_10289;
wire g65877_db;
wire g65877_sb;
wire TIMEBOOST_net_12330;
wire TIMEBOOST_net_3089;
wire g65878_sb;
wire g65879_da;
wire g65879_db;
wire g65879_sb;
wire TIMEBOOST_net_3953;
wire g65880_db;
wire g65880_sb;
wire TIMEBOOST_net_10290;
wire g65881_db;
wire g65881_sb;
wire TIMEBOOST_net_4628;
wire TIMEBOOST_net_14212;
wire g65882_sb;
wire TIMEBOOST_net_12875;
wire g65883_db;
wire g65883_sb;
wire TIMEBOOST_net_10678;
wire TIMEBOOST_net_14187;
wire g65884_sb;
wire TIMEBOOST_net_144;
wire TIMEBOOST_net_14815;
wire TIMEBOOST_net_145;
wire TIMEBOOST_net_14748;
wire TIMEBOOST_net_4302;
wire g65887_db;
wire g65887_sb;
wire TIMEBOOST_net_3513;
wire g65888_db;
wire g65888_sb;
wire TIMEBOOST_net_3327;
wire g65889_db;
wire g65889_sb;
wire TIMEBOOST_net_10486;
wire g65890_db;
wire g65890_sb;
wire TIMEBOOST_net_12443;
wire g65891_db;
wire g65891_sb;
wire TIMEBOOST_net_10662;
wire TIMEBOOST_net_12970;
wire g65892_sb;
wire TIMEBOOST_net_12368;
wire g65893_db;
wire g65893_sb;
wire TIMEBOOST_net_10487;
wire g65894_db;
wire g65894_sb;
wire TIMEBOOST_net_146;
wire TIMEBOOST_net_12626;
wire TIMEBOOST_net_3955;
wire g65896_db;
wire g65896_sb;
wire TIMEBOOST_net_4305;
wire TIMEBOOST_net_14469;
wire g65897_sb;
wire TIMEBOOST_net_3276;
wire TIMEBOOST_net_14425;
wire TIMEBOOST_net_13525;
wire TIMEBOOST_net_6402;
wire g65899_sb;
wire TIMEBOOST_net_4485;
wire TIMEBOOST_net_14605;
wire g65900_sb;
wire g65901_da;
wire g65901_db;
wire g65901_sb;
wire g65902_da;
wire g65902_db;
wire g65902_sb;
wire TIMEBOOST_net_9554;
wire g65903_db;
wire g65903_sb;
wire TIMEBOOST_net_9555;
wire g65904_db;
wire g65904_sb;
wire TIMEBOOST_net_349;
wire TIMEBOOST_net_4052;
wire g65905_sb;
wire TIMEBOOST_net_4630;
wire g65906_db;
wire g65906_sb;
wire TIMEBOOST_net_3018;
wire g65907_db;
wire g65907_sb;
wire TIMEBOOST_net_3956;
wire g65908_db;
wire g65908_sb;
wire TIMEBOOST_net_10339;
wire g65909_db;
wire g65909_sb;
wire TIMEBOOST_net_3957;
wire g65910_db;
wire g65910_sb;
wire TIMEBOOST_net_356;
wire TIMEBOOST_net_14346;
wire TIMEBOOST_net_14261;
wire g65912_db;
wire TIMEBOOST_net_3958;
wire g65913_db;
wire g65913_sb;
wire g65914_da;
wire g65914_db;
wire g65914_sb;
wire TIMEBOOST_net_10664;
wire g65915_db;
wire g65915_sb;
wire TIMEBOOST_net_12874;
wire g65916_db;
wire g65916_sb;
wire TIMEBOOST_net_170;
wire TIMEBOOST_net_14168;
wire TIMEBOOST_net_14369;
wire g65918_db;
wire g65919_da;
wire g65919_db;
wire g65919_sb;
wire TIMEBOOST_net_4486;
wire TIMEBOOST_net_14378;
wire g65920_sb;
wire TIMEBOOST_net_9916;
wire g65921_db;
wire g65921_sb;
wire TIMEBOOST_net_10667;
wire TIMEBOOST_net_12971;
wire TIMEBOOST_net_12434;
wire g65923_db;
wire g65923_sb;
wire g65924_da;
wire g65924_db;
wire g65924_sb;
wire TIMEBOOST_net_4542;
wire g65925_db;
wire TIMEBOOST_net_4543;
wire g65926_db;
wire TIMEBOOST_net_10674;
wire g65927_db;
wire TIMEBOOST_net_10675;
wire g65928_db;
wire TIMEBOOST_net_4546;
wire TIMEBOOST_net_12972;
wire TIMEBOOST_net_12335;
wire TIMEBOOST_net_14334;
wire TIMEBOOST_net_12873;
wire g65931_db;
wire g65931_sb;
wire g65932_p;
wire TIMEBOOST_net_147;
wire TIMEBOOST_net_12600;
wire TIMEBOOST_net_3190;
wire g65934_db;
wire g65934_sb;
wire TIMEBOOST_net_9556;
wire g65935_db;
wire g65935_sb;
wire TIMEBOOST_net_4487;
wire TIMEBOOST_net_14592;
wire g65936_sb;
wire g65937_p;
wire g65938_p;
wire g65939_p;
wire TIMEBOOST_net_10445;
wire g65940_db;
wire g65940_sb;
wire TIMEBOOST_net_1238;
wire g65941_db;
wire g65942_da;
wire g65942_db;
wire g65942_sb;
wire TIMEBOOST_net_9297;
wire TIMEBOOST_net_3959;
wire g65943_sb;
wire TIMEBOOST_net_12340;
wire TIMEBOOST_net_14417;
wire TIMEBOOST_net_12336;
wire g65945_db;
wire TIMEBOOST_net_4387;
wire g65946_db;
wire TIMEBOOST_net_12381;
wire g65947_db;
wire TIMEBOOST_net_4547;
wire TIMEBOOST_net_12973;
wire TIMEBOOST_net_4488;
wire TIMEBOOST_net_14358;
wire g65949_sb;
wire TIMEBOOST_net_165;
wire TIMEBOOST_net_12614;
wire TIMEBOOST_net_3019;
wire g65951_db;
wire g65951_sb;
wire TIMEBOOST_net_3960;
wire g65952_db;
wire g65952_sb;
wire TIMEBOOST_net_10340;
wire TIMEBOOST_net_14977;
wire g65953_sb;
wire TIMEBOOST_net_3961;
wire g65954_db;
wire g65954_sb;
wire TIMEBOOST_net_12615;
wire g65955_db;
wire TIMEBOOST_net_4548;
wire TIMEBOOST_net_12974;
wire TIMEBOOST_net_14766;
wire g65957_db;
wire g65957_sb;
wire TIMEBOOST_net_3741;
wire g65958_db;
wire g65958_sb;
wire TIMEBOOST_net_3021;
wire g65959_db;
wire TIMEBOOST_net_12631;
wire g65960_db;
wire g65960_sb;
wire TIMEBOOST_net_14292;
wire g65961_db;
wire g65962_da;
wire g65962_db;
wire g65962_sb;
wire TIMEBOOST_net_361;
wire g65963_db;
wire TIMEBOOST_net_3000;
wire g65964_db;
wire g65964_sb;
wire TIMEBOOST_net_4074;
wire g65965_db;
wire g65965_sb;
wire TIMEBOOST_net_4075;
wire g65966_db;
wire g65966_sb;
wire TIMEBOOST_net_4076;
wire g65967_db;
wire g65967_sb;
wire TIMEBOOST_net_13973;
wire g65968_db;
wire TIMEBOOST_net_10341;
wire g65969_db;
wire g65969_sb;
wire TIMEBOOST_net_10342;
wire TIMEBOOST_net_12716;
wire g65970_sb;
wire TIMEBOOST_net_4079;
wire TIMEBOOST_net_14994;
wire g65971_sb;
wire TIMEBOOST_net_9940;
wire TIMEBOOST_net_14627;
wire g65972_sb;
wire TIMEBOOST_net_12390;
wire TIMEBOOST_net_12658;
wire TIMEBOOST_net_90;
wire TIMEBOOST_net_12673;
wire TIMEBOOST_net_4549;
wire TIMEBOOST_net_12975;
wire TIMEBOOST_net_3962;
wire g65976_db;
wire g65976_sb;
wire TIMEBOOST_net_3963;
wire g65977_db;
wire g65977_sb;
wire TIMEBOOST_net_10291;
wire g65978_db;
wire g65978_sb;
wire g65983_p;
wire g65984_p;
wire TIMEBOOST_net_8;
wire TIMEBOOST_net_12857;
wire g65992_p;
wire g65993_p;
wire TIMEBOOST_net_9631;
wire g65994_db;
wire g65994_sb;
wire TIMEBOOST_net_149;
wire TIMEBOOST_net_3731;
wire TIMEBOOST_net_150;
wire g65996_db;
wire TIMEBOOST_net_9564;
wire g65997_db;
wire TIMEBOOST_net_12668;
wire g65998_db;
wire TIMEBOOST_net_121;
wire g65999_db;
wire TIMEBOOST_net_9529;
wire g66000_db;
wire TIMEBOOST_net_151;
wire TIMEBOOST_net_12567;
wire g66002_p;
wire g66003_p;
wire g66004_p;
wire g66005_p;
wire g66006_p;
wire g66007_p;
wire g66008_p;
wire g66009_p;
wire g66010_p;
wire g66011_p;
wire g66012_p;
wire g66013_p;
wire g66014_p;
wire g66015_p;
wire g66016_p;
wire g66066_p;
wire g66068_p;
wire g66072_p;
wire g66074_p;
wire g66075_p;
wire g66076_p;
wire g66077_p;
wire g66078_p;
wire g66079_p;
wire g66080_p;
wire g66081_p;
wire g66082_p;
wire g66083_p;
wire g66084_p;
wire g66085_p;
wire g66086_p;
wire g66087_p;
wire g66089_p;
wire g66090_p;
wire g66093_p;
wire g66094_p;
wire g66095_p;
wire g66096_p;
wire g66097_p;
wire g66098_p;
wire g66099_p;
wire g66100_p;
wire g66107_p;
wire g66108_p;
wire g66110_p;
wire g66113_p;
wire g66118_p;
wire g66121_p;
wire g66122_p;
wire g66124_p;
wire g66125_p;
wire g66127_p;
wire g66128_p;
wire g66129_p;
wire g66130_p;
wire g66132_p;
wire g66133_p;
wire g66134_p;
wire g66136_p;
wire g66138_p;
wire g66143_p;
wire g66145_p;
wire g66147_p;
wire g66153_p;
wire g66155_p;
wire g66160_p;
wire g66165_p;
wire g66176_p;
wire g66178_p;
wire g66184_p;
wire g66190_p;
wire g66194_p;
wire g66195_p;
wire g66197_p;
wire g66202_p;
wire g66215_p;
wire g66223_p;
wire g66232_p;
wire g66234_p;
wire g66237_p;
wire g66239_p;
wire g66248_p;
wire g66267_p;
wire g66269_p;
wire g66278_p;
wire g66286_p;
wire g66287_p;
wire g66290_dup_p;
wire g66291_p;
wire g66298_p;
wire g66299_p;
wire g66302_p;
wire g66303_p;
wire g66310_p;
wire g66315_p;
wire g66322_p;
wire g66323_p;
wire g66327_p;
wire g66336_p;
wire g66338_p;
wire g66357_p;
wire g66358_p;
wire TIMEBOOST_net_12908;
wire TIMEBOOST_net_12403;
wire g66397_sb;
wire TIMEBOOST_net_12907;
wire g66398_db;
wire g66398_sb;
wire TIMEBOOST_net_122;
wire TIMEBOOST_net_12395;
wire g66399_sb;
wire TIMEBOOST_net_3269;
wire g66400_db;
wire TIMEBOOST_net_13194;
wire TIMEBOOST_net_12404;
wire TIMEBOOST_net_9585;
wire TIMEBOOST_net_12405;
wire g66402_sb;
wire TIMEBOOST_net_9621;
wire TIMEBOOST_net_14635;
wire g66403_sb;
wire TIMEBOOST_net_13215;
wire g66404_db;
wire TIMEBOOST_net_3274;
wire TIMEBOOST_net_14644;
wire TIMEBOOST_net_13286;
wire TIMEBOOST_net_14645;
wire g66406_sb;
wire TIMEBOOST_net_13285;
wire TIMEBOOST_net_14835;
wire TIMEBOOST_net_13284;
wire g66408_db;
wire TIMEBOOST_net_12277;
wire TIMEBOOST_net_14834;
wire TIMEBOOST_net_3279;
wire g66410_db;
wire TIMEBOOST_net_14163;
wire g66411_db;
wire TIMEBOOST_net_124;
wire g66412_db;
wire TIMEBOOST_net_125;
wire g66413_db;
wire TIMEBOOST_net_126;
wire g66414_db;
wire TIMEBOOST_net_13189;
wire TIMEBOOST_net_14676;
wire g66415_sb;
wire TIMEBOOST_net_9630;
wire TIMEBOOST_net_14895;
wire TIMEBOOST_net_127;
wire g66417_db;
wire TIMEBOOST_net_3282;
wire TIMEBOOST_net_14731;
wire TIMEBOOST_net_128;
wire g66419_db;
wire TIMEBOOST_net_13188;
wire TIMEBOOST_net_13206;
wire TIMEBOOST_net_12883;
wire g66421_db;
wire TIMEBOOST_net_9633;
wire TIMEBOOST_net_13205;
wire TIMEBOOST_net_180;
wire g66423_db;
wire TIMEBOOST_net_9634;
wire TIMEBOOST_net_9675;
wire TIMEBOOST_net_129;
wire TIMEBOOST_net_15013;
wire TIMEBOOST_net_130;
wire g66426_db;
wire TIMEBOOST_net_131;
wire g66427_db;
wire TIMEBOOST_net_13332;
wire TIMEBOOST_net_9676;
wire TIMEBOOST_net_9576;
wire TIMEBOOST_net_14839;
wire TIMEBOOST_net_9636;
wire TIMEBOOST_net_14737;
wire g66433_da;
wire g66433_db;
wire g66433_sb;
wire TIMEBOOST_net_3733;
wire g66456_db;
wire g66456_sb;
wire TIMEBOOST_net_14998;
wire g66457_db;
wire g66457_sb;
wire g66458_p;
wire g66458_p0;
wire g66459_p0;
wire g66464_p;
wire g66464_p0;
wire g66465_p;
wire g66465_p0;
wire g66473_p;
wire g66475_p;
wire g66477_da;
wire g66477_db;
wire g66544_p;
wire g66547_p;
wire g66550_p;
wire g66577_p;
wire g66583_p;
wire g66584_p;
wire g66607_p;
wire g66620_p;
wire g66627_p;
wire g66628_p;
wire g66646_p;
wire g66649_p;
wire g66650_p;
wire g66652_p;
wire g66658_p;
wire g66662_p;
wire g66663_p;
wire g66669_p;
wire g66672_p;
wire g66714_p;
wire g66726_p;
wire g66728_p;
wire g66737_p;
wire g66738_p;
wire g66742_p;
wire g66752_p;
wire g66753_p;
wire g66759_p;
wire g66773_p;
wire g66777_p;
wire g66789_p;
wire g66805_p;
wire g66813_p;
wire g66825_p;
wire g66827_p;
wire g66854_p;
wire g66856_p;
wire g66866_p;
wire g66875_p;
wire g66876_p;
wire g66888_p;
wire g66889_p;
wire g66902_p;
wire g66911_p;
wire g66912_p;
wire g66913_p;
wire g66915_p;
wire g66917_p;
wire g66918_p;
wire g66921_p;
wire g66922_p;
wire g66923_p;
wire g66924_p;
wire g66925_p;
wire g66927_p;
wire g66929_p;
wire g66930_p;
wire g66931_p;
wire g66932_p;
wire g66933_p;
wire g66934_p;
wire g66935_p;
wire g66936_p;
wire g66937_p;
wire g66940_p;
wire g66941_p;
wire g66942_p;
wire g66944_p;
wire g66945_p;
wire g66946_p;
wire g66947_p;
wire g66948_p;
wire g66949_p;
wire g66951_p;
wire g66952_p;
wire g66953_p;
wire g66954_p;
wire g66955_p;
wire g66957_p;
wire g66959_p;
wire g66960_p;
wire g66963_p;
wire g66964_p;
wire g66965_p;
wire g66966_p;
wire g66968_p;
wire g66975_p;
wire g66978_p;
wire g66984_p;
wire g66985_p;
wire g66986_p;
wire g66987_p;
wire g66988_p;
wire g66989_p;
wire g66990_p;
wire g66997_p;
wire g67001_p;
wire g67003_p;
wire g67005_p;
wire g67006_p;
wire g67008_p;
wire g67010_p;
wire g67011_p;
wire g67014_p;
wire g67015_p;
wire g67017_p;
wire g67018_p;
wire g67019_p;
wire g67020_p;
wire g67021_p;
wire g67022_p;
wire g67023_p;
wire g67024_p;
wire g67025_p;
wire g67026_p;
wire g67029_p;
wire g67030_p;
wire g67031_p;
wire g67032_p;
wire g67033_p;
wire g67036_p;
wire TIMEBOOST_net_93;
wire g67040_db;
wire g67040_sb;
wire TIMEBOOST_net_94;
wire g67041_db;
wire TIMEBOOST_net_11;
wire g67042_db;
wire g67042_sb;
wire TIMEBOOST_net_12;
wire g67043_db;
wire g67044_da;
wire g67044_db;
wire g67044_sb;
wire g67045_da;
wire g67045_db;
wire g67046_da;
wire g67046_db;
wire g67046_sb;
wire TIMEBOOST_net_15196;
wire g67048_db;
wire g67048_sb;
wire TIMEBOOST_net_14997;
wire g67049_db;
wire g67049_sb;
wire TIMEBOOST_net_14673;
wire g67050_db;
wire TIMEBOOST_net_95;
wire g67051_db;
wire g67051_sb;
wire TIMEBOOST_net_84;
wire g67052_db;
wire TIMEBOOST_net_96;
wire g67053_db;
wire TIMEBOOST_net_49;
wire TIMEBOOST_net_9379;
wire TIMEBOOST_net_15017;
wire g67055_db;
wire TIMEBOOST_net_12854;
wire g67056_db;
wire TIMEBOOST_net_43;
wire TIMEBOOST_net_9386;
wire g67057_sb;
wire TIMEBOOST_net_44;
wire TIMEBOOST_net_12807;
wire TIMEBOOST_net_12710;
wire g67059_db;
wire TIMEBOOST_net_15200;
wire TIMEBOOST_net_12414;
wire TIMEBOOST_net_12705;
wire TIMEBOOST_net_9384;
wire TIMEBOOST_net_40;
wire TIMEBOOST_net_12412;
wire g67070_da;
wire g67070_db;
wire g67070_sb;
wire TIMEBOOST_net_85;
wire g67071_db;
wire TIMEBOOST_net_132;
wire TIMEBOOST_net_12700;
wire TIMEBOOST_net_12732;
wire g67073_db;
wire TIMEBOOST_net_14891;
wire g67074_db;
wire TIMEBOOST_net_14166;
wire g67075_db;
wire TIMEBOOST_net_9533;
wire TIMEBOOST_net_14693;
wire g67082_sb;
wire TIMEBOOST_net_2876;
wire g67083_db;
wire TIMEBOOST_net_100;
wire g67084_db;
wire TIMEBOOST_net_2877;
wire g67085_db;
wire TIMEBOOST_net_46;
wire TIMEBOOST_net_9387;
wire TIMEBOOST_net_41;
wire TIMEBOOST_net_12409;
wire TIMEBOOST_net_101;
wire g67088_db;
wire TIMEBOOST_net_102;
wire g67091_db;
wire TIMEBOOST_net_47;
wire TIMEBOOST_net_2888;
wire TIMEBOOST_net_103;
wire g67093_db;
wire TIMEBOOST_net_48;
wire g67094_db;
wire g67095_p;
wire g67096_p;
wire g67097_p;
wire g67098_p;
wire g67099_p;
wire g67100_p;
wire g67102_p;
wire g67103_p;
wire g67104_p;
wire g67105_p;
wire g67106_p;
wire g67107_p;
wire g67108_p;
wire g67109_p;
wire g67110_p;
wire g67111_p;
wire g67112_p;
wire g67113_p;
wire g67114_p;
wire g67115_p;
wire g67116_p;
wire g67117_p;
wire g67118_p;
wire g67119_p;
wire g67120_p;
wire g67122_p;
wire g67123_p;
wire g67125_p;
wire g67126_p;
wire g67127_p;
wire g67128_p;
wire g67129_p;
wire g67130_p;
wire g67131_p;
wire g67132_p;
wire g67133_p;
wire g67134_p;
wire g67135_p;
wire g67136_p;
wire g67138_p;
wire g67139_p;
wire g67140_p;
wire g67141_p;
wire g67142_p;
wire g67143_p;
wire TIMEBOOST_net_14671;
wire g67145_p;
wire g67146_p;
wire TIMEBOOST_net_12413;
wire g67148_p;
wire g67149_p;
wire g67150_p;
wire g67151_p;
wire g67152_p;
wire g67153_p;
wire g67154_p;
wire g67155_p;
wire g67156_p;
wire g67157_p;
wire g67311_p;
wire g67313_p;
wire g67324_p;
wire g67327_p;
wire g67329_p;
wire g67340_p;
wire g67353_p;
wire g67355_p;
wire g67360_p;
wire g67364_p;
wire g67369_p;
wire g67371_p;
wire g67386_p;
wire g67389_p;
wire g67390_p;
wire g67392_p;
wire g67394_p;
wire g67396_p;
wire g67397_p;
wire g67403_p;
wire g67405_p;
wire g67411_p;
wire g67421_p;
wire g67425_p;
wire g67430_p;
wire g67432_p;
wire g67434_p;
wire g67437_p;
wire g67446_p;
wire g67453_p;
wire g67457_p;
wire g67459_p;
wire g67463_p;
wire g67468_p;
wire g67489_p;
wire g67493_p;
wire g67495_p;
wire g67498_p;
wire g67502_p;
wire g67505_p;
wire g67506_p;
wire g67507_p;
wire g67514_p;
wire g67519_p;
wire g67523_p;
wire g67531_p;
wire g67534_p;
wire g67535_p;
wire g67536_p;
wire g67537_p;
wire g67538_p;
wire g67544_p;
wire g67545_p;
wire g67549_p;
wire g67559_p;
wire g67581_p;
wire g67582_p;
wire g67583_p;
wire g67592_p;
wire g67596_p;
wire g67600_p;
wire g67603_p;
wire g67605_p;
wire g67610_p;
wire g67613_p;
wire g67624_p;
wire g67625_p;
wire g67626_p;
wire g67631_p;
wire g67671_p;
wire g67672_p;
wire g67675_p;
wire g67680_p;
wire g67688_p;
wire g67689_p;
wire g67699_p;
wire g67707_p;
wire g67709_p;
wire g67712_p;
wire g67721_p;
wire g67722_p;
wire g67725_p;
wire g67731_p;
wire g67735_p;
wire g67739_p;
wire g67745_p;
wire g67746_p;
wire g67747_p;
wire g67754_p;
wire g67757_p;
wire g67758_p;
wire g67763_p;
wire g67765_p;
wire g67778_p;
wire g67783_p;
wire g67791_p;
wire g67799_p;
wire g67802_p;
wire g67804_p;
wire g67806_p;
wire g67807_p;
wire g67814_p;
wire g67828_p;
wire g68_p;
wire g70_p;
wire g73989_p;
wire g74028_p;
wire g74140_p;
wire g74153_p;
wire g74154_p;
wire g74162_dup_p;
wire g74174_p;
wire g74243_p;
wire g74245_p;
wire g74270_p;
wire g74283_p;
wire g74363_p;
wire g74408_p;
wire g74429_p;
wire g74434_da;
wire g74434_db;
wire g74434_sb;
wire g74470_p;
wire g74475_p;
wire g74553_p;
wire g74563_p;
wire g74576_p;
wire g74580_p;
wire g74628_p;
wire g74644_p;
wire g74660_p;
wire g74661_p;
wire g74689_p;
wire g74739_p;
wire g74749_p;
wire g74787_p;
wire g74859_p;
wire g74872_p;
wire g74879_p;
wire g74886_p;
wire g74920_p;
wire g74930_p;
wire g74961_p;
wire g74967_p;
wire g74981_p;
wire g74996_p;
wire TIMEBOOST_net_2864;
wire TIMEBOOST_net_2890;
wire g75024_sb;
wire g75059_p;
wire g75061_p;
wire g75067_p;
wire TIMEBOOST_net_13281;
wire g75072_db;
wire g75072_sb;
wire g75081_p;
wire g75084_p;
wire g75088_p;
wire g75126_p;
wire TIMEBOOST_net_9361;
wire g75160_db;
wire g75160_sb;
wire TIMEBOOST_net_13977;
wire g75162_db;
wire g75162_sb;
wire g75165_p;
wire g75174_p;
wire TIMEBOOST_net_12741;
wire TIMEBOOST_net_14020;
wire g75178_db;
wire g75181_da;
wire g75181_db;
wire g75200_p;
wire g75332_p;
wire g75413_db;
wire g75416_da;
wire g75416_db;
wire g75418_da;
wire g75418_db;
wire g75_p;
wire i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_29__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_31__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid;
wire n_0;
wire n_10002;
wire n_10007;
wire n_10010;
wire n_10014;
wire n_10017;
wire n_10020;
wire n_10023;
wire n_10026;
wire n_10029;
wire n_10032;
wire n_10035;
wire n_10038;
wire n_1004;
wire n_10041;
wire n_10048;
wire n_1005;
wire n_10051;
wire n_10054;
wire n_10057;
wire n_10060;
wire n_10063;
wire n_10066;
wire n_10069;
wire n_1007;
wire n_10075;
wire n_10078;
wire n_1008;
wire n_10081;
wire n_10084;
wire n_10087;
wire n_1009;
wire n_10090;
wire n_10093;
wire n_10096;
wire n_10099;
wire n_10102;
wire n_10105;
wire n_10106;
wire n_10109;
wire n_1011;
wire n_10112;
wire TIMEBOOST_net_9374;
wire n_10116;
wire TIMEBOOST_net_12083;
wire n_1012;
wire n_10120;
wire TIMEBOOST_net_9375;
wire n_10124;
wire n_10127;
wire TIMEBOOST_net_12135;
wire n_1013;
wire n_10131;
wire n_10134;
wire TIMEBOOST_net_12130;
wire TIMEBOOST_net_12075;
wire n_1014;
wire n_10141;
wire n_10143;
wire n_10144;
wire n_10147;
wire TIMEBOOST_net_9372;
wire n_1015;
wire n_10151;
wire n_10154;
wire n_10155;
wire n_10157;
wire n_1016;
wire n_10160;
wire n_10163;
wire TIMEBOOST_net_9438;
wire n_1017;
wire n_10170;
wire n_10173;
wire n_10176;
wire n_10179;
wire TIMEBOOST_net_12161;
wire n_10183;
wire n_10185;
wire n_10188;
wire n_1019;
wire TIMEBOOST_net_12155;
wire n_10193;
wire n_10195;
wire n_10198;
wire TIMEBOOST_net_12173;
wire n_10202;
wire n_10205;
wire TIMEBOOST_net_9373;
wire TIMEBOOST_net_12134;
wire n_10216;
wire n_10221;
wire TIMEBOOST_net_12133;
wire n_1023;
wire n_10230;
wire n_10232;
wire n_10235;
wire TIMEBOOST_net_12131;
wire TIMEBOOST_net_12158;
wire n_10244;
wire TIMEBOOST_net_12082;
wire TIMEBOOST_net_12132;
wire n_10252;
wire n_10254;
wire n_10256;
wire TIMEBOOST_net_12178;
wire n_10258;
wire n_10259;
wire n_10261;
wire TIMEBOOST_net_12174;
wire n_10268;
wire n_1027;
wire n_10270;
wire TIMEBOOST_net_12152;
wire n_10273;
wire TIMEBOOST_net_12166;
wire TIMEBOOST_net_12171;
wire TIMEBOOST_net_3764;
wire TIMEBOOST_net_12154;
wire TIMEBOOST_net_12153;
wire TIMEBOOST_net_12159;
wire n_1028;
wire n_10281;
wire n_10285;
wire n_10286;
wire n_10288;
wire n_10289;
wire n_10290;
wire n_10291;
wire n_10292;
wire n_10294;
wire n_10296;
wire n_10297;
wire n_10298;
wire n_10300;
wire n_10302;
wire n_10304;
wire n_10306;
wire n_10308;
wire n_1031;
wire n_10310;
wire n_10311;
wire n_10312;
wire n_10314;
wire n_10316;
wire n_10317;
wire n_10319;
wire n_10321;
wire n_10323;
wire n_10325;
wire n_10327;
wire n_10329;
wire n_1033;
wire n_10331;
wire n_10332;
wire n_10334;
wire n_10336;
wire n_10338;
wire n_1034;
wire n_10340;
wire n_10342;
wire n_10343;
wire n_10344;
wire n_10346;
wire n_10348;
wire n_10349;
wire n_1035;
wire n_10351;
wire n_10353;
wire n_10355;
wire n_10357;
wire n_10359;
wire n_1036;
wire n_10361;
wire n_10362;
wire n_10363;
wire n_10365;
wire n_10366;
wire n_10368;
wire n_1037;
wire n_10370;
wire n_10372;
wire n_10374;
wire n_10376;
wire n_10377;
wire n_10378;
wire n_1038;
wire n_10380;
wire n_10381;
wire n_10383;
wire n_10384;
wire n_10385;
wire n_10386;
wire n_10388;
wire n_1039;
wire n_10390;
wire n_10391;
wire n_10393;
wire n_10394;
wire n_10396;
wire n_10397;
wire n_10399;
wire n_104;
wire n_10400;
wire n_10401;
wire n_10402;
wire n_10404;
wire n_10405;
wire n_10407;
wire n_10408;
wire n_1041;
wire n_10410;
wire n_10411;
wire n_10412;
wire n_10413;
wire n_10414;
wire n_10416;
wire n_10417;
wire n_10418;
wire n_10419;
wire n_10421;
wire n_10423;
wire n_10424;
wire n_10426;
wire n_10428;
wire n_10430;
wire n_10432;
wire n_10433;
wire n_10434;
wire n_10436;
wire n_10438;
wire n_10439;
wire n_10440;
wire n_10441;
wire n_10443;
wire n_10444;
wire n_10445;
wire n_10446;
wire n_10447;
wire n_10449;
wire n_10450;
wire n_10451;
wire n_10453;
wire n_10455;
wire n_10457;
wire n_10459;
wire n_10460;
wire n_10462;
wire n_10463;
wire n_10464;
wire n_10465;
wire n_10467;
wire n_10469;
wire n_10470;
wire n_10473;
wire n_10474;
wire n_10476;
wire n_10477;
wire n_10478;
wire n_10479;
wire n_10481;
wire n_10483;
wire n_10485;
wire n_10487;
wire n_10489;
wire n_10491;
wire n_10493;
wire n_10495;
wire n_10497;
wire n_10499;
wire n_10501;
wire n_10503;
wire n_10506;
wire n_10508;
wire n_10509;
wire n_10511;
wire n_10513;
wire n_10515;
wire n_10518;
wire n_10521;
wire n_10524;
wire n_10527;
wire n_10530;
wire n_10533;
wire n_10541;
wire n_10544;
wire n_10547;
wire n_10553;
wire n_10554;
wire n_10556;
wire n_10559;
wire n_10560;
wire n_10561;
wire n_10564;
wire n_10566;
wire n_10569;
wire n_1057;
wire n_10572;
wire n_10575;
wire n_10576;
wire n_10577;
wire n_10579;
wire n_10584;
wire n_10588;
wire n_10592;
wire n_10595;
wire n_10596;
wire n_10599;
wire n_10602;
wire n_10605;
wire n_10608;
wire n_1061;
wire n_10611;
wire n_10614;
wire n_10617;
wire n_10622;
wire n_10624;
wire n_10627;
wire n_10630;
wire n_10631;
wire n_10634;
wire n_10637;
wire n_10638;
wire n_1064;
wire n_10641;
wire n_10644;
wire n_10647;
wire n_10650;
wire n_10653;
wire n_10656;
wire n_10659;
wire n_10660;
wire n_10661;
wire n_10662;
wire n_10669;
wire n_10672;
wire n_10675;
wire n_10676;
wire n_10679;
wire n_10680;
wire n_10681;
wire n_10682;
wire n_10685;
wire n_10688;
wire n_1069;
wire n_10691;
wire n_10693;
wire n_10696;
wire n_10699;
wire n_10702;
wire n_10705;
wire n_10708;
wire n_10711;
wire n_10715;
wire n_1072;
wire n_10728;
wire n_1073;
wire n_10731;
wire n_10734;
wire n_10738;
wire n_1074;
wire n_10741;
wire n_10744;
wire n_10747;
wire n_10750;
wire n_10753;
wire n_10754;
wire n_10755;
wire n_10758;
wire n_10763;
wire n_10764;
wire n_10765;
wire n_10768;
wire n_1077;
wire n_10771;
wire n_10774;
wire n_10777;
wire n_10780;
wire n_10781;
wire n_10782;
wire n_10784;
wire n_10785;
wire n_10787;
wire n_10788;
wire n_10789;
wire n_1079;
wire n_10791;
wire n_10792;
wire n_10793;
wire n_10795;
wire n_10797;
wire n_10799;
wire n_1080;
wire n_10800;
wire n_10802;
wire n_10803;
wire n_10804;
wire n_10806;
wire n_10807;
wire n_1081;
wire n_10810;
wire n_10812;
wire n_10813;
wire n_10815;
wire n_10817;
wire n_10819;
wire n_10820;
wire n_10821;
wire n_10823;
wire n_10825;
wire n_10828;
wire n_10829;
wire n_1083;
wire n_10832;
wire n_10833;
wire n_10834;
wire n_10835;
wire n_10836;
wire n_10838;
wire n_10839;
wire n_1084;
wire n_10841;
wire n_10843;
wire n_10845;
wire n_10847;
wire n_10848;
wire n_1085;
wire n_10851;
wire n_10853;
wire n_10855;
wire n_10856;
wire n_10859;
wire n_1086;
wire n_10860;
wire n_10864;
wire n_10865;
wire n_10866;
wire n_10867;
wire n_10870;
wire n_10873;
wire n_10875;
wire n_10876;
wire n_10877;
wire n_1088;
wire n_10880;
wire n_10881;
wire n_10882;
wire n_10885;
wire n_10889;
wire n_1089;
wire n_10890;
wire n_10891;
wire n_10892;
wire n_10895;
wire n_10898;
wire n_10901;
wire n_10902;
wire n_10903;
wire n_10904;
wire n_10905;
wire n_10906;
wire n_10907;
wire n_10908;
wire n_10909;
wire n_1091;
wire n_10912;
wire n_10913;
wire n_10916;
wire n_10917;
wire n_10918;
wire n_10919;
wire n_10922;
wire n_10923;
wire n_10927;
wire n_1093;
wire n_10930;
wire n_10931;
wire n_10932;
wire TIMEBOOST_net_12870;
wire n_10939;
wire n_1094;
wire n_10942;
wire n_10943;
wire n_10944;
wire n_10947;
wire n_1095;
wire n_10951;
wire n_10952;
wire n_10956;
wire n_1096;
wire n_10961;
wire n_10962;
wire n_10963;
wire n_10967;
wire n_10970;
wire n_10971;
wire n_10974;
wire n_10975;
wire n_10976;
wire n_10977;
wire n_10978;
wire n_1098;
wire n_10981;
wire n_10985;
wire n_10986;
wire n_10987;
wire n_1099;
wire n_10991;
wire n_10994;
wire n_11;
wire n_1100;
wire n_11002;
wire n_11005;
wire n_11008;
wire n_1101;
wire n_11013;
wire n_11014;
wire n_11019;
wire n_1103;
wire n_11034;
wire n_11036;
wire n_11037;
wire n_11038;
wire n_11039;
wire n_1104;
wire n_11040;
wire n_11041;
wire n_11042;
wire n_11043;
wire n_11044;
wire n_11046;
wire n_11047;
wire n_11048;
wire n_11049;
wire n_1105;
wire n_11050;
wire n_11051;
wire n_11053;
wire n_11054;
wire n_11055;
wire n_11056;
wire n_11057;
wire n_11058;
wire n_11059;
wire n_1106;
wire n_11060;
wire n_11061;
wire n_11062;
wire n_11063;
wire n_11064;
wire n_11065;
wire n_11066;
wire n_11067;
wire n_11069;
wire n_1107;
wire n_11070;
wire n_11071;
wire n_11072;
wire n_11073;
wire n_11075;
wire n_11076;
wire n_11077;
wire n_11078;
wire n_11079;
wire n_1108;
wire n_11081;
wire n_11083;
wire n_11084;
wire n_11085;
wire n_11086;
wire n_11087;
wire n_11088;
wire n_11089;
wire n_1109;
wire n_11090;
wire n_11091;
wire n_11092;
wire n_11093;
wire n_11094;
wire n_11095;
wire n_11096;
wire n_11097;
wire n_11099;
wire n_1110;
wire n_11100;
wire n_11101;
wire n_11102;
wire n_11104;
wire n_11106;
wire n_11107;
wire n_11108;
wire n_11109;
wire n_1111;
wire n_11110;
wire n_11111;
wire n_11113;
wire n_11115;
wire n_11118;
wire n_11119;
wire n_1112;
wire n_11120;
wire n_11121;
wire n_11122;
wire n_11123;
wire n_11124;
wire n_11125;
wire n_11126;
wire n_11129;
wire n_1113;
wire n_11130;
wire n_11131;
wire n_11132;
wire n_11134;
wire n_11135;
wire n_11136;
wire n_11137;
wire n_11138;
wire n_11139;
wire n_11140;
wire n_11142;
wire n_11143;
wire n_11144;
wire n_11145;
wire n_11146;
wire n_11147;
wire n_11148;
wire n_11149;
wire n_1115;
wire n_11152;
wire n_11153;
wire n_11155;
wire n_11157;
wire n_11158;
wire n_11159;
wire n_1116;
wire n_11161;
wire n_11162;
wire n_11164;
wire n_11165;
wire n_11167;
wire n_11169;
wire n_1117;
wire n_11171;
wire n_11173;
wire n_11174;
wire n_11175;
wire n_11177;
wire n_11178;
wire n_11179;
wire n_1118;
wire n_11180;
wire n_11181;
wire n_11182;
wire n_11184;
wire n_11186;
wire n_11187;
wire n_11188;
wire n_1119;
wire n_11190;
wire n_11191;
wire n_11193;
wire n_11194;
wire n_11196;
wire n_11198;
wire n_112;
wire n_1120;
wire n_11200;
wire n_11202;
wire n_11203;
wire n_11205;
wire n_11206;
wire n_11207;
wire n_11208;
wire n_11209;
wire n_11211;
wire n_11212;
wire n_11213;
wire n_11214;
wire n_11215;
wire n_11216;
wire n_11217;
wire n_11218;
wire n_11219;
wire n_1122;
wire n_11220;
wire n_11222;
wire n_11223;
wire n_11224;
wire n_11226;
wire n_11228;
wire n_11229;
wire n_1123;
wire n_11230;
wire n_11232;
wire n_11234;
wire n_11235;
wire n_11236;
wire n_11238;
wire n_11239;
wire n_1124;
wire n_11240;
wire n_11241;
wire n_11242;
wire n_11243;
wire n_11244;
wire n_11245;
wire n_11246;
wire n_11247;
wire n_11249;
wire n_1125;
wire n_11250;
wire n_11251;
wire n_11252;
wire n_11254;
wire n_11255;
wire n_11256;
wire n_11258;
wire n_11259;
wire n_1126;
wire n_11260;
wire n_11261;
wire n_11262;
wire n_11264;
wire n_11265;
wire n_11266;
wire n_11268;
wire n_11270;
wire n_11271;
wire n_11273;
wire n_11274;
wire n_11276;
wire n_11277;
wire n_11279;
wire n_11280;
wire n_11281;
wire n_11282;
wire n_11283;
wire n_11284;
wire n_11285;
wire n_11286;
wire n_11287;
wire n_11289;
wire n_11290;
wire n_11293;
wire n_11295;
wire n_11297;
wire n_11300;
wire n_11302;
wire n_11303;
wire n_11305;
wire n_11306;
wire n_11307;
wire n_11309;
wire n_11311;
wire n_11314;
wire n_11316;
wire n_11318;
wire n_11320;
wire n_11322;
wire n_11324;
wire n_11326;
wire n_11327;
wire n_11328;
wire n_1133;
wire n_11330;
wire n_11332;
wire n_11334;
wire n_11336;
wire n_11337;
wire n_11338;
wire n_1134;
wire n_11340;
wire n_11342;
wire n_11344;
wire n_11345;
wire n_11347;
wire n_11349;
wire n_11350;
wire n_11352;
wire n_11353;
wire n_11355;
wire n_11357;
wire n_11359;
wire n_11361;
wire n_11362;
wire n_11363;
wire n_11365;
wire n_11367;
wire n_11369;
wire n_11370;
wire n_11372;
wire n_11373;
wire n_11375;
wire n_11377;
wire n_11379;
wire n_11380;
wire n_11381;
wire n_11382;
wire n_11383;
wire n_11384;
wire n_11385;
wire n_11386;
wire n_11388;
wire n_11390;
wire n_11391;
wire n_11393;
wire n_11394;
wire n_11396;
wire n_11398;
wire n_11399;
wire n_11401;
wire n_11402;
wire n_11403;
wire n_11405;
wire n_11406;
wire n_11408;
wire n_11410;
wire n_11411;
wire n_11413;
wire n_11414;
wire n_11415;
wire n_11417;
wire n_11418;
wire n_11419;
wire n_11420;
wire n_11421;
wire n_11423;
wire n_11424;
wire n_11425;
wire n_11427;
wire n_11429;
wire n_11431;
wire n_11432;
wire n_11433;
wire n_11434;
wire n_11435;
wire n_11436;
wire n_11437;
wire n_11438;
wire n_11440;
wire n_11441;
wire n_11442;
wire n_11443;
wire n_11445;
wire n_11446;
wire n_11448;
wire n_11449;
wire n_11450;
wire n_11451;
wire n_11452;
wire n_11454;
wire n_11456;
wire n_11457;
wire n_11458;
wire n_11460;
wire n_11462;
wire n_11463;
wire n_11464;
wire n_11466;
wire n_11467;
wire n_11468;
wire n_11470;
wire n_11472;
wire n_11473;
wire n_11474;
wire n_11476;
wire n_11477;
wire n_11478;
wire n_11479;
wire n_11480;
wire n_11482;
wire n_11483;
wire n_11484;
wire n_11485;
wire n_11487;
wire n_11489;
wire n_11490;
wire n_11492;
wire n_11493;
wire n_11495;
wire n_11496;
wire n_11497;
wire n_11499;
wire n_11500;
wire n_11502;
wire n_11503;
wire n_11505;
wire n_11507;
wire n_11509;
wire n_11510;
wire n_11512;
wire n_11513;
wire n_11515;
wire n_11516;
wire n_11517;
wire n_11519;
wire n_11521;
wire n_11523;
wire n_11524;
wire n_11526;
wire n_11528;
wire n_11530;
wire n_11531;
wire n_11532;
wire n_11533;
wire n_11534;
wire n_11535;
wire n_11536;
wire n_11538;
wire n_11540;
wire n_11542;
wire n_11543;
wire n_11544;
wire n_11545;
wire n_11546;
wire n_11547;
wire n_11548;
wire n_11549;
wire n_11551;
wire n_11553;
wire n_11555;
wire n_11556;
wire n_11557;
wire n_11559;
wire n_11560;
wire n_11561;
wire n_11562;
wire n_11564;
wire n_11565;
wire n_11566;
wire n_11568;
wire n_11570;
wire n_11571;
wire n_11572;
wire n_11573;
wire n_11575;
wire n_11577;
wire n_11579;
wire n_11580;
wire n_11582;
wire n_11583;
wire n_11584;
wire n_11585;
wire n_11586;
wire n_11587;
wire n_11588;
wire n_11589;
wire n_1159;
wire n_11590;
wire n_11592;
wire n_11593;
wire n_11595;
wire n_11597;
wire n_11598;
wire n_11599;
wire n_1160;
wire n_11600;
wire n_11601;
wire n_11602;
wire n_11603;
wire n_11604;
wire n_11605;
wire n_11606;
wire n_11607;
wire n_11609;
wire n_1161;
wire n_11610;
wire n_11611;
wire n_11613;
wire n_11614;
wire n_11616;
wire n_11617;
wire n_11618;
wire n_1162;
wire n_11620;
wire n_11622;
wire n_11623;
wire n_11624;
wire n_11625;
wire n_11626;
wire n_11628;
wire n_11630;
wire n_11631;
wire n_11632;
wire n_11633;
wire n_11634;
wire n_11635;
wire n_11637;
wire n_11638;
wire n_11639;
wire n_1164;
wire n_11640;
wire n_11641;
wire n_11642;
wire n_11644;
wire n_11645;
wire n_11647;
wire n_11648;
wire n_1165;
wire n_11650;
wire n_11651;
wire n_11652;
wire n_11653;
wire n_11655;
wire n_11657;
wire n_11659;
wire n_1166;
wire n_11660;
wire n_11661;
wire n_11662;
wire n_11663;
wire n_11665;
wire n_11666;
wire n_11667;
wire n_11668;
wire n_11669;
wire n_1167;
wire n_11670;
wire n_11671;
wire n_11672;
wire n_11674;
wire n_11675;
wire n_11676;
wire n_11677;
wire n_11679;
wire n_1168;
wire n_11680;
wire n_11681;
wire n_11682;
wire n_11683;
wire n_11684;
wire n_11685;
wire n_11686;
wire n_11687;
wire n_11688;
wire n_11689;
wire n_1169;
wire n_11690;
wire n_11691;
wire n_11692;
wire n_11693;
wire n_11694;
wire n_11695;
wire n_11696;
wire n_11697;
wire n_11698;
wire n_11699;
wire n_1170;
wire n_11700;
wire n_11701;
wire n_11702;
wire n_11703;
wire n_11705;
wire n_11706;
wire n_11707;
wire n_11708;
wire n_11710;
wire n_11712;
wire n_11715;
wire n_11716;
wire n_11717;
wire n_11718;
wire n_11719;
wire n_11720;
wire n_11723;
wire n_11724;
wire n_11725;
wire n_11726;
wire n_11727;
wire n_11728;
wire n_1173;
wire n_11730;
wire n_11731;
wire n_11732;
wire n_11733;
wire n_11734;
wire n_11735;
wire n_11736;
wire n_11738;
wire n_11739;
wire n_1174;
wire n_11740;
wire n_11741;
wire n_1175;
wire n_1176;
wire n_11762;
wire n_11767;
wire n_1177;
wire n_11773;
wire n_11774;
wire n_11775;
wire n_11776;
wire n_11777;
wire n_11778;
wire n_1178;
wire n_11780;
wire n_11781;
wire n_11782;
wire n_11783;
wire n_11784;
wire n_11786;
wire n_11788;
wire n_11790;
wire n_11791;
wire n_11792;
wire n_11793;
wire n_11795;
wire n_11796;
wire TIMEBOOST_net_15104;
wire n_1180;
wire TIMEBOOST_net_12214;
wire TIMEBOOST_net_13410;
wire TIMEBOOST_net_12903;
wire TIMEBOOST_net_15065;
wire n_11805;
wire n_11806;
wire TIMEBOOST_net_12426;
wire TIMEBOOST_net_9505;
wire TIMEBOOST_net_15101;
wire TIMEBOOST_net_12439;
wire TIMEBOOST_net_12905;
wire TIMEBOOST_net_14629;
wire n_11814;
wire TIMEBOOST_net_9497;
wire n_11816;
wire TIMEBOOST_net_12418;
wire n_11818;
wire n_11819;
wire TIMEBOOST_net_15064;
wire TIMEBOOST_net_12438;
wire n_11822;
wire n_11823;
wire TIMEBOOST_net_12828;
wire TIMEBOOST_net_9495;
wire TIMEBOOST_net_12879;
wire TIMEBOOST_net_12829;
wire n_1183;
wire TIMEBOOST_net_9502;
wire n_11831;
wire TIMEBOOST_net_12428;
wire TIMEBOOST_net_12863;
wire TIMEBOOST_net_12441;
wire TIMEBOOST_net_15071;
wire n_11838;
wire n_11839;
wire n_11840;
wire n_11841;
wire TIMEBOOST_net_9515;
wire TIMEBOOST_net_12424;
wire n_11844;
wire n_11845;
wire n_11846;
wire n_11847;
wire n_11848;
wire n_11849;
wire n_1185;
wire n_11850;
wire n_11851;
wire n_11852;
wire n_11853;
wire n_11854;
wire n_11855;
wire n_11856;
wire n_11857;
wire n_11858;
wire n_11859;
wire n_1186;
wire n_11860;
wire n_11861;
wire n_11862;
wire n_11863;
wire n_11864;
wire n_11865;
wire n_11866;
wire n_11867;
wire n_11868;
wire n_11869;
wire n_1187;
wire n_11870;
wire n_11871;
wire n_11872;
wire n_11873;
wire n_11874;
wire n_11875;
wire n_11876;
wire n_11877;
wire n_11878;
wire n_1188;
wire n_11880;
wire n_11881;
wire n_11884;
wire n_11885;
wire TIMEBOOST_net_14783;
wire n_11887;
wire TIMEBOOST_net_12483;
wire TIMEBOOST_net_9443;
wire n_1189;
wire n_11890;
wire n_11891;
wire TIMEBOOST_net_15144;
wire n_11893;
wire TIMEBOOST_net_12866;
wire n_11895;
wire n_11896;
wire n_11897;
wire n_11898;
wire n_119;
wire n_1190;
wire n_11900;
wire TIMEBOOST_net_12410;
wire TIMEBOOST_net_15077;
wire n_11903;
wire TIMEBOOST_net_12904;
wire TIMEBOOST_net_15111;
wire TIMEBOOST_net_15137;
wire n_11907;
wire n_11908;
wire n_1191;
wire n_11910;
wire TIMEBOOST_net_9466;
wire n_11912;
wire n_11913;
wire n_11914;
wire n_11915;
wire n_11916;
wire TIMEBOOST_net_9513;
wire TIMEBOOST_net_12473;
wire TIMEBOOST_net_9491;
wire n_1192;
wire n_11920;
wire n_11921;
wire n_11923;
wire n_11924;
wire n_11925;
wire TIMEBOOST_net_15075;
wire n_11927;
wire n_11929;
wire n_1193;
wire n_11930;
wire n_11932;
wire n_11933;
wire n_11934;
wire TIMEBOOST_net_9521;
wire n_11937;
wire n_11938;
wire n_1194;
wire TIMEBOOST_net_9504;
wire TIMEBOOST_net_9520;
wire TIMEBOOST_net_9490;
wire TIMEBOOST_net_12458;
wire TIMEBOOST_net_15141;
wire TIMEBOOST_net_9512;
wire n_11948;
wire n_11949;
wire n_1195;
wire TIMEBOOST_net_9442;
wire n_11951;
wire n_11952;
wire n_11953;
wire n_11954;
wire TIMEBOOST_net_15139;
wire n_11956;
wire n_11957;
wire TIMEBOOST_net_9511;
wire TIMEBOOST_net_15066;
wire n_1196;
wire n_11960;
wire n_11961;
wire n_11962;
wire n_11964;
wire TIMEBOOST_net_15095;
wire TIMEBOOST_net_9496;
wire TIMEBOOST_net_12465;
wire n_11968;
wire n_1197;
wire n_11970;
wire TIMEBOOST_net_9510;
wire n_11972;
wire n_11973;
wire TIMEBOOST_net_15215;
wire n_11975;
wire n_11977;
wire n_11978;
wire TIMEBOOST_net_15142;
wire n_1198;
wire TIMEBOOST_net_15099;
wire TIMEBOOST_net_9441;
wire n_11984;
wire TIMEBOOST_net_9509;
wire n_11988;
wire n_1199;
wire n_11990;
wire n_11991;
wire n_11992;
wire TIMEBOOST_net_12894;
wire n_11995;
wire n_11996;
wire TIMEBOOST_net_15067;
wire TIMEBOOST_net_15110;
wire n_12;
wire n_1200;
wire n_12000;
wire n_12001;
wire n_12002;
wire n_12003;
wire n_12004;
wire TIMEBOOST_net_15096;
wire TIMEBOOST_net_9440;
wire n_12007;
wire n_12008;
wire n_12009;
wire n_1201;
wire n_12010;
wire n_12011;
wire TIMEBOOST_net_15130;
wire TIMEBOOST_net_9508;
wire TIMEBOOST_net_12572;
wire TIMEBOOST_net_12864;
wire TIMEBOOST_net_15195;
wire TIMEBOOST_net_15143;
wire n_1202;
wire n_12020;
wire TIMEBOOST_net_12718;
wire n_12022;
wire TIMEBOOST_net_12211;
wire n_12024;
wire TIMEBOOST_net_12464;
wire TIMEBOOST_net_15159;
wire n_12028;
wire TIMEBOOST_net_12210;
wire n_12031;
wire n_12032;
wire TIMEBOOST_net_9507;
wire n_12035;
wire n_12036;
wire n_12037;
wire n_12038;
wire n_1204;
wire n_12041;
wire TIMEBOOST_net_9465;
wire n_12044;
wire n_12045;
wire TIMEBOOST_net_15086;
wire n_12047;
wire n_12049;
wire TIMEBOOST_net_12773;
wire n_12051;
wire n_12052;
wire n_12053;
wire n_12054;
wire n_12055;
wire n_12056;
wire TIMEBOOST_net_12848;
wire n_12058;
wire TIMEBOOST_net_15087;
wire TIMEBOOST_net_12559;
wire n_12061;
wire TIMEBOOST_net_12193;
wire TIMEBOOST_net_12480;
wire TIMEBOOST_net_15092;
wire TIMEBOOST_net_12544;
wire n_12066;
wire TIMEBOOST_net_15080;
wire n_12068;
wire TIMEBOOST_net_15093;
wire n_1207;
wire n_12070;
wire TIMEBOOST_net_15124;
wire n_12072;
wire n_12073;
wire TIMEBOOST_net_12459;
wire n_12075;
wire TIMEBOOST_net_15136;
wire n_12078;
wire n_1208;
wire TIMEBOOST_net_15121;
wire n_12081;
wire TIMEBOOST_net_12550;
wire n_12084;
wire TIMEBOOST_net_12549;
wire TIMEBOOST_net_15120;
wire n_12088;
wire n_1209;
wire n_12090;
wire TIMEBOOST_net_15091;
wire TIMEBOOST_net_15090;
wire TIMEBOOST_net_12524;
wire TIMEBOOST_net_12557;
wire n_12097;
wire n_12099;
wire n_1210;
wire n_12100;
wire n_12101;
wire TIMEBOOST_net_15129;
wire TIMEBOOST_net_15089;
wire n_12104;
wire TIMEBOOST_net_15079;
wire TIMEBOOST_net_15193;
wire TIMEBOOST_net_15214;
wire TIMEBOOST_net_12556;
wire n_1211;
wire TIMEBOOST_net_15173;
wire TIMEBOOST_net_12199;
wire n_12112;
wire n_12113;
wire TIMEBOOST_net_15114;
wire n_12115;
wire n_12116;
wire n_12117;
wire TIMEBOOST_net_9481;
wire TIMEBOOST_net_15109;
wire TIMEBOOST_net_9485;
wire n_12122;
wire n_12124;
wire TIMEBOOST_net_12843;
wire n_12128;
wire n_12129;
wire n_1213;
wire n_12130;
wire n_12132;
wire n_12133;
wire n_12134;
wire n_12135;
wire n_12137;
wire n_12139;
wire n_12140;
wire n_12141;
wire n_12143;
wire n_12144;
wire n_12145;
wire n_12146;
wire n_12147;
wire n_12148;
wire n_1215;
wire n_12151;
wire n_12153;
wire n_12154;
wire n_12155;
wire n_12156;
wire n_12158;
wire n_12159;
wire n_1216;
wire n_12160;
wire n_12161;
wire n_12162;
wire n_12163;
wire n_12164;
wire n_12165;
wire n_12166;
wire n_12167;
wire n_12168;
wire n_12169;
wire n_1217;
wire n_12170;
wire n_12179;
wire n_1218;
wire TIMEBOOST_net_12501;
wire TIMEBOOST_net_12840;
wire TIMEBOOST_net_12191;
wire TIMEBOOST_net_14849;
wire TIMEBOOST_net_12578;
wire n_12186;
wire TIMEBOOST_net_15134;
wire TIMEBOOST_net_9506;
wire TIMEBOOST_net_12584;
wire n_1219;
wire TIMEBOOST_net_15078;
wire TIMEBOOST_net_12832;
wire TIMEBOOST_net_15072;
wire n_12194;
wire n_12195;
wire n_12196;
wire n_12197;
wire n_12198;
wire TIMEBOOST_net_15133;
wire n_1220;
wire n_12201;
wire n_12202;
wire n_12203;
wire TIMEBOOST_net_9498;
wire TIMEBOOST_net_12213;
wire n_12206;
wire n_12207;
wire n_12208;
wire n_1221;
wire TIMEBOOST_net_15122;
wire TIMEBOOST_net_12417;
wire n_12212;
wire TIMEBOOST_net_15105;
wire TIMEBOOST_net_12447;
wire n_12215;
wire TIMEBOOST_net_15076;
wire TIMEBOOST_net_12585;
wire n_12220;
wire TIMEBOOST_net_15145;
wire n_12222;
wire TIMEBOOST_net_15074;
wire n_12224;
wire TIMEBOOST_net_15119;
wire n_12227;
wire n_12228;
wire TIMEBOOST_net_9445;
wire TIMEBOOST_net_12583;
wire TIMEBOOST_net_15084;
wire TIMEBOOST_net_15128;
wire TIMEBOOST_net_12446;
wire n_12235;
wire n_12236;
wire n_12237;
wire n_12238;
wire TIMEBOOST_net_13855;
wire n_1224;
wire TIMEBOOST_net_15073;
wire n_12242;
wire n_12243;
wire n_12244;
wire n_12245;
wire n_12246;
wire n_12248;
wire n_1225;
wire n_12250;
wire TIMEBOOST_net_12437;
wire TIMEBOOST_net_15069;
wire TIMEBOOST_net_12525;
wire TIMEBOOST_net_14793;
wire n_12257;
wire n_12258;
wire n_12259;
wire n_1226;
wire TIMEBOOST_net_15100;
wire n_12264;
wire n_12266;
wire n_12267;
wire TIMEBOOST_net_15131;
wire TIMEBOOST_net_15068;
wire n_1227;
wire TIMEBOOST_net_15098;
wire n_12271;
wire TIMEBOOST_net_12587;
wire n_12273;
wire n_12274;
wire n_12275;
wire n_12276;
wire n_12277;
wire TIMEBOOST_net_12176;
wire n_1228;
wire n_12280;
wire n_12282;
wire n_12283;
wire TIMEBOOST_net_12896;
wire TIMEBOOST_net_15118;
wire n_12289;
wire n_1229;
wire n_12290;
wire TIMEBOOST_net_15108;
wire n_12292;
wire n_12293;
wire n_12294;
wire TIMEBOOST_net_15094;
wire TIMEBOOST_net_9494;
wire TIMEBOOST_net_12212;
wire n_123;
wire n_1230;
wire n_12300;
wire TIMEBOOST_net_12594;
wire TIMEBOOST_net_12440;
wire TIMEBOOST_net_15081;
wire TIMEBOOST_net_9493;
wire TIMEBOOST_net_12456;
wire n_12309;
wire n_1231;
wire n_12310;
wire TIMEBOOST_net_12208;
wire n_12313;
wire TIMEBOOST_net_15106;
wire TIMEBOOST_net_12425;
wire n_12318;
wire TIMEBOOST_net_12527;
wire TIMEBOOST_net_15070;
wire TIMEBOOST_net_15107;
wire TIMEBOOST_net_9492;
wire n_12323;
wire n_12325;
wire n_12326;
wire n_12327;
wire TIMEBOOST_net_12209;
wire TIMEBOOST_net_15103;
wire TIMEBOOST_net_12431;
wire n_12331;
wire TIMEBOOST_net_12175;
wire n_12334;
wire TIMEBOOST_net_12477;
wire TIMEBOOST_net_15117;
wire n_12337;
wire n_12338;
wire TIMEBOOST_net_15146;
wire TIMEBOOST_net_12767;
wire n_12341;
wire TIMEBOOST_net_15132;
wire TIMEBOOST_net_12768;
wire TIMEBOOST_net_12769;
wire n_12346;
wire n_12348;
wire TIMEBOOST_net_15198;
wire n_12351;
wire n_12352;
wire TIMEBOOST_net_12471;
wire TIMEBOOST_net_12457;
wire n_12356;
wire n_12357;
wire TIMEBOOST_net_15127;
wire TIMEBOOST_net_9475;
wire TIMEBOOST_net_15126;
wire n_12362;
wire n_12363;
wire n_12366;
wire TIMEBOOST_net_12470;
wire n_12369;
wire TIMEBOOST_net_15116;
wire n_12371;
wire n_12372;
wire TIMEBOOST_net_15147;
wire n_12374;
wire n_12375;
wire n_12376;
wire n_12378;
wire n_12379;
wire n_1238;
wire TIMEBOOST_net_12476;
wire n_12381;
wire n_12382;
wire n_12383;
wire TIMEBOOST_net_12558;
wire TIMEBOOST_net_12770;
wire n_12389;
wire TIMEBOOST_net_12468;
wire TIMEBOOST_net_9473;
wire n_12393;
wire TIMEBOOST_net_15125;
wire TIMEBOOST_net_9472;
wire TIMEBOOST_net_12489;
wire TIMEBOOST_net_12771;
wire TIMEBOOST_net_15115;
wire n_12402;
wire TIMEBOOST_net_15158;
wire TIMEBOOST_net_15199;
wire n_12406;
wire n_12408;
wire n_1241;
wire TIMEBOOST_net_12192;
wire TIMEBOOST_net_15157;
wire TIMEBOOST_net_12478;
wire n_12413;
wire TIMEBOOST_net_9470;
wire TIMEBOOST_net_15102;
wire n_12417;
wire TIMEBOOST_net_12488;
wire TIMEBOOST_net_12772;
wire TIMEBOOST_net_15154;
wire TIMEBOOST_net_15194;
wire n_12423;
wire TIMEBOOST_net_12564;
wire n_12425;
wire TIMEBOOST_net_9486;
wire n_12427;
wire n_12429;
wire n_12430;
wire TIMEBOOST_net_9484;
wire n_12433;
wire TIMEBOOST_net_12765;
wire TIMEBOOST_net_9483;
wire TIMEBOOST_net_12766;
wire TIMEBOOST_net_15113;
wire n_12439;
wire n_12440;
wire n_12441;
wire n_12442;
wire n_12446;
wire n_12447;
wire n_12448;
wire n_12449;
wire n_12450;
wire n_12451;
wire n_12452;
wire n_12453;
wire n_12454;
wire n_12455;
wire n_12457;
wire n_12459;
wire n_12460;
wire n_12461;
wire n_12462;
wire n_12463;
wire n_12464;
wire n_12465;
wire n_12466;
wire n_12468;
wire n_12469;
wire n_12471;
wire TIMEBOOST_net_2843;
wire n_12473;
wire n_12474;
wire n_12475;
wire n_12476;
wire n_12478;
wire n_12479;
wire n_1248;
wire n_12480;
wire n_12481;
wire n_12483;
wire n_12484;
wire n_12485;
wire n_12486;
wire n_12487;
wire n_12488;
wire n_12489;
wire n_12490;
wire n_12491;
wire n_12492;
wire n_12493;
wire n_12494;
wire n_12495;
wire n_12496;
wire n_12498;
wire n_12499;
wire n_12500;
wire n_12501;
wire n_12502;
wire n_12503;
wire n_12504;
wire n_12505;
wire n_12506;
wire n_12507;
wire n_12508;
wire n_12509;
wire n_1251;
wire n_12510;
wire n_12511;
wire n_12512;
wire n_12513;
wire n_12514;
wire n_12515;
wire n_12516;
wire n_12517;
wire n_12518;
wire n_12519;
wire n_1252;
wire n_12520;
wire n_12521;
wire n_12522;
wire n_12523;
wire n_12524;
wire n_12525;
wire n_12526;
wire n_12527;
wire n_12528;
wire n_12529;
wire n_1253;
wire n_12530;
wire n_12531;
wire n_12532;
wire n_12533;
wire n_12534;
wire n_12535;
wire n_12536;
wire n_12537;
wire n_12538;
wire n_12539;
wire n_12540;
wire n_12541;
wire n_12542;
wire n_12543;
wire n_12544;
wire n_12545;
wire n_12546;
wire n_12547;
wire n_12548;
wire n_12549;
wire n_12550;
wire n_12551;
wire n_12552;
wire n_12553;
wire n_12554;
wire n_12555;
wire n_12556;
wire n_12557;
wire n_12558;
wire n_12559;
wire n_12560;
wire n_12561;
wire n_12562;
wire n_12563;
wire n_12564;
wire n_12565;
wire n_12566;
wire n_12567;
wire n_12568;
wire n_12569;
wire n_12570;
wire n_12571;
wire n_12572;
wire n_12573;
wire n_12574;
wire n_12575;
wire n_12577;
wire n_12578;
wire n_12579;
wire n_1258;
wire n_12580;
wire n_12581;
wire n_12583;
wire n_12584;
wire n_12585;
wire n_12586;
wire n_12587;
wire n_12588;
wire n_12589;
wire n_1259;
wire n_12590;
wire n_12591;
wire n_12595;
wire n_12596;
wire n_12597;
wire n_12598;
wire n_12599;
wire n_1260;
wire n_12600;
wire n_12602;
wire n_12603;
wire n_12604;
wire n_12605;
wire n_12606;
wire n_12607;
wire n_1261;
wire n_12610;
wire n_12611;
wire n_12612;
wire n_12613;
wire n_12614;
wire n_12615;
wire n_12616;
wire n_12617;
wire n_12618;
wire n_12619;
wire n_12620;
wire n_12621;
wire n_12622;
wire n_12623;
wire n_12624;
wire n_12625;
wire n_12626;
wire n_12628;
wire n_12629;
wire n_1263;
wire n_12630;
wire n_12631;
wire n_12632;
wire n_12633;
wire n_12634;
wire n_12635;
wire n_12636;
wire n_12637;
wire n_12638;
wire n_12639;
wire n_1264;
wire n_12640;
wire n_12641;
wire n_12642;
wire n_12643;
wire n_12644;
wire n_12645;
wire n_12646;
wire n_12647;
wire n_12648;
wire n_12649;
wire n_1265;
wire n_12650;
wire n_12651;
wire n_12652;
wire n_12653;
wire n_12654;
wire n_12655;
wire n_12656;
wire n_12658;
wire n_12659;
wire n_1266;
wire n_12660;
wire n_12661;
wire n_12662;
wire n_12663;
wire n_12664;
wire n_12665;
wire n_12666;
wire n_12667;
wire n_12668;
wire n_12669;
wire n_12670;
wire n_12671;
wire n_12672;
wire n_12673;
wire n_12674;
wire n_12675;
wire n_12676;
wire n_12677;
wire n_12678;
wire n_12679;
wire n_12680;
wire n_12681;
wire n_12682;
wire n_12683;
wire n_12684;
wire n_12685;
wire n_12686;
wire n_12688;
wire n_12689;
wire n_1269;
wire n_12692;
wire n_12693;
wire n_12695;
wire n_12696;
wire n_12697;
wire n_12699;
wire n_1270;
wire n_12700;
wire n_12701;
wire n_12702;
wire n_12703;
wire n_12704;
wire n_12705;
wire n_12706;
wire n_12707;
wire n_12709;
wire n_12710;
wire n_12711;
wire n_12712;
wire n_12713;
wire n_12714;
wire n_12715;
wire n_12716;
wire n_12717;
wire n_1272;
wire n_12720;
wire n_12721;
wire n_12722;
wire n_12723;
wire n_12724;
wire n_12725;
wire n_12726;
wire n_12727;
wire n_12728;
wire n_12729;
wire n_1273;
wire n_12731;
wire n_12732;
wire n_12733;
wire n_12734;
wire n_12735;
wire n_12736;
wire n_12737;
wire n_12738;
wire n_1274;
wire n_12741;
wire n_12742;
wire n_12743;
wire n_12744;
wire n_12745;
wire n_12746;
wire n_12747;
wire n_12748;
wire n_12749;
wire n_1275;
wire n_12750;
wire n_12751;
wire n_12752;
wire n_12753;
wire n_12754;
wire n_12756;
wire n_12757;
wire n_12758;
wire n_12759;
wire n_1276;
wire n_12760;
wire n_12761;
wire n_12762;
wire n_12763;
wire n_12764;
wire n_12765;
wire n_12766;
wire n_12767;
wire n_12768;
wire n_12769;
wire n_1277;
wire n_12770;
wire n_12771;
wire n_12772;
wire n_12773;
wire n_12774;
wire n_12775;
wire n_12776;
wire n_12778;
wire n_12779;
wire n_12780;
wire n_12781;
wire n_12783;
wire n_12784;
wire n_12785;
wire n_12786;
wire n_12787;
wire n_12788;
wire n_12789;
wire n_1279;
wire n_12790;
wire n_12791;
wire n_12792;
wire n_12795;
wire n_12797;
wire n_12799;
wire n_1280;
wire n_12801;
wire n_12805;
wire n_12806;
wire n_12809;
wire n_1281;
wire n_12810;
wire n_12811;
wire n_12812;
wire n_12813;
wire n_12814;
wire n_12815;
wire n_12816;
wire n_12817;
wire n_12818;
wire n_12819;
wire n_1282;
wire n_12821;
wire n_12822;
wire n_12823;
wire n_12824;
wire n_12825;
wire n_12826;
wire n_12827;
wire n_12828;
wire n_12829;
wire n_1283;
wire n_12830;
wire n_12831;
wire n_12832;
wire n_12833;
wire n_12834;
wire n_12835;
wire n_12836;
wire n_12837;
wire n_12839;
wire n_1284;
wire n_12840;
wire n_12841;
wire n_12842;
wire n_12843;
wire n_12845;
wire n_12846;
wire n_12847;
wire n_12848;
wire n_12849;
wire n_1285;
wire n_12850;
wire n_12851;
wire n_12852;
wire n_12853;
wire n_12855;
wire n_12858;
wire n_12859;
wire n_1286;
wire n_12862;
wire n_12863;
wire n_12864;
wire n_12865;
wire n_12866;
wire n_12867;
wire n_12868;
wire n_12869;
wire n_1287;
wire n_12870;
wire n_12871;
wire n_12872;
wire n_12873;
wire n_12874;
wire n_12875;
wire n_12876;
wire n_12877;
wire n_12878;
wire n_12879;
wire n_1288;
wire n_12880;
wire n_12881;
wire n_12882;
wire n_12883;
wire n_12884;
wire n_12885;
wire n_12886;
wire n_12887;
wire n_12888;
wire n_12889;
wire n_1289;
wire n_12890;
wire n_12891;
wire n_12892;
wire n_12893;
wire n_12894;
wire n_12895;
wire n_12896;
wire n_12897;
wire n_12898;
wire n_12899;
wire n_1290;
wire n_12900;
wire n_12901;
wire n_12902;
wire n_12903;
wire n_12904;
wire n_12905;
wire n_12906;
wire n_12907;
wire n_12908;
wire n_1291;
wire n_12911;
wire n_12912;
wire n_12913;
wire n_12914;
wire n_12915;
wire n_12916;
wire n_12917;
wire n_12918;
wire n_12919;
wire n_12920;
wire n_12921;
wire n_12922;
wire n_12923;
wire n_12924;
wire n_12927;
wire n_12928;
wire n_12929;
wire n_1293;
wire n_12930;
wire n_12931;
wire n_12932;
wire n_12933;
wire n_12934;
wire n_12935;
wire n_12936;
wire n_12937;
wire n_12938;
wire n_12939;
wire n_1294;
wire n_12940;
wire n_12941;
wire n_12942;
wire n_12943;
wire n_12946;
wire n_12947;
wire n_12948;
wire n_12949;
wire n_12950;
wire n_12951;
wire n_12952;
wire n_12954;
wire n_12956;
wire n_12957;
wire n_12958;
wire n_12959;
wire n_12960;
wire n_12961;
wire n_12962;
wire n_12963;
wire n_12964;
wire n_12966;
wire n_12968;
wire n_12970;
wire n_12972;
wire n_12974;
wire n_12976;
wire n_12978;
wire n_12980;
wire n_12981;
wire n_12982;
wire n_12983;
wire n_12984;
wire n_12985;
wire n_12986;
wire n_12988;
wire n_1299;
wire n_12992;
wire n_12994;
wire TIMEBOOST_net_12703;
wire n_12998;
wire n_13000;
wire TIMEBOOST_net_12384;
wire TIMEBOOST_net_1170;
wire TIMEBOOST_net_4564;
wire TIMEBOOST_net_15014;
wire n_13010;
wire n_13012;
wire TIMEBOOST_net_727;
wire n_13018;
wire n_13020;
wire n_13022;
wire n_13026;
wire n_13027;
wire n_13028;
wire n_13034;
wire n_1304;
wire n_13041;
wire n_13042;
wire n_13043;
wire n_13044;
wire n_13045;
wire n_13046;
wire n_13047;
wire n_13048;
wire n_13049;
wire n_13050;
wire n_13051;
wire n_13052;
wire n_13053;
wire n_13054;
wire n_13055;
wire n_13056;
wire n_13057;
wire n_13058;
wire n_13059;
wire n_1306;
wire n_13060;
wire n_13061;
wire n_13063;
wire n_13064;
wire n_13065;
wire n_13066;
wire n_13067;
wire n_13068;
wire n_13073;
wire n_13074;
wire n_13075;
wire n_13076;
wire n_13077;
wire n_13078;
wire n_13079;
wire n_13080;
wire n_13081;
wire n_13082;
wire n_13083;
wire n_13084;
wire n_13085;
wire n_13086;
wire n_13087;
wire n_13088;
wire n_13089;
wire n_13090;
wire n_13091;
wire n_13093;
wire n_13094;
wire n_13095;
wire n_13097;
wire n_13098;
wire TIMEBOOST_net_12704;
wire n_13102;
wire n_13104;
wire n_13105;
wire n_13106;
wire TIMEBOOST_net_10924;
wire TIMEBOOST_net_893;
wire TIMEBOOST_net_890;
wire TIMEBOOST_net_856;
wire TIMEBOOST_net_12379;
wire TIMEBOOST_net_851;
wire n_13116;
wire n_13117;
wire n_13118;
wire n_13120;
wire n_13122;
wire n_13123;
wire n_13124;
wire n_13125;
wire n_13127;
wire n_13128;
wire n_13129;
wire n_13130;
wire n_13131;
wire n_13132;
wire n_13133;
wire n_13134;
wire n_13135;
wire n_13136;
wire n_13137;
wire n_13138;
wire n_13139;
wire n_13140;
wire n_13141;
wire n_13142;
wire n_13143;
wire n_13144;
wire n_13145;
wire n_13146;
wire TIMEBOOST_net_12698;
wire n_1315;
wire TIMEBOOST_net_10144;
wire TIMEBOOST_net_10945;
wire TIMEBOOST_net_865;
wire TIMEBOOST_net_12675;
wire n_1316;
wire TIMEBOOST_net_864;
wire n_13161;
wire n_13162;
wire n_13163;
wire n_13164;
wire n_13165;
wire n_13166;
wire n_13167;
wire n_13168;
wire n_13169;
wire n_1317;
wire n_13170;
wire n_13171;
wire n_13172;
wire n_13173;
wire n_13174;
wire n_13175;
wire n_13176;
wire n_13177;
wire n_13178;
wire n_13179;
wire n_1318;
wire n_13180;
wire n_13181;
wire n_13182;
wire n_13183;
wire n_13184;
wire n_13185;
wire n_13186;
wire TIMEBOOST_net_898;
wire TIMEBOOST_net_1202;
wire TIMEBOOST_net_897;
wire TIMEBOOST_net_13899;
wire TIMEBOOST_net_896;
wire TIMEBOOST_net_895;
wire TIMEBOOST_net_1201;
wire TIMEBOOST_net_13813;
wire TIMEBOOST_net_14983;
wire TIMEBOOST_net_14982;
wire TIMEBOOST_net_14763;
wire TIMEBOOST_net_1197;
wire TIMEBOOST_net_10770;
wire TIMEBOOST_net_1195;
wire TIMEBOOST_net_9660;
wire TIMEBOOST_net_891;
wire TIMEBOOST_net_1193;
wire TIMEBOOST_net_889;
wire TIMEBOOST_net_13335;
wire TIMEBOOST_net_888;
wire TIMEBOOST_net_9658;
wire TIMEBOOST_net_10823;
wire TIMEBOOST_net_1190;
wire TIMEBOOST_net_9657;
wire n_13218;
wire TIMEBOOST_net_887;
wire n_1322;
wire TIMEBOOST_net_1188;
wire n_13221;
wire TIMEBOOST_net_14220;
wire n_13223;
wire TIMEBOOST_net_1187;
wire TIMEBOOST_net_1186;
wire TIMEBOOST_net_9656;
wire n_13228;
wire TIMEBOOST_net_14059;
wire n_1323;
wire TIMEBOOST_net_862;
wire TIMEBOOST_net_861;
wire TIMEBOOST_net_860;
wire TIMEBOOST_net_859;
wire TIMEBOOST_net_858;
wire TIMEBOOST_net_857;
wire TIMEBOOST_net_14755;
wire TIMEBOOST_net_14828;
wire n_13249;
wire n_1325;
wire TIMEBOOST_net_12652;
wire TIMEBOOST_net_12380;
wire TIMEBOOST_net_855;
wire TIMEBOOST_net_12663;
wire n_1326;
wire TIMEBOOST_net_854;
wire TIMEBOOST_net_4130;
wire TIMEBOOST_net_12679;
wire n_1327;
wire TIMEBOOST_net_92;
wire n_13273;
wire TIMEBOOST_net_12717;
wire TIMEBOOST_net_9450;
wire TIMEBOOST_net_12678;
wire TIMEBOOST_net_12696;
wire TIMEBOOST_net_14641;
wire n_13286;
wire n_13287;
wire n_13289;
wire n_1329;
wire n_13290;
wire n_13291;
wire n_13292;
wire n_13295;
wire n_1330;
wire n_13302;
wire n_13303;
wire n_13304;
wire n_13305;
wire n_13306;
wire n_13308;
wire n_13309;
wire n_1331;
wire n_13310;
wire n_13311;
wire n_13313;
wire n_13314;
wire n_13315;
wire n_13317;
wire n_13318;
wire n_13319;
wire n_1332;
wire n_13320;
wire n_13321;
wire n_13323;
wire n_13325;
wire TIMEBOOST_net_1196;
wire n_13327;
wire n_13328;
wire n_13329;
wire n_1333;
wire TIMEBOOST_net_4131;
wire n_13332;
wire n_13333;
wire n_13334;
wire n_13335;
wire TIMEBOOST_net_13007;
wire n_13337;
wire n_13338;
wire n_13339;
wire n_1334;
wire n_13340;
wire n_13341;
wire n_13342;
wire n_1953;
wire TIMEBOOST_net_12966;
wire TIMEBOOST_net_13240;
wire n_13346;
wire TIMEBOOST_net_12958;
wire n_13348;
wire n_13349;
wire n_1335;
wire n_13350;
wire n_13353;
wire n_13354;
wire n_13355;
wire g64972_db;
wire n_13357;
wire n_13358;
wire n_13359;
wire n_13360;
wire n_13361;
wire n_13362;
wire n_13363;
wire n_13365;
wire n_13366;
wire n_13367;
wire n_13368;
wire n_13369;
wire n_1337;
wire n_13370;
wire n_13371;
wire n_13372;
wire n_13373;
wire n_13374;
wire n_13375;
wire n_13376;
wire n_13377;
wire n_13378;
wire n_13379;
wire n_1338;
wire n_13380;
wire n_13381;
wire n_13383;
wire n_13384;
wire n_13386;
wire n_13387;
wire n_13388;
wire n_13389;
wire n_13390;
wire n_13391;
wire n_13392;
wire n_13393;
wire n_13394;
wire n_13395;
wire n_13398;
wire n_13399;
wire n_1340;
wire n_13400;
wire n_13401;
wire n_13402;
wire n_13403;
wire n_13404;
wire n_13405;
wire n_13406;
wire n_13407;
wire n_13408;
wire n_13409;
wire n_1341;
wire n_13410;
wire n_13411;
wire n_13412;
wire n_13414;
wire n_13415;
wire n_13416;
wire n_13417;
wire n_13418;
wire n_13419;
wire n_1342;
wire n_13420;
wire n_13421;
wire n_13422;
wire n_13423;
wire n_13424;
wire n_13425;
wire n_13426;
wire n_13427;
wire n_13428;
wire n_13429;
wire n_1343;
wire n_13430;
wire n_13431;
wire n_13432;
wire n_13434;
wire n_13435;
wire TIMEBOOST_net_10593;
wire TIMEBOOST_net_14878;
wire TIMEBOOST_net_10509;
wire n_13439;
wire n_1344;
wire n_13441;
wire n_13442;
wire n_13444;
wire n_13445;
wire n_13446;
wire n_13447;
wire n_13448;
wire n_13449;
wire n_1345;
wire n_13450;
wire TIMEBOOST_net_10768;
wire n_13453;
wire n_13454;
wire n_13455;
wire TIMEBOOST_net_13972;
wire n_1346;
wire TIMEBOOST_net_10484;
wire n_13461;
wire n_13463;
wire n_13464;
wire TIMEBOOST_net_10485;
wire n_13467;
wire n_13468;
wire n_13469;
wire n_1347;
wire n_13470;
wire n_13474;
wire n_13475;
wire n_13479;
wire n_13481;
wire n_13482;
wire n_13483;
wire n_13484;
wire n_13485;
wire n_13486;
wire n_13487;
wire n_13488;
wire TIMEBOOST_net_13320;
wire n_1349;
wire n_13490;
wire n_13491;
wire n_13493;
wire n_13494;
wire n_13495;
wire n_13496;
wire n_13497;
wire n_13499;
wire n_135;
wire n_1350;
wire n_13500;
wire n_13502;
wire n_13503;
wire n_13504;
wire n_13505;
wire n_13506;
wire n_13508;
wire n_13509;
wire n_1351;
wire n_13511;
wire n_13512;
wire n_13513;
wire n_13514;
wire n_13515;
wire n_13516;
wire n_13517;
wire n_13518;
wire n_13519;
wire n_1352;
wire n_13520;
wire n_13521;
wire n_13522;
wire n_13523;
wire n_13524;
wire n_13525;
wire n_13526;
wire n_13527;
wire n_13528;
wire n_13529;
wire n_1353;
wire n_13530;
wire n_13531;
wire n_13532;
wire n_13533;
wire n_13534;
wire n_13535;
wire n_13536;
wire n_13537;
wire n_13538;
wire n_13539;
wire n_1354;
wire n_13540;
wire n_13541;
wire n_13543;
wire n_13544;
wire n_13546;
wire n_13547;
wire n_13548;
wire n_1355;
wire n_13550;
wire n_13552;
wire n_13553;
wire n_13554;
wire n_13555;
wire n_13556;
wire n_13557;
wire n_13558;
wire n_13559;
wire n_1356;
wire n_13560;
wire n_13561;
wire n_13562;
wire n_13563;
wire n_13564;
wire n_13565;
wire n_13566;
wire n_13568;
wire n_13569;
wire n_1357;
wire TIMEBOOST_net_15135;
wire n_13571;
wire n_13573;
wire n_13574;
wire n_13575;
wire n_13576;
wire n_13577;
wire n_13578;
wire n_13579;
wire n_1358;
wire n_13581;
wire n_13582;
wire n_13585;
wire n_13587;
wire n_1359;
wire n_13591;
wire n_13592;
wire TIMEBOOST_net_15123;
wire n_13595;
wire n_13597;
wire n_13599;
wire n_13601;
wire n_13603;
wire n_13605;
wire n_13607;
wire n_13608;
wire n_13609;
wire n_1361;
wire n_13611;
wire n_13613;
wire n_13614;
wire n_13616;
wire n_13617;
wire n_13618;
wire n_13619;
wire n_1362;
wire n_13620;
wire n_13621;
wire n_13622;
wire n_13623;
wire n_13624;
wire n_13625;
wire n_13627;
wire n_13628;
wire n_13629;
wire n_1363;
wire n_13631;
wire n_13632;
wire n_13634;
wire n_13635;
wire n_13636;
wire n_13638;
wire n_13640;
wire n_13641;
wire n_13642;
wire n_13643;
wire n_13645;
wire n_13646;
wire n_13647;
wire n_13648;
wire n_13649;
wire n_1365;
wire n_13650;
wire n_13651;
wire TIMEBOOST_net_10861;
wire n_13653;
wire n_13654;
wire TIMEBOOST_net_14933;
wire n_13657;
wire n_13658;
wire n_13659;
wire n_1366;
wire n_13661;
wire n_13662;
wire n_13663;
wire n_13664;
wire n_13666;
wire n_13667;
wire n_13668;
wire n_13670;
wire n_13671;
wire n_13672;
wire n_13673;
wire n_13674;
wire n_13678;
wire n_13679;
wire n_13680;
wire n_13681;
wire n_13682;
wire n_13685;
wire n_13686;
wire n_13687;
wire n_13688;
wire n_13689;
wire n_1369;
wire n_13691;
wire n_13692;
wire n_13693;
wire n_13694;
wire n_13695;
wire n_13696;
wire n_13697;
wire n_13698;
wire n_13701;
wire n_13703;
wire n_13704;
wire n_13705;
wire n_13709;
wire n_1371;
wire n_13710;
wire n_13711;
wire n_13712;
wire n_13715;
wire n_13716;
wire n_13717;
wire n_13719;
wire n_1372;
wire n_13720;
wire n_13721;
wire n_13722;
wire n_13724;
wire n_13725;
wire n_13727;
wire n_13728;
wire n_13729;
wire n_1373;
wire n_13731;
wire n_13732;
wire n_13734;
wire n_13735;
wire n_13736;
wire n_13738;
wire n_1374;
wire n_13740;
wire n_13741;
wire n_13743;
wire n_13744;
wire n_13745;
wire n_13747;
wire n_13748;
wire n_13749;
wire n_13750;
wire n_13752;
wire n_13753;
wire n_13754;
wire n_13755;
wire n_13756;
wire n_13757;
wire n_13758;
wire n_13759;
wire n_13760;
wire n_13761;
wire TIMEBOOST_net_12893;
wire n_13763;
wire n_13764;
wire n_13765;
wire n_13766;
wire n_13767;
wire n_13768;
wire n_1377;
wire n_13770;
wire n_13771;
wire n_13772;
wire TIMEBOOST_net_12849;
wire n_13774;
wire n_13775;
wire n_13776;
wire TIMEBOOST_net_12846;
wire TIMEBOOST_net_13137;
wire n_1378;
wire n_13780;
wire n_13781;
wire n_13783;
wire n_13784;
wire n_13785;
wire TIMEBOOST_net_1440;
wire n_13787;
wire n_13789;
wire n_1379;
wire n_13790;
wire n_13792;
wire n_13793;
wire n_13794;
wire n_13798;
wire n_13806;
wire n_13807;
wire n_13809;
wire n_1381;
wire n_13810;
wire n_13812;
wire n_13813;
wire n_13814;
wire n_13815;
wire n_13816;
wire n_13817;
wire n_13819;
wire n_1382;
wire n_13820;
wire n_13821;
wire n_13822;
wire n_13823;
wire n_13824;
wire n_13825;
wire n_13826;
wire n_13827;
wire n_13828;
wire n_13829;
wire n_1383;
wire n_13830;
wire n_13831;
wire n_1384;
wire n_13842;
wire n_13843;
wire n_13844;
wire TIMEBOOST_net_13496;
wire n_13846;
wire n_13847;
wire n_13849;
wire n_1385;
wire n_10139;
wire n_13854;
wire n_13856;
wire n_13857;
wire n_13859;
wire n_13862;
wire n_13863;
wire n_13865;
wire TIMEBOOST_net_6289;
wire n_13868;
wire TIMEBOOST_net_15252;
wire n_1387;
wire n_13871;
wire n_13873;
wire n_10275;
wire n_13875;
wire n_13878;
wire TIMEBOOST_net_12806;
wire n_1388;
wire n_10237;
wire n_10199;
wire n_10263;
wire TIMEBOOST_net_12805;
wire TIMEBOOST_net_12757;
wire n_13888;
wire n_10279;
wire n_1389;
wire n_13891;
wire n_10274;
wire n_14060;
wire TIMEBOOST_net_15224;
wire n_13899;
wire n_139;
wire n_1390;
wire n_13901;
wire n_13903;
wire TIMEBOOST_net_15227;
wire TIMEBOOST_net_12804;
wire n_13906;
wire n_13907;
wire n_13908;
wire n_1391;
wire n_13910;
wire n_13911;
wire n_13917;
wire n_13918;
wire n_13919;
wire n_1392;
wire n_13920;
wire n_13921;
wire n_13922;
wire n_13923;
wire n_13926;
wire TIMEBOOST_net_3737;
wire TIMEBOOST_net_12774;
wire n_1393;
wire n_13930;
wire TIMEBOOST_net_12603;
wire n_10278;
wire TIMEBOOST_net_15206;
wire TIMEBOOST_net_9463;
wire TIMEBOOST_net_3735;
wire n_13936;
wire n_13937;
wire n_13938;
wire TIMEBOOST_net_9462;
wire n_1394;
wire TIMEBOOST_net_12686;
wire TIMEBOOST_net_13000;
wire n_13942;
wire n_13943;
wire TIMEBOOST_net_12685;
wire TIMEBOOST_net_12723;
wire TIMEBOOST_net_12502;
wire n_13949;
wire n_1395;
wire TIMEBOOST_net_9461;
wire TIMEBOOST_net_12521;
wire n_13953;
wire n_13954;
wire TIMEBOOST_net_9460;
wire TIMEBOOST_net_9459;
wire n_13958;
wire n_1396;
wire n_13960;
wire n_10247;
wire TIMEBOOST_net_9458;
wire TIMEBOOST_net_9457;
wire TIMEBOOST_net_12522;
wire TIMEBOOST_net_12620;
wire n_1397;
wire n_10277;
wire n_13971;
wire n_13972;
wire n_13973;
wire n_13974;
wire TIMEBOOST_net_9456;
wire TIMEBOOST_net_12629;
wire TIMEBOOST_net_12764;
wire TIMEBOOST_net_12798;
wire n_1398;
wire n_13980;
wire TIMEBOOST_net_12169;
wire n_13982;
wire TIMEBOOST_net_12664;
wire TIMEBOOST_net_9416;
wire TIMEBOOST_net_12628;
wire n_13987;
wire n_10190;
wire n_1399;
wire n_13990;
wire n_13991;
wire n_13992;
wire n_13993;
wire n_13994;
wire n_13995;
wire n_13997;
wire n_13999;
wire n_14;
wire n_1400;
wire n_14000;
wire TIMEBOOST_net_9454;
wire n_14002;
wire n_14004;
wire n_14005;
wire n_14007;
wire TIMEBOOST_net_9410;
wire n_1401;
wire n_14011;
wire n_14013;
wire TIMEBOOST_net_9453;
wire n_14016;
wire TIMEBOOST_net_9406;
wire n_14018;
wire n_14019;
wire n_1402;
wire n_14020;
wire TIMEBOOST_net_9405;
wire n_14022;
wire TIMEBOOST_net_12682;
wire n_14024;
wire n_14025;
wire TIMEBOOST_net_9403;
wire n_14027;
wire n_14029;
wire n_1403;
wire TIMEBOOST_net_9400;
wire n_14033;
wire TIMEBOOST_net_15209;
wire n_14035;
wire TIMEBOOST_net_9396;
wire TIMEBOOST_net_9393;
wire n_1404;
wire TIMEBOOST_net_9392;
wire TIMEBOOST_net_15211;
wire TIMEBOOST_net_9407;
wire TIMEBOOST_net_12708;
wire TIMEBOOST_net_15257;
wire TIMEBOOST_net_12168;
wire TIMEBOOST_net_12946;
wire n_14049;
wire n_1405;
wire TIMEBOOST_net_12692;
wire n_14054;
wire n_14055;
wire n_14056;
wire n_1406;
wire TIMEBOOST_net_12167;
wire n_14061;
wire TIMEBOOST_net_12627;
wire TIMEBOOST_net_15256;
wire n_14069;
wire n_1407;
wire n_14070;
wire n_14072;
wire n_14073;
wire n_14074;
wire n_14075;
wire n_14076;
wire n_14077;
wire n_14078;
wire n_14079;
wire n_1408;
wire n_14080;
wire n_14081;
wire n_14082;
wire n_14083;
wire n_14084;
wire n_14085;
wire n_14086;
wire TIMEBOOST_net_11444;
wire n_14088;
wire n_1409;
wire n_14093;
wire n_14094;
wire TIMEBOOST_net_12799;
wire TIMEBOOST_net_9431;
wire n_14099;
wire n_1410;
wire n_14104;
wire TIMEBOOST_net_12616;
wire TIMEBOOST_net_12684;
wire TIMEBOOST_net_9429;
wire TIMEBOOST_net_12724;
wire n_1411;
wire n_14111;
wire TIMEBOOST_net_12725;
wire TIMEBOOST_net_12726;
wire TIMEBOOST_net_12660;
wire TIMEBOOST_net_12687;
wire TIMEBOOST_net_9425;
wire TIMEBOOST_net_12659;
wire n_1412;
wire TIMEBOOST_net_9424;
wire TIMEBOOST_net_9423;
wire TIMEBOOST_net_12735;
wire TIMEBOOST_net_12693;
wire TIMEBOOST_net_12739;
wire TIMEBOOST_net_12196;
wire n_14128;
wire n_1413;
wire TIMEBOOST_net_9420;
wire TIMEBOOST_net_9419;
wire TIMEBOOST_net_9418;
wire TIMEBOOST_net_9417;
wire n_1414;
wire n_14140;
wire n_14142;
wire n_14144;
wire n_1415;
wire TIMEBOOST_net_9414;
wire TIMEBOOST_net_9413;
wire TIMEBOOST_net_9412;
wire TIMEBOOST_net_9411;
wire n_1416;
wire TIMEBOOST_net_9409;
wire TIMEBOOST_net_6294;
wire TIMEBOOST_net_9378;
wire n_14166;
wire n_14167;
wire TIMEBOOST_net_12813;
wire n_1417;
wire n_14170;
wire n_14171;
wire n_14172;
wire n_14174;
wire TIMEBOOST_net_9391;
wire n_14177;
wire n_14178;
wire n_10250;
wire n_1418;
wire TIMEBOOST_net_9404;
wire n_10225;
wire TIMEBOOST_net_9402;
wire n_14185;
wire n_14186;
wire n_10213;
wire TIMEBOOST_net_9401;
wire n_1419;
wire TIMEBOOST_net_12638;
wire TIMEBOOST_net_12637;
wire TIMEBOOST_net_9390;
wire n_14194;
wire n_14195;
wire n_14197;
wire TIMEBOOST_net_9395;
wire TIMEBOOST_net_79;
wire TIMEBOOST_net_9394;
wire n_14201;
wire n_14202;
wire n_14203;
wire n_14205;
wire n_14207;
wire n_1421;
wire n_14211;
wire n_14212;
wire TIMEBOOST_net_12812;
wire TIMEBOOST_net_12811;
wire n_1422;
wire n_14220;
wire TIMEBOOST_net_9377;
wire n_14223;
wire n_14225;
wire n_14226;
wire TIMEBOOST_net_12810;
wire n_1423;
wire TIMEBOOST_net_12809;
wire TIMEBOOST_net_3648;
wire n_1424;
wire TIMEBOOST_net_12762;
wire n_14243;
wire n_14245;
wire TIMEBOOST_net_12808;
wire TIMEBOOST_net_9389;
wire n_1425;
wire n_14250;
wire n_14251;
wire n_14252;
wire n_14253;
wire n_14254;
wire n_14255;
wire n_14256;
wire n_14257;
wire n_14258;
wire n_1426;
wire n_14260;
wire n_14261;
wire n_14264;
wire n_14268;
wire n_14269;
wire n_14270;
wire n_14271;
wire n_14272;
wire n_14273;
wire n_14274;
wire n_14275;
wire n_14277;
wire n_1428;
wire n_14283;
wire n_14284;
wire n_14285;
wire n_14286;
wire n_1429;
wire n_14290;
wire n_14291;
wire n_14292;
wire n_14293;
wire n_14295;
wire n_14296;
wire n_14298;
wire n_143;
wire n_14300;
wire n_14301;
wire n_14302;
wire n_14303;
wire n_14304;
wire n_14305;
wire n_14306;
wire n_14307;
wire n_14308;
wire n_14309;
wire n_1431;
wire n_14310;
wire n_14311;
wire n_14312;
wire n_14313;
wire n_14314;
wire n_14315;
wire n_14316;
wire n_14317;
wire n_14318;
wire n_14319;
wire n_1432;
wire n_14320;
wire n_14321;
wire n_14322;
wire n_14323;
wire n_14324;
wire n_14325;
wire n_14326;
wire n_14327;
wire n_14328;
wire n_14329;
wire n_1433;
wire n_14330;
wire n_14331;
wire n_14332;
wire n_14333;
wire n_14334;
wire n_14335;
wire n_14336;
wire n_14337;
wire n_14338;
wire n_14339;
wire n_1434;
wire n_14340;
wire n_14341;
wire n_14342;
wire n_14343;
wire n_14344;
wire n_14345;
wire n_14346;
wire n_14347;
wire n_14348;
wire n_14349;
wire n_1435;
wire n_14350;
wire n_14351;
wire n_14352;
wire n_14353;
wire n_14354;
wire n_14355;
wire n_14356;
wire n_14357;
wire n_14358;
wire n_14359;
wire n_1436;
wire n_14360;
wire n_14361;
wire n_14362;
wire n_14363;
wire n_14364;
wire n_14365;
wire n_14366;
wire n_14367;
wire n_14368;
wire n_14369;
wire n_1437;
wire n_14370;
wire n_14371;
wire n_14372;
wire n_14373;
wire n_14374;
wire n_14375;
wire n_14376;
wire n_14377;
wire n_14378;
wire n_14379;
wire n_1438;
wire n_14380;
wire n_14381;
wire n_14382;
wire n_14383;
wire n_14384;
wire n_14385;
wire n_14386;
wire n_14387;
wire n_14388;
wire n_14389;
wire n_1439;
wire n_14390;
wire n_14391;
wire n_14392;
wire n_14393;
wire n_14394;
wire n_14396;
wire n_14397;
wire n_14399;
wire n_1440;
wire n_14401;
wire n_14402;
wire n_14403;
wire n_14407;
wire n_14408;
wire n_1441;
wire n_14410;
wire n_14413;
wire n_14414;
wire n_14415;
wire n_14416;
wire n_14419;
wire n_1442;
wire n_14420;
wire n_14421;
wire n_14422;
wire n_14426;
wire n_14427;
wire n_14428;
wire n_14429;
wire n_1443;
wire n_14430;
wire n_14431;
wire n_14432;
wire n_14433;
wire n_14434;
wire n_14435;
wire n_14436;
wire n_14437;
wire n_14438;
wire n_14439;
wire n_1444;
wire n_14440;
wire n_14441;
wire n_14442;
wire n_14443;
wire n_14444;
wire n_14445;
wire n_14446;
wire n_14447;
wire n_14448;
wire n_14449;
wire n_1445;
wire n_14451;
wire n_14454;
wire n_14456;
wire n_14457;
wire n_14458;
wire n_14459;
wire n_1446;
wire n_14460;
wire n_14461;
wire n_14462;
wire n_14467;
wire n_14468;
wire n_14469;
wire n_1447;
wire n_14471;
wire n_14472;
wire n_14473;
wire n_14474;
wire n_14475;
wire n_14476;
wire n_14477;
wire n_14478;
wire n_14479;
wire n_1448;
wire n_14480;
wire n_14481;
wire n_14482;
wire n_14483;
wire n_14484;
wire n_14485;
wire n_14486;
wire n_14487;
wire n_14489;
wire n_1449;
wire n_14490;
wire n_14491;
wire n_14493;
wire n_14494;
wire n_14495;
wire n_14497;
wire n_14498;
wire n_14499;
wire n_1450;
wire n_14500;
wire n_14504;
wire n_14505;
wire n_14507;
wire n_14508;
wire n_14510;
wire n_14511;
wire n_14512;
wire n_14513;
wire n_14514;
wire n_14515;
wire n_14517;
wire n_14518;
wire TIMEBOOST_net_13898;
wire n_1452;
wire n_14521;
wire n_14526;
wire TIMEBOOST_net_11839;
wire n_14528;
wire n_14529;
wire n_1453;
wire n_14530;
wire n_14531;
wire n_14532;
wire n_14534;
wire n_14535;
wire n_14536;
wire n_14539;
wire n_1454;
wire n_14541;
wire n_14543;
wire n_14544;
wire n_14545;
wire n_14547;
wire n_14548;
wire n_14549;
wire n_14550;
wire n_14551;
wire n_14554;
wire n_14556;
wire n_14557;
wire n_14558;
wire n_14559;
wire n_14560;
wire n_14563;
wire n_14564;
wire n_14565;
wire n_14566;
wire n_14567;
wire n_14569;
wire n_14570;
wire n_14571;
wire n_14572;
wire n_2153;
wire n_14577;
wire n_14578;
wire n_14579;
wire n_14580;
wire n_14582;
wire n_14583;
wire n_14585;
wire n_14586;
wire n_14588;
wire n_14589;
wire n_1459;
wire n_14590;
wire n_14591;
wire n_14592;
wire n_14593;
wire n_14594;
wire n_14595;
wire n_14596;
wire n_14597;
wire n_14598;
wire n_14599;
wire n_1460;
wire n_14601;
wire n_14602;
wire n_14603;
wire n_14604;
wire n_14605;
wire n_14607;
wire n_14608;
wire n_14609;
wire n_1461;
wire n_14610;
wire n_14611;
wire n_14612;
wire n_14613;
wire n_14614;
wire n_14615;
wire n_14616;
wire n_14617;
wire n_14618;
wire n_14619;
wire n_14620;
wire n_14621;
wire n_14622;
wire n_14623;
wire n_14624;
wire n_14625;
wire n_14626;
wire n_14627;
wire n_14628;
wire n_14629;
wire n_1463;
wire n_14630;
wire n_14631;
wire n_14632;
wire n_14633;
wire n_14634;
wire n_14635;
wire n_14636;
wire n_14637;
wire n_14638;
wire n_14639;
wire n_14640;
wire n_14641;
wire n_14642;
wire n_14643;
wire n_14644;
wire n_14645;
wire n_14646;
wire n_14648;
wire n_14649;
wire n_1465;
wire n_14650;
wire n_14651;
wire n_14652;
wire n_14653;
wire n_14654;
wire n_14655;
wire n_14656;
wire n_14657;
wire n_14658;
wire n_14659;
wire TIMEBOOST_net_907;
wire TIMEBOOST_net_13650;
wire n_14662;
wire n_14663;
wire n_14664;
wire n_14665;
wire n_14666;
wire n_14667;
wire n_14668;
wire n_14669;
wire n_1467;
wire n_14670;
wire n_14671;
wire TIMEBOOST_net_12827;
wire TIMEBOOST_net_12588;
wire n_14674;
wire TIMEBOOST_net_1225;
wire n_14676;
wire n_14678;
wire n_14679;
wire n_1468;
wire n_14680;
wire n_14681;
wire TIMEBOOST_net_710;
wire n_14683;
wire n_14685;
wire n_14686;
wire n_14687;
wire n_14688;
wire n_14689;
wire n_1469;
wire n_14690;
wire n_14691;
wire n_14693;
wire n_14694;
wire n_14695;
wire n_14696;
wire n_14697;
wire n_14698;
wire n_14699;
wire n_1470;
wire n_14700;
wire n_14701;
wire n_14702;
wire n_14703;
wire n_14705;
wire n_14706;
wire n_14708;
wire n_14709;
wire n_1471;
wire n_14710;
wire n_14711;
wire n_14713;
wire n_14715;
wire n_14717;
wire n_14719;
wire n_1472;
wire n_14721;
wire n_14722;
wire n_14723;
wire n_14724;
wire n_14725;
wire n_14726;
wire n_14727;
wire n_14728;
wire n_14730;
wire n_14731;
wire n_14733;
wire n_14734;
wire TIMEBOOST_net_14154;
wire n_14738;
wire n_1474;
wire n_14740;
wire n_14741;
wire n_14743;
wire n_14744;
wire n_14746;
wire TIMEBOOST_net_1448;
wire TIMEBOOST_net_14135;
wire n_14749;
wire n_1475;
wire TIMEBOOST_net_10331;
wire n_14751;
wire n_14753;
wire TIMEBOOST_net_4563;
wire n_14755;
wire n_14756;
wire n_14757;
wire n_14759;
wire n_1476;
wire n_14760;
wire n_14761;
wire n_14762;
wire n_14763;
wire n_14764;
wire n_14765;
wire n_14766;
wire n_14767;
wire n_14768;
wire n_14769;
wire n_1477;
wire n_14770;
wire n_14772;
wire n_14773;
wire n_14775;
wire n_14776;
wire n_14777;
wire n_14778;
wire n_1478;
wire n_14780;
wire n_14781;
wire n_14783;
wire n_14784;
wire n_14786;
wire n_14789;
wire n_1479;
wire n_14790;
wire n_14791;
wire n_14792;
wire n_14793;
wire n_14794;
wire n_14796;
wire n_14797;
wire n_14798;
wire n_14799;
wire n_148;
wire n_1480;
wire n_14800;
wire n_14802;
wire n_14803;
wire n_14804;
wire n_14805;
wire n_14806;
wire n_14807;
wire n_14808;
wire n_1481;
wire n_14810;
wire n_14811;
wire n_14812;
wire n_14813;
wire n_14814;
wire n_14815;
wire n_14816;
wire n_14817;
wire n_14818;
wire n_14819;
wire n_1482;
wire n_14821;
wire n_14822;
wire n_14824;
wire n_14825;
wire n_14826;
wire n_14828;
wire n_14829;
wire n_1483;
wire n_14830;
wire n_14832;
wire n_14833;
wire n_14834;
wire n_14836;
wire n_14837;
wire n_14838;
wire n_14839;
wire n_1484;
wire n_14840;
wire n_14841;
wire n_14842;
wire n_14844;
wire n_14845;
wire n_14846;
wire n_14847;
wire n_14848;
wire n_14849;
wire n_1485;
wire n_14850;
wire n_14851;
wire n_14852;
wire n_14853;
wire n_14854;
wire n_14855;
wire n_14856;
wire n_14858;
wire n_14859;
wire n_1486;
wire n_14860;
wire n_14861;
wire n_14862;
wire n_14863;
wire n_14864;
wire n_14865;
wire n_14866;
wire n_14867;
wire n_14869;
wire n_14871;
wire n_14873;
wire n_14875;
wire n_14877;
wire n_14879;
wire n_1488;
wire n_14880;
wire n_14881;
wire n_14883;
wire n_14884;
wire n_14885;
wire n_14887;
wire n_14888;
wire n_14889;
wire n_14890;
wire n_14891;
wire n_14892;
wire n_14893;
wire n_14894;
wire n_14895;
wire n_14896;
wire n_14897;
wire n_14898;
wire n_14899;
wire n_14900;
wire n_14901;
wire n_14902;
wire n_14903;
wire n_14904;
wire n_14905;
wire n_14906;
wire n_14907;
wire n_14908;
wire n_14909;
wire n_14910;
wire n_14911;
wire n_14912;
wire n_14913;
wire n_14914;
wire n_14915;
wire n_14916;
wire n_14917;
wire n_14918;
wire n_14919;
wire n_14920;
wire n_14921;
wire n_14922;
wire n_14923;
wire n_14924;
wire n_14925;
wire n_14926;
wire n_14927;
wire n_14928;
wire n_14929;
wire n_1493;
wire n_14930;
wire n_14931;
wire n_14932;
wire n_14933;
wire n_14934;
wire n_14939;
wire n_1495;
wire n_14956;
wire n_14957;
wire n_14960;
wire n_14961;
wire n_14963;
wire n_14965;
wire n_14967;
wire n_1497;
wire n_14971;
wire n_14981;
wire n_1499;
wire n_15;
wire n_150;
wire n_15001;
wire n_1501;
wire n_15014;
wire n_1502;
wire n_1503;
wire TIMEBOOST_net_175;
wire n_1504;
wire n_1505;
wire n_15054;
wire n_15055;
wire n_15065;
wire n_1507;
wire n_1508;
wire n_1509;
wire n_1510;
wire n_15117;
wire n_1512;
wire n_15125;
wire n_15128;
wire n_1513;
wire n_1514;
wire n_15142;
wire n_1515;
wire n_15187;
wire n_15188;
wire n_1519;
wire n_15196;
wire n_15197;
wire n_152;
wire n_15204;
wire n_15210;
wire n_15217;
wire n_1522;
wire n_1523;
wire n_15231;
wire n_1524;
wire n_15249;
wire n_15260;
wire n_15261;
wire n_15262;
wire n_15275;
wire n_15276;
wire n_15291;
wire n_15292;
wire n_15295;
wire n_15301;
wire n_15302;
wire n_15313;
wire n_15314;
wire TIMEBOOST_net_12080;
wire n_15317;
wire n_1532;
wire n_15324;
wire n_15325;
wire n_1533;
wire n_15330;
wire n_15331;
wire n_15347;
wire n_1535;
wire n_1536;
wire n_15365;
wire n_1537;
wire n_15370;
wire n_15371;
wire n_15372;
wire n_15373;
wire n_15376;
wire n_15377;
wire n_1538;
wire n_15385;
wire n_15388;
wire n_15389;
wire n_1539;
wire n_15390;
wire n_15397;
wire n_1540;
wire n_15401;
wire n_15402;
wire n_15403;
wire n_15405;
wire n_15406;
wire n_15407;
wire n_1541;
wire n_15414;
wire n_15417;
wire n_1542;
wire TIMEBOOST_net_82;
wire n_15434;
wire n_15435;
wire n_15436;
wire n_15438;
wire n_15439;
wire n_15440;
wire n_15441;
wire n_15442;
wire n_15444;
wire n_15445;
wire n_15446;
wire n_1545;
wire n_15453;
wire n_15456;
wire TIMEBOOST_net_11026;
wire n_15458;
wire n_1546;
wire n_15467;
wire n_1547;
wire n_15474;
wire n_1548;
wire n_1549;
wire n_1551;
wire n_15512;
wire n_15513;
wire n_15514;
wire n_15515;
wire n_15516;
wire n_15517;
wire n_15518;
wire TIMEBOOST_net_12713;
wire n_15527;
wire n_15528;
wire n_15529;
wire n_1553;
wire n_15533;
wire n_15534;
wire n_15537;
wire n_15538;
wire n_15539;
wire n_1554;
wire n_15540;
wire n_15549;
wire n_1555;
wire n_15551;
wire n_15552;
wire n_15553;
wire n_15558;
wire n_15560;
wire n_15562;
wire n_15565;
wire n_15566;
wire n_15567;
wire n_15568;
wire n_15569;
wire n_1557;
wire TIMEBOOST_net_14068;
wire TIMEBOOST_net_2878;
wire n_15581;
wire n_15584;
wire n_15585;
wire n_15586;
wire n_15587;
wire n_15589;
wire n_1559;
wire n_15590;
wire n_15591;
wire n_15592;
wire n_15593;
wire n_15594;
wire n_15598;
wire n_156;
wire n_15607;
wire n_1561;
wire n_15611;
wire n_15614;
wire n_1562;
wire TIMEBOOST_net_12982;
wire n_15638;
wire n_1564;
wire n_15645;
wire n_1565;
wire n_1567;
wire TIMEBOOST_net_13466;
wire n_15680;
wire n_15689;
wire n_1569;
wire n_15694;
wire n_15695;
wire TIMEBOOST_net_12939;
wire TIMEBOOST_net_10138;
wire n_15698;
wire n_15699;
wire TIMEBOOST_net_179;
wire n_1571;
wire n_1572;
wire TIMEBOOST_net_10139;
wire n_15729;
wire n_1573;
wire TIMEBOOST_net_13928;
wire n_15732;
wire n_15733;
wire n_15735;
wire n_15736;
wire TIMEBOOST_net_12598;
wire n_15738;
wire n_15739;
wire n_1574;
wire n_15741;
wire n_15744;
wire n_15746;
wire n_15748;
wire n_1575;
wire n_15754;
wire n_15755;
wire n_15756;
wire n_15757;
wire n_15758;
wire n_15759;
wire n_1576;
wire n_15760;
wire n_15762;
wire n_15769;
wire n_1577;
wire TIMEBOOST_net_3076;
wire n_1578;
wire n_15788;
wire n_1579;
wire n_15798;
wire n_1580;
wire n_15802;
wire n_15805;
wire n_15808;
wire n_1581;
wire n_15813;
wire n_15823;
wire n_15824;
wire n_1583;
wire n_1584;
wire n_1585;
wire n_15854;
wire n_15856;
wire n_15859;
wire n_1586;
wire n_1587;
wire n_1588;
wire n_1589;
wire n_1590;
wire n_15908;
wire TIMEBOOST_net_274;
wire n_1591;
wire n_15910;
wire n_15914;
wire n_15915;
wire n_15917;
wire n_15918;
wire n_15919;
wire n_1592;
wire n_15920;
wire TIMEBOOST_net_9637;
wire n_15922;
wire n_15923;
wire n_15924;
wire n_15927;
wire n_15928;
wire n_15929;
wire n_1593;
wire n_15931;
wire n_15932;
wire n_15935;
wire n_15936;
wire n_15937;
wire n_15939;
wire n_1594;
wire n_15940;
wire n_15941;
wire n_15942;
wire n_1595;
wire n_15958;
wire n_15959;
wire n_1596;
wire n_15960;
wire n_15969;
wire n_1597;
wire n_15979;
wire TIMEBOOST_net_15188;
wire n_15980;
wire n_15981;
wire n_15982;
wire n_15985;
wire n_15988;
wire n_1599;
wire n_15994;
wire n_15996;
wire n_15998;
wire n_15999;
wire n_160;
wire n_1600;
wire n_16000;
wire n_16001;
wire n_16002;
wire n_16003;
wire n_1601;
wire n_16015;
wire n_16016;
wire n_1602;
wire n_16021;
wire n_16022;
wire n_16027;
wire n_1603;
wire n_16030;
wire n_16033;
wire n_16034;
wire n_16036;
wire n_1604;
wire n_16046;
wire n_16047;
wire n_16048;
wire n_16049;
wire n_1605;
wire n_16052;
wire n_1606;
wire n_16066;
wire TIMEBOOST_net_12372;
wire n_1607;
wire n_16070;
wire n_16071;
wire n_16075;
wire n_16076;
wire n_1608;
wire n_16089;
wire n_1609;
wire n_1610;
wire n_16101;
wire n_16102;
wire n_16103;
wire n_16105;
wire n_1611;
wire n_1612;
wire n_1613;
wire n_16131;
wire n_1614;
wire TIMEBOOST_net_902;
wire n_1615;
wire n_16150;
wire n_16151;
wire n_16152;
wire n_16153;
wire n_16154;
wire n_16156;
wire n_16157;
wire TIMEBOOST_net_2032;
wire n_16159;
wire n_1616;
wire n_16160;
wire n_16161;
wire n_16162;
wire n_16163;
wire n_16164;
wire n_16165;
wire TIMEBOOST_net_12595;
wire n_16167;
wire n_16168;
wire n_16169;
wire TIMEBOOST_net_3009;
wire n_16170;
wire n_16173;
wire n_16175;
wire TIMEBOOST_net_14883;
wire n_16183;
wire n_1619;
wire n_16205;
wire n_16206;
wire n_16207;
wire n_16208;
wire n_16209;
wire n_1621;
wire n_16210;
wire n_16211;
wire n_16212;
wire n_16213;
wire n_16220;
wire n_16221;
wire n_16222;
wire n_16223;
wire n_16224;
wire n_16225;
wire n_16226;
wire n_16227;
wire n_16228;
wire n_16229;
wire n_1623;
wire n_16230;
wire n_16231;
wire n_16233;
wire n_16234;
wire n_16235;
wire n_16236;
wire n_16237;
wire n_16238;
wire n_16239;
wire n_1624;
wire n_16240;
wire n_16241;
wire n_16242;
wire n_16243;
wire n_16244;
wire n_16247;
wire n_16248;
wire n_16249;
wire n_1625;
wire n_16250;
wire n_16251;
wire n_16252;
wire n_16253;
wire n_16254;
wire n_16255;
wire n_16256;
wire n_16257;
wire n_16258;
wire n_16259;
wire n_1626;
wire n_16260;
wire n_16261;
wire n_16262;
wire n_16264;
wire n_16265;
wire n_16268;
wire n_16271;
wire n_16273;
wire n_16275;
wire n_1628;
wire n_16280;
wire n_16284;
wire n_16285;
wire n_16286;
wire n_16287;
wire n_16288;
wire n_16289;
wire n_1629;
wire n_16290;
wire n_16291;
wire n_16293;
wire n_16299;
wire n_1630;
wire n_16300;
wire n_16301;
wire n_16304;
wire n_16305;
wire n_16306;
wire n_16307;
wire n_16309;
wire n_1631;
wire n_16310;
wire n_16311;
wire n_16313;
wire n_16317;
wire n_1632;
wire n_16322;
wire n_16325;
wire n_16326;
wire n_1633;
wire n_16330;
wire n_16331;
wire n_16332;
wire n_16334;
wire n_16338;
wire n_1634;
wire n_1635;
wire n_16350;
wire n_16351;
wire n_16352;
wire n_16354;
wire n_16358;
wire n_16364;
wire n_16368;
wire n_16388;
wire n_16389;
wire n_1639;
wire n_16390;
wire n_16391;
wire TIMEBOOST_net_14950;
wire n_16393;
wire TIMEBOOST_net_12782;
wire n_16395;
wire n_16396;
wire n_16397;
wire n_16398;
wire n_16399;
wire n_1640;
wire n_16400;
wire n_16401;
wire n_16402;
wire n_16403;
wire n_16404;
wire n_16406;
wire n_16408;
wire n_16409;
wire n_1641;
wire n_16410;
wire n_16411;
wire n_16412;
wire n_16413;
wire n_1642;
wire n_16424;
wire n_16425;
wire n_16427;
wire n_16428;
wire n_16429;
wire TIMEBOOST_net_12081;
wire TIMEBOOST_net_12853;
wire n_16433;
wire n_16434;
wire n_16435;
wire n_16436;
wire n_16437;
wire n_16438;
wire n_16439;
wire TIMEBOOST_net_13223;
wire n_16441;
wire n_16442;
wire n_16444;
wire n_16445;
wire n_1645;
wire n_16451;
wire n_16452;
wire n_16455;
wire n_16456;
wire TIMEBOOST_net_12670;
wire TIMEBOOST_net_10947;
wire n_16459;
wire n_1646;
wire n_16460;
wire n_16462;
wire n_1647;
wire n_16474;
wire n_16475;
wire n_1648;
wire n_16485;
wire n_16486;
wire n_16487;
wire n_1649;
wire n_16490;
wire n_16491;
wire n_16492;
wire n_16493;
wire n_16494;
wire n_16495;
wire n_16496;
wire n_16497;
wire n_16499;
wire n_1650;
wire n_16501;
wire n_16503;
wire n_16504;
wire n_16507;
wire n_16511;
wire n_16512;
wire n_16513;
wire n_16516;
wire n_1652;
wire n_16520;
wire n_16521;
wire n_16523;
wire n_16524;
wire n_1653;
wire n_16533;
wire n_16534;
wire n_16535;
wire n_16536;
wire n_16537;
wire n_16538;
wire n_16539;
wire n_1654;
wire n_16540;
wire n_16541;
wire n_16542;
wire n_16543;
wire n_16544;
wire n_16547;
wire n_1655;
wire n_16550;
wire n_16552;
wire n_16553;
wire n_16554;
wire n_1656;
wire n_16560;
wire n_16564;
wire TIMEBOOST_net_11732;
wire n_16566;
wire n_1657;
wire n_16572;
wire n_16573;
wire n_16576;
wire n_16577;
wire n_16578;
wire n_16579;
wire n_1658;
wire n_16581;
wire n_16582;
wire n_16583;
wire n_16584;
wire n_16585;
wire n_16586;
wire n_16587;
wire n_16588;
wire n_16589;
wire n_1659;
wire n_16591;
wire n_16592;
wire n_16594;
wire n_16595;
wire n_16596;
wire n_16597;
wire n_16599;
wire n_1660;
wire n_16600;
wire n_16601;
wire n_16602;
wire n_16603;
wire TIMEBOOST_net_11692;
wire n_16605;
wire TIMEBOOST_net_12761;
wire TIMEBOOST_net_12763;
wire n_16610;
wire n_16611;
wire n_16612;
wire n_16613;
wire n_16614;
wire n_16615;
wire n_16616;
wire n_16617;
wire n_10180;
wire n_1662;
wire n_16622;
wire n_16623;
wire n_16624;
wire n_16625;
wire TIMEBOOST_net_12639;
wire n_16629;
wire n_1663;
wire n_16631;
wire n_16635;
wire n_16637;
wire n_1664;
wire n_1665;
wire n_16657;
wire n_1666;
wire n_1667;
wire n_1668;
wire n_16685;
wire n_1669;
wire n_16690;
wire n_16695;
wire n_16696;
wire n_16698;
wire n_1673;
wire n_16738;
wire n_1674;
wire n_16748;
wire n_1675;
wire n_16763;
wire n_1677;
wire n_16779;
wire n_1678;
wire n_1679;
wire n_16791;
wire n_16798;
wire n_168;
wire n_1680;
wire n_1681;
wire n_16810;
wire n_16816;
wire n_16818;
wire n_1683;
wire n_16834;
wire n_16835;
wire n_16836;
wire n_16837;
wire n_16838;
wire n_16839;
wire n_1684;
wire n_16840;
wire n_16841;
wire n_16842;
wire n_16843;
wire n_16844;
wire n_16845;
wire n_16848;
wire n_16849;
wire n_1685;
wire n_16850;
wire n_16851;
wire n_16852;
wire n_16853;
wire n_16854;
wire n_16855;
wire n_1686;
wire n_16860;
wire n_16864;
wire n_16867;
wire n_16871;
wire n_16876;
wire n_1688;
wire n_16888;
wire n_1689;
wire n_16891;
wire n_169;
wire n_1690;
wire n_16904;
wire n_16906;
wire n_16910;
wire n_16911;
wire n_16914;
wire n_16916;
wire n_1692;
wire n_1693;
wire n_16936;
wire n_1694;
wire n_16940;
wire n_16942;
wire n_16945;
wire n_16949;
wire n_1695;
wire n_16952;
wire n_1696;
wire n_16963;
wire n_16964;
wire n_16966;
wire n_16967;
wire n_1697;
wire n_16970;
wire n_16974;
wire TIMEBOOST_net_13805;
wire n_16977;
wire n_1698;
wire n_16980;
wire n_16981;
wire n_16984;
wire n_16985;
wire n_16986;
wire n_16987;
wire n_1699;
wire n_16992;
wire n_17;
wire n_1700;
wire n_1701;
wire n_17016;
wire n_17017;
wire TIMEBOOST_net_12683;
wire TIMEBOOST_net_12719;
wire n_1702;
wire TIMEBOOST_net_13239;
wire TIMEBOOST_net_9432;
wire n_17027;
wire n_17028;
wire n_17029;
wire n_17030;
wire n_17031;
wire n_17032;
wire n_17034;
wire n_17035;
wire n_17036;
wire n_17039;
wire n_1704;
wire n_17040;
wire n_17041;
wire n_17042;
wire n_17043;
wire n_17044;
wire n_17045;
wire n_17046;
wire n_17048;
wire n_17049;
wire n_17050;
wire n_17051;
wire TIMEBOOST_net_13465;
wire n_1708;
wire n_1709;
wire n_1714;
wire n_1715;
wire n_1716;
wire n_1717;
wire n_1718;
wire n_1719;
wire n_1721;
wire n_1722;
wire n_1724;
wire n_1737;
wire n_1739;
wire n_1740;
wire n_1742;
wire n_1743;
wire n_1746;
wire n_1748;
wire n_1750;
wire n_1752;
wire n_1754;
wire n_1755;
wire n_1756;
wire n_1758;
wire n_1759;
wire n_177;
wire n_1774;
wire n_1777;
wire n_1779;
wire n_1780;
wire n_1781;
wire n_1782;
wire n_1784;
wire n_1785;
wire n_1786;
wire n_1787;
wire n_1788;
wire n_1789;
wire n_1790;
wire n_1793;
wire n_1794;
wire n_1795;
wire n_1798;
wire n_1799;
wire n_18;
wire n_1800;
wire n_1802;
wire n_1803;
wire n_1804;
wire n_1805;
wire n_1806;
wire n_1808;
wire n_1809;
wire n_181;
wire n_1810;
wire n_1812;
wire n_1813;
wire n_1814;
wire n_1815;
wire n_1816;
wire n_1817;
wire n_1819;
wire n_1820;
wire n_1821;
wire n_1822;
wire n_1823;
wire n_1824;
wire n_1825;
wire n_1826;
wire n_1827;
wire n_1828;
wire n_1829;
wire n_1832;
wire n_1834;
wire n_1836;
wire n_1837;
wire n_1838;
wire n_1844;
wire n_1845;
wire TIMEBOOST_net_465;
wire n_1847;
wire n_1848;
wire n_1849;
wire n_1850;
wire n_1851;
wire n_1852;
wire n_1853;
wire n_1854;
wire n_1855;
wire n_1856;
wire TIMEBOOST_net_10397;
wire n_1858;
wire n_1859;
wire n_1860;
wire n_1861;
wire n_1862;
wire n_1863;
wire n_1864;
wire n_1865;
wire n_1866;
wire n_1867;
wire n_1868;
wire n_1869;
wire TIMEBOOST_net_13400;
wire n_1871;
wire TIMEBOOST_net_10396;
wire n_1873;
wire TIMEBOOST_net_464;
wire n_1875;
wire TIMEBOOST_net_13399;
wire n_1877;
wire TIMEBOOST_net_10395;
wire n_1879;
wire n_188;
wire TIMEBOOST_net_10394;
wire n_1881;
wire TIMEBOOST_net_463;
wire n_1883;
wire TIMEBOOST_net_462;
wire TIMEBOOST_net_461;
wire TIMEBOOST_net_459;
wire TIMEBOOST_net_457;
wire n_1888;
wire n_1889;
wire TIMEBOOST_net_3171;
wire TIMEBOOST_net_10393;
wire TIMEBOOST_net_12325;
wire n_1893;
wire n_1894;
wire n_1895;
wire n_1896;
wire n_1897;
wire n_1898;
wire n_1899;
wire n_1900;
wire TIMEBOOST_net_10532;
wire n_1902;
wire n_1903;
wire n_1904;
wire n_1906;
wire n_1907;
wire n_1908;
wire n_1909;
wire n_191;
wire TIMEBOOST_net_272;
wire TIMEBOOST_net_271;
wire n_1913;
wire n_1914;
wire TIMEBOOST_net_270;
wire n_1916;
wire n_1917;
wire n_1918;
wire n_1919;
wire n_1920;
wire n_1921;
wire n_1922;
wire n_1923;
wire TIMEBOOST_net_268;
wire n_1925;
wire TIMEBOOST_net_267;
wire n_1927;
wire n_1928;
wire n_1929;
wire n_193;
wire n_1930;
wire n_1931;
wire n_1932;
wire n_1933;
wire n_1934;
wire TIMEBOOST_net_10328;
wire n_1936;
wire n_1937;
wire TIMEBOOST_net_266;
wire TIMEBOOST_net_265;
wire n_1940;
wire TIMEBOOST_net_10327;
wire n_1943;
wire TIMEBOOST_net_217;
wire n_1945;
wire n_1946;
wire n_1947;
wire n_1948;
wire TIMEBOOST_net_10324;
wire TIMEBOOST_net_13655;
wire TIMEBOOST_net_13471;
wire TIMEBOOST_net_10322;
wire TIMEBOOST_net_10053;
wire n_1954;
wire n_1955;
wire n_1956;
wire n_1957;
wire n_1958;
wire n_1959;
wire n_1960;
wire n_1961;
wire n_1963;
wire n_1964;
wire n_1965;
wire n_1966;
wire n_1967;
wire n_1968;
wire n_1969;
wire n_1970;
wire n_1971;
wire n_1972;
wire n_1973;
wire n_1974;
wire n_1975;
wire n_1976;
wire n_1978;
wire n_1979;
wire n_1981;
wire n_1985;
wire n_1986;
wire n_1987;
wire n_1989;
wire n_1990;
wire n_1992;
wire n_1993;
wire n_1994;
wire n_1995;
wire TIMEBOOST_net_269;
wire n_1998;
wire n_1999;
wire n_2;
wire n_200;
wire n_2000;
wire n_2001;
wire n_2002;
wire n_2004;
wire n_2005;
wire n_2006;
wire n_2007;
wire n_2008;
wire n_2009;
wire n_2010;
wire n_2011;
wire n_2012;
wire n_2013;
wire n_2014;
wire TIMEBOOST_net_458;
wire n_2016;
wire n_2017;
wire n_2018;
wire n_2019;
wire n_202;
wire n_2022;
wire n_2023;
wire n_2024;
wire n_2027;
wire n_2028;
wire n_2029;
wire n_2031;
wire n_2032;
wire n_2033;
wire n_2034;
wire n_2035;
wire n_2036;
wire n_2037;
wire TIMEBOOST_net_460;
wire n_2039;
wire n_204;
wire n_2040;
wire n_2041;
wire n_2042;
wire n_2043;
wire n_2044;
wire n_2045;
wire n_2046;
wire n_2047;
wire n_2048;
wire n_2049;
wire n_205;
wire n_2051;
wire n_2052;
wire n_2053;
wire n_2054;
wire n_2055;
wire n_2057;
wire n_2058;
wire n_2059;
wire n_206;
wire n_2060;
wire n_2061;
wire n_2065;
wire n_2066;
wire n_2067;
wire n_2068;
wire n_2069;
wire n_207;
wire n_2070;
wire n_2071;
wire n_2072;
wire n_2074;
wire n_2075;
wire n_2076;
wire n_2077;
wire n_2078;
wire n_2079;
wire n_208;
wire n_2080;
wire n_2082;
wire n_2083;
wire n_2084;
wire n_2086;
wire n_2087;
wire n_2088;
wire n_2092;
wire n_2093;
wire n_2094;
wire n_21;
wire n_2100;
wire n_2101;
wire n_2102;
wire n_2103;
wire n_2104;
wire n_2105;
wire n_2106;
wire n_2108;
wire n_211;
wire n_2110;
wire n_2111;
wire n_2113;
wire n_2114;
wire n_2115;
wire n_2116;
wire n_2117;
wire n_2119;
wire n_2120;
wire n_2121;
wire n_2122;
wire n_2125;
wire n_2126;
wire n_2127;
wire n_2129;
wire n_213;
wire n_2131;
wire n_2132;
wire n_2134;
wire n_2135;
wire n_2136;
wire n_2137;
wire n_2138;
wire n_2140;
wire n_2146;
wire n_2147;
wire n_2150;
wire n_2151;
wire n_2152;
wire TIMEBOOST_net_10044;
wire n_2154;
wire TIMEBOOST_net_10326;
wire TIMEBOOST_net_10325;
wire TIMEBOOST_net_10323;
wire n_2159;
wire TIMEBOOST_net_9930;
wire n_2161;
wire n_2162;
wire n_2163;
wire n_2164;
wire n_2165;
wire n_2166;
wire n_2167;
wire n_2168;
wire n_2169;
wire n_2170;
wire n_2171;
wire n_2172;
wire n_2174;
wire n_2175;
wire n_2176;
wire n_2177;
wire n_2178;
wire n_2179;
wire n_2180;
wire n_2181;
wire TIMEBOOST_net_191;
wire n_2183;
wire n_2184;
wire n_2185;
wire n_2186;
wire n_2187;
wire n_2188;
wire n_2189;
wire TIMEBOOST_net_178;
wire n_2191;
wire n_2192;
wire n_2193;
wire n_2194;
wire n_2195;
wire TIMEBOOST_net_177;
wire n_2197;
wire n_2198;
wire n_2199;
wire n_22;
wire n_2200;
wire n_2201;
wire n_2202;
wire n_2203;
wire n_2204;
wire n_2205;
wire n_2206;
wire n_2207;
wire n_2208;
wire n_2209;
wire n_221;
wire n_2210;
wire n_2211;
wire n_2212;
wire n_2213;
wire n_2214;
wire n_2215;
wire n_2218;
wire n_2219;
wire n_2223;
wire n_2224;
wire n_2225;
wire n_2226;
wire n_2227;
wire n_2228;
wire n_2229;
wire n_2230;
wire n_2231;
wire n_2232;
wire n_2233;
wire n_2234;
wire n_2235;
wire n_2236;
wire n_2237;
wire n_2238;
wire n_2243;
wire n_2244;
wire n_2245;
wire n_2246;
wire n_2247;
wire n_2248;
wire n_2249;
wire n_2250;
wire n_2251;
wire n_2252;
wire n_2253;
wire n_2254;
wire n_2255;
wire n_2256;
wire n_2257;
wire n_2258;
wire n_2259;
wire n_2260;
wire n_2261;
wire n_2262;
wire n_2263;
wire n_2264;
wire n_2266;
wire TIMEBOOST_net_9531;
wire n_2269;
wire n_227;
wire n_2271;
wire n_2272;
wire n_2273;
wire n_2274;
wire n_2275;
wire n_2276;
wire n_2280;
wire n_2281;
wire n_2284;
wire n_2285;
wire n_2286;
wire n_2287;
wire n_2289;
wire n_2291;
wire n_2292;
wire n_2293;
wire n_2295;
wire n_2297;
wire n_2298;
wire n_2299;
wire n_23;
wire n_230;
wire n_2300;
wire n_2301;
wire n_2302;
wire n_2303;
wire n_2304;
wire n_2305;
wire n_2306;
wire n_2308;
wire n_231;
wire n_2311;
wire n_2313;
wire n_2314;
wire n_2315;
wire n_2316;
wire n_2319;
wire n_232;
wire n_2326;
wire n_2327;
wire n_2328;
wire n_2329;
wire n_233;
wire n_2331;
wire n_2337;
wire n_2339;
wire n_234;
wire n_2341;
wire n_2343;
wire n_2344;
wire n_2345;
wire n_2347;
wire n_2349;
wire n_235;
wire TIMEBOOST_net_14934;
wire n_2351;
wire n_2352;
wire n_2353;
wire n_2354;
wire TIMEBOOST_net_30;
wire n_2356;
wire n_2358;
wire n_2359;
wire n_236;
wire n_2361;
wire n_2362;
wire n_2363;
wire n_2364;
wire n_2366;
wire n_2367;
wire n_2369;
wire n_2370;
wire n_2371;
wire n_2372;
wire n_2373;
wire n_2374;
wire n_2376;
wire n_2377;
wire n_2378;
wire n_2379;
wire n_2380;
wire n_2386;
wire n_2387;
wire n_2388;
wire n_2389;
wire n_2390;
wire n_2392;
wire n_2395;
wire n_2396;
wire n_2397;
wire n_2398;
wire n_2399;
wire n_24;
wire n_2400;
wire n_2401;
wire n_2402;
wire n_2405;
wire n_2406;
wire n_2407;
wire n_2409;
wire n_2410;
wire n_2411;
wire n_2412;
wire n_2414;
wire n_2415;
wire n_2416;
wire n_2418;
wire n_2419;
wire n_242;
wire n_2420;
wire n_2421;
wire n_2422;
wire n_2423;
wire n_2424;
wire n_2425;
wire n_2426;
wire n_2427;
wire n_2428;
wire n_2429;
wire n_243;
wire n_2430;
wire n_2431;
wire n_2432;
wire n_2433;
wire n_2434;
wire n_2435;
wire n_2436;
wire n_2437;
wire n_2438;
wire TIMEBOOST_net_173;
wire n_2440;
wire n_2441;
wire n_2442;
wire n_2443;
wire n_2445;
wire n_2446;
wire n_2447;
wire n_2449;
wire n_245;
wire n_2451;
wire n_2453;
wire n_2455;
wire n_2456;
wire n_2457;
wire n_2458;
wire n_2459;
wire n_2460;
wire n_2461;
wire n_2462;
wire n_2463;
wire n_2464;
wire n_2468;
wire n_2469;
wire n_247;
wire n_2471;
wire n_2473;
wire n_2474;
wire n_2475;
wire n_2476;
wire n_2477;
wire n_2478;
wire n_2479;
wire n_2482;
wire n_2483;
wire n_2485;
wire n_2486;
wire n_2487;
wire n_2488;
wire n_249;
wire n_2490;
wire n_2491;
wire n_2492;
wire n_2493;
wire n_2494;
wire n_2496;
wire n_2497;
wire n_2498;
wire n_2499;
wire n_2500;
wire n_2501;
wire n_2502;
wire n_2503;
wire n_2504;
wire n_2505;
wire n_2507;
wire n_2508;
wire n_2509;
wire n_251;
wire n_2510;
wire n_2512;
wire n_2513;
wire n_2514;
wire n_2515;
wire n_2516;
wire n_2517;
wire n_2518;
wire n_2519;
wire n_2520;
wire n_2521;
wire n_2522;
wire n_2524;
wire n_2526;
wire n_2527;
wire n_2528;
wire n_2530;
wire n_2531;
wire n_2533;
wire n_2534;
wire n_2536;
wire n_2537;
wire n_2539;
wire n_2540;
wire n_2541;
wire n_2542;
wire n_2543;
wire n_2544;
wire n_2545;
wire n_2546;
wire n_2547;
wire n_255;
wire n_2552;
wire n_2553;
wire n_2555;
wire n_2556;
wire n_2557;
wire n_2558;
wire n_2559;
wire n_2560;
wire n_2562;
wire n_2564;
wire n_2566;
wire n_2567;
wire n_2568;
wire n_2569;
wire n_257;
wire n_2570;
wire n_2571;
wire n_2572;
wire n_2573;
wire n_2574;
wire n_2575;
wire n_2576;
wire n_2577;
wire n_2579;
wire n_2580;
wire n_2581;
wire n_2582;
wire n_2583;
wire n_2584;
wire n_2585;
wire n_2586;
wire n_2587;
wire n_2588;
wire n_2590;
wire n_2592;
wire n_2593;
wire n_2594;
wire n_2595;
wire n_2596;
wire n_2597;
wire n_2598;
wire n_2599;
wire n_26;
wire n_2600;
wire n_2601;
wire n_2602;
wire n_2603;
wire n_2604;
wire n_2605;
wire n_2606;
wire n_2608;
wire n_2609;
wire n_261;
wire n_2610;
wire n_2611;
wire n_2612;
wire n_2613;
wire n_2614;
wire n_2615;
wire n_2616;
wire n_2619;
wire n_2620;
wire n_2621;
wire TIMEBOOST_net_14724;
wire n_2623;
wire n_2624;
wire n_2625;
wire n_2626;
wire TIMEBOOST_net_10801;
wire n_2629;
wire n_263;
wire n_2630;
wire n_2631;
wire n_2632;
wire n_2633;
wire n_2634;
wire n_2635;
wire n_2636;
wire n_2637;
wire n_2638;
wire n_2639;
wire n_2640;
wire n_2641;
wire n_2643;
wire n_2644;
wire n_2645;
wire n_2646;
wire n_2648;
wire n_2649;
wire n_2651;
wire n_2652;
wire n_2653;
wire n_2654;
wire n_2655;
wire n_2656;
wire n_2657;
wire n_2658;
wire n_2659;
wire n_2660;
wire n_2661;
wire n_2662;
wire n_2663;
wire n_2664;
wire n_2665;
wire n_2666;
wire n_2667;
wire n_2668;
wire n_2669;
wire n_2670;
wire n_2671;
wire n_2672;
wire n_2673;
wire n_2674;
wire n_2675;
wire n_2676;
wire n_2677;
wire n_2678;
wire n_2679;
wire n_268;
wire n_2680;
wire n_2681;
wire n_2682;
wire n_2683;
wire n_2684;
wire n_2685;
wire n_2687;
wire n_2691;
wire n_2692;
wire n_2693;
wire n_2694;
wire n_2695;
wire n_2696;
wire n_2697;
wire n_2698;
wire n_2699;
wire n_27;
wire n_2700;
wire n_2701;
wire n_2702;
wire n_2705;
wire n_2706;
wire n_2707;
wire n_2708;
wire n_2709;
wire n_271;
wire n_2710;
wire n_2711;
wire n_2712;
wire n_2713;
wire n_2714;
wire n_2715;
wire n_2716;
wire n_2717;
wire n_2718;
wire n_2719;
wire n_272;
wire n_2720;
wire n_2721;
wire n_2722;
wire n_2723;
wire n_2725;
wire n_2726;
wire n_2727;
wire n_2728;
wire n_2729;
wire n_2730;
wire n_2731;
wire n_2732;
wire n_2734;
wire n_2735;
wire n_2738;
wire n_2739;
wire n_2740;
wire n_2742;
wire n_2744;
wire n_2745;
wire n_2746;
wire n_2747;
wire n_2748;
wire n_2750;
wire n_2751;
wire n_2752;
wire n_2753;
wire n_2754;
wire n_2755;
wire n_2756;
wire n_2757;
wire n_276;
wire n_2761;
wire n_2762;
wire n_2763;
wire n_2764;
wire n_2765;
wire n_2767;
wire n_2768;
wire n_2769;
wire n_277;
wire n_2770;
wire n_2774;
wire n_2775;
wire n_2776;
wire n_2777;
wire n_2778;
wire n_2779;
wire n_278;
wire n_2780;
wire n_2781;
wire n_2782;
wire n_2783;
wire n_2784;
wire n_2785;
wire n_2786;
wire n_2787;
wire n_2788;
wire n_2789;
wire n_279;
wire n_2790;
wire n_2792;
wire n_2793;
wire n_2794;
wire n_2795;
wire n_2797;
wire n_2799;
wire n_28;
wire n_2801;
wire n_2802;
wire n_2803;
wire n_2804;
wire n_2805;
wire n_2806;
wire n_2807;
wire n_2809;
wire n_2812;
wire n_2813;
wire n_2814;
wire n_2815;
wire n_2818;
wire n_2819;
wire n_282;
wire n_2820;
wire n_2821;
wire n_2822;
wire n_2823;
wire n_2824;
wire n_2825;
wire n_2826;
wire n_2828;
wire n_2829;
wire n_2830;
wire n_2831;
wire n_2833;
wire n_2834;
wire n_2835;
wire n_2836;
wire n_2838;
wire n_2839;
wire n_2840;
wire n_2841;
wire n_2842;
wire n_2843;
wire n_2844;
wire n_2846;
wire n_2847;
wire n_2848;
wire n_2849;
wire n_285;
wire n_2851;
wire n_2852;
wire n_2853;
wire n_2854;
wire n_2855;
wire n_2856;
wire n_2857;
wire n_2858;
wire n_2859;
wire n_2860;
wire n_2864;
wire n_2865;
wire n_2866;
wire n_2867;
wire n_2868;
wire n_2869;
wire n_287;
wire n_2870;
wire n_2871;
wire n_2872;
wire n_2873;
wire n_2874;
wire n_2876;
wire n_2877;
wire n_2878;
wire n_288;
wire n_2883;
wire n_2887;
wire n_2888;
wire n_2897;
wire TIMEBOOST_net_14151;
wire n_290;
wire n_2900;
wire n_2902;
wire n_2904;
wire n_2905;
wire n_2906;
wire n_2907;
wire n_2909;
wire n_2910;
wire n_2913;
wire n_2914;
wire n_2915;
wire n_2916;
wire n_2917;
wire n_2918;
wire n_2919;
wire n_292;
wire n_2920;
wire n_2921;
wire n_2922;
wire n_2924;
wire n_2925;
wire n_2926;
wire n_2927;
wire n_2929;
wire n_2930;
wire n_2931;
wire n_2932;
wire n_2933;
wire n_2934;
wire n_2935;
wire n_2937;
wire n_2938;
wire n_2939;
wire n_294;
wire n_2940;
wire n_2941;
wire n_2942;
wire n_2943;
wire n_2946;
wire n_2947;
wire n_2948;
wire n_2949;
wire n_2950;
wire n_2951;
wire n_2952;
wire n_2953;
wire n_2954;
wire n_2955;
wire n_2956;
wire n_2957;
wire n_2958;
wire n_2959;
wire n_2960;
wire n_2961;
wire n_2962;
wire n_2963;
wire n_2964;
wire n_2965;
wire n_2966;
wire n_2967;
wire n_2968;
wire n_2969;
wire n_297;
wire n_2970;
wire n_2971;
wire n_2972;
wire n_2973;
wire n_2979;
wire n_298;
wire n_2980;
wire n_2981;
wire n_2982;
wire n_2983;
wire n_2984;
wire n_2986;
wire n_2987;
wire n_2988;
wire n_2989;
wire n_2990;
wire n_2991;
wire n_2992;
wire n_2993;
wire n_2995;
wire n_2996;
wire n_2997;
wire n_2998;
wire n_2999;
wire n_300;
wire n_3000;
wire n_3001;
wire n_3004;
wire n_3005;
wire n_3006;
wire n_3007;
wire n_3008;
wire n_3013;
wire n_3014;
wire n_3015;
wire n_3016;
wire n_3017;
wire n_3018;
wire n_3019;
wire n_302;
wire n_3020;
wire n_3021;
wire n_3022;
wire n_3023;
wire n_3024;
wire n_3025;
wire n_3026;
wire n_3027;
wire n_3028;
wire n_303;
wire n_3030;
wire n_3031;
wire n_3032;
wire n_3033;
wire n_3034;
wire n_3036;
wire n_3037;
wire n_3039;
wire n_304;
wire n_3040;
wire n_3041;
wire n_3042;
wire n_3043;
wire n_3044;
wire n_3045;
wire n_3046;
wire n_3047;
wire n_3048;
wire n_3049;
wire n_3050;
wire n_3051;
wire n_3052;
wire n_3053;
wire n_3054;
wire n_3055;
wire n_3057;
wire n_3058;
wire n_3059;
wire n_306;
wire n_3060;
wire n_3061;
wire n_3062;
wire n_3064;
wire n_3066;
wire n_3068;
wire n_307;
wire n_3070;
wire n_3071;
wire n_3072;
wire n_3073;
wire n_3074;
wire n_3076;
wire n_3077;
wire n_3078;
wire n_3079;
wire n_3080;
wire n_3081;
wire n_3083;
wire n_3084;
wire n_3087;
wire n_3089;
wire n_3090;
wire n_3107;
wire n_3108;
wire n_3109;
wire n_3110;
wire n_3111;
wire n_3112;
wire n_3114;
wire n_3115;
wire n_3116;
wire n_3117;
wire n_3118;
wire n_3119;
wire n_3120;
wire n_3123;
wire n_3125;
wire n_3126;
wire TIMEBOOST_net_3096;
wire n_313;
wire n_3130;
wire n_3131;
wire n_3132;
wire n_3133;
wire n_3134;
wire n_3135;
wire n_3136;
wire n_3137;
wire n_3138;
wire n_3139;
wire n_3140;
wire n_3141;
wire n_3142;
wire n_3147;
wire n_3148;
wire n_3151;
wire n_3152;
wire n_3153;
wire n_3154;
wire n_3156;
wire n_3157;
wire n_3158;
wire n_3159;
wire n_3160;
wire n_3162;
wire n_3163;
wire n_3164;
wire n_3166;
wire n_3167;
wire n_3168;
wire n_3169;
wire n_317;
wire n_3170;
wire n_3171;
wire n_3172;
wire n_3173;
wire n_3174;
wire n_3175;
wire TIMEBOOST_net_10467;
wire n_3179;
wire n_3184;
wire n_3185;
wire n_3189;
wire n_319;
wire n_3190;
wire n_3191;
wire n_3192;
wire n_3193;
wire n_3194;
wire n_3195;
wire n_3196;
wire n_3197;
wire n_3198;
wire n_3199;
wire n_320;
wire n_3200;
wire n_3201;
wire n_3202;
wire n_3203;
wire n_3204;
wire n_3205;
wire n_3206;
wire n_3207;
wire n_3209;
wire n_321;
wire n_3210;
wire n_3211;
wire n_3212;
wire n_3213;
wire TIMEBOOST_net_10442;
wire n_3215;
wire n_3216;
wire n_3217;
wire n_3219;
wire n_3220;
wire n_3221;
wire n_3222;
wire n_3223;
wire n_3224;
wire n_3226;
wire n_3227;
wire n_3228;
wire n_3229;
wire n_323;
wire n_3231;
wire n_3232;
wire n_3233;
wire n_3235;
wire n_3236;
wire n_3237;
wire n_3238;
wire n_324;
wire n_3241;
wire n_3245;
wire n_3246;
wire n_3247;
wire n_3248;
wire n_325;
wire n_3250;
wire n_3251;
wire n_3252;
wire n_3254;
wire n_3255;
wire n_3256;
wire n_3257;
wire n_3258;
wire n_3259;
wire n_326;
wire n_3260;
wire n_3261;
wire n_3262;
wire n_3265;
wire n_3266;
wire n_3267;
wire n_3268;
wire n_3269;
wire n_3271;
wire n_3273;
wire n_3274;
wire n_3275;
wire n_3276;
wire n_3277;
wire n_3278;
wire n_3279;
wire n_3280;
wire n_3281;
wire n_3282;
wire TIMEBOOST_net_13643;
wire TIMEBOOST_net_14158;
wire n_3285;
wire TIMEBOOST_net_14157;
wire TIMEBOOST_net_11196;
wire TIMEBOOST_net_13630;
wire n_3289;
wire n_329;
wire n_3290;
wire n_3292;
wire n_3293;
wire n_3294;
wire n_3295;
wire n_3296;
wire n_3297;
wire n_3298;
wire n_3301;
wire n_3302;
wire n_3304;
wire n_3305;
wire n_3306;
wire n_331;
wire n_3310;
wire n_3313;
wire n_3314;
wire n_3315;
wire n_3316;
wire n_3317;
wire n_3318;
wire n_3319;
wire n_3320;
wire n_3321;
wire n_3323;
wire n_3324;
wire n_3325;
wire n_3326;
wire n_3327;
wire n_3329;
wire n_333;
wire n_3330;
wire n_3331;
wire n_3332;
wire n_3333;
wire n_3334;
wire n_3335;
wire n_3337;
wire n_3338;
wire n_3339;
wire n_3341;
wire n_3342;
wire n_3344;
wire n_3345;
wire n_3346;
wire n_3347;
wire TIMEBOOST_net_11173;
wire TIMEBOOST_net_11172;
wire n_335;
wire n_3350;
wire n_3351;
wire n_3352;
wire n_3353;
wire n_3354;
wire n_3355;
wire n_3356;
wire n_3357;
wire n_3358;
wire n_3359;
wire n_336;
wire TIMEBOOST_net_10633;
wire n_3361;
wire n_3363;
wire n_3364;
wire n_3365;
wire n_3366;
wire n_3367;
wire n_3368;
wire n_337;
wire n_3370;
wire n_3371;
wire n_3372;
wire n_3373;
wire n_3374;
wire n_3375;
wire n_3376;
wire n_3377;
wire n_3378;
wire n_3379;
wire n_3380;
wire n_3381;
wire n_3384;
wire n_3385;
wire n_3386;
wire n_3387;
wire n_3388;
wire n_3389;
wire n_3390;
wire n_3391;
wire n_3392;
wire n_3393;
wire n_3395;
wire n_3399;
wire n_34;
wire n_340;
wire n_3402;
wire n_3403;
wire n_3404;
wire n_3406;
wire n_3407;
wire n_3408;
wire n_3409;
wire n_341;
wire n_3410;
wire n_3413;
wire TIMEBOOST_net_10986;
wire n_3415;
wire n_3416;
wire n_3417;
wire n_3419;
wire n_342;
wire n_3420;
wire n_3421;
wire n_3422;
wire n_3423;
wire n_3424;
wire n_3425;
wire TIMEBOOST_net_11170;
wire TIMEBOOST_net_11171;
wire n_3428;
wire n_3429;
wire n_343;
wire n_3432;
wire n_3436;
wire n_3437;
wire n_3438;
wire n_3440;
wire n_3443;
wire n_3444;
wire n_3445;
wire n_3446;
wire n_3447;
wire n_3448;
wire n_3449;
wire n_345;
wire n_3450;
wire n_3452;
wire n_3453;
wire n_3454;
wire n_3455;
wire n_3456;
wire TIMEBOOST_net_11175;
wire TIMEBOOST_net_11174;
wire TIMEBOOST_net_13700;
wire n_3460;
wire TIMEBOOST_net_14084;
wire n_3462;
wire n_3463;
wire n_3464;
wire n_3465;
wire n_3466;
wire n_3467;
wire n_3468;
wire TIMEBOOST_net_11169;
wire TIMEBOOST_net_14085;
wire n_3471;
wire n_3472;
wire n_3474;
wire n_3475;
wire n_3476;
wire n_3477;
wire n_3478;
wire n_3479;
wire n_3480;
wire n_3481;
wire n_3482;
wire TIMEBOOST_net_11336;
wire n_3484;
wire n_3485;
wire n_3486;
wire n_3487;
wire n_3488;
wire n_3489;
wire n_349;
wire n_3490;
wire n_3491;
wire n_3492;
wire n_3493;
wire TIMEBOOST_net_11198;
wire TIMEBOOST_net_11039;
wire n_3496;
wire n_3497;
wire n_3498;
wire n_3499;
wire n_350;
wire n_3501;
wire n_3502;
wire n_3503;
wire n_3504;
wire n_3505;
wire TIMEBOOST_net_10527;
wire n_3507;
wire n_3508;
wire n_3509;
wire n_351;
wire n_3510;
wire TIMEBOOST_net_9806;
wire n_3512;
wire n_3513;
wire n_3514;
wire n_3515;
wire n_3516;
wire TIMEBOOST_net_10210;
wire n_3518;
wire n_3519;
wire n_3520;
wire n_3521;
wire n_3522;
wire n_3523;
wire n_3524;
wire n_3525;
wire n_3526;
wire n_3527;
wire TIMEBOOST_net_10428;
wire n_3529;
wire n_3530;
wire n_3531;
wire n_3533;
wire n_3534;
wire n_3535;
wire n_3536;
wire n_3537;
wire n_3538;
wire n_3539;
wire n_354;
wire n_3540;
wire TIMEBOOST_net_13358;
wire n_3542;
wire n_3543;
wire n_3544;
wire n_3545;
wire n_3546;
wire n_3547;
wire n_3548;
wire n_3549;
wire n_3550;
wire n_3551;
wire n_3552;
wire n_3553;
wire n_3554;
wire n_3555;
wire TIMEBOOST_net_10090;
wire n_3558;
wire n_3559;
wire n_3560;
wire n_3561;
wire n_3563;
wire n_3564;
wire n_3565;
wire n_3566;
wire n_3567;
wire n_3568;
wire n_3569;
wire n_357;
wire n_3570;
wire n_3571;
wire n_3572;
wire n_3573;
wire n_3574;
wire n_3575;
wire n_3576;
wire n_3577;
wire n_3578;
wire n_3579;
wire n_358;
wire n_3580;
wire n_3581;
wire n_3582;
wire n_3583;
wire n_3584;
wire n_3585;
wire n_3586;
wire n_3587;
wire n_3588;
wire n_3589;
wire TIMEBOOST_net_10441;
wire TIMEBOOST_net_10628;
wire n_3592;
wire n_3593;
wire n_3594;
wire n_3595;
wire n_3596;
wire n_3597;
wire n_3598;
wire n_3599;
wire n_36;
wire n_360;
wire n_3600;
wire n_3601;
wire n_3602;
wire n_3603;
wire n_3604;
wire n_3605;
wire n_3606;
wire n_3607;
wire n_3608;
wire n_3609;
wire n_3610;
wire n_3611;
wire n_3612;
wire n_3613;
wire n_3614;
wire n_3615;
wire n_3616;
wire n_3617;
wire n_3618;
wire n_3619;
wire n_362;
wire n_3620;
wire n_3621;
wire n_3622;
wire n_3623;
wire n_3624;
wire n_3625;
wire n_3626;
wire n_3627;
wire n_3628;
wire n_3629;
wire n_3630;
wire n_3631;
wire n_3632;
wire n_3633;
wire n_3634;
wire n_3635;
wire n_3636;
wire TIMEBOOST_net_9799;
wire n_3638;
wire n_3639;
wire n_364;
wire n_3640;
wire n_3641;
wire n_3642;
wire n_3643;
wire n_3644;
wire n_3645;
wire n_3646;
wire n_3647;
wire TIMEBOOST_net_493;
wire TIMEBOOST_net_10204;
wire n_3650;
wire n_3651;
wire TIMEBOOST_net_10101;
wire n_3653;
wire n_3654;
wire n_3655;
wire n_3656;
wire n_3657;
wire n_3658;
wire n_3659;
wire n_366;
wire n_3660;
wire n_3661;
wire n_3662;
wire n_3663;
wire n_3664;
wire n_3665;
wire n_3666;
wire n_3667;
wire n_3668;
wire n_3669;
wire n_3670;
wire n_3671;
wire n_3672;
wire n_3673;
wire n_3674;
wire n_3675;
wire n_3676;
wire n_3677;
wire n_3678;
wire n_3679;
wire n_3680;
wire n_3681;
wire n_3682;
wire n_3683;
wire n_3684;
wire n_3685;
wire n_3686;
wire n_3687;
wire n_3688;
wire TIMEBOOST_net_12913;
wire n_369;
wire n_3690;
wire n_3691;
wire n_3692;
wire n_3693;
wire n_3694;
wire n_3695;
wire n_3696;
wire n_3697;
wire n_3698;
wire n_3699;
wire n_370;
wire n_3700;
wire n_3701;
wire n_3702;
wire n_3703;
wire n_3704;
wire n_3705;
wire n_3706;
wire n_3707;
wire n_3708;
wire n_3709;
wire n_3710;
wire n_3711;
wire n_3712;
wire n_3713;
wire n_3714;
wire n_3715;
wire n_3716;
wire n_3717;
wire n_3718;
wire n_3719;
wire n_372;
wire n_3720;
wire n_3721;
wire n_3722;
wire n_3723;
wire n_3724;
wire n_3725;
wire n_3726;
wire n_3727;
wire n_3728;
wire n_3729;
wire n_373;
wire n_3730;
wire n_3731;
wire n_3732;
wire n_3733;
wire n_3734;
wire n_3735;
wire n_3736;
wire n_3737;
wire n_3738;
wire n_3739;
wire n_374;
wire n_3740;
wire n_3741;
wire n_3742;
wire n_3743;
wire n_3744;
wire n_3745;
wire n_3746;
wire n_3747;
wire n_3748;
wire n_3749;
wire n_375;
wire n_3750;
wire n_3751;
wire n_3752;
wire n_3753;
wire n_3754;
wire n_3755;
wire n_3756;
wire n_3757;
wire n_3758;
wire n_3759;
wire n_376;
wire n_3760;
wire n_3761;
wire n_3762;
wire n_3763;
wire n_3764;
wire n_3765;
wire TIMEBOOST_net_9925;
wire n_3767;
wire n_3768;
wire n_3769;
wire n_377;
wire n_3770;
wire n_3771;
wire n_3772;
wire n_3773;
wire n_3774;
wire n_3775;
wire n_3776;
wire n_3777;
wire n_3778;
wire n_3779;
wire n_378;
wire n_3780;
wire n_3781;
wire n_3782;
wire n_3783;
wire n_3784;
wire n_3785;
wire TIMEBOOST_net_10531;
wire n_3787;
wire n_3788;
wire n_3789;
wire n_3790;
wire n_3791;
wire n_3792;
wire n_3793;
wire n_3794;
wire n_3795;
wire n_3796;
wire n_3797;
wire n_3798;
wire n_3799;
wire n_38;
wire n_3800;
wire n_3805;
wire n_3806;
wire n_3807;
wire n_3808;
wire n_3809;
wire n_3810;
wire n_3811;
wire n_3812;
wire TIMEBOOST_net_10100;
wire n_3814;
wire n_3815;
wire TIMEBOOST_net_10062;
wire TIMEBOOST_net_10061;
wire TIMEBOOST_net_10060;
wire TIMEBOOST_net_10059;
wire n_382;
wire n_3820;
wire TIMEBOOST_net_10056;
wire TIMEBOOST_net_10099;
wire n_3823;
wire TIMEBOOST_net_12994;
wire TIMEBOOST_net_10055;
wire TIMEBOOST_net_10098;
wire n_3827;
wire TIMEBOOST_net_10301;
wire TIMEBOOST_net_10097;
wire n_3830;
wire n_3831;
wire n_3832;
wire n_3833;
wire TIMEBOOST_net_10054;
wire TIMEBOOST_net_10096;
wire TIMEBOOST_net_13421;
wire TIMEBOOST_net_13420;
wire TIMEBOOST_net_10095;
wire n_3839;
wire n_384;
wire TIMEBOOST_net_13417;
wire TIMEBOOST_net_15176;
wire TIMEBOOST_net_10052;
wire TIMEBOOST_net_10051;
wire TIMEBOOST_net_10050;
wire TIMEBOOST_net_10094;
wire TIMEBOOST_net_10151;
wire TIMEBOOST_net_10093;
wire n_3848;
wire TIMEBOOST_net_10049;
wire n_385;
wire TIMEBOOST_net_10476;
wire n_3851;
wire TIMEBOOST_net_10525;
wire TIMEBOOST_net_10468;
wire TIMEBOOST_net_10463;
wire TIMEBOOST_net_10523;
wire TIMEBOOST_net_10522;
wire TIMEBOOST_net_10466;
wire TIMEBOOST_net_10465;
wire TIMEBOOST_net_13196;
wire n_386;
wire TIMEBOOST_net_10521;
wire TIMEBOOST_net_10462;
wire n_3862;
wire TIMEBOOST_net_13497;
wire n_3864;
wire TIMEBOOST_net_10520;
wire TIMEBOOST_net_10519;
wire n_3867;
wire TIMEBOOST_net_10168;
wire TIMEBOOST_net_10563;
wire n_3870;
wire n_3871;
wire n_3872;
wire TIMEBOOST_net_13248;
wire n_3874;
wire n_3875;
wire n_3876;
wire TIMEBOOST_net_10479;
wire n_3878;
wire n_3880;
wire n_3881;
wire TIMEBOOST_net_10298;
wire TIMEBOOST_net_13184;
wire TIMEBOOST_net_10518;
wire TIMEBOOST_net_13198;
wire n_3887;
wire TIMEBOOST_net_13133;
wire TIMEBOOST_net_10297;
wire n_389;
wire n_3890;
wire TIMEBOOST_net_13132;
wire TIMEBOOST_net_10296;
wire n_3893;
wire TIMEBOOST_net_13107;
wire TIMEBOOST_net_10092;
wire TIMEBOOST_net_10295;
wire n_3897;
wire n_3898;
wire TIMEBOOST_net_10294;
wire TIMEBOOST_net_10561;
wire TIMEBOOST_net_10517;
wire TIMEBOOST_net_10235;
wire n_3903;
wire TIMEBOOST_net_10560;
wire TIMEBOOST_net_13197;
wire TIMEBOOST_net_10516;
wire n_3907;
wire n_3908;
wire n_3909;
wire n_391;
wire n_3910;
wire TIMEBOOST_net_10645;
wire TIMEBOOST_net_13775;
wire TIMEBOOST_net_13422;
wire TIMEBOOST_net_10408;
wire TIMEBOOST_net_10464;
wire n_3916;
wire n_3917;
wire n_3918;
wire TIMEBOOST_net_10058;
wire TIMEBOOST_net_13590;
wire TIMEBOOST_net_13419;
wire TIMEBOOST_net_10406;
wire TIMEBOOST_net_13418;
wire TIMEBOOST_net_13424;
wire TIMEBOOST_net_10515;
wire n_3926;
wire TIMEBOOST_net_13423;
wire n_3928;
wire n_3929;
wire n_393;
wire TIMEBOOST_net_492;
wire n_3931;
wire TIMEBOOST_net_13414;
wire TIMEBOOST_net_10514;
wire TIMEBOOST_net_13413;
wire n_3935;
wire TIMEBOOST_net_13481;
wire TIMEBOOST_net_10478;
wire n_3938;
wire n_3939;
wire n_3940;
wire TIMEBOOST_net_10477;
wire n_3942;
wire n_3943;
wire TIMEBOOST_net_13416;
wire TIMEBOOST_net_14628;
wire TIMEBOOST_net_10414;
wire TIMEBOOST_net_10621;
wire TIMEBOOST_net_10620;
wire n_3949;
wire n_395;
wire TIMEBOOST_net_9882;
wire TIMEBOOST_net_10613;
wire TIMEBOOST_net_10415;
wire n_3953;
wire n_3954;
wire TIMEBOOST_net_10630;
wire n_3956;
wire TIMEBOOST_net_10614;
wire TIMEBOOST_net_10612;
wire TIMEBOOST_net_10439;
wire n_396;
wire TIMEBOOST_net_10604;
wire TIMEBOOST_net_10420;
wire TIMEBOOST_net_9881;
wire TIMEBOOST_net_10538;
wire TIMEBOOST_net_13673;
wire n_3965;
wire TIMEBOOST_net_9880;
wire TIMEBOOST_net_12625;
wire TIMEBOOST_net_9879;
wire TIMEBOOST_net_9804;
wire n_397;
wire n_3970;
wire n_3971;
wire n_3972;
wire TIMEBOOST_net_9878;
wire n_3974;
wire TIMEBOOST_net_10438;
wire TIMEBOOST_net_10437;
wire TIMEBOOST_net_12749;
wire TIMEBOOST_net_13828;
wire TIMEBOOST_net_9875;
wire n_398;
wire TIMEBOOST_net_494;
wire n_3981;
wire n_3982;
wire TIMEBOOST_net_10423;
wire n_3984;
wire n_3985;
wire n_3986;
wire TIMEBOOST_net_10419;
wire n_3988;
wire TIMEBOOST_net_9874;
wire TIMEBOOST_net_10249;
wire TIMEBOOST_net_10248;
wire TIMEBOOST_net_10418;
wire n_3993;
wire n_3994;
wire TIMEBOOST_net_10629;
wire TIMEBOOST_net_12787;
wire n_3997;
wire TIMEBOOST_net_12788;
wire n_3999;
wire n_40;
wire TIMEBOOST_net_13671;
wire TIMEBOOST_net_13182;
wire n_4002;
wire n_4003;
wire n_4004;
wire n_4005;
wire n_4006;
wire n_4007;
wire n_4008;
wire n_4009;
wire n_401;
wire n_4010;
wire n_4011;
wire n_4012;
wire n_4013;
wire n_4014;
wire n_4015;
wire TIMEBOOST_net_10627;
wire TIMEBOOST_net_9871;
wire TIMEBOOST_net_9870;
wire n_4019;
wire n_4020;
wire n_4021;
wire TIMEBOOST_net_13818;
wire TIMEBOOST_net_10625;
wire n_4024;
wire TIMEBOOST_net_10417;
wire n_4026;
wire n_4027;
wire TIMEBOOST_net_10416;
wire TIMEBOOST_net_10411;
wire n_4030;
wire TIMEBOOST_net_10436;
wire n_4032;
wire n_4033;
wire TIMEBOOST_net_12624;
wire TIMEBOOST_net_10409;
wire TIMEBOOST_net_9868;
wire TIMEBOOST_net_10605;
wire TIMEBOOST_net_13819;
wire TIMEBOOST_net_13767;
wire n_404;
wire TIMEBOOST_net_13820;
wire TIMEBOOST_net_13776;
wire n_4042;
wire n_4043;
wire n_4044;
wire TIMEBOOST_net_10624;
wire TIMEBOOST_net_10609;
wire TIMEBOOST_net_10410;
wire TIMEBOOST_net_10615;
wire TIMEBOOST_net_10435;
wire n_405;
wire TIMEBOOST_net_10412;
wire TIMEBOOST_net_10434;
wire TIMEBOOST_net_13800;
wire TIMEBOOST_net_10618;
wire TIMEBOOST_net_13573;
wire TIMEBOOST_net_10606;
wire n_4056;
wire TIMEBOOST_net_10413;
wire n_4058;
wire TIMEBOOST_net_13574;
wire n_4060;
wire n_4061;
wire TIMEBOOST_net_10433;
wire TIMEBOOST_net_10617;
wire n_4064;
wire TIMEBOOST_net_10422;
wire TIMEBOOST_net_10616;
wire TIMEBOOST_net_10610;
wire n_4068;
wire TIMEBOOST_net_10623;
wire n_407;
wire TIMEBOOST_net_12623;
wire TIMEBOOST_net_10622;
wire n_4072;
wire TIMEBOOST_net_10619;
wire TIMEBOOST_net_10607;
wire TIMEBOOST_net_10603;
wire TIMEBOOST_net_10421;
wire TIMEBOOST_net_12285;
wire n_4078;
wire n_408;
wire n_4080;
wire n_4084;
wire n_4085;
wire n_4086;
wire n_4088;
wire n_409;
wire n_4090;
wire n_4092;
wire n_4093;
wire n_4095;
wire n_4096;
wire n_4097;
wire n_4098;
wire n_4100;
wire n_4101;
wire n_4102;
wire n_4103;
wire n_4104;
wire n_4105;
wire n_4106;
wire n_4107;
wire n_4108;
wire n_4109;
wire n_411;
wire n_4111;
wire n_4112;
wire n_4113;
wire n_4114;
wire n_4115;
wire n_4119;
wire n_412;
wire TIMEBOOST_net_868;
wire n_4123;
wire n_4125;
wire n_413;
wire n_4130;
wire n_4131;
wire n_4132;
wire n_4134;
wire n_4135;
wire n_4136;
wire n_4137;
wire n_4138;
wire n_4140;
wire n_4142;
wire n_4143;
wire n_4144;
wire n_4145;
wire n_4146;
wire n_4149;
wire n_4151;
wire n_4152;
wire n_4153;
wire n_4154;
wire n_4155;
wire n_4156;
wire n_4157;
wire n_4158;
wire TIMEBOOST_net_14898;
wire n_416;
wire n_4160;
wire n_4161;
wire n_4162;
wire n_4163;
wire n_4165;
wire n_4167;
wire n_4168;
wire n_4169;
wire n_4170;
wire n_4171;
wire n_4172;
wire n_4177;
wire TIMEBOOST_net_320;
wire n_4188;
wire n_419;
wire n_4190;
wire TIMEBOOST_net_11698;
wire n_4192;
wire TIMEBOOST_net_11329;
wire n_4194;
wire TIMEBOOST_net_11696;
wire n_4196;
wire n_4197;
wire n_4198;
wire n_4199;
wire n_42;
wire n_420;
wire n_4200;
wire n_4201;
wire n_4202;
wire TIMEBOOST_net_11222;
wire n_4204;
wire n_4205;
wire n_4206;
wire n_4207;
wire n_4208;
wire n_4209;
wire n_4210;
wire n_4211;
wire n_4212;
wire n_4213;
wire n_4214;
wire n_4216;
wire TIMEBOOST_net_11258;
wire n_4219;
wire n_4220;
wire n_4221;
wire n_4222;
wire n_4223;
wire n_4224;
wire n_4225;
wire n_4226;
wire n_4227;
wire n_4228;
wire n_4229;
wire TIMEBOOST_net_10821;
wire n_4231;
wire n_4232;
wire n_4233;
wire n_4234;
wire n_4235;
wire n_4236;
wire n_4237;
wire n_4238;
wire n_4239;
wire n_424;
wire n_4240;
wire n_4241;
wire TIMEBOOST_net_10383;
wire n_4243;
wire n_4244;
wire n_4245;
wire n_4246;
wire TIMEBOOST_net_10211;
wire TIMEBOOST_net_13784;
wire n_4249;
wire n_425;
wire n_4250;
wire n_4251;
wire n_4252;
wire TIMEBOOST_net_10382;
wire n_4254;
wire n_4255;
wire n_4256;
wire n_4257;
wire n_4258;
wire n_4259;
wire n_4260;
wire n_4261;
wire n_4262;
wire n_4263;
wire TIMEBOOST_net_10250;
wire n_4265;
wire n_4266;
wire n_4267;
wire n_4269;
wire n_4270;
wire n_4271;
wire n_4272;
wire n_4273;
wire n_4274;
wire n_4275;
wire n_4276;
wire n_4277;
wire n_4278;
wire n_4279;
wire n_4280;
wire n_4281;
wire n_4282;
wire n_4283;
wire n_4284;
wire TIMEBOOST_net_13306;
wire TIMEBOOST_net_10351;
wire n_4287;
wire n_4288;
wire n_4289;
wire n_4290;
wire n_4291;
wire n_4292;
wire n_4293;
wire n_4295;
wire n_4296;
wire n_4297;
wire n_4298;
wire n_4299;
wire n_430;
wire n_4300;
wire n_4301;
wire n_4302;
wire n_4303;
wire n_4304;
wire n_4305;
wire n_4306;
wire n_4307;
wire n_4308;
wire n_4309;
wire n_4310;
wire n_4311;
wire n_4312;
wire n_4313;
wire n_4314;
wire n_4315;
wire n_4316;
wire n_4317;
wire n_4318;
wire n_4319;
wire n_432;
wire n_4320;
wire n_4321;
wire n_4322;
wire n_4323;
wire n_4324;
wire n_4325;
wire n_4326;
wire n_4327;
wire n_4328;
wire n_4329;
wire n_433;
wire n_4330;
wire n_4331;
wire n_4332;
wire n_4333;
wire n_4334;
wire n_4335;
wire n_4336;
wire n_4337;
wire n_4338;
wire n_4339;
wire n_434;
wire n_4340;
wire n_4341;
wire n_4342;
wire n_4343;
wire n_4344;
wire n_4345;
wire n_4346;
wire n_4347;
wire TIMEBOOST_net_15186;
wire n_4349;
wire n_4350;
wire n_4351;
wire n_4352;
wire n_4353;
wire n_4354;
wire n_4355;
wire n_4356;
wire n_4357;
wire n_4358;
wire n_4359;
wire n_436;
wire TIMEBOOST_net_15187;
wire n_4361;
wire n_4362;
wire n_4363;
wire n_4364;
wire n_4365;
wire n_4366;
wire n_4367;
wire n_4368;
wire n_4369;
wire n_4370;
wire n_4371;
wire n_4372;
wire n_4373;
wire n_4374;
wire n_4375;
wire n_4376;
wire n_4377;
wire n_4378;
wire n_4379;
wire n_4380;
wire n_4381;
wire n_4382;
wire n_4383;
wire n_4384;
wire n_4385;
wire n_4386;
wire n_4387;
wire n_4388;
wire n_4389;
wire n_439;
wire n_4390;
wire n_4391;
wire n_4392;
wire n_4393;
wire n_4394;
wire n_4395;
wire n_4396;
wire n_4397;
wire n_4398;
wire n_4399;
wire n_440;
wire n_4400;
wire n_4401;
wire n_4402;
wire n_4403;
wire n_4404;
wire n_4405;
wire TIMEBOOST_net_9927;
wire n_4407;
wire n_4408;
wire n_4409;
wire n_4410;
wire n_4411;
wire n_4412;
wire TIMEBOOST_net_14621;
wire TIMEBOOST_net_9926;
wire n_4415;
wire n_4416;
wire n_4417;
wire n_4418;
wire n_4419;
wire n_4420;
wire n_4421;
wire n_4422;
wire n_4423;
wire n_4424;
wire n_4425;
wire n_4426;
wire n_4427;
wire n_4428;
wire n_4429;
wire n_4430;
wire n_4431;
wire n_4432;
wire n_4433;
wire n_4434;
wire n_4435;
wire n_4436;
wire n_4437;
wire n_4438;
wire n_4439;
wire n_4440;
wire n_4441;
wire n_4442;
wire n_4443;
wire n_4444;
wire n_4445;
wire n_4446;
wire n_4447;
wire n_4448;
wire n_4449;
wire n_4450;
wire n_4451;
wire n_4452;
wire n_4453;
wire n_4454;
wire n_4455;
wire n_4456;
wire n_4457;
wire n_4458;
wire n_4459;
wire n_4460;
wire n_4461;
wire n_4462;
wire n_4463;
wire n_4464;
wire n_4465;
wire n_4466;
wire n_4467;
wire n_4468;
wire n_4469;
wire n_447;
wire n_4470;
wire n_4471;
wire n_4472;
wire n_4473;
wire n_4474;
wire n_4475;
wire n_4476;
wire n_4477;
wire n_4478;
wire n_4479;
wire n_4480;
wire n_4481;
wire n_4482;
wire n_4483;
wire n_4484;
wire n_4485;
wire n_4486;
wire n_4487;
wire n_4488;
wire n_4489;
wire n_4490;
wire n_4491;
wire n_4492;
wire n_4493;
wire TIMEBOOST_net_13602;
wire n_4495;
wire n_4496;
wire n_4497;
wire n_4498;
wire n_4499;
wire n_4500;
wire n_4501;
wire n_4502;
wire n_4503;
wire n_4504;
wire n_4505;
wire n_4506;
wire n_4507;
wire n_4508;
wire n_4509;
wire n_4510;
wire n_4511;
wire n_4512;
wire n_4513;
wire n_4514;
wire n_4515;
wire TIMEBOOST_net_13398;
wire TIMEBOOST_net_10085;
wire n_4518;
wire n_4519;
wire n_4520;
wire n_4521;
wire TIMEBOOST_net_10321;
wire n_4523;
wire n_4524;
wire n_4525;
wire n_4527;
wire n_4528;
wire n_4532;
wire n_4533;
wire n_4534;
wire n_4535;
wire n_4536;
wire n_4537;
wire n_454;
wire n_4591;
wire TIMEBOOST_net_10149;
wire n_4593;
wire n_4594;
wire n_4595;
wire TIMEBOOST_net_4815;
wire TIMEBOOST_net_4115;
wire n_4598;
wire TIMEBOOST_net_10732;
wire n_46;
wire n_4601;
wire n_4603;
wire n_4605;
wire n_4607;
wire n_4608;
wire n_4609;
wire n_4610;
wire TIMEBOOST_net_10246;
wire n_4612;
wire TIMEBOOST_net_10444;
wire n_4614;
wire n_4616;
wire n_4617;
wire n_4618;
wire n_4619;
wire n_4621;
wire n_4623;
wire n_4625;
wire n_4627;
wire n_4628;
wire n_4629;
wire n_4630;
wire n_4631;
wire n_4632;
wire n_4633;
wire n_4634;
wire n_4635;
wire n_4636;
wire n_4637;
wire n_4638;
wire n_4639;
wire n_4641;
wire n_4642;
wire n_4644;
wire n_4645;
wire n_4646;
wire n_4647;
wire n_4649;
wire n_4652;
wire n_4654;
wire n_4655;
wire n_4656;
wire n_4658;
wire n_4659;
wire n_4660;
wire n_4661;
wire n_4662;
wire n_4663;
wire n_4664;
wire n_4666;
wire n_4667;
wire n_4668;
wire n_4669;
wire n_4670;
wire n_4671;
wire n_4672;
wire n_4673;
wire n_4674;
wire n_4675;
wire TIMEBOOST_net_222;
wire n_4677;
wire n_4678;
wire n_4679;
wire n_4680;
wire n_4681;
wire n_4683;
wire n_4685;
wire n_4686;
wire TIMEBOOST_net_11697;
wire n_4688;
wire TIMEBOOST_net_11694;
wire n_4691;
wire n_4692;
wire n_4693;
wire n_4694;
wire n_4695;
wire n_4696;
wire n_4697;
wire TIMEBOOST_net_11607;
wire n_4699;
wire n_47;
wire n_4700;
wire n_4702;
wire n_4703;
wire n_4704;
wire TIMEBOOST_net_13994;
wire TIMEBOOST_net_11328;
wire n_4707;
wire n_4708;
wire n_471;
wire TIMEBOOST_net_11580;
wire n_4711;
wire n_4712;
wire n_4713;
wire n_4714;
wire n_4715;
wire TIMEBOOST_net_259;
wire n_4717;
wire n_4718;
wire n_4719;
wire n_4720;
wire n_4721;
wire n_4722;
wire TIMEBOOST_net_10137;
wire TIMEBOOST_net_10169;
wire n_4725;
wire n_4726;
wire n_4727;
wire n_4728;
wire n_4729;
wire n_4730;
wire TIMEBOOST_net_10562;
wire n_4732;
wire n_4733;
wire n_4734;
wire n_4735;
wire n_4736;
wire n_4737;
wire n_4739;
wire n_4740;
wire n_4741;
wire n_4743;
wire n_4744;
wire n_4746;
wire TIMEBOOST_net_883;
wire TIMEBOOST_net_10581;
wire TIMEBOOST_net_14118;
wire TIMEBOOST_net_9343;
wire TIMEBOOST_net_882;
wire TIMEBOOST_net_9342;
wire TIMEBOOST_net_10592;
wire TIMEBOOST_net_490;
wire TIMEBOOST_net_489;
wire TIMEBOOST_net_3739;
wire TIMEBOOST_net_9311;
wire TIMEBOOST_net_10583;
wire TIMEBOOST_net_881;
wire TIMEBOOST_net_10582;
wire TIMEBOOST_net_487;
wire TIMEBOOST_net_880;
wire TIMEBOOST_net_10822;
wire TIMEBOOST_net_879;
wire TIMEBOOST_net_485;
wire TIMEBOOST_net_484;
wire TIMEBOOST_net_9344;
wire TIMEBOOST_net_10591;
wire TIMEBOOST_net_483;
wire TIMEBOOST_net_10590;
wire TIMEBOOST_net_12727;
wire TIMEBOOST_net_10589;
wire TIMEBOOST_net_10588;
wire TIMEBOOST_net_10587;
wire TIMEBOOST_net_10586;
wire TIMEBOOST_net_10585;
wire TIMEBOOST_net_878;
wire n_4778;
wire TIMEBOOST_net_10584;
wire n_4780;
wire n_4781;
wire n_4782;
wire n_4783;
wire n_4784;
wire n_4785;
wire n_4786;
wire n_4792;
wire n_4793;
wire n_4795;
wire n_4796;
wire n_4797;
wire n_4798;
wire n_4799;
wire n_4800;
wire n_4802;
wire n_4803;
wire n_4806;
wire n_4807;
wire n_4808;
wire n_4809;
wire n_4811;
wire n_4812;
wire n_4813;
wire n_4814;
wire n_4815;
wire n_4816;
wire n_4818;
wire n_4819;
wire n_4820;
wire n_4822;
wire n_4823;
wire n_4824;
wire n_4825;
wire n_4826;
wire n_4828;
wire n_4830;
wire n_4831;
wire n_4832;
wire n_4833;
wire n_4834;
wire n_4835;
wire n_4836;
wire n_4837;
wire n_4838;
wire n_4839;
wire n_4840;
wire n_4841;
wire n_4842;
wire n_4843;
wire n_4844;
wire n_4845;
wire n_4846;
wire n_4847;
wire n_4848;
wire n_4849;
wire n_4851;
wire n_4853;
wire n_4855;
wire n_4856;
wire n_4857;
wire n_4858;
wire n_4859;
wire n_4860;
wire n_4861;
wire n_4862;
wire n_4863;
wire n_4864;
wire n_4866;
wire n_4867;
wire n_4868;
wire n_4869;
wire n_4870;
wire n_4871;
wire n_4872;
wire n_4873;
wire n_4874;
wire TIMEBOOST_net_14508;
wire n_4877;
wire n_4878;
wire n_4879;
wire n_4880;
wire n_4881;
wire n_4883;
wire n_4884;
wire TIMEBOOST_net_11643;
wire n_4886;
wire TIMEBOOST_net_11693;
wire TIMEBOOST_net_11207;
wire n_4889;
wire n_4890;
wire n_4891;
wire n_4892;
wire TIMEBOOST_net_13908;
wire n_4894;
wire n_4895;
wire n_4896;
wire n_4897;
wire n_4899;
wire n_4900;
wire n_4901;
wire n_4902;
wire n_4903;
wire n_4904;
wire n_4905;
wire n_4906;
wire n_4907;
wire n_4908;
wire n_4909;
wire n_4911;
wire n_4912;
wire n_4913;
wire n_4914;
wire n_4915;
wire n_4917;
wire n_4918;
wire n_4920;
wire n_4922;
wire n_4924;
wire n_4926;
wire n_4928;
wire n_4930;
wire n_4932;
wire n_4934;
wire n_4936;
wire n_4939;
wire n_4941;
wire n_4943;
wire n_4945;
wire n_4947;
wire n_4949;
wire n_4951;
wire n_4953;
wire n_4955;
wire n_4957;
wire n_4959;
wire n_4961;
wire n_4963;
wire n_4965;
wire n_4968;
wire n_497;
wire n_4970;
wire n_4973;
wire n_4975;
wire n_4978;
wire n_4980;
wire n_4982;
wire n_4984;
wire n_4986;
wire n_4988;
wire n_4991;
wire n_4993;
wire n_4996;
wire n_4999;
wire n_50;
wire n_5001;
wire n_5003;
wire n_5006;
wire n_5009;
wire n_5012;
wire n_5014;
wire n_5016;
wire n_5018;
wire n_5021;
wire n_5023;
wire n_5025;
wire n_5027;
wire n_5029;
wire n_5031;
wire n_5033;
wire n_5036;
wire n_5038;
wire n_504;
wire n_5040;
wire n_5042;
wire n_5044;
wire n_5046;
wire n_5048;
wire n_5050;
wire n_5052;
wire n_5054;
wire n_5056;
wire n_5058;
wire n_5060;
wire n_5062;
wire n_5064;
wire n_5066;
wire n_5068;
wire n_5071;
wire n_5074;
wire n_5076;
wire n_5078;
wire n_5080;
wire n_5082;
wire n_5084;
wire n_5086;
wire n_5088;
wire n_5090;
wire n_5092;
wire n_5094;
wire n_5096;
wire n_5098;
wire n_5100;
wire n_5102;
wire n_5104;
wire n_5106;
wire n_5108;
wire n_5110;
wire n_5112;
wire n_5114;
wire n_5116;
wire n_5118;
wire n_512;
wire n_5120;
wire n_5122;
wire n_5124;
wire n_5126;
wire n_5128;
wire n_513;
wire n_5130;
wire n_5132;
wire n_5134;
wire n_5136;
wire n_5138;
wire n_5140;
wire n_5143;
wire n_5146;
wire n_5149;
wire n_5151;
wire n_5153;
wire n_5156;
wire n_5158;
wire n_5161;
wire n_5163;
wire n_5166;
wire n_5168;
wire n_5170;
wire n_5172;
wire n_5174;
wire n_5176;
wire n_5179;
wire n_518;
wire n_5181;
wire n_5183;
wire n_5185;
wire n_5188;
wire n_519;
wire n_5190;
wire n_5192;
wire n_5194;
wire n_5196;
wire n_5198;
wire n_520;
wire n_5200;
wire n_5203;
wire n_5205;
wire n_5207;
wire n_521;
wire n_5210;
wire n_5212;
wire n_5214;
wire n_5216;
wire n_5218;
wire n_522;
wire n_5221;
wire n_5223;
wire n_5225;
wire n_5227;
wire n_5228;
wire n_5229;
wire n_523;
wire n_5230;
wire TIMEBOOST_net_11354;
wire n_5232;
wire n_5235;
wire n_5237;
wire n_524;
wire n_5240;
wire n_5242;
wire n_5244;
wire n_5246;
wire n_5248;
wire n_525;
wire n_5251;
wire n_5253;
wire n_5255;
wire n_5258;
wire n_526;
wire n_5260;
wire n_5263;
wire n_5265;
wire n_5267;
wire n_5269;
wire n_527;
wire n_5272;
wire n_5275;
wire n_5277;
wire n_5279;
wire n_528;
wire n_5281;
wire n_5283;
wire n_5285;
wire n_5288;
wire n_529;
wire n_5290;
wire n_5293;
wire n_5296;
wire n_5298;
wire n_530;
wire n_5300;
wire n_5303;
wire n_5305;
wire n_5308;
wire n_531;
wire n_5311;
wire n_5313;
wire n_5315;
wire n_5318;
wire n_532;
wire n_5320;
wire n_5323;
wire n_5325;
wire n_5327;
wire n_533;
wire n_5330;
wire n_5332;
wire n_5335;
wire n_5337;
wire n_5339;
wire n_534;
wire n_5342;
wire n_5345;
wire n_5347;
wire n_5349;
wire n_535;
wire n_5351;
wire n_5354;
wire n_5356;
wire n_5358;
wire n_536;
wire n_5361;
wire n_5363;
wire n_5366;
wire n_5368;
wire n_5371;
wire n_5373;
wire n_5376;
wire n_5378;
wire n_538;
wire n_5380;
wire n_5383;
wire n_5386;
wire n_5388;
wire n_539;
wire n_5391;
wire n_5393;
wire n_5396;
wire n_5399;
wire n_540;
wire n_5402;
wire n_5404;
wire n_5406;
wire n_5409;
wire n_541;
wire n_5412;
wire n_5414;
wire n_5416;
wire n_5418;
wire n_5421;
wire n_5424;
wire n_5427;
wire n_5429;
wire n_5431;
wire n_5433;
wire n_5435;
wire n_5438;
wire n_544;
wire n_5441;
wire n_5444;
wire n_5446;
wire n_5448;
wire n_545;
wire n_5450;
wire n_5452;
wire n_5454;
wire n_5456;
wire n_5458;
wire n_546;
wire n_5461;
wire n_5463;
wire n_5465;
wire n_5467;
wire n_547;
wire n_5470;
wire n_5472;
wire n_5474;
wire n_5476;
wire n_5478;
wire n_5481;
wire n_5483;
wire n_5486;
wire n_5489;
wire n_549;
wire n_5491;
wire n_5493;
wire n_5495;
wire n_5497;
wire n_5499;
wire n_550;
wire n_5501;
wire n_5503;
wire n_5505;
wire n_5507;
wire n_5509;
wire n_551;
wire n_5511;
wire n_5513;
wire n_5515;
wire n_5517;
wire n_5519;
wire n_5521;
wire n_5523;
wire n_5526;
wire n_5528;
wire n_5531;
wire n_5534;
wire n_5537;
wire n_5539;
wire n_554;
wire n_5541;
wire n_5543;
wire n_5545;
wire n_5546;
wire n_5547;
wire n_5548;
wire n_5549;
wire n_5552;
wire n_5553;
wire n_5554;
wire n_5555;
wire n_5556;
wire n_5557;
wire n_5558;
wire n_5559;
wire n_5561;
wire n_5563;
wire n_5565;
wire n_5566;
wire n_5567;
wire n_5568;
wire n_5569;
wire n_5570;
wire n_5571;
wire n_5572;
wire n_5573;
wire n_5574;
wire n_5575;
wire n_5576;
wire n_5577;
wire n_5578;
wire n_5579;
wire n_558;
wire n_5580;
wire n_5581;
wire n_5582;
wire n_5583;
wire n_5585;
wire n_5587;
wire n_5588;
wire n_5589;
wire n_559;
wire n_5591;
wire n_5592;
wire n_5593;
wire n_5594;
wire n_5595;
wire n_5597;
wire n_5598;
wire n_560;
wire n_5600;
wire n_5601;
wire n_5603;
wire n_5604;
wire n_5606;
wire n_5607;
wire n_5608;
wire n_5609;
wire n_561;
wire n_5611;
wire n_5612;
wire n_5614;
wire n_5616;
wire n_5617;
wire n_5618;
wire n_5619;
wire n_562;
wire n_5620;
wire n_5622;
wire n_5623;
wire n_5625;
wire n_5626;
wire n_5627;
wire n_5628;
wire n_563;
wire n_5630;
wire n_5631;
wire n_5632;
wire n_5633;
wire n_5634;
wire n_5635;
wire n_5636;
wire n_5637;
wire n_5638;
wire n_5639;
wire n_564;
wire n_5640;
wire n_5641;
wire n_5642;
wire n_5643;
wire n_5644;
wire TIMEBOOST_net_13937;
wire n_5646;
wire n_5648;
wire n_5649;
wire n_565;
wire n_5650;
wire n_5651;
wire n_5652;
wire n_5654;
wire n_5655;
wire n_5656;
wire n_5657;
wire n_5658;
wire n_566;
wire n_5660;
wire n_5662;
wire n_5663;
wire n_5664;
wire n_5666;
wire n_5668;
wire n_5669;
wire n_567;
wire n_5670;
wire n_5672;
wire n_5673;
wire n_5675;
wire n_5676;
wire n_5678;
wire n_5679;
wire n_568;
wire n_5681;
wire n_5682;
wire n_5684;
wire n_5686;
wire n_5687;
wire n_5688;
wire n_5689;
wire n_5691;
wire n_5694;
wire n_5696;
wire n_5699;
wire n_57;
wire n_5701;
wire n_5702;
wire n_5703;
wire n_5704;
wire n_5705;
wire n_5707;
wire n_5708;
wire n_5709;
wire n_5710;
wire n_5712;
wire n_5713;
wire n_5716;
wire n_5717;
wire n_5718;
wire n_5722;
wire n_5723;
wire n_5724;
wire n_5725;
wire n_5728;
wire TIMEBOOST_net_11647;
wire n_573;
wire n_5730;
wire n_5731;
wire n_5732;
wire n_5733;
wire n_5735;
wire n_5736;
wire n_5737;
wire n_5739;
wire n_574;
wire n_5740;
wire n_5741;
wire n_5742;
wire n_5743;
wire n_5744;
wire n_5745;
wire n_5747;
wire n_5748;
wire TIMEBOOST_net_13483;
wire n_5750;
wire n_5751;
wire TIMEBOOST_net_11645;
wire n_5753;
wire n_5754;
wire n_5755;
wire n_5757;
wire n_5758;
wire TIMEBOOST_net_11358;
wire n_5763;
wire n_5766;
wire n_5768;
wire n_5769;
wire n_5770;
wire n_5772;
wire n_5774;
wire n_5776;
wire n_5778;
wire n_5780;
wire n_5782;
wire n_5784;
wire n_5786;
wire n_5788;
wire n_5790;
wire n_5792;
wire n_5794;
wire n_5796;
wire n_5798;
wire n_580;
wire n_5800;
wire n_5802;
wire n_5804;
wire n_5806;
wire n_5808;
wire n_581;
wire n_5810;
wire n_5812;
wire n_5814;
wire n_5816;
wire n_5819;
wire n_582;
wire n_5822;
wire n_5824;
wire n_5827;
wire n_583;
wire n_5830;
wire n_5833;
wire n_5836;
wire n_5838;
wire n_584;
wire n_5840;
wire n_5842;
wire n_5844;
wire n_5846;
wire n_5848;
wire n_585;
wire n_5850;
wire n_5852;
wire n_5854;
wire n_5856;
wire n_5858;
wire n_586;
wire n_5860;
wire n_5862;
wire n_5864;
wire n_5866;
wire n_5868;
wire n_587;
wire n_5870;
wire n_5872;
wire n_5874;
wire n_5876;
wire n_5878;
wire n_588;
wire n_5880;
wire n_5882;
wire n_5884;
wire n_5886;
wire n_5888;
wire n_5890;
wire n_5892;
wire n_5894;
wire n_5896;
wire n_5898;
wire n_5900;
wire n_5902;
wire n_5904;
wire n_5906;
wire n_5908;
wire n_5910;
wire n_5912;
wire n_5914;
wire n_5916;
wire n_5918;
wire n_592;
wire n_5920;
wire n_5922;
wire n_5924;
wire n_5926;
wire n_5928;
wire n_593;
wire n_5930;
wire n_5932;
wire n_5934;
wire n_5936;
wire n_5938;
wire n_594;
wire n_5940;
wire n_5942;
wire n_5944;
wire n_5946;
wire n_5948;
wire n_595;
wire n_5950;
wire n_5952;
wire n_5954;
wire n_5956;
wire n_5958;
wire n_596;
wire n_5960;
wire n_5962;
wire n_5964;
wire n_5966;
wire n_5967;
wire n_5969;
wire n_597;
wire n_5971;
wire n_5973;
wire n_5975;
wire n_5977;
wire n_5979;
wire n_598;
wire n_5981;
wire n_5983;
wire n_5985;
wire n_5987;
wire n_5989;
wire n_599;
wire n_5991;
wire n_5993;
wire n_5995;
wire n_5997;
wire n_5999;
wire n_6;
wire n_600;
wire n_6001;
wire n_6003;
wire n_6005;
wire n_6007;
wire n_6009;
wire n_601;
wire n_6011;
wire n_6013;
wire n_6015;
wire n_6017;
wire n_6019;
wire n_602;
wire n_6021;
wire n_6023;
wire n_6025;
wire n_6027;
wire n_6029;
wire n_603;
wire n_6031;
wire n_6033;
wire n_6035;
wire n_6037;
wire n_6039;
wire n_604;
wire n_6040;
wire n_6041;
wire n_6043;
wire n_6045;
wire n_6047;
wire n_6049;
wire n_605;
wire n_6051;
wire n_6053;
wire n_6054;
wire n_6056;
wire n_6058;
wire n_606;
wire n_6060;
wire n_6061;
wire n_6063;
wire n_6065;
wire n_6067;
wire n_6069;
wire n_607;
wire n_6071;
wire n_6073;
wire n_6075;
wire n_6077;
wire n_6079;
wire n_6081;
wire n_6083;
wire n_6085;
wire n_6087;
wire n_6089;
wire n_609;
wire n_6091;
wire n_6093;
wire n_6095;
wire n_6097;
wire n_6099;
wire n_61;
wire n_610;
wire n_6101;
wire n_6103;
wire n_6105;
wire n_6107;
wire n_6109;
wire n_611;
wire n_6111;
wire n_6112;
wire n_6115;
wire n_6117;
wire n_6119;
wire n_612;
wire n_6121;
wire n_6123;
wire n_6125;
wire n_6127;
wire n_6129;
wire n_613;
wire n_6132;
wire n_6135;
wire n_6136;
wire n_6138;
wire n_614;
wire n_6140;
wire n_6142;
wire n_6144;
wire n_6146;
wire n_6148;
wire n_615;
wire n_6150;
wire n_6152;
wire n_6154;
wire n_6156;
wire n_6158;
wire n_616;
wire n_6160;
wire n_6162;
wire n_6164;
wire n_6166;
wire n_6168;
wire n_617;
wire n_6171;
wire n_6173;
wire n_6175;
wire n_6177;
wire n_6179;
wire n_6181;
wire n_6184;
wire n_6186;
wire n_6189;
wire n_6191;
wire n_6193;
wire n_6195;
wire n_6196;
wire n_6199;
wire n_620;
wire n_6200;
wire n_6201;
wire n_6204;
wire n_6206;
wire n_6208;
wire n_621;
wire n_6211;
wire n_6213;
wire n_6216;
wire n_6218;
wire n_622;
wire n_6221;
wire n_6223;
wire n_6226;
wire n_6228;
wire n_623;
wire n_6230;
wire n_6231;
wire n_6232;
wire n_6234;
wire n_6235;
wire n_6238;
wire n_624;
wire n_6240;
wire n_6243;
wire n_6246;
wire n_6249;
wire n_625;
wire n_6252;
wire n_6254;
wire n_6257;
wire n_6259;
wire n_626;
wire n_6261;
wire n_6264;
wire n_6266;
wire n_6268;
wire n_627;
wire n_6271;
wire n_6273;
wire n_6276;
wire n_6278;
wire n_6281;
wire n_6284;
wire n_6286;
wire n_6287;
wire n_6289;
wire n_629;
wire n_6292;
wire n_6295;
wire n_6297;
wire n_6298;
wire n_6301;
wire n_6303;
wire n_6305;
wire n_6308;
wire n_6311;
wire n_6313;
wire n_6315;
wire n_6318;
wire n_6319;
wire n_6321;
wire n_6323;
wire n_6325;
wire n_6327;
wire n_6329;
wire n_6331;
wire n_6333;
wire n_6334;
wire n_6335;
wire n_6337;
wire n_6338;
wire n_6340;
wire n_6342;
wire n_6344;
wire n_6345;
wire n_6347;
wire n_6348;
wire n_6350;
wire n_6353;
wire n_6355;
wire n_6356;
wire n_6358;
wire n_6361;
wire n_6364;
wire n_6366;
wire n_6369;
wire n_6371;
wire n_6372;
wire n_6373;
wire n_6374;
wire n_6376;
wire n_6379;
wire n_6382;
wire n_6384;
wire n_6386;
wire n_6388;
wire n_639;
wire n_6390;
wire n_6391;
wire n_6393;
wire n_6395;
wire n_6398;
wire n_640;
wire n_6400;
wire n_6402;
wire n_6405;
wire n_6407;
wire n_641;
wire n_6410;
wire n_6413;
wire n_6415;
wire n_6417;
wire n_642;
wire n_6420;
wire n_6423;
wire n_6425;
wire n_6427;
wire n_643;
wire n_6430;
wire n_6431;
wire n_6433;
wire n_6435;
wire n_6436;
wire n_6438;
wire n_6440;
wire n_6443;
wire n_6446;
wire n_6448;
wire n_645;
wire n_6451;
wire n_6453;
wire n_6456;
wire n_6458;
wire n_646;
wire n_6461;
wire n_6463;
wire n_6465;
wire n_6468;
wire n_6470;
wire n_6473;
wire n_6475;
wire n_6477;
wire n_648;
wire n_6480;
wire n_6483;
wire n_6485;
wire n_6488;
wire n_649;
wire n_6490;
wire n_6493;
wire n_6495;
wire n_6498;
wire n_65;
wire n_650;
wire n_6501;
wire n_6504;
wire n_6506;
wire n_6509;
wire n_6512;
wire n_6514;
wire n_6516;
wire n_6518;
wire n_652;
wire n_6521;
wire n_6523;
wire n_6526;
wire n_6528;
wire n_653;
wire n_6530;
wire n_6532;
wire n_6534;
wire n_6536;
wire n_6538;
wire n_6541;
wire n_6543;
wire n_6546;
wire n_6548;
wire n_655;
wire n_6550;
wire n_6553;
wire n_6554;
wire n_6556;
wire n_6558;
wire n_656;
wire n_6561;
wire n_6563;
wire n_6566;
wire n_6567;
wire n_6569;
wire n_657;
wire n_6572;
wire n_6575;
wire n_6578;
wire n_658;
wire n_6580;
wire n_6582;
wire n_6585;
wire n_6587;
wire n_6589;
wire n_659;
wire n_6592;
wire n_6594;
wire n_6596;
wire n_6598;
wire n_660;
wire n_6601;
wire n_6603;
wire n_6605;
wire n_6607;
wire n_661;
wire n_6610;
wire n_6613;
wire n_6615;
wire n_6617;
wire n_662;
wire n_6620;
wire n_6621;
wire n_6623;
wire n_6624;
wire n_6626;
wire n_6629;
wire n_663;
wire n_6631;
wire n_6634;
wire n_6636;
wire n_6639;
wire n_664;
wire n_6641;
wire n_6644;
wire n_6645;
wire n_6647;
wire n_6649;
wire n_665;
wire n_6651;
wire n_6654;
wire n_6657;
wire n_6659;
wire n_666;
wire n_6662;
wire n_6665;
wire n_6668;
wire n_667;
wire n_6670;
wire n_6672;
wire n_6674;
wire n_6676;
wire n_6678;
wire n_668;
wire n_6680;
wire n_6682;
wire n_6684;
wire n_6686;
wire n_6689;
wire n_669;
wire n_6691;
wire n_6693;
wire n_6695;
wire n_6697;
wire n_6699;
wire n_67;
wire n_670;
wire n_6701;
wire n_6703;
wire n_6705;
wire n_6707;
wire n_6709;
wire n_671;
wire n_6712;
wire n_6714;
wire n_6716;
wire n_6718;
wire n_672;
wire n_6720;
wire n_6722;
wire n_6724;
wire n_6726;
wire n_6729;
wire n_673;
wire n_6731;
wire n_6733;
wire n_6735;
wire n_6738;
wire n_674;
wire n_6741;
wire n_6743;
wire n_6745;
wire n_6747;
wire n_6749;
wire n_675;
wire n_6752;
wire n_6754;
wire n_6757;
wire n_6759;
wire n_676;
wire n_6761;
wire n_6763;
wire n_6766;
wire n_6768;
wire n_677;
wire n_6770;
wire n_6772;
wire n_6774;
wire n_6776;
wire n_6778;
wire n_678;
wire n_6781;
wire n_6783;
wire n_6785;
wire n_6788;
wire n_6789;
wire n_6791;
wire n_6793;
wire n_6795;
wire n_6797;
wire n_6799;
wire n_6801;
wire n_6804;
wire n_6806;
wire n_6809;
wire n_681;
wire n_6812;
wire n_6814;
wire n_6816;
wire n_6819;
wire n_6821;
wire n_6824;
wire n_6826;
wire n_6828;
wire n_6830;
wire n_6833;
wire n_6835;
wire n_6837;
wire n_6840;
wire n_6842;
wire n_6845;
wire n_6847;
wire n_6849;
wire n_6851;
wire n_6853;
wire n_6855;
wire n_6857;
wire n_6859;
wire n_6861;
wire n_6863;
wire n_6865;
wire n_6867;
wire n_6868;
wire n_6869;
wire n_6871;
wire n_6872;
wire n_6875;
wire n_6876;
wire n_6878;
wire n_6880;
wire n_6883;
wire n_6885;
wire n_6886;
wire n_6887;
wire n_6889;
wire n_689;
wire n_6892;
wire n_6895;
wire n_6897;
wire n_6898;
wire n_6900;
wire n_6902;
wire n_6903;
wire n_6905;
wire n_6908;
wire n_691;
wire n_6910;
wire n_6911;
wire n_6913;
wire n_6915;
wire n_6917;
wire n_6919;
wire n_692;
wire n_6920;
wire n_6922;
wire n_6924;
wire n_6926;
wire n_6929;
wire n_6932;
wire n_6934;
wire n_6935;
wire n_6937;
wire n_6940;
wire n_6941;
wire n_6942;
wire n_6943;
wire n_6944;
wire n_6946;
wire n_6948;
wire n_695;
wire n_6951;
wire n_6953;
wire n_6956;
wire n_6958;
wire n_696;
wire n_6961;
wire n_6963;
wire n_6965;
wire n_6967;
wire n_6969;
wire n_6971;
wire n_6973;
wire n_6975;
wire n_6977;
wire n_6978;
wire n_6980;
wire n_6982;
wire n_6983;
wire n_6984;
wire n_6985;
wire n_6986;
wire n_6987;
wire TIMEBOOST_net_12960;
wire n_6989;
wire n_6991;
wire n_6992;
wire n_6993;
wire n_6994;
wire n_6995;
wire n_6996;
wire n_6997;
wire n_6998;
wire n_6999;
wire n_700;
wire n_7000;
wire n_7001;
wire n_7002;
wire n_7003;
wire n_7004;
wire n_7005;
wire n_7006;
wire n_7007;
wire n_7008;
wire n_7009;
wire n_7010;
wire n_7011;
wire n_7012;
wire n_7013;
wire n_7014;
wire n_7015;
wire n_7016;
wire n_7018;
wire n_7019;
wire n_7027;
wire n_7028;
wire n_7029;
wire n_703;
wire n_7030;
wire n_7031;
wire n_7032;
wire n_7033;
wire n_7038;
wire n_7039;
wire n_7040;
wire n_7043;
wire n_7044;
wire n_7045;
wire n_7046;
wire n_7047;
wire n_7048;
wire n_7049;
wire n_705;
wire n_7050;
wire n_7051;
wire n_7052;
wire n_7053;
wire n_7054;
wire n_7055;
wire n_7056;
wire n_7057;
wire n_7058;
wire n_7059;
wire n_7060;
wire n_7061;
wire n_7062;
wire n_7063;
wire n_7064;
wire n_7065;
wire n_7066;
wire n_7067;
wire n_7068;
wire n_7069;
wire n_707;
wire n_7070;
wire n_7071;
wire n_7072;
wire n_7073;
wire n_7074;
wire n_7075;
wire TIMEBOOST_net_14833;
wire n_7078;
wire n_7079;
wire n_708;
wire n_7080;
wire n_7081;
wire n_7082;
wire n_7083;
wire n_7084;
wire g52462_da;
wire g52468_da;
wire TIMEBOOST_net_4415;
wire TIMEBOOST_net_12968;
wire n_709;
wire n_7091;
wire n_7092;
wire n_7093;
wire n_7094;
wire n_7095;
wire n_7096;
wire n_7102;
wire n_7108;
wire n_711;
wire n_7110;
wire n_7112;
wire n_7114;
wire n_7115;
wire n_7117;
wire n_7119;
wire n_7121;
wire n_7122;
wire n_7123;
wire n_7125;
wire n_7126;
wire n_7128;
wire n_713;
wire n_7130;
wire n_7132;
wire n_7134;
wire n_7135;
wire n_7136;
wire n_7137;
wire n_7139;
wire n_7141;
wire n_7143;
wire n_7145;
wire n_7147;
wire n_7149;
wire n_715;
wire n_7151;
wire n_7153;
wire n_7155;
wire n_7157;
wire n_7159;
wire n_716;
wire n_7161;
wire n_7163;
wire n_7165;
wire n_7168;
wire n_7171;
wire n_7174;
wire n_7177;
wire n_7180;
wire n_7182;
wire n_7185;
wire n_7187;
wire n_7189;
wire n_7191;
wire n_7193;
wire n_7195;
wire n_7197;
wire n_72;
wire n_7200;
wire n_7203;
wire n_7205;
wire n_7207;
wire n_7209;
wire n_721;
wire n_7210;
wire n_7211;
wire n_7212;
wire n_7213;
wire n_7214;
wire n_7215;
wire n_7216;
wire n_7217;
wire TIMEBOOST_net_10407;
wire TIMEBOOST_net_10512;
wire n_722;
wire n_7220;
wire TIMEBOOST_net_13576;
wire TIMEBOOST_net_10431;
wire TIMEBOOST_net_10626;
wire n_7227;
wire n_7228;
wire n_7229;
wire n_7231;
wire n_7232;
wire n_7233;
wire n_7234;
wire n_7235;
wire n_7236;
wire n_7237;
wire n_7238;
wire n_7239;
wire n_7240;
wire n_7241;
wire n_7242;
wire n_7243;
wire n_7244;
wire n_7245;
wire n_7246;
wire n_7247;
wire n_7248;
wire n_7249;
wire n_725;
wire n_7250;
wire n_7251;
wire n_7252;
wire n_7253;
wire n_7254;
wire n_7255;
wire n_7256;
wire n_7257;
wire n_7258;
wire n_7259;
wire n_7260;
wire n_7261;
wire n_7262;
wire n_7263;
wire n_7264;
wire n_7265;
wire n_7266;
wire n_7267;
wire n_7268;
wire n_7269;
wire n_727;
wire n_7270;
wire n_7271;
wire n_7272;
wire n_7273;
wire n_7274;
wire n_7275;
wire n_7276;
wire n_7277;
wire n_7278;
wire n_7279;
wire n_7280;
wire n_7281;
wire n_7282;
wire n_7283;
wire n_7284;
wire n_7285;
wire n_7286;
wire n_7287;
wire n_7288;
wire n_7289;
wire n_729;
wire n_7290;
wire n_7291;
wire n_7293;
wire n_7294;
wire n_7295;
wire n_7296;
wire n_7297;
wire n_7298;
wire n_730;
wire n_7300;
wire n_7307;
wire n_7308;
wire n_7309;
wire n_731;
wire n_7310;
wire n_7311;
wire n_7312;
wire n_7313;
wire n_7315;
wire n_7316;
wire n_7317;
wire TIMEBOOST_net_11140;
wire n_7320;
wire n_7321;
wire n_7322;
wire n_7324;
wire n_7325;
wire n_7326;
wire TIMEBOOST_net_722;
wire n_7329;
wire n_733;
wire n_7330;
wire TIMEBOOST_net_721;
wire n_7333;
wire TIMEBOOST_net_13981;
wire TIMEBOOST_net_11588;
wire TIMEBOOST_net_10909;
wire n_7338;
wire n_7339;
wire n_734;
wire n_7341;
wire TIMEBOOST_net_11653;
wire n_7350;
wire n_736;
wire n_7362;
wire n_7364;
wire n_7366;
wire n_7368;
wire n_7369;
wire n_737;
wire n_7371;
wire n_7373;
wire n_7374;
wire n_7375;
wire n_7377;
wire n_7379;
wire n_738;
wire n_7381;
wire n_7383;
wire n_7385;
wire n_7386;
wire n_7387;
wire n_7388;
wire n_739;
wire n_7390;
wire n_7392;
wire n_7393;
wire n_7396;
wire n_7397;
wire n_7398;
wire n_7399;
wire n_74;
wire n_740;
wire n_7400;
wire n_7401;
wire n_7404;
wire n_7405;
wire n_7406;
wire n_7407;
wire n_7408;
wire n_7409;
wire n_741;
wire n_7410;
wire n_7411;
wire n_7412;
wire n_7413;
wire n_7414;
wire n_7415;
wire n_7416;
wire n_7417;
wire n_7418;
wire n_7419;
wire n_742;
wire n_7420;
wire n_7421;
wire n_7422;
wire n_7423;
wire n_7424;
wire n_7425;
wire n_7426;
wire n_7427;
wire n_7428;
wire n_7429;
wire n_743;
wire n_7430;
wire n_7431;
wire n_7432;
wire n_7433;
wire n_7434;
wire n_7435;
wire n_7436;
wire n_7437;
wire n_7438;
wire n_7439;
wire n_744;
wire n_7440;
wire n_7442;
wire n_7443;
wire n_7444;
wire n_7445;
wire n_7446;
wire n_7447;
wire n_7448;
wire n_7449;
wire n_745;
wire n_7450;
wire n_7451;
wire n_7452;
wire n_7453;
wire n_7454;
wire n_7455;
wire n_7456;
wire n_7457;
wire n_7458;
wire n_7459;
wire n_746;
wire n_7460;
wire n_7461;
wire n_7462;
wire n_7463;
wire n_7464;
wire n_7465;
wire n_7466;
wire n_7467;
wire n_7468;
wire n_7469;
wire n_747;
wire n_7470;
wire TIMEBOOST_net_14569;
wire n_7472;
wire n_7473;
wire n_7474;
wire n_7475;
wire n_7476;
wire n_7477;
wire n_7478;
wire n_7479;
wire n_748;
wire n_7480;
wire n_7481;
wire n_7482;
wire n_7483;
wire n_7484;
wire n_7485;
wire n_7486;
wire n_7487;
wire n_7488;
wire n_7489;
wire n_7490;
wire n_7491;
wire n_7492;
wire n_7493;
wire n_7494;
wire n_7495;
wire n_7496;
wire n_7497;
wire n_7498;
wire n_7499;
wire n_75;
wire n_7500;
wire n_7504;
wire n_7505;
wire n_7508;
wire n_7509;
wire n_7510;
wire n_7511;
wire n_7512;
wire n_7513;
wire n_7514;
wire n_7515;
wire n_7516;
wire n_7517;
wire n_7518;
wire n_7519;
wire n_7521;
wire n_7522;
wire n_7523;
wire n_7524;
wire n_7525;
wire n_7527;
wire n_7528;
wire n_7529;
wire n_7530;
wire n_7531;
wire n_7532;
wire n_7534;
wire n_7535;
wire n_7538;
wire n_7539;
wire n_7540;
wire n_7541;
wire n_7542;
wire n_7543;
wire n_7544;
wire n_7547;
wire n_7548;
wire n_7550;
wire n_7551;
wire n_7552;
wire n_7557;
wire n_7558;
wire n_7559;
wire n_7560;
wire n_7561;
wire n_7562;
wire n_7564;
wire n_7565;
wire n_7567;
wire n_7568;
wire n_7569;
wire n_7571;
wire n_7574;
wire n_7575;
wire n_7576;
wire n_7577;
wire n_7578;
wire n_7579;
wire n_7580;
wire n_7581;
wire n_7582;
wire n_7583;
wire n_7584;
wire n_7585;
wire n_7586;
wire n_7587;
wire n_7588;
wire n_7589;
wire n_7590;
wire n_7591;
wire n_7592;
wire n_7593;
wire n_7594;
wire n_7595;
wire n_7596;
wire n_7597;
wire n_7598;
wire n_7599;
wire n_76;
wire n_7600;
wire n_7601;
wire n_7602;
wire n_7603;
wire n_7604;
wire n_7605;
wire n_7606;
wire n_7607;
wire n_7608;
wire n_7609;
wire n_7610;
wire n_7611;
wire n_7612;
wire n_7613;
wire n_7614;
wire n_7615;
wire n_7616;
wire n_7617;
wire n_7618;
wire n_7619;
wire n_7620;
wire n_7621;
wire n_7622;
wire n_7624;
wire n_7625;
wire n_7626;
wire n_7627;
wire n_7628;
wire n_7629;
wire n_763;
wire n_7630;
wire n_7631;
wire n_7632;
wire n_7633;
wire n_7634;
wire n_7635;
wire n_7636;
wire n_7637;
wire n_7638;
wire n_7639;
wire n_7640;
wire n_7642;
wire n_7643;
wire n_7645;
wire n_7646;
wire n_7647;
wire n_7648;
wire n_7649;
wire n_7650;
wire n_7651;
wire n_7652;
wire n_7653;
wire n_7654;
wire n_7655;
wire n_7656;
wire n_7657;
wire n_7658;
wire n_7661;
wire n_7663;
wire n_7664;
wire n_7665;
wire n_7666;
wire n_7667;
wire n_7669;
wire n_7671;
wire n_7672;
wire n_7673;
wire n_7677;
wire n_7679;
wire n_7681;
wire n_7683;
wire n_7684;
wire n_7685;
wire n_7687;
wire n_7689;
wire n_7692;
wire n_7694;
wire n_7695;
wire n_7697;
wire n_7698;
wire n_7699;
wire n_7701;
wire n_7702;
wire n_7704;
wire n_7705;
wire n_7706;
wire n_7707;
wire n_7708;
wire n_7709;
wire TIMEBOOST_net_11188;
wire n_7711;
wire n_7712;
wire n_7714;
wire n_7715;
wire n_7716;
wire n_7717;
wire n_7718;
wire n_7719;
wire n_7720;
wire n_7721;
wire n_7722;
wire n_7723;
wire n_7724;
wire n_7725;
wire n_7726;
wire TIMEBOOST_net_319;
wire TIMEBOOST_net_318;
wire n_7731;
wire n_7733;
wire n_7734;
wire n_7735;
wire n_7737;
wire n_7738;
wire n_7739;
wire n_7740;
wire n_7742;
wire n_7743;
wire n_7744;
wire n_7745;
wire n_7746;
wire n_7747;
wire n_7749;
wire n_7750;
wire n_7751;
wire n_7752;
wire n_7753;
wire n_7754;
wire n_7755;
wire n_7756;
wire n_7757;
wire n_7759;
wire n_7760;
wire n_7761;
wire n_7762;
wire n_7764;
wire n_7766;
wire n_7767;
wire n_7768;
wire n_7769;
wire n_7771;
wire n_7773;
wire n_7774;
wire n_7776;
wire n_7777;
wire n_7779;
wire n_7780;
wire n_7781;
wire n_7782;
wire n_7783;
wire n_7785;
wire n_7786;
wire n_7787;
wire n_7788;
wire n_7789;
wire n_779;
wire n_7790;
wire n_7791;
wire n_7792;
wire n_7793;
wire n_7794;
wire n_7795;
wire n_7796;
wire n_7797;
wire n_7798;
wire n_7799;
wire n_7800;
wire n_7801;
wire n_7802;
wire n_7803;
wire n_7804;
wire n_7805;
wire n_7806;
wire n_7807;
wire n_7808;
wire n_7809;
wire n_7810;
wire n_7811;
wire n_7812;
wire n_7813;
wire n_7814;
wire n_7815;
wire n_7816;
wire n_7817;
wire n_7818;
wire n_7819;
wire n_7820;
wire n_7821;
wire n_7822;
wire n_7823;
wire n_7824;
wire n_7826;
wire n_7828;
wire n_783;
wire n_7830;
wire n_7833;
wire n_7835;
wire n_7836;
wire n_7838;
wire n_784;
wire n_7840;
wire n_7842;
wire n_7844;
wire n_7845;
wire n_7847;
wire n_7849;
wire n_785;
wire n_7851;
wire n_7853;
wire n_7855;
wire n_7857;
wire n_7859;
wire n_7861;
wire n_7863;
wire n_7865;
wire n_7867;
wire n_7869;
wire n_7871;
wire n_7873;
wire n_7875;
wire n_7877;
wire n_7879;
wire n_7881;
wire n_7883;
wire n_7885;
wire n_7887;
wire n_7889;
wire n_7891;
wire n_7893;
wire n_7895;
wire n_7897;
wire n_7899;
wire n_790;
wire n_7901;
wire n_7903;
wire n_7905;
wire n_7907;
wire n_7909;
wire n_791;
wire n_7911;
wire n_7913;
wire n_7915;
wire n_7917;
wire n_7919;
wire n_7921;
wire n_7923;
wire n_7925;
wire n_7927;
wire n_7929;
wire n_7931;
wire n_7933;
wire n_7935;
wire n_7937;
wire n_7939;
wire n_7941;
wire n_7943;
wire n_7945;
wire n_7947;
wire n_7949;
wire n_7951;
wire n_7953;
wire n_7955;
wire n_7957;
wire n_7959;
wire n_7961;
wire n_7963;
wire n_7965;
wire n_7967;
wire n_7969;
wire n_7971;
wire n_7973;
wire n_7975;
wire n_7977;
wire n_7979;
wire n_798;
wire n_7981;
wire n_7983;
wire n_7985;
wire n_7987;
wire n_7989;
wire n_7991;
wire n_7993;
wire n_7995;
wire n_7997;
wire n_7999;
wire n_8001;
wire n_8003;
wire n_8005;
wire n_8007;
wire n_8009;
wire n_8012;
wire n_8014;
wire n_8017;
wire n_8019;
wire n_802;
wire n_8021;
wire n_8024;
wire n_8027;
wire n_8030;
wire n_8032;
wire n_8034;
wire n_8036;
wire n_8039;
wire n_8041;
wire n_8044;
wire n_8047;
wire n_8049;
wire n_8052;
wire n_8054;
wire n_8056;
wire n_8059;
wire n_8060;
wire n_8062;
wire n_8064;
wire n_8066;
wire n_8068;
wire n_8069;
wire n_8071;
wire n_8073;
wire n_8076;
wire n_8079;
wire n_808;
wire n_8082;
wire n_8084;
wire n_8087;
wire n_8089;
wire n_8092;
wire n_8094;
wire n_8097;
wire n_8100;
wire n_8102;
wire n_8105;
wire n_8107;
wire n_8109;
wire n_8111;
wire n_8114;
wire n_8116;
wire n_8118;
wire n_8119;
wire n_812;
wire n_8121;
wire n_8123;
wire n_8125;
wire n_8128;
wire n_813;
wire n_8130;
wire n_8132;
wire n_8135;
wire n_8137;
wire n_8139;
wire n_8140;
wire n_8142;
wire n_8144;
wire n_8147;
wire n_815;
wire n_8150;
wire n_8152;
wire n_8154;
wire n_8157;
wire n_8159;
wire n_816;
wire n_8161;
wire n_8163;
wire n_8166;
wire n_8168;
wire n_817;
wire n_8171;
wire n_8173;
wire n_8175;
wire n_8176;
wire n_8178;
wire n_8180;
wire n_8182;
wire n_8184;
wire n_8186;
wire n_8189;
wire n_819;
wire n_8191;
wire n_8193;
wire n_8196;
wire n_8198;
wire n_8200;
wire n_8203;
wire n_8205;
wire n_8208;
wire n_8210;
wire n_8213;
wire n_8215;
wire n_8218;
wire n_8220;
wire n_8223;
wire n_8226;
wire n_8229;
wire n_8231;
wire n_8232;
wire n_8234;
wire n_8236;
wire n_8239;
wire n_824;
wire n_8241;
wire n_8244;
wire n_8246;
wire n_8248;
wire n_8251;
wire n_8253;
wire n_8255;
wire n_8258;
wire n_826;
wire n_8260;
wire n_8262;
wire n_8264;
wire n_8267;
wire n_8269;
wire n_8271;
wire n_8272;
wire n_8274;
wire n_8277;
wire n_8279;
wire n_8281;
wire n_8283;
wire n_8285;
wire n_8288;
wire n_829;
wire n_8291;
wire n_8293;
wire n_8295;
wire n_8297;
wire n_8299;
wire n_83;
wire n_8302;
wire n_8304;
wire n_8307;
wire n_8309;
wire n_8311;
wire n_8313;
wire n_8316;
wire n_8319;
wire n_832;
wire n_8321;
wire n_8323;
wire n_8325;
wire n_8327;
wire n_8329;
wire n_833;
wire n_8331;
wire n_8333;
wire n_8335;
wire n_8337;
wire n_8339;
wire n_8341;
wire n_8344;
wire n_8346;
wire n_8349;
wire n_8351;
wire n_8353;
wire n_8355;
wire n_8358;
wire n_836;
wire n_8360;
wire n_8362;
wire n_8364;
wire n_8366;
wire n_8368;
wire n_837;
wire n_8371;
wire n_8373;
wire n_8376;
wire n_8379;
wire n_838;
wire n_8382;
wire n_8384;
wire n_8387;
wire n_8389;
wire n_839;
wire n_8391;
wire n_8393;
wire n_8395;
wire n_8397;
wire n_84;
wire n_840;
wire n_8400;
wire n_8402;
wire n_8404;
wire n_8406;
wire n_8407;
wire n_8409;
wire n_841;
wire n_8411;
wire n_8413;
wire n_8415;
wire n_8417;
wire n_8419;
wire n_842;
wire n_8421;
wire n_8423;
wire n_8426;
wire n_8428;
wire n_843;
wire n_8430;
wire n_8431;
wire n_8432;
wire n_8433;
wire n_8434;
wire n_8436;
wire n_8437;
wire n_8438;
wire n_8439;
wire n_844;
wire n_8440;
wire n_8441;
wire n_8442;
wire n_8444;
wire n_8445;
wire n_8446;
wire n_8447;
wire n_8448;
wire n_8449;
wire n_845;
wire n_8450;
wire n_8451;
wire n_8452;
wire n_8453;
wire n_8454;
wire n_8455;
wire n_8456;
wire n_8457;
wire n_8458;
wire n_8459;
wire n_8460;
wire n_8461;
wire n_8462;
wire n_8463;
wire n_8464;
wire n_8465;
wire n_8466;
wire n_8467;
wire n_8468;
wire n_8469;
wire n_847;
wire n_8470;
wire n_8472;
wire n_8474;
wire n_8476;
wire n_8477;
wire n_8478;
wire n_8480;
wire n_8481;
wire n_8482;
wire n_8483;
wire n_8484;
wire n_8485;
wire n_8486;
wire n_8487;
wire n_8488;
wire n_8489;
wire n_849;
wire TIMEBOOST_net_14012;
wire n_8492;
wire n_8493;
wire n_8494;
wire n_8495;
wire n_8496;
wire n_8498;
wire n_85;
wire n_850;
wire TIMEBOOST_net_11731;
wire n_8501;
wire n_8502;
wire n_8503;
wire n_8504;
wire n_8505;
wire n_8506;
wire n_8508;
wire n_8509;
wire n_851;
wire n_8510;
wire n_8511;
wire n_8512;
wire n_8513;
wire n_8514;
wire n_8515;
wire n_8516;
wire n_8517;
wire n_8518;
wire n_8519;
wire n_852;
wire n_8520;
wire n_8521;
wire n_8522;
wire n_8523;
wire n_8524;
wire n_8525;
wire n_8526;
wire n_8527;
wire n_8528;
wire n_8529;
wire n_853;
wire n_8530;
wire n_8531;
wire TIMEBOOST_net_10982;
wire n_8535;
wire n_8538;
wire TIMEBOOST_net_1154;
wire n_8540;
wire n_8541;
wire n_8542;
wire n_8547;
wire n_8548;
wire n_8549;
wire n_855;
wire n_8550;
wire n_8551;
wire n_8552;
wire n_8553;
wire n_8554;
wire n_8555;
wire n_8556;
wire n_8557;
wire n_8558;
wire n_8559;
wire n_8560;
wire n_8561;
wire n_8562;
wire n_8563;
wire n_8564;
wire n_8565;
wire n_8566;
wire n_8567;
wire n_8568;
wire n_8569;
wire n_8570;
wire n_8571;
wire n_8572;
wire n_8573;
wire n_8574;
wire n_8575;
wire n_8576;
wire n_8579;
wire n_858;
wire TIMEBOOST_net_1172;
wire n_8582;
wire n_8583;
wire n_8585;
wire n_8588;
wire n_8589;
wire n_8590;
wire n_8591;
wire n_8595;
wire n_8596;
wire n_8597;
wire n_8598;
wire n_8601;
wire n_8602;
wire n_8603;
wire n_8604;
wire n_8605;
wire n_8606;
wire n_8607;
wire n_8609;
wire n_861;
wire n_8611;
wire n_8613;
wire n_8615;
wire n_8616;
wire n_8617;
wire n_8618;
wire n_8619;
wire n_8620;
wire n_8621;
wire n_8622;
wire n_8623;
wire n_8624;
wire n_8625;
wire n_8626;
wire n_8627;
wire n_8628;
wire n_8629;
wire n_863;
wire n_8630;
wire n_8631;
wire n_8632;
wire n_8633;
wire n_8634;
wire n_8635;
wire n_8636;
wire n_8637;
wire n_8638;
wire n_864;
wire n_8640;
wire n_8641;
wire n_8642;
wire n_8643;
wire n_8644;
wire n_8645;
wire n_8646;
wire n_8647;
wire n_8648;
wire n_8649;
wire n_865;
wire n_8650;
wire n_8651;
wire n_8652;
wire n_8653;
wire n_8655;
wire n_8656;
wire n_8657;
wire n_8658;
wire n_8659;
wire n_866;
wire n_8660;
wire n_8661;
wire n_8662;
wire n_8664;
wire n_8665;
wire n_8668;
wire n_8669;
wire n_867;
wire n_8672;
wire n_8673;
wire n_8674;
wire n_8675;
wire n_8676;
wire n_8677;
wire n_8678;
wire n_868;
wire n_8680;
wire n_8682;
wire n_8686;
wire n_8687;
wire n_8688;
wire n_869;
wire n_8692;
wire n_8693;
wire n_8694;
wire n_8695;
wire n_8697;
wire n_8699;
wire n_870;
wire n_8701;
wire n_8703;
wire n_8705;
wire n_8707;
wire n_8708;
wire n_8709;
wire n_871;
wire n_8711;
wire n_8712;
wire n_8713;
wire n_8714;
wire n_8716;
wire n_8717;
wire n_872;
wire n_8721;
wire n_8723;
wire n_8724;
wire n_8725;
wire n_8726;
wire n_8727;
wire n_8728;
wire n_8730;
wire n_8731;
wire n_8732;
wire n_8733;
wire n_8734;
wire TIMEBOOST_net_11897;
wire TIMEBOOST_net_11896;
wire n_874;
wire TIMEBOOST_net_11895;
wire TIMEBOOST_net_11894;
wire TIMEBOOST_net_11768;
wire TIMEBOOST_net_11915;
wire TIMEBOOST_net_2899;
wire n_8745;
wire TIMEBOOST_net_12484;
wire n_8747;
wire TIMEBOOST_net_14352;
wire n_8749;
wire n_875;
wire n_8750;
wire n_8751;
wire n_8752;
wire TIMEBOOST_net_5199;
wire n_8757;
wire n_8759;
wire n_876;
wire n_8760;
wire n_8765;
wire n_877;
wire n_878;
wire n_8780;
wire n_8782;
wire n_8784;
wire n_879;
wire n_8790;
wire n_8792;
wire n_8794;
wire n_8796;
wire n_880;
wire n_8800;
wire n_8801;
wire n_881;
wire n_8818;
wire n_8819;
wire n_882;
wire n_8820;
wire n_883;
wire n_8831;
wire n_8832;
wire TIMEBOOST_net_14098;
wire n_884;
wire TIMEBOOST_net_14023;
wire n_8842;
wire n_8843;
wire n_8846;
wire n_8847;
wire n_8848;
wire n_8849;
wire n_885;
wire n_8850;
wire n_8851;
wire n_8852;
wire n_8853;
wire n_8854;
wire n_8855;
wire n_8857;
wire n_8859;
wire n_886;
wire n_8860;
wire n_8861;
wire n_8863;
wire n_8864;
wire n_8866;
wire n_8867;
wire n_887;
wire n_8871;
wire n_8872;
wire n_8874;
wire n_8875;
wire n_8876;
wire n_8877;
wire n_8879;
wire n_888;
wire n_8880;
wire n_8884;
wire n_8887;
wire n_8888;
wire n_8889;
wire n_889;
wire n_8890;
wire n_8892;
wire n_8896;
wire n_8897;
wire n_8898;
wire n_8899;
wire n_890;
wire n_8900;
wire n_8902;
wire n_8904;
wire n_8906;
wire n_8908;
wire n_891;
wire n_8910;
wire n_8912;
wire n_8914;
wire n_8916;
wire n_8917;
wire n_8919;
wire n_892;
wire n_8920;
wire n_8921;
wire n_8924;
wire n_8926;
wire n_8927;
wire n_8928;
wire n_893;
wire n_8932;
wire n_8934;
wire n_8935;
wire n_8939;
wire n_894;
wire n_8940;
wire n_8941;
wire n_8943;
wire n_8944;
wire n_8945;
wire n_8946;
wire n_8947;
wire n_8949;
wire n_895;
wire n_8950;
wire TIMEBOOST_net_13310;
wire TIMEBOOST_net_13307;
wire n_8953;
wire n_8954;
wire n_8955;
wire n_8957;
wire n_8959;
wire n_896;
wire n_8960;
wire n_8961;
wire n_8962;
wire n_8963;
wire n_8964;
wire n_8965;
wire n_8966;
wire n_8967;
wire n_8968;
wire n_8969;
wire n_897;
wire n_8970;
wire n_8971;
wire n_8973;
wire n_8975;
wire n_8977;
wire n_8979;
wire n_898;
wire n_8981;
wire n_8983;
wire n_8986;
wire n_8989;
wire n_899;
wire n_8990;
wire n_8991;
wire n_8992;
wire n_8993;
wire n_8994;
wire n_8995;
wire n_8996;
wire n_8997;
wire n_8998;
wire n_8999;
wire n_9;
wire n_900;
wire n_9000;
wire n_9001;
wire n_9002;
wire n_9003;
wire n_9004;
wire n_9005;
wire n_9006;
wire n_9007;
wire n_9008;
wire n_9009;
wire n_901;
wire n_9010;
wire n_9011;
wire n_9012;
wire n_9013;
wire n_9014;
wire n_9015;
wire n_9016;
wire n_9017;
wire n_9018;
wire n_9019;
wire n_902;
wire n_9020;
wire n_9021;
wire n_9022;
wire n_9023;
wire n_9024;
wire n_9025;
wire n_9026;
wire n_9027;
wire n_9028;
wire n_9029;
wire n_903;
wire n_9030;
wire n_9031;
wire n_9032;
wire n_9033;
wire n_9034;
wire n_9035;
wire n_9036;
wire n_9037;
wire n_9038;
wire n_9039;
wire n_904;
wire n_9040;
wire n_9041;
wire n_9042;
wire n_9043;
wire n_9044;
wire n_9045;
wire n_9046;
wire n_9047;
wire n_9048;
wire n_9049;
wire n_905;
wire n_9050;
wire n_9051;
wire n_9052;
wire TIMEBOOST_net_13432;
wire n_9054;
wire n_9055;
wire n_9056;
wire n_9057;
wire n_9058;
wire n_9059;
wire n_906;
wire TIMEBOOST_net_12743;
wire n_9061;
wire n_9062;
wire n_9063;
wire n_9064;
wire n_9065;
wire n_9066;
wire n_9067;
wire TIMEBOOST_net_12742;
wire n_9069;
wire n_907;
wire n_9070;
wire n_9071;
wire n_9072;
wire n_9073;
wire n_9074;
wire n_9075;
wire n_9076;
wire n_9077;
wire n_9078;
wire n_9079;
wire n_908;
wire n_9080;
wire n_9081;
wire n_9082;
wire n_9083;
wire n_9084;
wire n_9085;
wire n_9086;
wire n_9087;
wire n_9088;
wire n_9089;
wire n_909;
wire n_9090;
wire n_9091;
wire n_9092;
wire n_9093;
wire n_9094;
wire n_9095;
wire n_9096;
wire n_9097;
wire n_9098;
wire n_9099;
wire n_910;
wire n_9100;
wire n_9101;
wire n_9102;
wire n_9103;
wire n_9104;
wire n_9105;
wire n_9106;
wire n_9107;
wire n_9108;
wire n_9109;
wire n_911;
wire n_9110;
wire n_9111;
wire n_9112;
wire n_9113;
wire n_9114;
wire n_9115;
wire n_9116;
wire n_9117;
wire n_9118;
wire n_9119;
wire n_912;
wire n_9120;
wire n_9121;
wire n_9122;
wire n_9123;
wire n_9124;
wire n_9125;
wire n_9126;
wire n_9127;
wire n_9128;
wire n_9129;
wire n_913;
wire n_9130;
wire n_9131;
wire n_9132;
wire n_9133;
wire n_9134;
wire n_9135;
wire n_9136;
wire n_9137;
wire n_9138;
wire n_9139;
wire n_914;
wire n_9140;
wire n_9141;
wire n_9142;
wire n_9143;
wire n_9144;
wire n_9145;
wire n_9146;
wire n_915;
wire n_9152;
wire n_9153;
wire n_9154;
wire n_9155;
wire n_916;
wire n_9160;
wire n_9163;
wire n_9168;
wire n_917;
wire n_9170;
wire n_9171;
wire n_9172;
wire n_9173;
wire n_9174;
wire n_9175;
wire n_9176;
wire n_9177;
wire n_9178;
wire n_9179;
wire n_918;
wire n_9180;
wire n_9181;
wire n_9182;
wire n_9183;
wire n_9184;
wire n_9185;
wire n_9187;
wire n_9188;
wire n_9189;
wire n_919;
wire n_9191;
wire n_9192;
wire n_9194;
wire n_9197;
wire n_9198;
wire n_9199;
wire n_920;
wire n_9200;
wire n_9201;
wire n_9202;
wire n_9203;
wire n_9204;
wire n_9205;
wire n_9206;
wire n_9207;
wire n_9208;
wire n_9209;
wire n_921;
wire n_9210;
wire n_9214;
wire n_9215;
wire n_9216;
wire n_9217;
wire n_9218;
wire n_9219;
wire n_922;
wire n_9220;
wire n_9221;
wire n_9222;
wire n_9223;
wire n_9224;
wire n_9225;
wire n_9226;
wire n_9227;
wire n_9228;
wire n_9229;
wire n_923;
wire n_9230;
wire n_9231;
wire n_9232;
wire n_9233;
wire n_9234;
wire n_9235;
wire n_9236;
wire n_9237;
wire n_9238;
wire n_9239;
wire n_924;
wire n_9241;
wire n_925;
wire n_9256;
wire n_926;
wire n_9260;
wire n_9261;
wire n_9262;
wire n_9265;
wire n_9269;
wire n_927;
wire n_9270;
wire n_9271;
wire n_9272;
wire n_9274;
wire n_9276;
wire n_9277;
wire n_928;
wire n_9280;
wire n_9283;
wire n_9284;
wire n_9285;
wire n_9286;
wire n_9287;
wire n_929;
wire n_9290;
wire n_9293;
wire n_9294;
wire n_9295;
wire n_9296;
wire n_9297;
wire n_9298;
wire n_9299;
wire n_930;
wire n_9301;
wire n_9303;
wire n_9305;
wire n_9306;
wire n_9307;
wire n_9309;
wire n_931;
wire n_9311;
wire n_9312;
wire n_9315;
wire n_9319;
wire n_9320;
wire n_9321;
wire n_9322;
wire n_9325;
wire n_9328;
wire n_9329;
wire n_9330;
wire n_9331;
wire n_9332;
wire n_9334;
wire n_9335;
wire n_9336;
wire n_9338;
wire n_9340;
wire n_9341;
wire n_9342;
wire n_9343;
wire n_9345;
wire n_9346;
wire n_9348;
wire n_9350;
wire n_9353;
wire n_9355;
wire n_9358;
wire n_9361;
wire n_9363;
wire n_9366;
wire n_9368;
wire n_937;
wire n_9371;
wire n_9372;
wire n_9374;
wire n_9377;
wire n_9379;
wire n_938;
wire n_9381;
wire n_9383;
wire n_9385;
wire n_9387;
wire n_9389;
wire n_939;
wire n_9391;
wire n_9393;
wire n_9396;
wire n_9398;
wire n_940;
wire n_9400;
wire n_9402;
wire n_9404;
wire n_9405;
wire n_9406;
wire n_9407;
wire n_9408;
wire n_9409;
wire n_941;
wire n_9410;
wire n_9411;
wire TIMEBOOST_net_13829;
wire n_9413;
wire n_9414;
wire n_9415;
wire n_9416;
wire n_9418;
wire n_9419;
wire n_9420;
wire n_9421;
wire n_9423;
wire n_9424;
wire n_9425;
wire n_9426;
wire n_9427;
wire n_9428;
wire n_943;
wire n_9430;
wire n_9431;
wire n_9432;
wire n_9433;
wire n_9434;
wire n_9435;
wire n_9436;
wire n_9437;
wire n_9438;
wire n_9439;
wire n_944;
wire n_9440;
wire n_9441;
wire n_9442;
wire n_9443;
wire n_9444;
wire n_9445;
wire n_9446;
wire n_9447;
wire n_9448;
wire n_9449;
wire n_945;
wire n_9450;
wire n_9451;
wire n_9452;
wire n_9453;
wire n_9454;
wire n_9455;
wire n_9456;
wire n_9457;
wire n_9458;
wire n_9459;
wire n_946;
wire n_9460;
wire n_9461;
wire n_9462;
wire n_9463;
wire n_9464;
wire n_9465;
wire n_9466;
wire n_9467;
wire n_9468;
wire n_9469;
wire n_947;
wire n_9470;
wire n_9471;
wire n_9472;
wire n_9473;
wire n_9474;
wire n_9475;
wire n_9476;
wire n_9477;
wire n_9478;
wire n_9479;
wire n_948;
wire n_9480;
wire n_9481;
wire n_9482;
wire n_9483;
wire n_9484;
wire n_9485;
wire n_9486;
wire n_9487;
wire n_9488;
wire n_9489;
wire n_9490;
wire n_9491;
wire n_9492;
wire n_9493;
wire n_9494;
wire n_9495;
wire n_9496;
wire n_9497;
wire n_9498;
wire n_9499;
wire n_95;
wire n_950;
wire n_9500;
wire n_9501;
wire n_9502;
wire n_9503;
wire n_9504;
wire n_9505;
wire n_9506;
wire n_9507;
wire n_9508;
wire n_9509;
wire n_951;
wire n_9510;
wire n_9511;
wire n_9512;
wire n_9513;
wire n_9514;
wire n_9515;
wire n_9516;
wire n_9517;
wire n_9518;
wire n_9519;
wire n_952;
wire n_9520;
wire n_9521;
wire n_9522;
wire n_9523;
wire n_9524;
wire n_9525;
wire n_9526;
wire n_9527;
wire n_9528;
wire n_9529;
wire n_9530;
wire n_9531;
wire n_9532;
wire n_9534;
wire n_9535;
wire n_9537;
wire n_9538;
wire n_9539;
wire n_9540;
wire n_9541;
wire n_9542;
wire n_9543;
wire n_9544;
wire n_9545;
wire n_9546;
wire n_9547;
wire n_9548;
wire n_9549;
wire n_9550;
wire n_9551;
wire n_9552;
wire n_9553;
wire n_9554;
wire n_9555;
wire n_9556;
wire n_9557;
wire n_9558;
wire n_9559;
wire n_956;
wire n_9560;
wire n_9561;
wire n_9562;
wire n_9563;
wire n_9564;
wire n_9565;
wire n_9567;
wire n_9568;
wire n_9569;
wire n_957;
wire n_9570;
wire n_9571;
wire n_9572;
wire n_9573;
wire n_9575;
wire n_9576;
wire n_9578;
wire n_9579;
wire n_9580;
wire n_9582;
wire n_9583;
wire n_9584;
wire n_9585;
wire n_9586;
wire n_9588;
wire n_9589;
wire n_959;
wire n_9590;
wire n_9591;
wire n_9592;
wire n_9593;
wire n_9594;
wire n_9596;
wire n_9598;
wire n_960;
wire n_9600;
wire n_9602;
wire n_9604;
wire n_9605;
wire n_9607;
wire n_9608;
wire n_961;
wire n_9610;
wire n_9612;
wire n_9613;
wire n_9615;
wire n_9617;
wire n_9619;
wire n_9621;
wire n_9622;
wire n_9623;
wire n_9624;
wire n_9625;
wire n_9626;
wire n_9627;
wire n_9629;
wire n_963;
wire n_9631;
wire n_9633;
wire n_9635;
wire n_9637;
wire n_9639;
wire n_964;
wire n_9640;
wire n_9642;
wire n_9643;
wire n_9645;
wire n_9647;
wire n_9648;
wire n_9649;
wire n_965;
wire n_9651;
wire n_9653;
wire n_9655;
wire n_9657;
wire n_9658;
wire n_9659;
wire n_9660;
wire n_9661;
wire n_9662;
wire n_9663;
wire n_9665;
wire n_9666;
wire n_9667;
wire n_9668;
wire n_9669;
wire n_9670;
wire n_9671;
wire n_9673;
wire TIMEBOOST_net_13379;
wire n_9676;
wire n_9677;
wire n_9678;
wire n_9680;
wire n_9682;
wire n_9683;
wire n_9684;
wire n_9685;
wire n_9686;
wire n_9687;
wire n_9689;
wire n_969;
wire n_9690;
wire n_9691;
wire n_9692;
wire n_9693;
wire n_9694;
wire n_9696;
wire n_9697;
wire n_9698;
wire TIMEBOOST_net_13120;
wire n_9701;
wire n_9702;
wire n_9703;
wire n_9704;
wire n_9705;
wire n_9706;
wire n_9707;
wire n_9708;
wire n_9709;
wire n_971;
wire n_9710;
wire n_9711;
wire n_9712;
wire n_9713;
wire n_9714;
wire n_9715;
wire n_9716;
wire n_9717;
wire n_9718;
wire n_9719;
wire n_9720;
wire n_9721;
wire n_9722;
wire n_9723;
wire n_9724;
wire n_9725;
wire n_9726;
wire n_9727;
wire n_9728;
wire n_9729;
wire n_973;
wire n_9731;
wire n_9732;
wire n_9733;
wire n_9734;
wire n_9735;
wire n_9737;
wire n_9738;
wire n_9740;
wire n_9741;
wire n_9742;
wire n_9744;
wire n_9745;
wire n_9746;
wire n_9747;
wire n_9748;
wire TIMEBOOST_net_9382;
wire n_9750;
wire n_9751;
wire n_9752;
wire n_9753;
wire n_9754;
wire n_9756;
wire n_9757;
wire n_9759;
wire n_976;
wire n_9761;
wire TIMEBOOST_net_13106;
wire n_9765;
wire n_9767;
wire n_9768;
wire n_977;
wire n_9770;
wire n_9771;
wire n_9773;
wire n_9775;
wire n_9776;
wire n_9777;
wire n_9779;
wire n_978;
wire TIMEBOOST_net_13125;
wire n_9783;
wire n_9785;
wire n_9786;
wire n_9787;
wire n_9788;
wire n_9789;
wire n_9790;
wire n_9791;
wire n_9793;
wire n_9794;
wire n_9796;
wire n_9798;
wire n_980;
wire n_9800;
wire n_9802;
wire n_9804;
wire n_9805;
wire n_9807;
wire n_9808;
wire n_9810;
wire n_9811;
wire n_9813;
wire n_9814;
wire n_9816;
wire n_9818;
wire n_982;
wire n_9820;
wire n_9822;
wire n_9823;
wire n_9824;
wire n_9825;
wire n_9826;
wire n_9827;
wire n_9828;
wire n_9829;
wire n_983;
wire n_9830;
wire n_9831;
wire n_9832;
wire n_9833;
wire n_9834;
wire n_9835;
wire n_9836;
wire n_9837;
wire n_9838;
wire n_9839;
wire n_9840;
wire n_9841;
wire n_9842;
wire n_9843;
wire n_9844;
wire n_9845;
wire n_9846;
wire n_9847;
wire n_9848;
wire n_9849;
wire n_9850;
wire n_9851;
wire n_9852;
wire n_9853;
wire n_9854;
wire n_9855;
wire n_9856;
wire n_9857;
wire n_9858;
wire n_9859;
wire n_9860;
wire n_9861;
wire n_9862;
wire n_9863;
wire n_9864;
wire n_9865;
wire n_9866;
wire n_9867;
wire n_9868;
wire n_9869;
wire n_987;
wire n_9870;
wire n_9871;
wire n_9872;
wire n_9873;
wire n_9874;
wire n_9875;
wire n_9876;
wire n_9877;
wire n_9878;
wire n_9879;
wire n_988;
wire n_9880;
wire n_9881;
wire n_9882;
wire n_9883;
wire n_9884;
wire n_9885;
wire n_9886;
wire n_9887;
wire n_9888;
wire n_9889;
wire n_9890;
wire n_9891;
wire n_9892;
wire n_9893;
wire TIMEBOOST_net_13759;
wire n_9895;
wire n_9896;
wire n_9897;
wire n_9898;
wire n_9899;
wire n_990;
wire n_9901;
wire n_9902;
wire n_9903;
wire n_9904;
wire n_9906;
wire n_9908;
wire n_9910;
wire n_9912;
wire n_9914;
wire n_9916;
wire n_9918;
wire n_992;
wire n_9920;
wire n_9922;
wire n_9924;
wire n_9926;
wire n_9928;
wire n_993;
wire n_9931;
wire n_9932;
wire n_994;
wire n_9941;
wire n_9942;
wire n_9947;
wire n_9950;
wire n_9953;
wire n_9956;
wire n_996;
wire n_9962;
wire n_9968;
wire n_9971;
wire n_9975;
wire n_9976;
wire n_9979;
wire n_998;
wire n_9982;
wire n_9988;
wire n_999;
wire n_9991;
wire n_9992;
wire n_9993;
wire n_9997;
wire out_bckp_irdy_out;
wire out_bckp_perr_en_out;
wire output_backup_devsel_out_reg_Q;
wire output_backup_par_en_out_reg_Q;
wire output_backup_par_out_reg_Q;
wire output_backup_perr_out_reg_Q;
wire output_backup_serr_en_out_reg_Q;
wire output_backup_stop_out_reg_Q;
wire output_backup_tar_ad_en_out_reg_Q;
wire output_backup_trdy_out_reg_Q;
wire parchk_pci_ad_out_in;
wire parchk_pci_ad_out_in_1168;
wire parchk_pci_ad_out_in_1169;
wire parchk_pci_ad_out_in_1170;
wire parchk_pci_ad_out_in_1171;
wire parchk_pci_ad_out_in_1172;
wire parchk_pci_ad_out_in_1173;
wire parchk_pci_ad_out_in_1174;
wire parchk_pci_ad_out_in_1175;
wire parchk_pci_ad_out_in_1176;
wire parchk_pci_ad_out_in_1177;
wire parchk_pci_ad_out_in_1178;
wire parchk_pci_ad_out_in_1179;
wire parchk_pci_ad_out_in_1180;
wire parchk_pci_ad_out_in_1181;
wire parchk_pci_ad_out_in_1182;
wire parchk_pci_ad_out_in_1183;
wire parchk_pci_ad_out_in_1184;
wire parchk_pci_ad_out_in_1185;
wire parchk_pci_ad_out_in_1186;
wire parchk_pci_ad_out_in_1187;
wire parchk_pci_ad_out_in_1188;
wire parchk_pci_ad_out_in_1189;
wire parchk_pci_ad_out_in_1190;
wire parchk_pci_ad_out_in_1191;
wire parchk_pci_ad_out_in_1192;
wire parchk_pci_ad_out_in_1193;
wire parchk_pci_ad_out_in_1194;
wire parchk_pci_ad_out_in_1195;
wire parchk_pci_ad_out_in_1196;
wire parchk_pci_ad_out_in_1197;
wire parchk_pci_ad_out_in_1198;
wire parchk_pci_ad_reg_in;
wire parchk_pci_ad_reg_in_1205;
wire parchk_pci_ad_reg_in_1206;
wire parchk_pci_ad_reg_in_1207;
wire parchk_pci_ad_reg_in_1208;
wire parchk_pci_ad_reg_in_1209;
wire parchk_pci_ad_reg_in_1210;
wire parchk_pci_ad_reg_in_1211;
wire parchk_pci_ad_reg_in_1212;
wire parchk_pci_ad_reg_in_1213;
wire parchk_pci_ad_reg_in_1214;
wire parchk_pci_ad_reg_in_1215;
wire parchk_pci_ad_reg_in_1216;
wire parchk_pci_ad_reg_in_1217;
wire parchk_pci_ad_reg_in_1218;
wire parchk_pci_ad_reg_in_1219;
wire parchk_pci_ad_reg_in_1220;
wire parchk_pci_ad_reg_in_1221;
wire parchk_pci_ad_reg_in_1222;
wire parchk_pci_ad_reg_in_1223;
wire parchk_pci_ad_reg_in_1224;
wire parchk_pci_ad_reg_in_1225;
wire parchk_pci_ad_reg_in_1226;
wire parchk_pci_ad_reg_in_1227;
wire parchk_pci_ad_reg_in_1228;
wire parchk_pci_ad_reg_in_1229;
wire parchk_pci_ad_reg_in_1230;
wire parchk_pci_ad_reg_in_1231;
wire parchk_pci_ad_reg_in_1232;
wire parchk_pci_ad_reg_in_1233;
wire parchk_pci_ad_reg_in_1235;
wire parchk_pci_cbe_en_in;
wire parchk_pci_cbe_out_in;
wire parchk_pci_cbe_out_in_1202;
wire parchk_pci_cbe_out_in_1203;
wire parchk_pci_cbe_out_in_1204;
wire parchk_pci_cbe_reg_in;
wire parchk_pci_cbe_reg_in_1236;
wire parchk_pci_cbe_reg_in_1237;
wire parchk_pci_cbe_reg_in_1238;
wire parchk_pci_frame_en_in;
wire parchk_pci_frame_reg_in;
wire parchk_pci_irdy_en_in;
wire parchk_pci_par_en_in;
wire parchk_pci_perr_out_in;
wire parchk_pci_serr_en_in;
wire parchk_pci_serr_out_in;
wire parchk_pci_trdy_en_in;
wire parchk_pci_trdy_reg_in;
wire parity_checker_check_for_serr_on_second;
wire parity_checker_check_for_serr_on_second_reg_Q;
wire parity_checker_check_perr;
wire parity_checker_check_perr_reg_Q;
wire parity_checker_frame_and_irdy_en_prev;
wire parity_checker_frame_and_irdy_en_prev_prev;
wire parity_checker_frame_dec2;
wire parity_checker_master_perr_report;
wire parity_checker_master_perr_report_reg_Q;
wire parity_checker_pci_perr_en_reg;
wire parity_checker_perr_sampled;
wire pci_inti_conf_int_in;
wire pci_resi_conf_soft_res_in;
wire pci_target_unit_del_sync_addr_in;
wire pci_target_unit_del_sync_addr_in_204;
wire pci_target_unit_del_sync_addr_in_205;
wire pci_target_unit_del_sync_addr_in_206;
wire pci_target_unit_del_sync_addr_in_207;
wire pci_target_unit_del_sync_addr_in_208;
wire pci_target_unit_del_sync_addr_in_209;
wire pci_target_unit_del_sync_addr_in_210;
wire pci_target_unit_del_sync_addr_in_211;
wire pci_target_unit_del_sync_addr_in_212;
wire pci_target_unit_del_sync_addr_in_213;
wire pci_target_unit_del_sync_addr_in_214;
wire pci_target_unit_del_sync_addr_in_215;
wire pci_target_unit_del_sync_addr_in_216;
wire pci_target_unit_del_sync_addr_in_217;
wire pci_target_unit_del_sync_addr_in_218;
wire pci_target_unit_del_sync_addr_in_219;
wire pci_target_unit_del_sync_addr_in_220;
wire pci_target_unit_del_sync_addr_in_221;
wire pci_target_unit_del_sync_addr_in_222;
wire pci_target_unit_del_sync_addr_in_223;
wire pci_target_unit_del_sync_addr_in_224;
wire pci_target_unit_del_sync_addr_in_225;
wire pci_target_unit_del_sync_addr_in_226;
wire pci_target_unit_del_sync_addr_in_227;
wire pci_target_unit_del_sync_addr_in_228;
wire pci_target_unit_del_sync_addr_in_229;
wire pci_target_unit_del_sync_addr_in_230;
wire pci_target_unit_del_sync_addr_in_231;
wire pci_target_unit_del_sync_addr_in_232;
wire pci_target_unit_del_sync_addr_in_233;
wire pci_target_unit_del_sync_addr_in_234;
wire pci_target_unit_del_sync_bc_in;
wire pci_target_unit_del_sync_bc_in_201;
wire pci_target_unit_del_sync_bc_in_202;
wire pci_target_unit_del_sync_bc_in_203;
wire pci_target_unit_del_sync_be_out_reg_0__Q;
wire pci_target_unit_del_sync_be_out_reg_1__Q;
wire pci_target_unit_del_sync_be_out_reg_2__Q;
wire pci_target_unit_del_sync_be_out_reg_3__Q;
wire pci_target_unit_del_sync_comp_cycle_count_0_;
wire pci_target_unit_del_sync_comp_cycle_count_10_;
wire pci_target_unit_del_sync_comp_cycle_count_11_;
wire pci_target_unit_del_sync_comp_cycle_count_12_;
wire pci_target_unit_del_sync_comp_cycle_count_13_;
wire pci_target_unit_del_sync_comp_cycle_count_14_;
wire pci_target_unit_del_sync_comp_cycle_count_15_;
wire pci_target_unit_del_sync_comp_cycle_count_1_;
wire pci_target_unit_del_sync_comp_cycle_count_2_;
wire pci_target_unit_del_sync_comp_cycle_count_3_;
wire pci_target_unit_del_sync_comp_cycle_count_4_;
wire pci_target_unit_del_sync_comp_cycle_count_5_;
wire pci_target_unit_del_sync_comp_cycle_count_6_;
wire pci_target_unit_del_sync_comp_cycle_count_7_;
wire pci_target_unit_del_sync_comp_cycle_count_8_;
wire pci_target_unit_del_sync_comp_cycle_count_9_;
wire pci_target_unit_del_sync_comp_cycle_count_reg_16__Q;
wire pci_target_unit_del_sync_comp_done_reg_clr;
wire pci_target_unit_del_sync_comp_done_reg_clr_reg_Q;
wire pci_target_unit_del_sync_comp_done_reg_main;
wire pci_target_unit_del_sync_comp_done_reg_main_reg_Q;
wire pci_target_unit_del_sync_comp_flush_out_reg_Q;
wire pci_target_unit_del_sync_comp_in;
wire pci_target_unit_del_sync_comp_rty_exp_clr;
wire pci_target_unit_del_sync_comp_rty_exp_clr_reg_Q;
wire pci_target_unit_del_sync_comp_rty_exp_reg;
wire pci_target_unit_del_sync_req_comp_pending;
wire pci_target_unit_del_sync_req_comp_pending_sample;
wire pci_target_unit_del_sync_req_comp_pending_sample_reg_Q;
wire pci_target_unit_del_sync_req_done_reg;
wire pci_target_unit_del_sync_req_rty_exp_clr;
wire pci_target_unit_del_sync_req_rty_exp_clr_reg_Q;
wire pci_target_unit_del_sync_req_rty_exp_reg;
wire pci_target_unit_del_sync_req_sync_sync_data_out_reg_0__Q;
wire pci_target_unit_del_sync_sync_comp_done;
wire pci_target_unit_del_sync_sync_comp_req_pending;
wire pci_target_unit_del_sync_sync_comp_rty_exp_clr;
wire pci_target_unit_del_sync_sync_req_comp_pending;
wire pci_target_unit_del_sync_sync_req_rty_exp;
wire pci_target_unit_fifos_inGreyCount_0_;
wire pci_target_unit_fifos_inGreyCount_reg_0__Q;
wire pci_target_unit_fifos_inGreyCount_reg_1__Q;
wire pci_target_unit_fifos_outGreyCount_0_;
wire pci_target_unit_fifos_outGreyCount_reg_0__Q;
wire pci_target_unit_fifos_outGreyCount_reg_1__Q;
wire pci_target_unit_fifos_pcir_control_in_192;
wire pci_target_unit_fifos_pcir_data_in;
wire pci_target_unit_fifos_pcir_data_in_158;
wire pci_target_unit_fifos_pcir_data_in_159;
wire pci_target_unit_fifos_pcir_data_in_160;
wire pci_target_unit_fifos_pcir_data_in_161;
wire pci_target_unit_fifos_pcir_data_in_162;
wire pci_target_unit_fifos_pcir_data_in_163;
wire pci_target_unit_fifos_pcir_data_in_164;
wire pci_target_unit_fifos_pcir_data_in_165;
wire pci_target_unit_fifos_pcir_data_in_166;
wire pci_target_unit_fifos_pcir_data_in_167;
wire pci_target_unit_fifos_pcir_data_in_168;
wire pci_target_unit_fifos_pcir_data_in_169;
wire pci_target_unit_fifos_pcir_data_in_170;
wire pci_target_unit_fifos_pcir_data_in_171;
wire pci_target_unit_fifos_pcir_data_in_172;
wire pci_target_unit_fifos_pcir_data_in_173;
wire pci_target_unit_fifos_pcir_data_in_174;
wire pci_target_unit_fifos_pcir_data_in_175;
wire pci_target_unit_fifos_pcir_data_in_176;
wire pci_target_unit_fifos_pcir_data_in_177;
wire pci_target_unit_fifos_pcir_data_in_178;
wire pci_target_unit_fifos_pcir_data_in_179;
wire pci_target_unit_fifos_pcir_data_in_180;
wire pci_target_unit_fifos_pcir_data_in_181;
wire pci_target_unit_fifos_pcir_data_in_182;
wire pci_target_unit_fifos_pcir_data_in_183;
wire pci_target_unit_fifos_pcir_data_in_184;
wire pci_target_unit_fifos_pcir_data_in_185;
wire pci_target_unit_fifos_pcir_data_in_186;
wire pci_target_unit_fifos_pcir_data_in_187;
wire pci_target_unit_fifos_pcir_data_in_188;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_1_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_2__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_1__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_39;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_40;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_0_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_1_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_2_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_0__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_1__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_2__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_0__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_1__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_2__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_0_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_1_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_2_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_100;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_101;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__Q;
wire pci_target_unit_fifos_pcir_flush_in;
wire pci_target_unit_fifos_pcir_wenable_in;
wire pci_target_unit_fifos_pcir_whole_waddr;
wire pci_target_unit_fifos_pcir_whole_waddr_94;
wire pci_target_unit_fifos_pciw_addr_data_in;
wire pci_target_unit_fifos_pciw_addr_data_in_121;
wire pci_target_unit_fifos_pciw_addr_data_in_122;
wire pci_target_unit_fifos_pciw_addr_data_in_123;
wire pci_target_unit_fifos_pciw_addr_data_in_124;
wire pci_target_unit_fifos_pciw_addr_data_in_125;
wire pci_target_unit_fifos_pciw_addr_data_in_126;
wire pci_target_unit_fifos_pciw_addr_data_in_127;
wire pci_target_unit_fifos_pciw_addr_data_in_128;
wire pci_target_unit_fifos_pciw_addr_data_in_129;
wire pci_target_unit_fifos_pciw_addr_data_in_130;
wire pci_target_unit_fifos_pciw_addr_data_in_131;
wire pci_target_unit_fifos_pciw_addr_data_in_132;
wire pci_target_unit_fifos_pciw_addr_data_in_133;
wire pci_target_unit_fifos_pciw_addr_data_in_134;
wire pci_target_unit_fifos_pciw_addr_data_in_135;
wire pci_target_unit_fifos_pciw_addr_data_in_136;
wire pci_target_unit_fifos_pciw_addr_data_in_137;
wire pci_target_unit_fifos_pciw_addr_data_in_138;
wire pci_target_unit_fifos_pciw_addr_data_in_139;
wire pci_target_unit_fifos_pciw_addr_data_in_140;
wire pci_target_unit_fifos_pciw_addr_data_in_141;
wire pci_target_unit_fifos_pciw_addr_data_in_142;
wire pci_target_unit_fifos_pciw_addr_data_in_143;
wire pci_target_unit_fifos_pciw_addr_data_in_144;
wire pci_target_unit_fifos_pciw_addr_data_in_145;
wire pci_target_unit_fifos_pciw_addr_data_in_146;
wire pci_target_unit_fifos_pciw_addr_data_in_147;
wire pci_target_unit_fifos_pciw_addr_data_in_148;
wire pci_target_unit_fifos_pciw_addr_data_in_149;
wire pci_target_unit_fifos_pciw_addr_data_in_150;
wire pci_target_unit_fifos_pciw_addr_data_in_151;
wire pci_target_unit_fifos_pciw_cbe_in;
wire pci_target_unit_fifos_pciw_cbe_in_152;
wire pci_target_unit_fifos_pciw_cbe_in_153;
wire pci_target_unit_fifos_pciw_cbe_in_154;
wire pci_target_unit_fifos_pciw_control_in;
wire pci_target_unit_fifos_pciw_control_in_155;
wire pci_target_unit_fifos_pciw_control_in_156;
wire pci_target_unit_fifos_pciw_control_in_157;
wire pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_74;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_75;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_0__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_1__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_2__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_0__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_1__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_2__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus2;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_94;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_95;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_2_;
wire pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_0__153;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_1__192;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_2__231;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_3__270;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__Q;
wire pci_target_unit_fifos_pciw_inTransactionCount_0_;
wire pci_target_unit_fifos_pciw_inTransactionCount_1_;
wire pci_target_unit_fifos_pciw_inTransactionCount_reg_1__Q;
wire pci_target_unit_fifos_pciw_outTransactionCount_1_;
wire pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q;
wire pci_target_unit_fifos_pciw_outTransactionCount_reg_1__Q;
wire pci_target_unit_fifos_pciw_wenable_in;
wire pci_target_unit_fifos_pciw_whole_waddr;
wire pci_target_unit_fifos_pciw_whole_waddr_47;
wire pci_target_unit_fifos_wb_clk_inGreyCount_0_;
wire pci_target_unit_fifos_wb_clk_inGreyCount_1_;
wire pci_target_unit_fifos_wb_clk_sync_inGreyCount;
wire pci_target_unit_fifos_wb_clk_sync_inGreyCount_36;
wire pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg_Q;
wire pci_target_unit_pci_target_if_keep_desconnect_wo_data_set;
wire pci_target_unit_pci_target_if_norm_address_reg_0__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_1__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_2__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_3__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_4__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_5__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_6__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_7__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_8__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_9__Q;
wire pci_target_unit_pci_target_if_norm_prf_en;
wire pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_77;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_0__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_10__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_11__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_12__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_13__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_14__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_15__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_16__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_17__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_18__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_19__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_1__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_20__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_21__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_22__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_23__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_24__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_25__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_26__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_27__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_28__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_29__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_2__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_30__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_31__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_3__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_4__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_5__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_6__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_7__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_8__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_9__Q;
wire pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_0__Q;
wire pci_target_unit_pci_target_if_same_read_reg;
wire pci_target_unit_pci_target_if_target_rd_completed;
wire pci_target_unit_pci_target_sm_backoff;
wire pci_target_unit_pci_target_sm_bckp_trdy_reg_reg_Q;
wire pci_target_unit_pci_target_sm_cnf_progress;
wire pci_target_unit_pci_target_sm_master_will_request_read;
wire pci_target_unit_pci_target_sm_n_2;
wire pci_target_unit_pci_target_sm_n_3;
wire pci_target_unit_pci_target_sm_previous_frame;
wire pci_target_unit_pci_target_sm_rd_from_fifo;
wire pci_target_unit_pci_target_sm_rd_progress;
wire pci_target_unit_pci_target_sm_rd_request;
wire pci_target_unit_pci_target_sm_rd_request_reg_Q;
wire pci_target_unit_pci_target_sm_read_completed_reg;
wire pci_target_unit_pci_target_sm_read_completed_reg_reg_Q;
wire pci_target_unit_pci_target_sm_same_read_reg;
wire pci_target_unit_pci_target_sm_state_backoff_reg_reg_Q;
wire pci_target_unit_pci_target_sm_state_transfere_reg;
wire pci_target_unit_pci_target_sm_state_transfere_reg_reg_Q;
wire pci_target_unit_pci_target_sm_wr_progress;
wire pci_target_unit_pci_target_sm_wr_to_fifo;
wire pci_target_unit_pcit_if_comp_flush_in;
wire pci_target_unit_pcit_if_pcir_fifo_control_in_637;
wire pci_target_unit_pcit_if_pcir_fifo_data_in;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_766;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_767;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_768;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_769;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_770;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_771;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_772;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_773;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_774;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_775;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_776;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_777;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_778;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_779;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_780;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_781;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_782;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_783;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_784;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_785;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_786;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_787;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_788;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_789;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_790;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_791;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_792;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_793;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_794;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_795;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_796;
wire pci_target_unit_pcit_if_req_req_pending_in;
wire pci_target_unit_pcit_if_strd_addr_in;
wire pci_target_unit_pcit_if_strd_addr_in_686;
wire pci_target_unit_pcit_if_strd_addr_in_687;
wire pci_target_unit_pcit_if_strd_addr_in_688;
wire pci_target_unit_pcit_if_strd_addr_in_689;
wire pci_target_unit_pcit_if_strd_addr_in_690;
wire pci_target_unit_pcit_if_strd_addr_in_691;
wire pci_target_unit_pcit_if_strd_addr_in_692;
wire pci_target_unit_pcit_if_strd_addr_in_693;
wire pci_target_unit_pcit_if_strd_addr_in_694;
wire pci_target_unit_pcit_if_strd_addr_in_695;
wire pci_target_unit_pcit_if_strd_addr_in_696;
wire pci_target_unit_pcit_if_strd_addr_in_697;
wire pci_target_unit_pcit_if_strd_addr_in_698;
wire pci_target_unit_pcit_if_strd_addr_in_699;
wire pci_target_unit_pcit_if_strd_addr_in_700;
wire pci_target_unit_pcit_if_strd_addr_in_701;
wire pci_target_unit_pcit_if_strd_addr_in_702;
wire pci_target_unit_pcit_if_strd_addr_in_703;
wire pci_target_unit_pcit_if_strd_addr_in_704;
wire pci_target_unit_pcit_if_strd_addr_in_705;
wire pci_target_unit_pcit_if_strd_addr_in_706;
wire pci_target_unit_pcit_if_strd_addr_in_707;
wire pci_target_unit_pcit_if_strd_addr_in_708;
wire pci_target_unit_pcit_if_strd_addr_in_709;
wire pci_target_unit_pcit_if_strd_addr_in_710;
wire pci_target_unit_pcit_if_strd_addr_in_711;
wire pci_target_unit_pcit_if_strd_addr_in_712;
wire pci_target_unit_pcit_if_strd_addr_in_713;
wire pci_target_unit_pcit_if_strd_addr_in_714;
wire pci_target_unit_pcit_if_strd_addr_in_715;
wire pci_target_unit_pcit_if_strd_addr_in_716;
wire pci_target_unit_pcit_if_strd_bc_in;
wire pci_target_unit_pcit_if_strd_bc_in_717;
wire pci_target_unit_pcit_if_strd_bc_in_718;
wire pci_target_unit_pcit_if_strd_bc_in_719;
wire pci_target_unit_wbm_sm_pci_tar_burst_ok;
wire pci_target_unit_wbm_sm_pci_tar_read_request;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_50;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_51;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_52;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_53;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_54;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_55;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_56;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_57;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_58;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_59;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_60;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_61;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_62;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_63;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_64;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_65;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_66;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_67;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_68;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_69;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_70;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_71;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_72;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_73;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_74;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_75;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_76;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_77;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_78;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_79;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_80;
wire pci_target_unit_wbm_sm_pciw_fifo_cbe_in;
wire pci_target_unit_wbm_sm_pciw_fifo_cbe_in_81;
wire pci_target_unit_wbm_sm_pciw_fifo_cbe_in_82;
wire pci_target_unit_wbm_sm_pciw_fifo_cbe_in_83;
wire pci_target_unit_wbm_sm_pciw_fifo_control_in;
wire pci_target_unit_wbm_sm_pciw_fifo_control_in_84;
wire pci_target_unit_wbm_sm_pciw_fifo_control_in_85;
wire pci_target_unit_wbm_sm_pciw_fifo_control_in_86;
wire pci_target_unit_wishbone_master_addr_into_cnt_reg;
wire pci_target_unit_wishbone_master_bc_register_reg_0__Q;
wire pci_target_unit_wishbone_master_bc_register_reg_1__Q;
wire pci_target_unit_wishbone_master_bc_register_reg_2__Q;
wire pci_target_unit_wishbone_master_bc_register_reg_3__Q;
wire pci_target_unit_wishbone_master_burst_chopped;
wire pci_target_unit_wishbone_master_burst_chopped_delayed;
wire pci_target_unit_wishbone_master_burst_chopped_delayed_reg_Q;
wire pci_target_unit_wishbone_master_c_state_0_;
wire pci_target_unit_wishbone_master_c_state_1_;
wire pci_target_unit_wishbone_master_c_state_2_;
wire pci_target_unit_wishbone_master_first_data_is_burst_reg;
wire pci_target_unit_wishbone_master_first_wb_data_access;
wire pci_target_unit_wishbone_master_read_bound;
wire pci_target_unit_wishbone_master_read_count_0_;
wire pci_target_unit_wishbone_master_read_count_1_;
wire pci_target_unit_wishbone_master_read_count_reg_2__Q;
wire pci_target_unit_wishbone_master_reset_rty_cnt;
wire pci_target_unit_wishbone_master_reset_rty_cnt_reg_Q;
wire pci_target_unit_wishbone_master_retried;
wire pci_target_unit_wishbone_master_rty_counter_0_;
wire pci_target_unit_wishbone_master_rty_counter_1_;
wire pci_target_unit_wishbone_master_rty_counter_3_;
wire pci_target_unit_wishbone_master_rty_counter_4_;
wire pci_target_unit_wishbone_master_rty_counter_5_;
wire pci_target_unit_wishbone_master_rty_counter_6_;
wire pci_target_unit_wishbone_master_rty_counter_7_;
wire pci_target_unit_wishbone_master_wb_cyc_o_reg_Q;
wire pciu_am1_in;
wire pciu_am1_in_518;
wire pciu_am1_in_519;
wire pciu_am1_in_520;
wire pciu_am1_in_521;
wire pciu_am1_in_522;
wire pciu_am1_in_523;
wire pciu_am1_in_524;
wire pciu_am1_in_525;
wire pciu_am1_in_526;
wire pciu_am1_in_527;
wire pciu_am1_in_528;
wire pciu_am1_in_529;
wire pciu_am1_in_530;
wire pciu_am1_in_531;
wire pciu_am1_in_532;
wire pciu_am1_in_533;
wire pciu_am1_in_534;
wire pciu_am1_in_535;
wire pciu_am1_in_536;
wire pciu_am1_in_537;
wire pciu_am1_in_538;
wire pciu_am1_in_539;
wire pciu_am1_in_540;
wire pciu_bar0_in;
wire pciu_bar0_in_361;
wire pciu_bar0_in_362;
wire pciu_bar0_in_363;
wire pciu_bar0_in_364;
wire pciu_bar0_in_365;
wire pciu_bar0_in_366;
wire pciu_bar0_in_367;
wire pciu_bar0_in_368;
wire pciu_bar0_in_369;
wire pciu_bar0_in_370;
wire pciu_bar0_in_371;
wire pciu_bar0_in_372;
wire pciu_bar0_in_373;
wire pciu_bar0_in_374;
wire pciu_bar0_in_375;
wire pciu_bar0_in_376;
wire pciu_bar0_in_377;
wire pciu_bar0_in_378;
wire pciu_bar0_in_379;
wire pciu_bar1_in;
wire pciu_bar1_in_380;
wire pciu_bar1_in_381;
wire pciu_bar1_in_382;
wire pciu_bar1_in_383;
wire pciu_bar1_in_384;
wire pciu_bar1_in_385;
wire pciu_bar1_in_386;
wire pciu_bar1_in_387;
wire pciu_bar1_in_388;
wire pciu_bar1_in_389;
wire pciu_bar1_in_390;
wire pciu_bar1_in_391;
wire pciu_bar1_in_392;
wire pciu_bar1_in_393;
wire pciu_bar1_in_394;
wire pciu_bar1_in_395;
wire pciu_bar1_in_396;
wire pciu_bar1_in_397;
wire pciu_bar1_in_398;
wire pciu_bar1_in_399;
wire pciu_bar1_in_400;
wire pciu_bar1_in_401;
wire pciu_bar1_in_402;
wire pciu_cache_line_size_in_775;
wire pciu_cache_line_size_in_776;
wire pciu_cache_line_size_in_777;
wire pciu_cache_lsize_not_zero_in;
wire pciu_pciif_bckp_stop_in;
wire pciu_pciif_idsel_reg_in;
wire pciu_pciif_stop_reg_in;
wire pciu_pref_en_in_320;
wire wbm_cyc_o_1378;
wire wbs_ack_o_1307;
wire wbs_err_o_1309;
wire wbs_rty_o_1308;
wire wbs_wbb3_2_wbb2_dat_o_i;
wire wbs_wbb3_2_wbb2_dat_o_i_100;
wire wbs_wbb3_2_wbb2_dat_o_i_101;
wire wbs_wbb3_2_wbb2_dat_o_i_102;
wire wbs_wbb3_2_wbb2_dat_o_i_103;
wire wbs_wbb3_2_wbb2_dat_o_i_104;
wire wbs_wbb3_2_wbb2_dat_o_i_105;
wire wbs_wbb3_2_wbb2_dat_o_i_106;
wire wbs_wbb3_2_wbb2_dat_o_i_107;
wire wbs_wbb3_2_wbb2_dat_o_i_108;
wire wbs_wbb3_2_wbb2_dat_o_i_109;
wire wbs_wbb3_2_wbb2_dat_o_i_110;
wire wbs_wbb3_2_wbb2_dat_o_i_111;
wire wbs_wbb3_2_wbb2_dat_o_i_112;
wire wbs_wbb3_2_wbb2_dat_o_i_113;
wire wbs_wbb3_2_wbb2_dat_o_i_114;
wire wbs_wbb3_2_wbb2_dat_o_i_115;
wire wbs_wbb3_2_wbb2_dat_o_i_116;
wire wbs_wbb3_2_wbb2_dat_o_i_117;
wire wbs_wbb3_2_wbb2_dat_o_i_118;
wire wbs_wbb3_2_wbb2_dat_o_i_119;
wire wbs_wbb3_2_wbb2_dat_o_i_120;
wire wbs_wbb3_2_wbb2_dat_o_i_121;
wire wbs_wbb3_2_wbb2_dat_o_i_122;
wire wbs_wbb3_2_wbb2_dat_o_i_123;
wire wbs_wbb3_2_wbb2_dat_o_i_124;
wire wbs_wbb3_2_wbb2_dat_o_i_125;
wire wbs_wbb3_2_wbb2_dat_o_i_126;
wire wbs_wbb3_2_wbb2_dat_o_i_127;
wire wbs_wbb3_2_wbb2_dat_o_i_128;
wire wbs_wbb3_2_wbb2_dat_o_i_129;
wire wbs_wbb3_2_wbb2_dat_o_i_130;
wire wbu_addr_in;
wire wbu_addr_in_250;
wire wbu_addr_in_251;
wire wbu_addr_in_252;
wire wbu_addr_in_253;
wire wbu_addr_in_254;
wire wbu_addr_in_255;
wire wbu_addr_in_256;
wire wbu_addr_in_257;
wire wbu_addr_in_258;
wire wbu_addr_in_259;
wire wbu_addr_in_260;
wire wbu_addr_in_261;
wire wbu_addr_in_262;
wire wbu_addr_in_263;
wire wbu_addr_in_264;
wire wbu_addr_in_265;
wire wbu_addr_in_266;
wire wbu_addr_in_267;
wire wbu_addr_in_268;
wire wbu_addr_in_269;
wire wbu_addr_in_270;
wire wbu_addr_in_271;
wire wbu_addr_in_272;
wire wbu_addr_in_273;
wire wbu_addr_in_274;
wire wbu_addr_in_275;
wire wbu_addr_in_276;
wire wbu_addr_in_277;
wire wbu_addr_in_278;
wire wbu_addr_in_279;
wire wbu_addr_in_280;
wire wbu_am1_in;
wire wbu_am2_in;
wire wbu_bar1_in;
wire wbu_bar2_in;
wire wbu_cache_line_size_in_206;
wire wbu_cache_line_size_in_207;
wire wbu_cache_line_size_in_208;
wire wbu_cache_line_size_in_209;
wire wbu_cache_line_size_in_210;
wire wbu_cache_line_size_in_211;
wire wbu_latency_tim_val_in;
wire wbu_latency_tim_val_in_243;
wire wbu_latency_tim_val_in_244;
wire wbu_latency_tim_val_in_245;
wire wbu_latency_tim_val_in_246;
wire wbu_latency_tim_val_in_247;
wire wbu_latency_tim_val_in_248;
wire wbu_latency_tim_val_in_249;
wire wbu_map_in_131;
wire wbu_map_in_132;
wire wbu_mrl_en_in_141;
wire wbu_mrl_en_in_142;
wire wbu_pci_drcomp_pending_in;
wire wbu_pciif_devsel_reg_in;
wire wbu_pciif_frame_out_in;
wire wbu_pref_en_in_136;
wire wbu_pref_en_in_137;
wire wbu_sel_in;
wire wbu_sel_in_312;
wire wbu_sel_in_313;
wire wbu_sel_in_314;
wire wbu_wb_init_complete_in;
wire wbu_we_in;
wire wishbone_slave_unit_del_sync_addr_out_reg_0__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_10__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_11__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_12__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_13__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_14__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_15__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_16__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_17__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_18__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_19__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_1__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_20__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_21__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_22__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_23__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_24__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_25__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_26__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_27__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_28__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_29__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_2__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_30__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_31__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_3__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_4__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_5__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_6__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_7__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_8__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_9__Q;
wire wishbone_slave_unit_del_sync_bc_out_reg_0__Q;
wire wishbone_slave_unit_del_sync_bc_out_reg_1__Q;
wire wishbone_slave_unit_del_sync_bc_out_reg_2__Q;
wire wishbone_slave_unit_del_sync_bc_out_reg_3__Q;
wire wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_0_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_10_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_11_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_12_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_1_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_2_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_3_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_4_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_5_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_6_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_7_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_8_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_9_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_10__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_11__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_12__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_8__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_9__Q;
wire wishbone_slave_unit_del_sync_comp_done_reg_clr;
wire wishbone_slave_unit_del_sync_comp_done_reg_clr_reg_Q;
wire wishbone_slave_unit_del_sync_comp_done_reg_main;
wire wishbone_slave_unit_del_sync_comp_flush_out;
wire wishbone_slave_unit_del_sync_comp_req_pending_reg_Q;
wire wishbone_slave_unit_del_sync_comp_rty_exp_clr;
wire wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg_Q;
wire wishbone_slave_unit_del_sync_comp_rty_exp_reg;
wire wishbone_slave_unit_del_sync_req_comp_pending;
wire wishbone_slave_unit_del_sync_req_comp_pending_sample;
wire wishbone_slave_unit_del_sync_req_comp_pending_sample_reg_Q;
wire wishbone_slave_unit_del_sync_req_done_reg;
wire wishbone_slave_unit_del_sync_req_done_reg_reg_Q;
wire wishbone_slave_unit_del_sync_req_rty_exp_clr;
wire wishbone_slave_unit_del_sync_req_rty_exp_clr_reg_Q;
wire wishbone_slave_unit_del_sync_req_rty_exp_reg;
wire wishbone_slave_unit_del_sync_sync_comp_done;
wire wishbone_slave_unit_del_sync_sync_comp_req_pending;
wire wishbone_slave_unit_del_sync_sync_comp_rty_exp_clr;
wire wishbone_slave_unit_del_sync_sync_req_comp_pending;
wire wishbone_slave_unit_del_sync_sync_req_rty_exp;
wire wishbone_slave_unit_del_sync_we_out_reg_Q;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_100;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_101;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_70;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_71;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_72;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_73;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_74;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_75;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_76;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_77;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_78;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_79;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_80;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_81;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_82;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_83;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_84;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_85;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_86;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_87;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_88;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_89;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_90;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_91;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_92;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_93;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_94;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_95;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_96;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_97;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_98;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_99;
wire wishbone_slave_unit_fifos_inGreyCount_0_;
wire wishbone_slave_unit_fifos_inGreyCount_reg_0__Q;
wire wishbone_slave_unit_fifos_inGreyCount_reg_1__Q;
wire wishbone_slave_unit_fifos_inGreyCount_reg_2__Q;
wire wishbone_slave_unit_fifos_outGreyCount_0_;
wire wishbone_slave_unit_fifos_outGreyCount_1_;
wire wishbone_slave_unit_fifos_outGreyCount_2_;
wire wishbone_slave_unit_fifos_pci_clk_inGreyCount_0_;
wire wishbone_slave_unit_fifos_pci_clk_inGreyCount_1_;
wire wishbone_slave_unit_fifos_pci_clk_inGreyCount_2_;
wire wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_2__Q;
wire wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount;
wire wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_49;
wire wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_50;
wire wishbone_slave_unit_fifos_wbr_be_in;
wire wishbone_slave_unit_fifos_wbr_be_in_264;
wire wishbone_slave_unit_fifos_wbr_be_in_265;
wire wishbone_slave_unit_fifos_wbr_be_in_266;
wire wishbone_slave_unit_fifos_wbr_control_in;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_0_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_1_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_1_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_3_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_45;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_46;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_47;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_0_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_1_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_2_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_3_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_0_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_1_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_2_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_3_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_0_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__43;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__46;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__47;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__51;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__56;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__59;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__62;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__67;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__70;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_11__466;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__484;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__487;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13_;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__509;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__522;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__531;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__532;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__536;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__544;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_14__583;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_15__622;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_2__6;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__177;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__178;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__183;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__236;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__237;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__238;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__243;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__247;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__248;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__249;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__258;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__260;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__265;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__271;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_7__310;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__330;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__342;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__358;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__359;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__360;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__363;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__365;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__374;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__376;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__377;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__379;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__380;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__9__Q;
wire wishbone_slave_unit_fifos_wbr_whole_waddr;
wire wishbone_slave_unit_fifos_wbr_whole_waddr_104;
wire wishbone_slave_unit_fifos_wbr_whole_waddr_105;
wire wishbone_slave_unit_fifos_wbr_whole_waddr_106;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_70;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_71;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_72;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus1;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_93;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_94;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_95;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_11__465;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_13__543;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_14__582;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_15__621;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_4__213;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_6__252;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__291;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__309;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__Q;
wire wishbone_slave_unit_fifos_wbw_inTransactionCount_0_;
wire wishbone_slave_unit_fifos_wbw_inTransactionCount_1_;
wire wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_0__Q;
wire wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_1__Q;
wire wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q;
wire wishbone_slave_unit_fifos_wbw_outTransactionCount_0_;
wire wishbone_slave_unit_fifos_wbw_outTransactionCount_1_;
wire wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_0__Q;
wire wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_1__Q;
wire wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q;
wire wishbone_slave_unit_fifos_wbw_whole_waddr;
wire wishbone_slave_unit_fifos_wbw_whole_waddr_55;
wire wishbone_slave_unit_fifos_wbw_whole_waddr_56;
wire wishbone_slave_unit_fifos_wbw_whole_waddr_57;
wire wishbone_slave_unit_pci_initiator_if_current_byte_address;
wire wishbone_slave_unit_pci_initiator_if_current_byte_address_36;
wire wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q;
wire wishbone_slave_unit_pci_initiator_if_data_source;
wire wishbone_slave_unit_pci_initiator_if_del_read_req;
wire wishbone_slave_unit_pci_initiator_if_del_write_req;
wire wishbone_slave_unit_pci_initiator_if_err_recovery;
wire wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__Q;
wire wishbone_slave_unit_pci_initiator_if_posted_write_req;
wire wishbone_slave_unit_pci_initiator_if_read_bound;
wire wishbone_slave_unit_pci_initiator_if_read_count_0_;
wire wishbone_slave_unit_pci_initiator_if_read_count_1_;
wire wishbone_slave_unit_pci_initiator_if_read_count_2_;
wire wishbone_slave_unit_pci_initiator_if_read_count_3_;
wire wishbone_slave_unit_pci_initiator_if_read_count_reg_3__Q;
wire wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg_Q;
wire wishbone_slave_unit_pci_initiator_if_write_req_int;
wire wishbone_slave_unit_pci_initiator_sm_cur_state_0_;
wire wishbone_slave_unit_pci_initiator_sm_cur_state_1_;
wire wishbone_slave_unit_pci_initiator_sm_cur_state_2_;
wire wishbone_slave_unit_pci_initiator_sm_cur_state_3_;
wire wishbone_slave_unit_pci_initiator_sm_decode_count_0_;
wire wishbone_slave_unit_pci_initiator_sm_decode_count_1_;
wire wishbone_slave_unit_pci_initiator_sm_decode_count_2_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_0_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_1_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_2_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_3_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_4_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_5_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_6_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_7_;
wire wishbone_slave_unit_pci_initiator_sm_mabort1;
wire wishbone_slave_unit_pci_initiator_sm_mabort2;
wire wishbone_slave_unit_pci_initiator_sm_rdata_selector;
wire wishbone_slave_unit_pci_initiator_sm_rdata_selector_14;
wire wishbone_slave_unit_pci_initiator_sm_timeout;
wire wishbone_slave_unit_pci_initiator_sm_transfer;
wire wishbone_slave_unit_pcim_if_del_bc_in;
wire wishbone_slave_unit_pcim_if_del_bc_in_382;
wire wishbone_slave_unit_pcim_if_del_bc_in_383;
wire wishbone_slave_unit_pcim_if_del_burst_in;
wire wishbone_slave_unit_pcim_if_del_req_in;
wire wishbone_slave_unit_pcim_if_del_we_in;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_384;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_385;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_386;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_387;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_388;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_389;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_390;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_391;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_392;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_393;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_394;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_395;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_396;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_397;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_398;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_399;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_400;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_401;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_402;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_403;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_404;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_405;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_406;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_407;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_408;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_409;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_410;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_411;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_412;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_413;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_414;
wire wishbone_slave_unit_pcim_if_wbw_cbe_in;
wire wishbone_slave_unit_pcim_if_wbw_cbe_in_416;
wire wishbone_slave_unit_pcim_if_wbw_cbe_in_417;
wire wishbone_slave_unit_pcim_sm_be_in_557;
wire wishbone_slave_unit_pcim_sm_be_in_558;
wire wishbone_slave_unit_pcim_sm_be_in_559;
wire wishbone_slave_unit_pcim_sm_data_in;
wire wishbone_slave_unit_pcim_sm_data_in_635;
wire wishbone_slave_unit_pcim_sm_data_in_636;
wire wishbone_slave_unit_pcim_sm_data_in_637;
wire wishbone_slave_unit_pcim_sm_data_in_638;
wire wishbone_slave_unit_pcim_sm_data_in_639;
wire wishbone_slave_unit_pcim_sm_data_in_640;
wire wishbone_slave_unit_pcim_sm_data_in_641;
wire wishbone_slave_unit_pcim_sm_data_in_642;
wire wishbone_slave_unit_pcim_sm_data_in_643;
wire wishbone_slave_unit_pcim_sm_data_in_644;
wire wishbone_slave_unit_pcim_sm_data_in_645;
wire wishbone_slave_unit_pcim_sm_data_in_646;
wire wishbone_slave_unit_pcim_sm_data_in_647;
wire wishbone_slave_unit_pcim_sm_data_in_648;
wire wishbone_slave_unit_pcim_sm_data_in_649;
wire wishbone_slave_unit_pcim_sm_data_in_650;
wire wishbone_slave_unit_pcim_sm_data_in_651;
wire wishbone_slave_unit_pcim_sm_data_in_652;
wire wishbone_slave_unit_pcim_sm_data_in_653;
wire wishbone_slave_unit_pcim_sm_data_in_654;
wire wishbone_slave_unit_pcim_sm_data_in_655;
wire wishbone_slave_unit_pcim_sm_data_in_656;
wire wishbone_slave_unit_pcim_sm_data_in_657;
wire wishbone_slave_unit_pcim_sm_data_in_658;
wire wishbone_slave_unit_pcim_sm_data_in_659;
wire wishbone_slave_unit_pcim_sm_data_in_660;
wire wishbone_slave_unit_pcim_sm_data_in_661;
wire wishbone_slave_unit_pcim_sm_data_in_662;
wire wishbone_slave_unit_pcim_sm_data_in_663;
wire wishbone_slave_unit_pcim_sm_data_in_664;
wire wishbone_slave_unit_pcim_sm_data_in_665;
wire wishbone_slave_unit_pcim_sm_last_in;
wire wishbone_slave_unit_pcim_sm_rdy_in;
wire wishbone_slave_unit_wbs_sm_del_req_pending_in;
wire wishbone_slave_unit_wbs_sm_wbr_control_in;
wire wishbone_slave_unit_wbs_sm_wbr_control_in_190;
wire wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg_Q;
wire wishbone_slave_unit_wishbone_slave_c_state;
wire wishbone_slave_unit_wishbone_slave_c_state_1;
wire wishbone_slave_unit_wishbone_slave_c_state_2;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_0__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_10__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_11__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_12__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_13__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_14__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_15__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_16__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_17__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_18__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_19__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_1__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_20__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_21__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_22__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_23__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_24__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_25__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_26__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_27__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_28__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_29__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_2__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_30__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_31__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_32__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_33__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_34__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_35__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_3__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_4__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_5__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_6__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_7__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_8__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_9__Q;
wire wishbone_slave_unit_wishbone_slave_del_addr_hit;
wire wishbone_slave_unit_wishbone_slave_del_completion_allow;
wire wishbone_slave_unit_wishbone_slave_do_del_request;
wire wishbone_slave_unit_wishbone_slave_img_hit_0_;
wire wishbone_slave_unit_wishbone_slave_img_hit_1_;
wire wishbone_slave_unit_wishbone_slave_img_hit_2_;
wire wishbone_slave_unit_wishbone_slave_img_hit_3_;
wire wishbone_slave_unit_wishbone_slave_img_hit_4_;
wire wishbone_slave_unit_wishbone_slave_img_wallow;
wire wishbone_slave_unit_wishbone_slave_map;
wire wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q;
wire wishbone_slave_unit_wishbone_slave_pref_en_reg_Q;
wire wishbone_slave_unit_wishbone_slave_wb_conf_hit;
wire wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg_Q;
wire TIMEBOOST_net_0;
wire TIMEBOOST_net_1;
wire TIMEBOOST_net_2;
wire TIMEBOOST_net_3;
wire TIMEBOOST_net_4;
wire TIMEBOOST_net_5;

// Start cells
in01f04 FE_OCPC1822_n_16560 ( .a(n_16560), .o(FE_OCPN1822_n_16560) );
in01f08 FE_OCPC1823_n_16560 ( .a(FE_OCPN1822_n_16560), .o(FE_OCPN1823_n_16560) );
in01f04 FE_OCPC1824_n_12030 ( .a(FE_OCP_RBN2284_FE_RN_494_0), .o(FE_OCPN1824_n_12030) );
in01f08 FE_OCPC1825_n_12030 ( .a(FE_OCPN1824_n_12030), .o(FE_OCPN1825_n_12030) );
in01f08 FE_OCPC1827_n_14995 ( .a(FE_OCP_RBN1922_n_10273), .o(FE_OCPN1827_n_14995) );
in01f01 FE_OCPC1831_n_16949 ( .a(n_16949), .o(FE_OCPN1831_n_16949) );
in01m02 FE_OCPC1832_n_16949 ( .a(FE_OCPN1831_n_16949), .o(FE_OCPN1832_n_16949) );
in01f02 FE_OCPC1833_n_11884 ( .a(n_11884), .o(FE_OCPN1833_n_11884) );
in01f04 FE_OCPC1834_n_11884 ( .a(FE_OCPN1833_n_11884), .o(FE_OCPN1834_n_11884) );
in01f01 FE_OCPC1835_n_16798 ( .a(n_16798), .o(FE_OCPN1835_n_16798) );
in01f04 FE_OCPC1836_n_16798 ( .a(FE_OCPN1835_n_16798), .o(FE_OCPN1836_n_16798) );
in01f01 FE_OCPC1837_n_1238 ( .a(n_1238), .o(FE_OCPN1837_n_1238) );
in01s02 FE_OCPC1838_n_1238 ( .a(FE_OCPN1837_n_1238), .o(FE_OCPN1838_n_1238) );
in01m02 FE_OCPC1839_n_1238 ( .a(FE_OCPN1837_n_1238), .o(FE_OCPN1839_n_1238) );
in01f01 FE_OCPC1840_n_16089 ( .a(n_16089), .o(FE_OCPN1840_n_16089) );
in01f04 FE_OCPC1841_n_16089 ( .a(FE_OCPN1840_n_16089), .o(FE_OCPN1841_n_16089) );
in01f08 FE_OCPC1842_n_16033 ( .a(n_16033), .o(FE_OCPN1842_n_16033) );
in01f08 FE_OCPC1843_n_16033 ( .a(FE_OCPN1842_n_16033), .o(FE_OCPN1843_n_16033) );
in01f02 FE_OCPC1844_n_16427 ( .a(n_16427), .o(FE_OCPN1844_n_16427) );
in01f03 FE_OCPC1845_n_16427 ( .a(FE_OCPN1844_n_16427), .o(TIMEBOOST_net_5) );
in01f01 FE_OCPC1846_n_14981 ( .a(n_14981), .o(FE_OCPN1846_n_14981) );
in01f06 FE_OCPC1847_n_14981 ( .a(FE_OCPN1846_n_14981), .o(FE_OCPN1847_n_14981) );
in01f08 FE_OCPC1848_n_15998 ( .a(n_15998), .o(FE_OCPN1848_n_15998) );
in01f02 FE_OCPC1849_n_15998 ( .a(FE_OCPN1848_n_15998), .o(FE_OCPN1849_n_15998) );
in01f06 FE_OCPC1850_n_15998 ( .a(FE_OCPN1848_n_15998), .o(FE_OCPN1850_n_15998) );
in01f10 FE_OCPC1851_n_16538 ( .a(n_16538), .o(FE_OCPN1851_n_16538) );
in01f10 FE_OCPC1852_n_16538 ( .a(FE_OCPN1851_n_16538), .o(FE_OCPN1852_n_16538) );
in01m10 FE_OCPC1853_n_2071 ( .a(n_2071), .o(FE_OCPN1853_n_2071) );
in01m08 FE_OCPC1854_n_2071 ( .a(FE_OCPN1853_n_2071), .o(FE_OCPN1854_n_2071) );
in01s01 FE_OCPC1855_n_2071 ( .a(FE_OCPN1853_n_2071), .o(FE_OCPN1855_n_2071) );
in01f03 FE_OCPC1856_FE_OFN1774_n_13800 ( .a(FE_OFN1774_n_13800), .o(FE_OCPN1856_FE_OFN1774_n_13800) );
in01f06 FE_OCPC1860_FE_OFN468_n_15534 ( .a(FE_OFN2137_n_15534), .o(FE_OCPN1860_FE_OFN468_n_15534) );
in01f08 FE_OCPC1861_FE_OFN468_n_15534 ( .a(FE_OCPN1860_FE_OFN468_n_15534), .o(FE_OCPN1861_FE_OFN468_n_15534) );
in01f02 FE_OCPC1862_FE_OFN474_n_16992 ( .a(FE_OFN2142_n_16992), .o(FE_OCPN1862_FE_OFN474_n_16992) );
in01f04 FE_OCPC1863_FE_OFN474_n_16992 ( .a(FE_OCPN1862_FE_OFN474_n_16992), .o(FE_OCPN1863_FE_OFN474_n_16992) );
in01f01 FE_OCPC1865_n_12377 ( .a(n_12381), .o(FE_OCPN1865_n_12377) );
in01f04 FE_OCPC1866_n_12377 ( .a(n_12381), .o(FE_OCPN1866_n_12377) );
in01f08 FE_OCPC1871_FE_OFN474_n_16992 ( .a(FE_OFN2142_n_16992), .o(FE_OCPN1871_FE_OFN474_n_16992) );
in01f04 FE_OCPC1872_FE_OFN474_n_16992 ( .a(FE_OCPN1871_FE_OFN474_n_16992), .o(FE_OCPN1872_FE_OFN474_n_16992) );
in01f08 FE_OCPC1873_FE_OFN474_n_16992 ( .a(FE_OCPN1871_FE_OFN474_n_16992), .o(FE_OCPN1873_FE_OFN474_n_16992) );
in01f03 FE_OCPC1875_n_14526 ( .a(n_16460), .o(FE_OCPN1875_n_14526) );
in01f06 FE_OCPC1876_n_13903 ( .a(n_13903), .o(FE_OCPN1876_n_13903) );
in01f06 FE_OCPC1877_n_13903 ( .a(FE_OCPN1876_n_13903), .o(FE_OCPN1877_n_13903) );
in01f04 FE_OCPC1878_FE_OFN470_n_10588 ( .a(FE_OFN2131_n_10588), .o(FE_OCPN1878_FE_OFN470_n_10588) );
in01f04 FE_OCPC1879_FE_OFN470_n_10588 ( .a(FE_OCPN1878_FE_OFN470_n_10588), .o(FE_OCPN1879_FE_OFN470_n_10588) );
in01f04 FE_OCPC1880_n_9991 ( .a(n_9991), .o(FE_OCPN1880_n_9991) );
in01f06 FE_OCPC1881_n_9991 ( .a(FE_OCPN1880_n_9991), .o(FE_OCPN1881_n_9991) );
in01f02 FE_OCPC1882_n_9991 ( .a(FE_OCPN1880_n_9991), .o(FE_OCPN1882_n_9991) );
in01f06 FE_OCPC1883_n_15566 ( .a(n_15566), .o(FE_OCPN1883_n_15566) );
in01f10 FE_OCPC1884_n_15566 ( .a(FE_OCPN1883_n_15566), .o(FE_OCPN1884_n_15566) );
in01f02 FE_OCPC1885_FE_OFN1508_n_15587 ( .a(FE_OFN1508_n_15587), .o(FE_OCPN1885_FE_OFN1508_n_15587) );
in01f04 FE_OCPC1886_FE_OFN1508_n_15587 ( .a(FE_OCPN1885_FE_OFN1508_n_15587), .o(FE_OCPN1886_FE_OFN1508_n_15587) );
in01f08 FE_OCPC1887_FE_OFN473_n_16992 ( .a(FE_OFN2139_n_16992), .o(FE_OCPN1887_FE_OFN473_n_16992) );
in01f08 FE_OCPC1888_FE_OFN473_n_16992 ( .a(FE_OCPN1887_FE_OFN473_n_16992), .o(FE_OCPN1888_FE_OFN473_n_16992) );
in01f01 FE_OCPC1889_n_16553 ( .a(n_16553), .o(FE_OCPN1889_n_16553) );
in01f02 FE_OCPC1890_n_16553 ( .a(FE_OCPN1889_n_16553), .o(FE_OCPN1890_n_16553) );
in01f04 FE_OCPC1891_FE_OFN1727_n_9975 ( .a(FE_OFN1727_n_9975), .o(FE_OCPN1891_FE_OFN1727_n_9975) );
in01f06 FE_OCPC1892_FE_OFN1727_n_9975 ( .a(FE_OCPN1891_FE_OFN1727_n_9975), .o(FE_OCPN1892_FE_OFN1727_n_9975) );
in01f04 FE_OCPC1895_FE_OFN1559_n_12042 ( .a(FE_OFN1559_n_12042), .o(FE_OCPN1895_FE_OFN1559_n_12042) );
in01f06 FE_OCPC1897_n_3231 ( .a(n_3231), .o(FE_OCPN1897_n_3231) );
in01f08 FE_OCPC1898_n_3231 ( .a(FE_OCPN1897_n_3231), .o(FE_OCPN1898_n_3231) );
in01f04 FE_OCPC1899_n_16810 ( .a(n_16810), .o(FE_OCPN1899_n_16810) );
in01f02 FE_OCPC1900_n_16810 ( .a(FE_OCPN1899_n_16810), .o(FE_OCPN1900_n_16810) );
in01f02 FE_OCPC1901_n_16810 ( .a(FE_OCPN1899_n_16810), .o(FE_OCPN1901_n_16810) );
in01f02 FE_OCPC1902_FE_OFN1061_n_16720 ( .a(FE_OFN1061_n_16720), .o(FE_OCPN1902_FE_OFN1061_n_16720) );
in01f02 FE_OCPC1903_FE_OFN1061_n_16720 ( .a(FE_OCPN1902_FE_OFN1061_n_16720), .o(FE_OCPN1903_FE_OFN1061_n_16720) );
in01f02 FE_OCPC1904_n_8927 ( .a(n_8927), .o(FE_OCPN1904_n_8927) );
in01f06 FE_OCPC1905_n_8927 ( .a(FE_OCPN1904_n_8927), .o(FE_OCPN1905_n_8927) );
in01f02 FE_OCPC1907_n_11767 ( .a(FE_OCP_RBN1970_n_11767), .o(FE_OCPN1907_n_11767) );
in01f08 FE_OCPC1908_n_16497 ( .a(FE_OFN2127_n_16497), .o(FE_OCPN1908_n_16497) );
in01f10 FE_OCPC1909_n_16497 ( .a(FE_OCPN1908_n_16497), .o(FE_OCPN1909_n_16497) );
in01f06 FE_OCPC1910_FE_OFN1152_n_13249 ( .a(FE_OFN1152_n_13249), .o(FE_OCPN1910_FE_OFN1152_n_13249) );
in01f08 FE_OCPC1911_FE_OFN1152_n_13249 ( .a(FE_OCPN1910_FE_OFN1152_n_13249), .o(FE_OCPN1911_FE_OFN1152_n_13249) );
in01f02 FE_OCPC1912_FE_OFN1150_n_13249 ( .a(FE_OFN1150_n_13249), .o(FE_OCPN1912_FE_OFN1150_n_13249) );
in01f02 FE_OCPC1913_FE_OFN1150_n_13249 ( .a(FE_OCPN1912_FE_OFN1150_n_13249), .o(FE_OCPN1913_FE_OFN1150_n_13249) );
in01f06 FE_OCPC1914_FE_OFN1522_n_10892 ( .a(FE_OFN1522_n_10892), .o(FE_OCPN1914_FE_OFN1522_n_10892) );
in01f08 FE_OCPC1915_FE_OFN1522_n_10892 ( .a(FE_OCPN1914_FE_OFN1522_n_10892), .o(FE_OCPN1915_FE_OFN1522_n_10892) );
in01f02 FE_OCPC2014_n_10195 ( .a(n_10195), .o(FE_OCPN2014_n_10195) );
in01f04 FE_OCPC2015_n_10195 ( .a(FE_OCPN2014_n_10195), .o(FE_OCPN2015_n_10195) );
in01f06 FE_OCPC2217_n_13997 ( .a(n_13997), .o(FE_OCPN2217_n_13997) );
in01f08 FE_OCPC2218_n_13997 ( .a(FE_OCPN2217_n_13997), .o(FE_OCPN2218_n_13997) );
in01f02 FE_OCPC2219_n_13997 ( .a(FE_OCPN2217_n_13997), .o(FE_OCPN2219_n_13997) );
in01f02 FE_OCPUNCOC1951_FE_OFN697_n_16760 ( .a(FE_OFN697_n_16760), .o(FE_OCPUNCON1951_FE_OFN697_n_16760) );
in01f08 FE_OCPUNCOC1952_FE_OFN697_n_16760 ( .a(FE_OCPUNCON1951_FE_OFN697_n_16760), .o(FE_OCPUNCON1952_FE_OFN697_n_16760) );
in01m06 FE_OCP_DRV_C1949_n_8660 ( .a(FE_OCP_DRV_N2262_n_8660), .o(FE_OCP_DRV_N1949_n_8660) );
in01f08 FE_OCP_DRV_C1950_n_8660 ( .a(FE_OCP_DRV_N1949_n_8660), .o(FE_OCP_DRV_N1950_n_8660) );
in01f02 FE_OCP_DRV_C2261_n_8660 ( .a(n_8660), .o(FE_OCP_DRV_N2261_n_8660) );
in01f04 FE_OCP_DRV_C2262_n_8660 ( .a(FE_OCP_DRV_N2261_n_8660), .o(FE_OCP_DRV_N2262_n_8660) );
in01s01 FE_OCP_RBC1917_wbs_cti_i_1_ ( .a(FE_OCP_RBN1918_wbs_cti_i_1_), .o(FE_OCP_RBN1917_wbs_cti_i_1_) );
in01f80 FE_OCP_RBC1918_wbs_cti_i_1_ ( .a(wbs_cti_i_1_), .o(FE_OCP_RBN1918_wbs_cti_i_1_) );
in01f02 FE_OCP_RBC1921_n_10273 ( .a(n_10273), .o(FE_OCP_RBN1921_n_10273) );
in01f06 FE_OCP_RBC1922_n_10273 ( .a(FE_OCP_RBN1921_n_10273), .o(FE_OCP_RBN1922_n_10273) );
in01f02 FE_OCP_RBC1923_n_10273 ( .a(FE_OCP_RBN1921_n_10273), .o(FE_OCP_RBN1923_n_10273) );
in01f01 FE_OCP_RBC1924_n_10273 ( .a(FE_OCP_RBN1923_n_10273), .o(FE_OCP_RBN1924_n_10273) );
in01f02 FE_OCP_RBC1925_n_10259 ( .a(n_10259), .o(FE_OCP_RBN1925_n_10259) );
in01f02 FE_OCP_RBC1926_n_10259 ( .a(FE_OCP_RBN1925_n_10259), .o(FE_OCP_RBN1926_n_10259) );
in01f02 FE_OCP_RBC1927_n_10259 ( .a(FE_OCP_RBN1925_n_10259), .o(FE_OCP_RBN1927_n_10259) );
in01f04 FE_OCP_RBC1928_n_10259 ( .a(FE_OCP_RBN1925_n_10259), .o(FE_OCP_RBN1928_n_10259) );
in01f10 FE_OCP_RBC1929_parchk_pci_trdy_reg_in ( .a(parchk_pci_trdy_reg_in), .o(FE_OCP_RBN1929_parchk_pci_trdy_reg_in) );
in01f08 FE_OCP_RBC1930_parchk_pci_trdy_reg_in ( .a(FE_OCP_RBN1929_parchk_pci_trdy_reg_in), .o(FE_OCP_RBN1930_parchk_pci_trdy_reg_in) );
in01f04 FE_OCP_RBC1932_FE_OFN1515_n_10538 ( .a(FE_OCP_RBN1966_FE_RN_459_0), .o(FE_OCP_RBN1932_FE_OFN1515_n_10538) );
in01f02 FE_OCP_RBC1933_FE_OFN1515_n_10538 ( .a(FE_OCP_RBN1966_FE_RN_459_0), .o(FE_OCP_RBN1933_FE_OFN1515_n_10538) );
in01f02 FE_OCP_RBC1934_FE_OFN1515_n_10538 ( .a(FE_OCP_RBN1966_FE_RN_459_0), .o(FE_OCP_RBN1934_FE_OFN1515_n_10538) );
in01f02 FE_OCP_RBC1954_FE_RN_462_0 ( .a(FE_RN_462_0), .o(FE_OCP_RBN1954_FE_RN_462_0) );
in01f02 FE_OCP_RBC1955_n_16981 ( .a(n_16981), .o(FE_OCP_RBN1955_n_16981) );
in01f04 FE_OCP_RBC1956_n_16981 ( .a(n_16981), .o(FE_OCP_RBN1956_n_16981) );
in01f02 FE_OCP_RBC1961_FE_OFN1591_n_13741 ( .a(FE_OFN1591_n_13741), .o(FE_OCP_RBN1961_FE_OFN1591_n_13741) );
in01f02 FE_OCP_RBC1962_FE_OFN1591_n_13741 ( .a(FE_OFN1591_n_13741), .o(FE_OCP_RBN1962_FE_OFN1591_n_13741) );
in01f02 FE_OCP_RBC1963_FE_OFN1591_n_13741 ( .a(FE_OFN1591_n_13741), .o(FE_OCP_RBN1963_FE_OFN1591_n_13741) );
in01f04 FE_OCP_RBC1964_FE_OFN1591_n_13741 ( .a(FE_OCP_RBN1963_FE_OFN1591_n_13741), .o(FE_OCP_RBN1964_FE_OFN1591_n_13741) );
in01f02 FE_OCP_RBC1965_FE_RN_459_0 ( .a(FE_RN_459_0), .o(FE_OCP_RBN1965_FE_RN_459_0) );
in01f02 FE_OCP_RBC1966_FE_RN_459_0 ( .a(FE_OCP_RBN1965_FE_RN_459_0), .o(FE_OCP_RBN1966_FE_RN_459_0) );
in01f04 FE_OCP_RBC1967_FE_RN_459_0 ( .a(FE_OCP_RBN1965_FE_RN_459_0), .o(FE_OCP_RBN1967_FE_RN_459_0) );
in01f06 FE_OCP_RBC1968_FE_OFN1532_n_10143 ( .a(FE_OFN1532_n_10143), .o(FE_OCP_RBN1968_FE_OFN1532_n_10143) );
in01f06 FE_OCP_RBC1969_FE_OFN1532_n_10143 ( .a(FE_OFN1532_n_10143), .o(FE_OCP_RBN1969_FE_OFN1532_n_10143) );
in01f02 FE_OCP_RBC1970_n_11767 ( .a(n_11767), .o(FE_OCP_RBN1970_n_11767) );
in01f02 FE_OCP_RBC1971_n_11767 ( .a(FE_OCP_RBN1970_n_11767), .o(FE_OCP_RBN1971_n_11767) );
in01f02 FE_OCP_RBC1972_n_11767 ( .a(FE_OCP_RBN1970_n_11767), .o(FE_OCP_RBN1972_n_11767) );
in01f06 FE_OCP_RBC1973_n_12381 ( .a(n_12381), .o(FE_OCP_RBN1973_n_12381) );
in01f01 FE_OCP_RBC1974_n_12381 ( .a(n_12381), .o(FE_OCP_RBN1974_n_12381) );
in01f01 FE_OCP_RBC1975_n_12381 ( .a(n_12381), .o(FE_OCP_RBN1975_n_12381) );
in01f04 FE_OCP_RBC1976_n_12381 ( .a(n_12381), .o(FE_OCP_RBN1976_n_12381) );
in01f01 FE_OCP_RBC1977_n_10273 ( .a(FE_OCP_RBN1922_n_10273), .o(FE_OCP_RBN1977_n_10273) );
in01f01 FE_OCP_RBC1978_n_10273 ( .a(FE_OCP_RBN1922_n_10273), .o(FE_OCP_RBN1978_n_10273) );
in01f04 FE_OCP_RBC1979_n_10273 ( .a(FE_OCP_RBN1922_n_10273), .o(FE_OCP_RBN1979_n_10273) );
in01f02 FE_OCP_RBC1980_n_10273 ( .a(FE_OCP_RBN1922_n_10273), .o(FE_OCP_RBN1980_n_10273) );
in01f01 FE_OCP_RBC1981_FE_OFN1591_n_13741 ( .a(FE_OCP_RBN1964_FE_OFN1591_n_13741), .o(FE_OCP_RBN1981_FE_OFN1591_n_13741) );
in01f01 FE_OCP_RBC1983_FE_OFN1591_n_13741 ( .a(FE_OCP_RBN1964_FE_OFN1591_n_13741), .o(FE_OCP_RBN1983_FE_OFN1591_n_13741) );
in01f02 FE_OCP_RBC1984_FE_OFN1591_n_13741 ( .a(FE_OCP_RBN1964_FE_OFN1591_n_13741), .o(FE_OCP_RBN1984_FE_OFN1591_n_13741) );
in01f04 FE_OCP_RBC1985_FE_OFN1591_n_13741 ( .a(FE_OCP_RBN1964_FE_OFN1591_n_13741), .o(FE_OCP_RBN1985_FE_OFN1591_n_13741) );
in01f08 FE_OCP_RBC1994_n_13971 ( .a(n_13971), .o(FE_OCP_RBN1994_n_13971) );
in01f04 FE_OCP_RBC1995_n_13971 ( .a(FE_OCP_RBN1994_n_13971), .o(FE_OCP_RBN1995_n_13971) );
in01f04 FE_OCP_RBC1996_n_13971 ( .a(FE_OCP_RBN1994_n_13971), .o(FE_OCP_RBN1996_n_13971) );
in01f08 FE_OCP_RBC1997_n_13971 ( .a(FE_OCP_RBN1994_n_13971), .o(FE_OCP_RBN1997_n_13971) );
in01f04 FE_OCP_RBC1998_n_13971 ( .a(FE_OCP_RBN1994_n_13971), .o(FE_OCP_RBN1998_n_13971) );
in01f02 FE_OCP_RBC1999_n_13971 ( .a(FE_OCP_RBN1994_n_13971), .o(FE_OCP_RBN1999_n_13971) );
in01m02 FE_OCP_RBC2000_n_1403 ( .a(n_1403), .o(FE_OCP_RBN2000_n_1403) );
in01f02 FE_OCP_RBC2003_FE_OFN1026_n_16760 ( .a(FE_OFN1026_n_16760), .o(FE_OCP_RBN2003_FE_OFN1026_n_16760) );
in01f01 FE_OCP_RBC2004_FE_OFN1026_n_16760 ( .a(FE_OFN1026_n_16760), .o(FE_OCP_RBN2004_FE_OFN1026_n_16760) );
in01f06 FE_OCP_RBC2005_FE_RN_459_0 ( .a(FE_OCP_RBN1967_FE_RN_459_0), .o(FE_OCP_RBN2005_FE_RN_459_0) );
in01f04 FE_OCP_RBC2006_FE_RN_459_0 ( .a(FE_OCP_RBN1967_FE_RN_459_0), .o(FE_OCP_RBN2006_FE_RN_459_0) );
in01f01 FE_OCP_RBC2007_n_16698 ( .a(n_16698), .o(FE_OCP_RBN2007_n_16698) );
in01f06 FE_OCP_RBC2008_n_16698 ( .a(n_16698), .o(FE_OCP_RBN2008_n_16698) );
in01f06 FE_OCP_RBC2009_n_16698 ( .a(FE_OCP_RBN2008_n_16698), .o(FE_OCP_RBN2009_n_16698) );
in01f06 FE_OCP_RBC2010_n_16698 ( .a(FE_OCP_RBN2008_n_16698), .o(FE_OCP_RBN2010_n_16698) );
in01f06 FE_OCP_RBC2011_n_16698 ( .a(FE_OCP_RBN2008_n_16698), .o(FE_OCP_RBN2011_n_16698) );
in01f04 FE_OCP_RBC2012_n_16698 ( .a(FE_OCP_RBN2008_n_16698), .o(FE_OCP_RBN2012_n_16698) );
in01f04 FE_OCP_RBC2013_FE_OCPN1895_FE_OFN1559_n_12042 ( .a(FE_OCPN1895_FE_OFN1559_n_12042), .o(FE_OCP_RBN2013_FE_OCPN1895_FE_OFN1559_n_12042) );
in01f04 FE_OCP_RBC2016_n_16970 ( .a(n_16970), .o(FE_OCP_RBN2016_n_16970) );
in01f01 FE_OCP_RBC2017_n_16970 ( .a(n_16970), .o(FE_OCP_RBN2017_n_16970) );
in01f02 FE_OCP_RBC2018_n_16970 ( .a(n_16970), .o(FE_OCP_RBN2018_n_16970) );
in01f01 FE_OCP_RBC2019_n_16970 ( .a(n_16970), .o(FE_OCP_RBN2019_n_16970) );
in01f01 FE_OCP_RBC2220_n_15347 ( .a(n_15347), .o(FE_OCP_RBN2220_n_15347) );
in01f02 FE_OCP_RBC2221_n_15347 ( .a(n_15347), .o(FE_OCP_RBN2221_n_15347) );
in01f03 FE_OCP_RBC2222_n_15347 ( .a(n_15347), .o(FE_OCP_RBN2222_n_15347) );
in01f06 FE_OCP_RBC2223_n_15347 ( .a(n_15347), .o(FE_OCP_RBN2223_n_15347) );
in01f02 FE_OCP_RBC2224_n_16322 ( .a(n_16322), .o(FE_OCP_RBN2224_n_16322) );
in01f03 FE_OCP_RBC2225_n_16322 ( .a(n_16322), .o(FE_OCP_RBN2225_n_16322) );
in01f02 FE_OCP_RBC2226_g75174_p ( .a(g75174_p), .o(FE_OCP_RBN2226_g75174_p) );
in01f02 FE_OCP_RBC2227_g75174_p ( .a(g75174_p), .o(FE_OCP_RBN2227_g75174_p) );
in01f02 FE_OCP_RBC2228_n_15969 ( .a(n_15969), .o(FE_OCP_RBN2228_n_15969) );
in01f04 FE_OCP_RBC2229_n_15969 ( .a(FE_OCP_RBN2228_n_15969), .o(FE_OCP_RBN2229_n_15969) );
in01f04 FE_OCP_RBC2231_FE_RN_390_0 ( .a(FE_RN_390_0), .o(FE_OCP_RBN2231_FE_RN_390_0) );
in01f02 FE_OCP_RBC2232_n_16273 ( .a(n_16273), .o(FE_OCP_RBN2232_n_16273) );
in01f02 FE_OCP_RBC2233_n_16273 ( .a(n_16273), .o(FE_OCP_RBN2233_n_16273) );
in01f01 FE_OCP_RBC2237_g74749_p ( .a(g74749_p), .o(FE_OCP_RBN2237_g74749_p) );
in01f04 FE_OCP_RBC2238_g74749_p ( .a(g74749_p), .o(FE_OCP_RBN2238_g74749_p) );
in01f02 FE_OCP_RBC2239_g74749_p ( .a(g74749_p), .o(FE_OCP_RBN2239_g74749_p) );
in01s01 FE_OCP_RBC2265_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_ ( .a(FE_OCP_RBN2269_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_), .o(FE_OCP_RBN2265_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_) );
in01f80 FE_OCP_RBC2269_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_ ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_), .o(FE_OCP_RBN2269_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_) );
in01f10 FE_OCP_RBC2270_g75061_p ( .a(g75061_p), .o(FE_OCP_RBN2270_g75061_p) );
in01f04 FE_OCP_RBC2271_g75061_p ( .a(g75061_p), .o(FE_OCP_RBN2271_g75061_p) );
in01f01 FE_OCP_RBC2272_n_10268 ( .a(n_10268), .o(FE_OCP_RBN2272_n_10268) );
in01f02 FE_OCP_RBC2273_n_10268 ( .a(n_10268), .o(FE_OCP_RBN2273_n_10268) );
in01f04 FE_OCP_RBC2274_n_10268 ( .a(FE_OCP_RBN2273_n_10268), .o(FE_OCP_RBN2274_n_10268) );
in01f02 FE_OCP_RBC2275_n_10268 ( .a(FE_OCP_RBN2273_n_10268), .o(FE_OCP_RBN2275_n_10268) );
in01f20 FE_OCP_RBC2277_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_ ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_), .o(FE_OCP_RBN2277_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_) );
in01f02 FE_OCP_RBC2278_n_16974 ( .a(n_16974), .o(FE_OCP_RBN2278_n_16974) );
in01f01 FE_OCP_RBC2279_n_16974 ( .a(n_16974), .o(FE_OCP_RBN2279_n_16974) );
in01f02 FE_OCP_RBC2280_g74996_p ( .a(g74996_p), .o(FE_OCP_RBN2280_g74996_p) );
in01f02 FE_OCP_RBC2281_g74996_p ( .a(g74996_p), .o(FE_OCP_RBN2281_g74996_p) );
in01f02 FE_OCP_RBC2282_g74996_p ( .a(g74996_p), .o(FE_OCP_RBN2282_g74996_p) );
in01f02 FE_OCP_RBC2283_g74996_p ( .a(g74996_p), .o(FE_OCP_RBN2283_g74996_p) );
in01f02 FE_OCP_RBC2284_FE_RN_494_0 ( .a(FE_RN_494_0), .o(FE_OCP_RBN2284_FE_RN_494_0) );
in01f04 FE_OCP_RBC2285_FE_RN_494_0 ( .a(FE_RN_494_0), .o(FE_OCP_RBN2285_FE_RN_494_0) );
in01f08 FE_OCP_RBC2286_FE_RN_494_0 ( .a(FE_OCP_RBN2285_FE_RN_494_0), .o(FE_OCP_RBN2286_FE_RN_494_0) );
in01s01 FE_OCP_RBC2289_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_ ( .a(FE_OCP_RBN2290_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .o(FE_OCP_RBN2289_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_) );
in01f20 FE_OCP_RBC2290_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_ ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .o(FE_OCP_RBN2290_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_) );
in01f06 FE_OCP_RBC2291_FE_OFN1575_n_12028 ( .a(FE_OFN1575_n_12028), .o(FE_OCP_RBN2291_FE_OFN1575_n_12028) );
in01f06 FE_OCP_RBC2292_FE_OFN1575_n_12028 ( .a(FE_OFN1575_n_12028), .o(FE_OCP_RBN2292_FE_OFN1575_n_12028) );
in01f04 FE_OCP_RBC2293_FE_OFN1581_n_12306 ( .a(FE_OFN1581_n_12306), .o(FE_OCP_RBN2293_FE_OFN1581_n_12306) );
in01m08 FE_OFC1001_n_15978 ( .a(FE_OFN997_n_15978), .o(FE_OFN1001_n_15978) );
in01s04 FE_OFC1002_n_2047 ( .a(n_2047), .o(FE_OFN1002_n_2047) );
in01s06 FE_OFC1003_n_2047 ( .a(FE_OFN1002_n_2047), .o(FE_OFN1003_n_2047) );
in01f06 FE_OFC1004_n_16288 ( .a(n_16288), .o(FE_OFN1004_n_16288) );
in01f08 FE_OFC1005_n_16288 ( .a(FE_OFN1004_n_16288), .o(FE_OFN1005_n_16288) );
in01f10 FE_OFC1006_n_16288 ( .a(FE_OFN1004_n_16288), .o(FE_OFN1006_n_16288) );
in01s01 FE_OFC1007_n_4734 ( .a(n_4734), .o(FE_OFN1007_n_4734) );
in01s03 FE_OFC1008_n_4734 ( .a(n_4734), .o(FE_OFN1008_n_4734) );
in01s02 FE_OFC1009_n_4734 ( .a(n_4734), .o(FE_OFN1009_n_4734) );
in01s03 FE_OFC1010_n_4734 ( .a(FE_OFN1008_n_4734), .o(FE_OFN1010_n_4734) );
in01s06 FE_OFC1011_n_4734 ( .a(FE_OFN1008_n_4734), .o(FE_OFN1011_n_4734) );
in01s03 FE_OFC1012_n_4734 ( .a(FE_OFN1009_n_4734), .o(FE_OFN1012_n_4734) );
in01s03 FE_OFC1013_n_4734 ( .a(FE_OFN1009_n_4734), .o(FE_OFN1013_n_4734) );
in01s06 FE_OFC1014_n_2053 ( .a(n_2053), .o(FE_OFN1014_n_2053) );
in01s03 FE_OFC1015_n_2053 ( .a(FE_OFN1014_n_2053), .o(FE_OFN1015_n_2053) );
in01s08 FE_OFC1016_n_2053 ( .a(FE_OFN1014_n_2053), .o(FE_OFN1016_n_2053) );
in01s03 FE_OFC1017_n_2053 ( .a(FE_OFN1014_n_2053), .o(FE_OFN1017_n_2053) );
in01m06 FE_OFC1018_n_11877 ( .a(n_11877), .o(FE_OFN1018_n_11877) );
in01m02 FE_OFC1019_n_11877 ( .a(n_11877), .o(FE_OFN1019_n_11877) );
in01m04 FE_OFC1020_n_11877 ( .a(n_11877), .o(FE_OFN1020_n_11877) );
in01m08 FE_OFC1021_n_11877 ( .a(FE_OFN1018_n_11877), .o(FE_OFN1021_n_11877) );
in01m08 FE_OFC1022_n_11877 ( .a(FE_OFN1018_n_11877), .o(FE_OFN1022_n_11877) );
in01m04 FE_OFC1023_n_11877 ( .a(FE_OFN1019_n_11877), .o(FE_OFN1023_n_11877) );
in01m02 FE_OFC1024_n_11877 ( .a(FE_OFN1019_n_11877), .o(FE_OFN1024_n_11877) );
in01m06 FE_OFC1025_n_11877 ( .a(FE_OFN1020_n_11877), .o(FE_OFN1025_n_11877) );
in01m02 FE_OFC1028_n_4732 ( .a(n_4732), .o(FE_OFN1028_n_4732) );
in01s02 FE_OFC1029_n_4732 ( .a(n_4732), .o(FE_OFN1029_n_4732) );
in01s02 FE_OFC1030_n_4732 ( .a(n_4732), .o(FE_OFN1030_n_4732) );
in01s03 FE_OFC1031_n_4732 ( .a(FE_OFN1028_n_4732), .o(FE_OFN1031_n_4732) );
in01s03 FE_OFC1032_n_4732 ( .a(FE_OFN1029_n_4732), .o(FE_OFN1032_n_4732) );
in01s03 FE_OFC1033_n_4732 ( .a(FE_OFN1030_n_4732), .o(FE_OFN1033_n_4732) );
in01s03 FE_OFC1034_n_4732 ( .a(FE_OFN1030_n_4732), .o(FE_OFN1034_n_4732) );
in01s01 FE_OFC1035_n_4732 ( .a(FE_OFN1028_n_4732), .o(FE_OFN1035_n_4732) );
in01s02 FE_OFC1036_n_4732 ( .a(FE_OFN1028_n_4732), .o(FE_OFN1036_n_4732) );
in01s03 FE_OFC1037_n_4732 ( .a(FE_OFN1029_n_4732), .o(FE_OFN1037_n_4732) );
in01s03 FE_OFC1038_n_2037 ( .a(n_2037), .o(FE_OFN1038_n_2037) );
in01s01 FE_OFC1039_n_2037 ( .a(n_2037), .o(FE_OFN1039_n_2037) );
in01s01 FE_OFC1040_n_2037 ( .a(n_2037), .o(FE_OFN1040_n_2037) );
in01s06 FE_OFC1041_n_2037 ( .a(FE_OFN1038_n_2037), .o(FE_OFN1041_n_2037) );
in01s06 FE_OFC1042_n_2037 ( .a(FE_OFN1038_n_2037), .o(FE_OFN1042_n_2037) );
in01s06 FE_OFC1043_n_2037 ( .a(FE_OFN1039_n_2037), .o(FE_OFN1043_n_2037) );
in01s06 FE_OFC1044_n_2037 ( .a(FE_OFN1040_n_2037), .o(FE_OFN1044_n_2037) );
in01s03 FE_OFC1045_n_16657 ( .a(n_16657), .o(FE_OFN1045_n_16657) );
in01s08 FE_OFC1046_n_16657 ( .a(FE_OFN1045_n_16657), .o(FE_OFN1046_n_16657) );
in01s04 FE_OFC1047_n_16657 ( .a(n_16657), .o(FE_OFN1047_n_16657) );
in01s03 FE_OFC1048_n_16657 ( .a(n_16657), .o(FE_OFN1048_n_16657) );
in01s06 FE_OFC1049_n_16657 ( .a(FE_OFN1048_n_16657), .o(FE_OFN1049_n_16657) );
in01s02 FE_OFC1050_n_16657 ( .a(FE_OFN1047_n_16657), .o(FE_OFN1050_n_16657) );
in01s08 FE_OFC1051_n_16657 ( .a(FE_OFN1047_n_16657), .o(FE_OFN1051_n_16657) );
in01s02 FE_OFC1052_n_4727 ( .a(n_4727), .o(FE_OFN1052_n_4727) );
in01s03 FE_OFC1053_n_4727 ( .a(n_4727), .o(FE_OFN1053_n_4727) );
in01m02 FE_OFC1054_n_4727 ( .a(n_4727), .o(FE_OFN1054_n_4727) );
in01s06 FE_OFC1055_n_4727 ( .a(FE_OFN1053_n_4727), .o(FE_OFN1055_n_4727) );
in01s06 FE_OFC1056_n_4727 ( .a(FE_OFN1053_n_4727), .o(FE_OFN1056_n_4727) );
in01s03 FE_OFC1057_n_4727 ( .a(FE_OFN1054_n_4727), .o(FE_OFN1057_n_4727) );
in01s01 FE_OFC1058_n_4727 ( .a(FE_OFN1054_n_4727), .o(FE_OFN1058_n_4727) );
in01s02 FE_OFC1059_n_4727 ( .a(FE_OFN1054_n_4727), .o(FE_OFN1059_n_4727) );
in01f02 FE_OFC1061_n_16720 ( .a(FE_OFN1060_n_16720), .o(TIMEBOOST_net_3) );
in01f06 FE_OFC1062_n_15808 ( .a(n_15808), .o(FE_OFN1062_n_15808) );
in01f10 FE_OFC1063_n_15808 ( .a(FE_OFN1062_n_15808), .o(FE_OFN1063_n_15808) );
in01f06 FE_OFC1064_n_15808 ( .a(n_15808), .o(FE_OFN1064_n_15808) );
in01f04 FE_OFC1065_n_15808 ( .a(FE_OFN1064_n_15808), .o(FE_OFN1065_n_15808) );
in01f06 FE_OFC1066_n_15808 ( .a(FE_OFN1064_n_15808), .o(FE_OFN1066_n_15808) );
in01f08 FE_OFC1067_n_15729 ( .a(n_15729), .o(FE_OFN1067_n_15729) );
in01f06 FE_OFC1068_n_15729 ( .a(FE_OFN1067_n_15729), .o(FE_OFN1068_n_15729) );
in01f08 FE_OFC1069_n_15729 ( .a(FE_OFN1067_n_15729), .o(FE_OFN1069_n_15729) );
in01f06 FE_OFC1070_n_15729 ( .a(FE_OFN1067_n_15729), .o(FE_OFN1070_n_15729) );
in01f04 FE_OFC1071_n_15729 ( .a(FE_OFN1067_n_15729), .o(FE_OFN1071_n_15729) );
in01s01 FE_OFC1072_n_4740 ( .a(n_4740), .o(FE_OFN1072_n_4740) );
in01s04 FE_OFC1073_n_4740 ( .a(n_4740), .o(FE_OFN1073_n_4740) );
in01s04 FE_OFC1074_n_4740 ( .a(FE_OFN1073_n_4740), .o(FE_OFN1074_n_4740) );
in01s04 FE_OFC1075_n_4740 ( .a(FE_OFN1073_n_4740), .o(FE_OFN1075_n_4740) );
in01s04 FE_OFC1076_n_4740 ( .a(FE_OFN1073_n_4740), .o(FE_OFN1076_n_4740) );
in01s04 FE_OFC1077_n_4740 ( .a(FE_OFN1073_n_4740), .o(FE_OFN1077_n_4740) );
in01m02 FE_OFC1078_n_4778 ( .a(n_4778), .o(FE_OFN1078_n_4778) );
in01s08 FE_OFC1079_n_4778 ( .a(FE_OFN1078_n_4778), .o(FE_OFN1079_n_4778) );
in01f04 FE_OFC1080_n_13221 ( .a(n_13221), .o(FE_OFN1080_n_13221) );
in01f08 FE_OFC1081_n_13221 ( .a(n_13221), .o(FE_OFN1081_n_13221) );
in01f06 FE_OFC1082_n_13221 ( .a(FE_OFN1080_n_13221), .o(FE_OFN1082_n_13221) );
in01f04 FE_OFC1083_n_13221 ( .a(FE_OFN1080_n_13221), .o(FE_OFN1083_n_13221) );
in01m08 FE_OFC1084_n_13221 ( .a(FE_OFN1081_n_13221), .o(FE_OFN1084_n_13221) );
in01f08 FE_OFC1085_n_13221 ( .a(FE_OFN1081_n_13221), .o(FE_OFN1085_n_13221) );
in01m01 FE_OFC1086_g64577_p ( .a(g64577_p), .o(FE_OFN1086_g64577_p) );
in01f06 FE_OFC1087_g64577_p ( .a(g64577_p), .o(FE_OFN1087_g64577_p) );
in01f02 FE_OFC1088_g64577_p ( .a(g64577_p), .o(FE_OFN1088_g64577_p) );
in01f02 FE_OFC1089_g64577_p ( .a(g64577_p), .o(FE_OFN1089_g64577_p) );
in01s02 FE_OFC1090_g64577_p ( .a(FE_OFN1086_g64577_p), .o(FE_OFN1090_g64577_p) );
in01m04 FE_OFC1091_g64577_p ( .a(FE_OFN1087_g64577_p), .o(FE_OFN1091_g64577_p) );
in01m08 FE_OFC1092_g64577_p ( .a(FE_OFN1087_g64577_p), .o(FE_OFN1092_g64577_p) );
in01m02 FE_OFC1093_g64577_p ( .a(FE_OFN1087_g64577_p), .o(FE_OFN1093_g64577_p) );
in01s01 FE_OFC1094_g64577_p ( .a(FE_OFN1087_g64577_p), .o(TIMEBOOST_net_1) );
in01m02 FE_OFC1095_g64577_p ( .a(FE_OFN1089_g64577_p), .o(FE_OFN1095_g64577_p) );
in01s02 FE_OFC1096_g64577_p ( .a(FE_OFN1089_g64577_p), .o(FE_OFN1096_g64577_p) );
in01m06 FE_OFC1097_g64577_p ( .a(FE_OFN1089_g64577_p), .o(FE_OFN1097_g64577_p) );
in01s02 FE_OFC1098_g64577_p ( .a(FE_OFN1090_g64577_p), .o(FE_OFN1098_g64577_p) );
in01s02 FE_OFC1099_g64577_p ( .a(FE_OFN1090_g64577_p), .o(FE_OFN1099_g64577_p) );
in01s02 FE_OFC1100_g64577_p ( .a(FE_OFN1088_g64577_p), .o(FE_OFN1100_g64577_p) );
in01s06 FE_OFC1101_g64577_p ( .a(FE_OFN1091_g64577_p), .o(FE_OFN1101_g64577_p) );
in01m06 FE_OFC1102_g64577_p ( .a(FE_OFN1091_g64577_p), .o(FE_OFN1102_g64577_p) );
in01s02 FE_OFC1103_g64577_p ( .a(FE_OFN1088_g64577_p), .o(FE_OFN1103_g64577_p) );
in01m03 FE_OFC1104_g64577_p ( .a(FE_OFN1088_g64577_p), .o(FE_OFN1104_g64577_p) );
in01s10 FE_OFC1105_g64577_p ( .a(FE_OFN1092_g64577_p), .o(FE_OFN1105_g64577_p) );
in01m08 FE_OFC1106_g64577_p ( .a(FE_OFN1088_g64577_p), .o(FE_OFN1106_g64577_p) );
in01s02 FE_OFC1107_g64577_p ( .a(FE_OFN1088_g64577_p), .o(FE_OFN1107_g64577_p) );
in01s06 FE_OFC1108_g64577_p ( .a(FE_OFN1096_g64577_p), .o(FE_OFN1108_g64577_p) );
in01s08 FE_OFC1109_g64577_p ( .a(FE_OFN1097_g64577_p), .o(FE_OFN1109_g64577_p) );
in01m06 FE_OFC1110_g64577_p ( .a(FE_OFN1093_g64577_p), .o(FE_OFN1110_g64577_p) );
in01s02 FE_OFC1111_g64577_p ( .a(FE_OFN1093_g64577_p), .o(FE_OFN1111_g64577_p) );
in01s06 FE_OFC1112_g64577_p ( .a(FE_OFN1102_g64577_p), .o(FE_OFN1112_g64577_p) );
in01s02 FE_OFC1113_g64577_p ( .a(FE_OFN1103_g64577_p), .o(FE_OFN1113_g64577_p) );
in01s02 FE_OFC1114_g64577_p ( .a(FE_OFN1103_g64577_p), .o(FE_OFN1114_g64577_p) );
in01s06 FE_OFC1115_g64577_p ( .a(FE_OFN1101_g64577_p), .o(FE_OFN1115_g64577_p) );
in01s06 FE_OFC1116_g64577_p ( .a(FE_OFN1102_g64577_p), .o(FE_OFN1116_g64577_p) );
in01s10 FE_OFC1117_g64577_p ( .a(FE_OFN1105_g64577_p), .o(FE_OFN1117_g64577_p) );
in01s06 FE_OFC1118_g64577_p ( .a(FE_OFN1108_g64577_p), .o(FE_OFN1118_g64577_p) );
in01s08 FE_OFC1119_g64577_p ( .a(FE_OFN1109_g64577_p), .o(FE_OFN1119_g64577_p) );
in01s08 FE_OFC1120_g64577_p ( .a(FE_OFN1109_g64577_p), .o(FE_OFN1120_g64577_p) );
in01s06 FE_OFC1121_g64577_p ( .a(FE_OFN1101_g64577_p), .o(FE_OFN1121_g64577_p) );
in01s06 FE_OFC1122_g64577_p ( .a(FE_OFN1102_g64577_p), .o(FE_OFN1122_g64577_p) );
in01s06 FE_OFC1123_g64577_p ( .a(FE_OFN1102_g64577_p), .o(FE_OFN1123_g64577_p) );
in01s06 FE_OFC1124_g64577_p ( .a(FE_OFN1105_g64577_p), .o(FE_OFN1124_g64577_p) );
in01s10 FE_OFC1125_g64577_p ( .a(FE_OFN1105_g64577_p), .o(FE_OFN1125_g64577_p) );
in01s06 FE_OFC1126_g64577_p ( .a(FE_OFN1110_g64577_p), .o(FE_OFN1126_g64577_p) );
in01s02 FE_OFC1127_g64577_p ( .a(FE_OFN1111_g64577_p), .o(FE_OFN1127_g64577_p) );
in01s03 FE_OFC1128_g64577_p ( .a(FE_OFN1111_g64577_p), .o(FE_OFN1128_g64577_p) );
in01s06 FE_OFC1129_g64577_p ( .a(FE_OFN1108_g64577_p), .o(FE_OFN1129_g64577_p) );
in01s06 FE_OFC1130_g64577_p ( .a(FE_OFN1101_g64577_p), .o(FE_OFN1130_g64577_p) );
in01s06 FE_OFC1131_g64577_p ( .a(FE_OFN1101_g64577_p), .o(FE_OFN1131_g64577_p) );
in01s06 FE_OFC1132_g64577_p ( .a(FE_OFN1110_g64577_p), .o(FE_OFN1132_g64577_p) );
in01s06 FE_OFC1133_g64577_p ( .a(FE_OFN1110_g64577_p), .o(FE_OFN1133_g64577_p) );
in01s06 FE_OFC1134_g64577_p ( .a(FE_OFN1113_g64577_p), .o(FE_OFN1134_g64577_p) );
in01s06 FE_OFC1135_g64577_p ( .a(FE_OFN1114_g64577_p), .o(FE_OFN1135_g64577_p) );
in01s06 FE_OFC1136_g64577_p ( .a(FE_OFN1108_g64577_p), .o(FE_OFN1136_g64577_p) );
in01s06 FE_OFC1137_g64577_p ( .a(FE_OFN1108_g64577_p), .o(FE_OFN1137_g64577_p) );
in01s03 FE_OFC1138_g64577_p ( .a(FE_OFN1107_g64577_p), .o(FE_OFN1138_g64577_p) );
in01s03 FE_OFC1139_g64577_p ( .a(FE_OFN1138_g64577_p), .o(FE_OFN1139_g64577_p) );
in01s03 FE_OFC1140_g64577_p ( .a(FE_OFN1138_g64577_p), .o(FE_OFN1140_g64577_p) );
in01f06 FE_OFC1141_n_15261 ( .a(n_15261), .o(FE_OFN1141_n_15261) );
in01f06 FE_OFC1142_n_15261 ( .a(FE_OFN1141_n_15261), .o(FE_OFN1142_n_15261) );
in01f06 FE_OFC1143_n_15261 ( .a(FE_OFN1141_n_15261), .o(FE_OFN1143_n_15261) );
in01m06 FE_OFC1144_n_15261 ( .a(FE_OFN1141_n_15261), .o(FE_OFN1144_n_15261) );
in01f08 FE_OFC1145_n_15261 ( .a(FE_OFN1141_n_15261), .o(FE_OFN1145_n_15261) );
in01f10 FE_OFC1146_n_13249 ( .a(n_13249), .o(FE_OFN1146_n_13249) );
in01f04 FE_OFC1147_n_13249 ( .a(FE_OFN1146_n_13249), .o(FE_OFN1147_n_13249) );
in01f08 FE_OFC1148_n_13249 ( .a(FE_OFN1146_n_13249), .o(FE_OFN1148_n_13249) );
in01f04 FE_OFC1149_n_13249 ( .a(FE_OFN1146_n_13249), .o(FE_OFN1149_n_13249) );
in01f08 FE_OFC1150_n_13249 ( .a(FE_OFN1146_n_13249), .o(FE_OFN1150_n_13249) );
in01f08 FE_OFC1151_n_13249 ( .a(FE_OFN1146_n_13249), .o(FE_OFN1151_n_13249) );
in01m04 FE_OFC1152_n_13249 ( .a(FE_OFN1146_n_13249), .o(FE_OFN1152_n_13249) );
in01f06 FE_OFC1153_n_3464 ( .a(n_3464), .o(FE_OFN1153_n_3464) );
in01m04 FE_OFC1154_n_3464 ( .a(FE_OFN1153_n_3464), .o(FE_OFN1154_n_3464) );
in01f08 FE_OFC1155_n_3464 ( .a(FE_OFN1153_n_3464), .o(FE_OFN1155_n_3464) );
in01m02 FE_OFC1156_n_7498 ( .a(n_7498), .o(FE_OFN1156_n_7498) );
in01m06 FE_OFC1157_n_15325 ( .a(n_15325), .o(FE_OFN1157_n_15325) );
in01m08 FE_OFC1158_n_15325 ( .a(FE_OFN1157_n_15325), .o(FE_OFN1158_n_15325) );
in01s10 FE_OFC1159_n_15325 ( .a(FE_OFN1157_n_15325), .o(FE_OFN1159_n_15325) );
in01m01 FE_OFC1160_n_5615 ( .a(n_5592), .o(FE_OFN1160_n_5615) );
in01m02 FE_OFC1161_n_5615 ( .a(n_5592), .o(FE_OFN1161_n_5615) );
in01s02 FE_OFC1162_n_5615 ( .a(n_5592), .o(FE_OFN1162_n_5615) );
in01s04 FE_OFC1163_n_5615 ( .a(FE_OFN1160_n_5615), .o(FE_OFN1163_n_5615) );
in01m04 FE_OFC1164_n_5615 ( .a(FE_OFN1161_n_5615), .o(FE_OFN1164_n_5615) );
in01s02 FE_OFC1165_n_5615 ( .a(FE_OFN1161_n_5615), .o(FE_OFN1165_n_5615) );
in01s06 FE_OFC1166_n_5615 ( .a(FE_OFN1162_n_5615), .o(FE_OFN1166_n_5615) );
in01f08 FE_OFC1167_n_5592 ( .a(n_5592), .o(FE_OFN1167_n_5592) );
in01s04 FE_OFC1168_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1168_n_5592) );
in01m04 FE_OFC1169_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1169_n_5592) );
in01s04 FE_OFC1170_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1170_n_5592) );
in01s06 FE_OFC1171_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1171_n_5592) );
in01m02 FE_OFC1172_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1172_n_5592) );
in01m08 FE_OFC1173_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1173_n_5592) );
in01s06 FE_OFC1174_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1174_n_5592) );
in01f02 FE_OFC1175_n_3476 ( .a(n_3476), .o(FE_OFN1175_n_3476) );
in01f03 FE_OFC1176_n_3476 ( .a(n_3476), .o(FE_OFN1176_n_3476) );
in01f02 FE_OFC1177_n_3476 ( .a(n_3476), .o(FE_OFN1177_n_3476) );
in01f02 FE_OFC1178_n_3476 ( .a(n_3476), .o(FE_OFN1178_n_3476) );
in01m06 FE_OFC1179_n_3476 ( .a(FE_OFN1178_n_3476), .o(FE_OFN1179_n_3476) );
in01m06 FE_OFC1180_n_3476 ( .a(FE_OFN1175_n_3476), .o(FE_OFN1180_n_3476) );
in01f04 FE_OFC1181_n_3476 ( .a(FE_OFN1175_n_3476), .o(FE_OFN1181_n_3476) );
in01m06 FE_OFC1182_n_3476 ( .a(FE_OFN1176_n_3476), .o(FE_OFN1182_n_3476) );
in01m06 FE_OFC1183_n_3476 ( .a(FE_OFN1176_n_3476), .o(FE_OFN1183_n_3476) );
in01m06 FE_OFC1184_n_3476 ( .a(FE_OFN1177_n_3476), .o(FE_OFN1184_n_3476) );
in01m06 FE_OFC1185_n_3476 ( .a(FE_OFN1177_n_3476), .o(FE_OFN1185_n_3476) );
in01m04 FE_OFC1186_n_3476 ( .a(FE_OFN1178_n_3476), .o(FE_OFN1186_n_3476) );
in01f02 FE_OFC1187_n_5742 ( .a(n_5742), .o(FE_OFN1187_n_5742) );
in01f03 FE_OFC1188_n_5742 ( .a(FE_OFN1187_n_5742), .o(FE_OFN1188_n_5742) );
in01f06 FE_OFC1189_n_5742 ( .a(FE_OFN1187_n_5742), .o(FE_OFN1189_n_5742) );
in01m02 FE_OFC1190_n_6935 ( .a(n_6935), .o(FE_OFN1190_n_6935) );
in01f08 FE_OFC1191_n_6935 ( .a(n_6935), .o(FE_OFN1191_n_6935) );
in01f10 FE_OFC1192_n_6935 ( .a(FE_OFN1191_n_6935), .o(FE_OFN1192_n_6935) );
in01m04 FE_OFC1193_n_6935 ( .a(FE_OFN1190_n_6935), .o(FE_OFN1193_n_6935) );
in01m02 FE_OFC1194_n_6935 ( .a(FE_OFN1190_n_6935), .o(FE_OFN1194_n_6935) );
in01m01 FE_OFC1195_n_4090 ( .a(n_4090), .o(FE_OFN1195_n_4090) );
in01s01 FE_OFC1196_n_4090 ( .a(FE_OFN1195_n_4090), .o(FE_OFN1196_n_4090) );
in01s02 FE_OFC1197_n_4090 ( .a(FE_OFN1195_n_4090), .o(FE_OFN1197_n_4090) );
in01m01 FE_OFC1198_n_4090 ( .a(n_4090), .o(FE_OFN1198_n_4090) );
in01m01 FE_OFC1199_n_4090 ( .a(n_4090), .o(FE_OFN1199_n_4090) );
in01s04 FE_OFC1200_n_4090 ( .a(FE_OFN1198_n_4090), .o(FE_OFN1200_n_4090) );
in01s02 FE_OFC1201_n_4090 ( .a(n_4090), .o(FE_OFN1201_n_4090) );
in01s06 FE_OFC1202_n_4090 ( .a(FE_OFN1201_n_4090), .o(FE_OFN1202_n_4090) );
in01s02 FE_OFC1203_n_4090 ( .a(FE_OFN1199_n_4090), .o(FE_OFN1203_n_4090) );
in01s02 FE_OFC1204_n_4090 ( .a(FE_OFN1199_n_4090), .o(FE_OFN1204_n_4090) );
in01s04 FE_OFC1205_n_6356 ( .a(n_6356), .o(FE_OFN1205_n_6356) );
in01s04 FE_OFC1206_n_6356 ( .a(FE_OFN1205_n_6356), .o(FE_OFN1206_n_6356) );
in01s04 FE_OFC1207_n_6356 ( .a(FE_OFN1205_n_6356), .o(FE_OFN1207_n_6356) );
in01s04 FE_OFC1208_n_6356 ( .a(FE_OFN1205_n_6356), .o(FE_OFN1208_n_6356) );
in01s02 FE_OFC1209_n_4151 ( .a(n_4151), .o(FE_OFN1209_n_4151) );
in01s04 FE_OFC1210_n_4151 ( .a(n_4151), .o(FE_OFN1210_n_4151) );
in01s02 FE_OFC1211_n_4151 ( .a(n_4151), .o(FE_OFN1211_n_4151) );
in01s06 FE_OFC1212_n_4151 ( .a(FE_OFN1210_n_4151), .o(FE_OFN1212_n_4151) );
in01s06 FE_OFC1213_n_4151 ( .a(FE_OFN1210_n_4151), .o(FE_OFN1213_n_4151) );
in01s06 FE_OFC1214_n_4151 ( .a(FE_OFN1209_n_4151), .o(FE_OFN1214_n_4151) );
in01s03 FE_OFC1215_n_4151 ( .a(FE_OFN1211_n_4151), .o(FE_OFN1215_n_4151) );
in01s01 FE_OFC1216_n_4151 ( .a(FE_OFN1211_n_4151), .o(FE_OFN1216_n_4151) );
in01s04 FE_OFC1217_n_6886 ( .a(n_6886), .o(FE_OFN1217_n_6886) );
in01s04 FE_OFC1218_n_6886 ( .a(FE_OFN1217_n_6886), .o(FE_OFN1218_n_6886) );
in01s08 FE_OFC1219_n_6886 ( .a(FE_OFN1217_n_6886), .o(FE_OFN1219_n_6886) );
in01m08 FE_OFC1220_n_6391 ( .a(n_6391), .o(FE_OFN1220_n_6391) );
in01m08 FE_OFC1221_n_6391 ( .a(FE_OFN1220_n_6391), .o(FE_OFN1221_n_6391) );
in01m06 FE_OFC1222_n_6391 ( .a(FE_OFN1220_n_6391), .o(FE_OFN1222_n_6391) );
in01m06 FE_OFC1223_n_6391 ( .a(FE_OFN1220_n_6391), .o(FE_OFN1223_n_6391) );
in01m02 FE_OFC1224_n_6391 ( .a(FE_OFN1220_n_6391), .o(FE_OFN1224_n_6391) );
in01s02 FE_OFC1225_n_6391 ( .a(FE_OFN1220_n_6391), .o(FE_OFN1225_n_6391) );
in01m01 FE_OFC1226_n_6391 ( .a(FE_OFN1220_n_6391), .o(FE_OFN1226_n_6391) );
in01m08 FE_OFC1227_n_6391 ( .a(FE_OFN1221_n_6391), .o(FE_OFN1227_n_6391) );
in01m06 FE_OFC1228_n_6391 ( .a(FE_OFN1221_n_6391), .o(FE_OFN1228_n_6391) );
in01s06 FE_OFC1229_n_6391 ( .a(FE_OFN1222_n_6391), .o(FE_OFN1229_n_6391) );
in01s08 FE_OFC1230_n_6391 ( .a(FE_OFN1227_n_6391), .o(FE_OFN1230_n_6391) );
in01s08 FE_OFC1231_n_6391 ( .a(FE_OFN1227_n_6391), .o(FE_OFN1231_n_6391) );
in01s08 FE_OFC1232_n_6391 ( .a(FE_OFN1227_n_6391), .o(FE_OFN1232_n_6391) );
in01s08 FE_OFC1233_n_6391 ( .a(FE_OFN1228_n_6391), .o(FE_OFN1233_n_6391) );
in01s10 FE_OFC1234_n_6391 ( .a(FE_OFN1229_n_6391), .o(FE_OFN1234_n_6391) );
in01s08 FE_OFC1235_n_6391 ( .a(FE_OFN1228_n_6391), .o(FE_OFN1235_n_6391) );
in01s08 FE_OFC1236_n_6391 ( .a(FE_OFN1228_n_6391), .o(FE_OFN1236_n_6391) );
in01s01 FE_OFC1237_n_4092 ( .a(n_4092), .o(FE_OFN1237_n_4092) );
in01s04 FE_OFC1238_n_4092 ( .a(n_4092), .o(FE_OFN1238_n_4092) );
in01s02 FE_OFC1239_n_4092 ( .a(n_4092), .o(FE_OFN1239_n_4092) );
in01s02 FE_OFC1240_n_4092 ( .a(n_4092), .o(FE_OFN1240_n_4092) );
in01s06 FE_OFC1241_n_4092 ( .a(FE_OFN1238_n_4092), .o(FE_OFN1241_n_4092) );
in01s04 FE_OFC1242_n_4092 ( .a(FE_OFN1238_n_4092), .o(FE_OFN1242_n_4092) );
in01s06 FE_OFC1243_n_4092 ( .a(FE_OFN1240_n_4092), .o(FE_OFN1243_n_4092) );
in01s06 FE_OFC1244_n_4092 ( .a(FE_OFN1239_n_4092), .o(FE_OFN1244_n_4092) );
in01m06 FE_OFC1245_n_4093 ( .a(n_4093), .o(FE_OFN1245_n_4093) );
in01s02 FE_OFC1246_n_4093 ( .a(FE_OFN1245_n_4093), .o(FE_OFN1246_n_4093) );
in01s02 FE_OFC1247_n_4093 ( .a(FE_OFN1245_n_4093), .o(FE_OFN1247_n_4093) );
in01s06 FE_OFC1248_n_4093 ( .a(FE_OFN1245_n_4093), .o(FE_OFN1248_n_4093) );
in01s06 FE_OFC1249_n_4093 ( .a(FE_OFN1245_n_4093), .o(FE_OFN1249_n_4093) );
in01s06 FE_OFC1250_n_4093 ( .a(FE_OFN1245_n_4093), .o(FE_OFN1250_n_4093) );
in01s02 FE_OFC1251_n_4143 ( .a(n_4143), .o(FE_OFN1251_n_4143) );
in01s01 FE_OFC1252_n_4143 ( .a(FE_OFN1251_n_4143), .o(FE_OFN1252_n_4143) );
in01s04 FE_OFC1253_n_4143 ( .a(FE_OFN1251_n_4143), .o(FE_OFN1253_n_4143) );
in01s02 FE_OFC1254_n_4143 ( .a(n_4143), .o(FE_OFN1254_n_4143) );
in01s02 FE_OFC1255_n_4143 ( .a(n_4143), .o(FE_OFN1255_n_4143) );
in01s02 FE_OFC1256_n_4143 ( .a(n_4143), .o(FE_OFN1256_n_4143) );
in01s01 FE_OFC1257_n_4143 ( .a(FE_OFN1254_n_4143), .o(FE_OFN1257_n_4143) );
in01s04 FE_OFC1258_n_4143 ( .a(FE_OFN1254_n_4143), .o(FE_OFN1258_n_4143) );
in01s01 FE_OFC1259_n_4143 ( .a(FE_OFN1255_n_4143), .o(FE_OFN1259_n_4143) );
in01s04 FE_OFC1260_n_4143 ( .a(FE_OFN1255_n_4143), .o(FE_OFN1260_n_4143) );
in01s06 FE_OFC1261_n_4143 ( .a(FE_OFN1256_n_4143), .o(FE_OFN1261_n_4143) );
in01s02 FE_OFC1262_n_4095 ( .a(n_4095), .o(FE_OFN1262_n_4095) );
in01s02 FE_OFC1263_n_4095 ( .a(n_4095), .o(FE_OFN1263_n_4095) );
in01s04 FE_OFC1264_n_4095 ( .a(FE_OFN1262_n_4095), .o(FE_OFN1264_n_4095) );
in01s02 FE_OFC1265_n_4095 ( .a(FE_OFN1262_n_4095), .o(FE_OFN1265_n_4095) );
in01s02 FE_OFC1266_n_4095 ( .a(n_4095), .o(FE_OFN1266_n_4095) );
in01s02 FE_OFC1267_n_4095 ( .a(n_4095), .o(FE_OFN1267_n_4095) );
in01s06 FE_OFC1268_n_4095 ( .a(FE_OFN1263_n_4095), .o(FE_OFN1268_n_4095) );
in01s06 FE_OFC1269_n_4095 ( .a(FE_OFN1267_n_4095), .o(FE_OFN1269_n_4095) );
in01s06 FE_OFC1270_n_4095 ( .a(FE_OFN1266_n_4095), .o(FE_OFN1270_n_4095) );
in01m06 FE_OFC1271_n_4096 ( .a(n_4096), .o(FE_OFN1271_n_4096) );
in01s08 FE_OFC1272_n_4096 ( .a(FE_OFN1271_n_4096), .o(FE_OFN1272_n_4096) );
in01s02 FE_OFC1273_n_4096 ( .a(FE_OFN1271_n_4096), .o(FE_OFN1273_n_4096) );
in01s04 FE_OFC1274_n_4096 ( .a(FE_OFN1271_n_4096), .o(FE_OFN1274_n_4096) );
in01s04 FE_OFC1275_n_4096 ( .a(FE_OFN1271_n_4096), .o(FE_OFN1275_n_4096) );
in01s06 FE_OFC1276_n_4096 ( .a(FE_OFN1271_n_4096), .o(FE_OFN1276_n_4096) );
in01s02 FE_OFC1277_n_4097 ( .a(n_4097), .o(FE_OFN1277_n_4097) );
in01s04 FE_OFC1278_n_4097 ( .a(FE_OFN1277_n_4097), .o(FE_OFN1278_n_4097) );
in01s02 FE_OFC1279_n_4097 ( .a(FE_OFN1277_n_4097), .o(FE_OFN1279_n_4097) );
in01s02 FE_OFC1280_n_4097 ( .a(n_4097), .o(FE_OFN1280_n_4097) );
in01s04 FE_OFC1281_n_4097 ( .a(n_4097), .o(FE_OFN1281_n_4097) );
in01s01 FE_OFC1282_n_4097 ( .a(FE_OFN1280_n_4097), .o(FE_OFN1282_n_4097) );
in01s06 FE_OFC1283_n_4097 ( .a(FE_OFN1280_n_4097), .o(FE_OFN1283_n_4097) );
in01s06 FE_OFC1284_n_4097 ( .a(FE_OFN1281_n_4097), .o(FE_OFN1284_n_4097) );
in01s06 FE_OFC1285_n_4097 ( .a(FE_OFN1281_n_4097), .o(FE_OFN1285_n_4097) );
in01m01 FE_OFC1286_n_4098 ( .a(n_4098), .o(FE_OFN1286_n_4098) );
in01s01 FE_OFC1287_n_4098 ( .a(n_4098), .o(FE_OFN1287_n_4098) );
in01s04 FE_OFC1288_n_4098 ( .a(FE_OFN1286_n_4098), .o(FE_OFN1288_n_4098) );
in01s02 FE_OFC1289_n_4098 ( .a(FE_OFN1287_n_4098), .o(FE_OFN1289_n_4098) );
in01m02 FE_OFC1290_n_4098 ( .a(n_4098), .o(FE_OFN1290_n_4098) );
in01s02 FE_OFC1291_n_4098 ( .a(n_4098), .o(FE_OFN1291_n_4098) );
in01s02 FE_OFC1292_n_4098 ( .a(n_4098), .o(FE_OFN1292_n_4098) );
in01s06 FE_OFC1293_n_4098 ( .a(FE_OFN1290_n_4098), .o(FE_OFN1293_n_4098) );
in01s06 FE_OFC1294_n_4098 ( .a(FE_OFN1291_n_4098), .o(FE_OFN1294_n_4098) );
in01s06 FE_OFC1295_n_4098 ( .a(FE_OFN1292_n_4098), .o(FE_OFN1295_n_4098) );
in01m01 FE_OFC1296_n_5763 ( .a(n_5763), .o(FE_OFN1296_n_5763) );
in01m02 FE_OFC1297_n_5763 ( .a(n_5763), .o(FE_OFN1297_n_5763) );
in01m01 FE_OFC1298_n_5763 ( .a(n_5763), .o(FE_OFN1298_n_5763) );
in01s04 FE_OFC1299_n_5763 ( .a(FE_OFN1297_n_5763), .o(FE_OFN1299_n_5763) );
in01s04 FE_OFC1300_n_5763 ( .a(FE_OFN1298_n_5763), .o(FE_OFN1300_n_5763) );
in01s06 FE_OFC1301_n_5763 ( .a(FE_OFN1297_n_5763), .o(FE_OFN1301_n_5763) );
in01s06 FE_OFC1302_n_5763 ( .a(FE_OFN1296_n_5763), .o(FE_OFN1302_n_5763) );
in01f03 FE_OFC1303_n_13124 ( .a(n_13124), .o(FE_OFN1303_n_13124) );
in01f04 FE_OFC1304_n_13124 ( .a(FE_OFN1303_n_13124), .o(FE_OFN1304_n_13124) );
in01f03 FE_OFC1305_n_13124 ( .a(FE_OFN1303_n_13124), .o(FE_OFN1305_n_13124) );
in01f02 FE_OFC1306_n_13124 ( .a(FE_OFN1303_n_13124), .o(FE_OFN1306_n_13124) );
in01s10 FE_OFC1307_n_6624 ( .a(n_6624), .o(FE_OFN1307_n_6624) );
in01s10 FE_OFC1308_n_6624 ( .a(n_6624), .o(FE_OFN1308_n_6624) );
in01m10 FE_OFC1309_n_6624 ( .a(n_6624), .o(FE_OFN1309_n_6624) );
in01s08 FE_OFC1310_n_6624 ( .a(FE_OFN1308_n_6624), .o(FE_OFN1310_n_6624) );
in01s10 FE_OFC1311_n_6624 ( .a(FE_OFN1307_n_6624), .o(FE_OFN1311_n_6624) );
in01s06 FE_OFC1312_n_6624 ( .a(FE_OFN1307_n_6624), .o(FE_OFN1312_n_6624) );
in01s08 FE_OFC1313_n_6624 ( .a(FE_OFN1308_n_6624), .o(FE_OFN1313_n_6624) );
in01s08 FE_OFC1314_n_6624 ( .a(FE_OFN1308_n_6624), .o(FE_OFN1314_n_6624) );
in01m08 FE_OFC1315_n_6624 ( .a(FE_OFN1308_n_6624), .o(FE_OFN1315_n_6624) );
in01s10 FE_OFC1316_n_6624 ( .a(FE_OFN1309_n_6624), .o(FE_OFN1316_n_6624) );
in01m10 FE_OFC1317_n_6624 ( .a(FE_OFN1309_n_6624), .o(FE_OFN1317_n_6624) );
in01m04 FE_OFC1318_n_6436 ( .a(n_6436), .o(FE_OFN1318_n_6436) );
in01m02 FE_OFC1319_n_6436 ( .a(FE_OFN1318_n_6436), .o(FE_OFN1319_n_6436) );
in01m06 FE_OFC1320_n_6436 ( .a(FE_OFN1318_n_6436), .o(FE_OFN1320_n_6436) );
in01s08 FE_OFC1321_n_6436 ( .a(n_6436), .o(FE_OFN1321_n_6436) );
in01s06 FE_OFC1322_n_6436 ( .a(FE_OFN1321_n_6436), .o(FE_OFN1322_n_6436) );
in01s08 FE_OFC1323_n_6436 ( .a(FE_OFN1321_n_6436), .o(FE_OFN1323_n_6436) );
in01f04 FE_OFC1324_n_13547 ( .a(n_13547), .o(FE_OFN1324_n_13547) );
in01f03 FE_OFC1325_n_13547 ( .a(n_13547), .o(FE_OFN1325_n_13547) );
in01m06 FE_OFC1326_n_13547 ( .a(FE_OFN1324_n_13547), .o(FE_OFN1326_n_13547) );
in01m08 FE_OFC1327_n_13547 ( .a(FE_OFN1324_n_13547), .o(FE_OFN1327_n_13547) );
in01f04 FE_OFC1328_n_13547 ( .a(n_13547), .o(FE_OFN1328_n_13547) );
in01f01 FE_OFC1329_n_13547 ( .a(n_13547), .o(FE_OFN1329_n_13547) );
in01f06 FE_OFC1330_n_13547 ( .a(FE_OFN1325_n_13547), .o(FE_OFN1330_n_13547) );
in01m08 FE_OFC1331_n_13547 ( .a(FE_OFN1328_n_13547), .o(FE_OFN1331_n_13547) );
in01m04 FE_OFC1332_n_13547 ( .a(FE_OFN1328_n_13547), .o(FE_OFN1332_n_13547) );
in01f02 FE_OFC1333_n_13547 ( .a(FE_OFN1329_n_13547), .o(FE_OFN1333_n_13547) );
in01f02 FE_OFC1334_n_13720 ( .a(n_13720), .o(FE_OFN1334_n_13720) );
in01f02 FE_OFC1335_n_13720 ( .a(FE_OFN1334_n_13720), .o(FE_OFN1335_n_13720) );
in01f02 FE_OFC1336_n_16439 ( .a(n_16439), .o(FE_OFN1336_n_16439) );
in01f06 FE_OFC1337_n_16439 ( .a(FE_OFN1336_n_16439), .o(FE_OFN1337_n_16439) );
in01f06 FE_OFC1338_n_8567 ( .a(n_8567), .o(FE_OFN1338_n_8567) );
in01s04 FE_OFC1339_n_8567 ( .a(n_8567), .o(FE_OFN1339_n_8567) );
in01f02 FE_OFC1340_n_8567 ( .a(n_8567), .o(FE_OFN1340_n_8567) );
in01f04 FE_OFC1341_n_8567 ( .a(FE_OFN1339_n_8567), .o(FE_OFN1341_n_8567) );
in01f06 FE_OFC1342_n_8567 ( .a(FE_OFN1339_n_8567), .o(FE_OFN1342_n_8567) );
in01f04 FE_OFC1343_n_8567 ( .a(FE_OFN1340_n_8567), .o(FE_OFN1343_n_8567) );
in01f04 FE_OFC1344_n_8567 ( .a(FE_OFN1340_n_8567), .o(FE_OFN1344_n_8567) );
in01f06 FE_OFC1345_n_8567 ( .a(FE_OFN1338_n_8567), .o(FE_OFN1345_n_8567) );
in01s02 FE_OFC1346_n_8567 ( .a(FE_OFN1338_n_8567), .o(FE_OFN1346_n_8567) );
in01f02 FE_OFC1347_n_8567 ( .a(FE_OFN1338_n_8567), .o(FE_OFN1347_n_8567) );
in01f08 FE_OFC1348_n_8567 ( .a(FE_OFN1338_n_8567), .o(FE_OFN1348_n_8567) );
in01f02 FE_OFC1349_n_8567 ( .a(FE_OFN1338_n_8567), .o(FE_OFN1349_n_8567) );
in01f08 FE_OFC1350_n_8567 ( .a(FE_OFN1341_n_8567), .o(FE_OFN1350_n_8567) );
in01f08 FE_OFC1351_n_8567 ( .a(FE_OFN1342_n_8567), .o(FE_OFN1351_n_8567) );
in01f08 FE_OFC1352_n_8567 ( .a(FE_OFN1343_n_8567), .o(FE_OFN1352_n_8567) );
in01f08 FE_OFC1353_n_8567 ( .a(FE_OFN1343_n_8567), .o(FE_OFN1353_n_8567) );
in01f04 FE_OFC1354_n_8567 ( .a(FE_OFN1346_n_8567), .o(FE_OFN1354_n_8567) );
in01f06 FE_OFC1355_n_8567 ( .a(FE_OFN1347_n_8567), .o(FE_OFN1355_n_8567) );
in01f02 FE_OFC1356_n_8567 ( .a(FE_OFN1347_n_8567), .o(FE_OFN1356_n_8567) );
in01f08 FE_OFC1357_n_8567 ( .a(FE_OFN1348_n_8567), .o(FE_OFN1357_n_8567) );
in01f04 FE_OFC1358_n_8567 ( .a(FE_OFN1341_n_8567), .o(FE_OFN1358_n_8567) );
in01f02 FE_OFC1359_n_8567 ( .a(FE_OFN1345_n_8567), .o(FE_OFN1359_n_8567) );
in01f08 FE_OFC1360_n_8567 ( .a(FE_OFN1345_n_8567), .o(FE_OFN1360_n_8567) );
in01f08 FE_OFC1361_n_8567 ( .a(FE_OFN1348_n_8567), .o(FE_OFN1361_n_8567) );
in01f08 FE_OFC1362_n_8567 ( .a(FE_OFN1348_n_8567), .o(FE_OFN1362_n_8567) );
in01f08 FE_OFC1363_n_8567 ( .a(FE_OFN1342_n_8567), .o(FE_OFN1363_n_8567) );
in01f02 FE_OFC1364_n_8567 ( .a(FE_OFN1342_n_8567), .o(FE_OFN1364_n_8567) );
in01f02 FE_OFC1365_n_8567 ( .a(FE_OFN1344_n_8567), .o(FE_OFN1365_n_8567) );
in01f06 FE_OFC1366_n_8567 ( .a(FE_OFN1344_n_8567), .o(FE_OFN1366_n_8567) );
in01f08 FE_OFC1367_n_8567 ( .a(FE_OFN1345_n_8567), .o(FE_OFN1367_n_8567) );
in01f08 FE_OFC1368_n_8567 ( .a(FE_OFN1351_n_8567), .o(FE_OFN1368_n_8567) );
in01f08 FE_OFC1369_n_8567 ( .a(FE_OFN1352_n_8567), .o(FE_OFN1369_n_8567) );
in01f08 FE_OFC1370_n_8567 ( .a(FE_OFN1353_n_8567), .o(FE_OFN1370_n_8567) );
in01s02 FE_OFC1371_n_8567 ( .a(FE_OFN1345_n_8567), .o(FE_OFN1371_n_8567) );
in01f04 FE_OFC1372_n_8567 ( .a(FE_OFN1354_n_8567), .o(FE_OFN1372_n_8567) );
in01f06 FE_OFC1373_n_8567 ( .a(FE_OFN1354_n_8567), .o(FE_OFN1373_n_8567) );
in01f08 FE_OFC1374_n_8567 ( .a(FE_OFN1356_n_8567), .o(FE_OFN1374_n_8567) );
in01f08 FE_OFC1376_n_8567 ( .a(FE_OFN1357_n_8567), .o(FE_OFN1376_n_8567) );
in01f08 FE_OFC1377_n_8567 ( .a(FE_OFN1350_n_8567), .o(FE_OFN1377_n_8567) );
in01f06 FE_OFC1378_n_8567 ( .a(FE_OFN1358_n_8567), .o(FE_OFN1378_n_8567) );
in01f02 FE_OFC1379_n_8567 ( .a(FE_OFN1358_n_8567), .o(FE_OFN1379_n_8567) );
in01f06 FE_OFC1380_n_8567 ( .a(FE_OFN1351_n_8567), .o(FE_OFN1380_n_8567) );
in01f06 FE_OFC1381_n_8567 ( .a(FE_OFN1352_n_8567), .o(FE_OFN1381_n_8567) );
in01f08 FE_OFC1382_n_8567 ( .a(FE_OFN1353_n_8567), .o(FE_OFN1382_n_8567) );
in01f06 FE_OFC1383_n_8567 ( .a(FE_OFN1359_n_8567), .o(FE_OFN1383_n_8567) );
in01f08 FE_OFC1384_n_8567 ( .a(FE_OFN1360_n_8567), .o(FE_OFN1384_n_8567) );
in01f06 FE_OFC1385_n_8567 ( .a(FE_OFN1355_n_8567), .o(FE_OFN1385_n_8567) );
in01f02 FE_OFC1386_n_8567 ( .a(FE_OFN1355_n_8567), .o(FE_OFN1386_n_8567) );
in01f08 FE_OFC1387_n_8567 ( .a(FE_OFN1355_n_8567), .o(FE_OFN1387_n_8567) );
in01f06 FE_OFC1388_n_8567 ( .a(FE_OFN1355_n_8567), .o(FE_OFN1388_n_8567) );
in01f08 FE_OFC1389_n_8567 ( .a(FE_OFN1357_n_8567), .o(FE_OFN1389_n_8567) );
in01f06 FE_OFC1390_n_8567 ( .a(FE_OFN1362_n_8567), .o(FE_OFN1390_n_8567) );
in01f08 FE_OFC1391_n_8567 ( .a(FE_OFN1350_n_8567), .o(FE_OFN1391_n_8567) );
in01f06 FE_OFC1392_n_8567 ( .a(FE_OFN1351_n_8567), .o(FE_OFN1392_n_8567) );
in01f10 FE_OFC1394_n_8567 ( .a(FE_OFN1363_n_8567), .o(FE_OFN1394_n_8567) );
in01f08 FE_OFC1396_n_8567 ( .a(FE_OFN1364_n_8567), .o(FE_OFN1396_n_8567) );
in01f06 FE_OFC1397_n_8567 ( .a(FE_OFN1352_n_8567), .o(FE_OFN1397_n_8567) );
in01f08 FE_OFC1398_n_8567 ( .a(FE_OFN1352_n_8567), .o(FE_OFN1398_n_8567) );
in01f08 FE_OFC1399_n_8567 ( .a(FE_OFN1353_n_8567), .o(FE_OFN1399_n_8567) );
in01f08 FE_OFC1400_n_8567 ( .a(FE_OFN1353_n_8567), .o(FE_OFN1400_n_8567) );
in01f06 FE_OFC1401_n_8567 ( .a(FE_OFN1365_n_8567), .o(FE_OFN1401_n_8567) );
in01f08 FE_OFC1402_n_8567 ( .a(FE_OFN1366_n_8567), .o(FE_OFN1402_n_8567) );
in01f08 FE_OFC1403_n_8567 ( .a(FE_OFN1366_n_8567), .o(FE_OFN1403_n_8567) );
in01f08 FE_OFC1404_n_8567 ( .a(FE_OFN1367_n_8567), .o(FE_OFN1404_n_8567) );
in01f08 FE_OFC1405_n_8567 ( .a(FE_OFN1360_n_8567), .o(FE_OFN1405_n_8567) );
in01f08 FE_OFC1406_n_8567 ( .a(FE_OFN1357_n_8567), .o(FE_OFN1406_n_8567) );
in01f08 FE_OFC1407_n_8567 ( .a(FE_OFN1357_n_8567), .o(FE_OFN1407_n_8567) );
in01f08 FE_OFC1408_n_8567 ( .a(FE_OFN1361_n_8567), .o(FE_OFN1408_n_8567) );
in01f06 FE_OFC1409_n_8567 ( .a(FE_OFN1362_n_8567), .o(FE_OFN1409_n_8567) );
in01f06 FE_OFC1410_n_8567 ( .a(FE_OFN1362_n_8567), .o(FE_OFN1410_n_8567) );
in01f08 FE_OFC1411_n_8567 ( .a(FE_OFN1350_n_8567), .o(FE_OFN1411_n_8567) );
in01f06 FE_OFC1412_n_8567 ( .a(FE_OFN1351_n_8567), .o(FE_OFN1412_n_8567) );
in01f06 FE_OFC1413_n_8567 ( .a(FE_OFN1351_n_8567), .o(FE_OFN1413_n_8567) );
in01f08 FE_OFC1414_n_8567 ( .a(FE_OFN1367_n_8567), .o(FE_OFN1414_n_8567) );
in01f08 FE_OFC1415_n_8567 ( .a(FE_OFN1367_n_8567), .o(FE_OFN1415_n_8567) );
in01f08 FE_OFC1416_n_8567 ( .a(FE_OFN1360_n_8567), .o(FE_OFN1416_n_8567) );
in01f08 FE_OFC1417_n_8567 ( .a(FE_OFN1360_n_8567), .o(FE_OFN1417_n_8567) );
in01f06 FE_OFC1419_n_8567 ( .a(FE_OFN1371_n_8567), .o(FE_OFN1419_n_8567) );
in01f08 FE_OFC1420_n_8567 ( .a(FE_OFN1350_n_8567), .o(FE_OFN1420_n_8567) );
in01f08 FE_OFC1421_n_8567 ( .a(FE_OFN1350_n_8567), .o(FE_OFN1421_n_8567) );
in01f06 FE_OFC1422_n_8567 ( .a(FE_OFN1361_n_8567), .o(FE_OFN1422_n_8567) );
in01f06 FE_OFC1423_n_8567 ( .a(FE_OFN1361_n_8567), .o(FE_OFN1423_n_8567) );
in01f08 FE_OFC1424_n_8567 ( .a(FE_OFN1361_n_8567), .o(FE_OFN1424_n_8567) );
in01f06 FE_OFC1425_n_8567 ( .a(FE_OFN1361_n_8567), .o(FE_OFN1425_n_8567) );
in01f04 FE_OFC1426_n_8567 ( .a(FE_OFN1379_n_8567), .o(FE_OFN1426_n_8567) );
in01f06 FE_OFC1427_n_8567 ( .a(FE_OFN1426_n_8567), .o(FE_OFN1427_n_8567) );
in01f04 FE_OFC1428_n_8567 ( .a(FE_OFN1426_n_8567), .o(FE_OFN1428_n_8567) );
in01f04 FE_OFC1429_n_16779 ( .a(n_16779), .o(FE_OFN1429_n_16779) );
in01f04 FE_OFC1430_n_16779 ( .a(n_16779), .o(FE_OFN1430_n_16779) );
in01f02 FE_OFC1431_n_16779 ( .a(FE_OFN1429_n_16779), .o(FE_OFN1431_n_16779) );
in01f08 FE_OFC1432_n_16779 ( .a(FE_OFN1429_n_16779), .o(FE_OFN1432_n_16779) );
in01f06 FE_OFC1433_n_16779 ( .a(FE_OFN1430_n_16779), .o(FE_OFN1433_n_16779) );
in01m01 FE_OFC1434_n_9372 ( .a(n_9372), .o(FE_OFN1434_n_9372) );
in01f10 FE_OFC1435_n_9372 ( .a(n_9372), .o(FE_OFN1435_n_9372) );
in01m08 FE_OFC1436_n_9372 ( .a(FE_OFN1435_n_9372), .o(FE_OFN1436_n_9372) );
in01m06 FE_OFC1437_n_9372 ( .a(FE_OFN1435_n_9372), .o(FE_OFN1437_n_9372) );
in01f08 FE_OFC1438_n_9372 ( .a(FE_OFN1435_n_9372), .o(FE_OFN1438_n_9372) );
in01f08 FE_OFC1439_n_9372 ( .a(FE_OFN1435_n_9372), .o(FE_OFN1439_n_9372) );
in01f08 FE_OFC1440_n_9372 ( .a(FE_OFN1435_n_9372), .o(FE_OFN1440_n_9372) );
in01m06 FE_OFC1441_n_9372 ( .a(FE_OFN1435_n_9372), .o(FE_OFN1441_n_9372) );
in01f04 FE_OFC1442_n_11125 ( .a(n_11125), .o(FE_OFN1442_n_11125) );
in01f04 FE_OFC1443_n_11125 ( .a(n_11125), .o(FE_OFN1443_n_11125) );
in01f04 FE_OFC1444_n_11125 ( .a(FE_OFN1442_n_11125), .o(FE_OFN1444_n_11125) );
in01f10 FE_OFC1445_n_11125 ( .a(FE_OFN1443_n_11125), .o(FE_OFN1445_n_11125) );
in01f08 FE_OFC1446_n_11125 ( .a(FE_OFN1442_n_11125), .o(FE_OFN1446_n_11125) );
in01f04 FE_OFC1447_n_9163 ( .a(n_9163), .o(FE_OFN1447_n_9163) );
in01f01 FE_OFC1448_n_9163 ( .a(n_9163), .o(FE_OFN1448_n_9163) );
in01f03 FE_OFC1449_n_9163 ( .a(FE_OFN1448_n_9163), .o(FE_OFN1449_n_9163) );
in01f02 FE_OFC1450_n_9163 ( .a(FE_OFN1448_n_9163), .o(FE_OFN1450_n_9163) );
in01f06 FE_OFC1451_n_10588 ( .a(n_10588), .o(FE_OFN1451_n_10588) );
in01f02 FE_OFC1452_n_10588 ( .a(n_10588), .o(FE_OFN1452_n_10588) );
in01f06 FE_OFC1453_n_10588 ( .a(FE_OFN1452_n_10588), .o(FE_OFN1453_n_10588) );
in01f06 FE_OFC1454_n_11138 ( .a(n_11138), .o(FE_OFN1454_n_11138) );
in01f06 FE_OFC1455_n_11138 ( .a(FE_OFN1454_n_11138), .o(FE_OFN1455_n_11138) );
in01f06 FE_OFC1456_n_11138 ( .a(FE_OFN1454_n_11138), .o(FE_OFN1456_n_11138) );
in01f06 FE_OFC1457_n_11138 ( .a(FE_OFN1454_n_11138), .o(FE_OFN1457_n_11138) );
in01f06 FE_OFC1458_n_11138 ( .a(FE_OFN1454_n_11138), .o(FE_OFN1458_n_11138) );
in01f06 FE_OFC1459_n_11795 ( .a(n_11795), .o(FE_OFN1459_n_11795) );
in01f08 FE_OFC1460_n_11795 ( .a(FE_OFN1459_n_11795), .o(FE_OFN1460_n_11795) );
in01f04 FE_OFC1461_n_11795 ( .a(FE_OFN1459_n_11795), .o(FE_OFN1461_n_11795) );
in01f06 FE_OFC1462_n_11795 ( .a(FE_OFN1459_n_11795), .o(FE_OFN1462_n_11795) );
in01f04 FE_OFC1463_n_10789 ( .a(n_10789), .o(FE_OFN1463_n_10789) );
in01f04 FE_OFC1464_n_10789 ( .a(n_10789), .o(FE_OFN1464_n_10789) );
in01f06 FE_OFC1465_n_10789 ( .a(FE_OFN1463_n_10789), .o(FE_OFN1465_n_10789) );
in01f06 FE_OFC1466_n_10789 ( .a(FE_OFN1464_n_10789), .o(FE_OFN1466_n_10789) );
in01f06 FE_OFC1467_n_10789 ( .a(FE_OFN1464_n_10789), .o(FE_OFN1467_n_10789) );
in01f06 FE_OFC1468_n_10789 ( .a(FE_OFN1463_n_10789), .o(FE_OFN1468_n_10789) );
in01f03 FE_OFC1469_g52675_p ( .a(g52675_p), .o(FE_OFN1469_g52675_p) );
in01s01 FE_OFC146_g65530_p ( .a(g65530_p), .o(FE_OFN146_g65530_p) );
in01f04 FE_OFC1470_g52675_p ( .a(FE_OFN1469_g52675_p), .o(FE_OFN1470_g52675_p) );
in01f03 FE_OFC1471_g52675_p ( .a(FE_OFN1469_g52675_p), .o(FE_OFN1471_g52675_p) );
in01f03 FE_OFC1472_g52675_p ( .a(FE_OFN1469_g52675_p), .o(FE_OFN1472_g52675_p) );
in01f04 FE_OFC1473_n_16637 ( .a(n_16637), .o(FE_OFN1473_n_16637) );
in01f04 FE_OFC1474_n_16637 ( .a(n_16637), .o(FE_OFN1474_n_16637) );
in01f06 FE_OFC1475_n_16637 ( .a(n_16637), .o(FE_OFN1475_n_16637) );
in01f06 FE_OFC1477_n_16637 ( .a(FE_OFN1473_n_16637), .o(FE_OFN1477_n_16637) );
in01f08 FE_OFC1478_n_16637 ( .a(FE_OFN1474_n_16637), .o(FE_OFN1478_n_16637) );
in01f08 FE_OFC1479_n_16637 ( .a(FE_OFN1475_n_16637), .o(FE_OFN1479_n_16637) );
in01s01 FE_OFC147_g65530_p ( .a(FE_OFN146_g65530_p), .o(FE_OFN147_g65530_p) );
in01f03 FE_OFC1480_n_15534 ( .a(n_15534), .o(FE_OFN1480_n_15534) );
in01f04 FE_OFC1481_n_15534 ( .a(n_15534), .o(FE_OFN1481_n_15534) );
in01f02 FE_OFC1483_n_15534 ( .a(n_15534), .o(FE_OFN1483_n_15534) );
in01f06 FE_OFC1484_n_15534 ( .a(FE_OFN1480_n_15534), .o(FE_OFN1484_n_15534) );
in01f06 FE_OFC1485_n_15534 ( .a(FE_OFN1483_n_15534), .o(FE_OFN1485_n_15534) );
in01f08 FE_OFC1486_n_16992 ( .a(n_16992), .o(FE_OFN1486_n_16992) );
in01f04 FE_OFC1487_n_9320 ( .a(n_9320), .o(FE_OFN1487_n_9320) );
in01f02 FE_OFC1488_n_9320 ( .a(n_9320), .o(FE_OFN1488_n_9320) );
in01f06 FE_OFC1489_n_9320 ( .a(FE_OFN1487_n_9320), .o(FE_OFN1489_n_9320) );
in01f06 FE_OFC1490_n_9320 ( .a(FE_OFN1487_n_9320), .o(FE_OFN1490_n_9320) );
in01f01 FE_OFC1491_n_9320 ( .a(FE_OFN1487_n_9320), .o(FE_OFN1491_n_9320) );
in01f06 FE_OFC1492_n_9320 ( .a(FE_OFN1490_n_9320), .o(FE_OFN1492_n_9320) );
in01f08 FE_OFC1493_n_9320 ( .a(FE_OFN1492_n_9320), .o(FE_OFN1493_n_9320) );
in01f04 FE_OFC1495_n_15558 ( .a(n_15558), .o(FE_OFN1495_n_15558) );
in01f01 FE_OFC1496_n_15558 ( .a(n_15558), .o(FE_OFN1496_n_15558) );
in01f02 FE_OFC1497_n_15558 ( .a(n_15558), .o(FE_OFN1497_n_15558) );
in01f06 FE_OFC1498_n_15558 ( .a(FE_OFN1495_n_15558), .o(FE_OFN1498_n_15558) );
in01f06 FE_OFC1499_n_15558 ( .a(FE_OFN1495_n_15558), .o(FE_OFN1499_n_15558) );
in01f02 FE_OFC1500_n_15558 ( .a(FE_OFN1496_n_15558), .o(FE_OFN1500_n_15558) );
in01f02 FE_OFC1501_n_15558 ( .a(FE_OFN1496_n_15558), .o(FE_OFN1501_n_15558) );
in01f06 FE_OFC1502_n_15558 ( .a(FE_OFN1497_n_15558), .o(FE_OFN1502_n_15558) );
in01f08 FE_OFC1505_n_15768 ( .a(FE_OFN1503_n_15768), .o(FE_OFN1505_n_15768) );
in01f01 FE_OFC1506_n_15768 ( .a(FE_OFN1503_n_15768), .o(FE_OFN1506_n_15768) );
in01f06 FE_OFC1507_n_15587 ( .a(n_15587), .o(FE_OFN1507_n_15587) );
in01f06 FE_OFC1508_n_15587 ( .a(FE_OFN1507_n_15587), .o(FE_OFN1508_n_15587) );
in01f06 FE_OFC1509_n_15587 ( .a(FE_OFN1507_n_15587), .o(FE_OFN1509_n_15587) );
in01f04 FE_OFC1510_n_15587 ( .a(FE_OFN1507_n_15587), .o(FE_OFN1510_n_15587) );
in01f04 FE_OFC1511_n_15587 ( .a(FE_OFN1507_n_15587), .o(FE_OFN1511_n_15587) );
in01f04 FE_OFC1513_n_14987 ( .a(FE_OCP_RBN1923_n_10273), .o(FE_OFN1513_n_14987) );
in01f02 FE_OFC1514_n_10538 ( .a(FE_OCP_RBN1965_FE_RN_459_0), .o(FE_OFN1514_n_10538) );
in01f04 FE_OFC1519_n_10892 ( .a(n_10892), .o(FE_OFN1519_n_10892) );
in01f03 FE_OFC1520_n_10892 ( .a(n_10892), .o(FE_OFN1520_n_10892) );
in01f02 FE_OFC1521_n_10892 ( .a(FE_OFN1519_n_10892), .o(FE_OFN1521_n_10892) );
in01f08 FE_OFC1522_n_10892 ( .a(FE_OFN1519_n_10892), .o(FE_OFN1522_n_10892) );
in01f06 FE_OFC1523_n_10892 ( .a(FE_OFN1520_n_10892), .o(FE_OFN1523_n_10892) );
in01f02 FE_OFC1524_n_10853 ( .a(n_10853), .o(FE_OFN1524_n_10853) );
in01f03 FE_OFC1525_n_10853 ( .a(n_10853), .o(FE_OFN1525_n_10853) );
in01f04 FE_OFC1526_n_10853 ( .a(n_10853), .o(FE_OFN1526_n_10853) );
in01f04 FE_OFC1527_n_10853 ( .a(FE_OFN1524_n_10853), .o(FE_OFN1527_n_10853) );
in01f06 FE_OFC1528_n_10853 ( .a(FE_OFN1526_n_10853), .o(FE_OFN1528_n_10853) );
in01f06 FE_OFC1529_n_10853 ( .a(FE_OFN1525_n_10853), .o(FE_OFN1529_n_10853) );
in01f06 FE_OFC1530_n_10853 ( .a(FE_OFN1526_n_10853), .o(FE_OFN1530_n_10853) );
in01f02 FE_OFC1531_n_10143 ( .a(n_10143), .o(FE_OFN1531_n_10143) );
in01f06 FE_OFC1532_n_10143 ( .a(n_10143), .o(FE_OFN1532_n_10143) );
in01f02 FE_OFC1533_n_10143 ( .a(n_10143), .o(FE_OFN1533_n_10143) );
in01f02 FE_OFC1535_n_10143 ( .a(FE_OFN1533_n_10143), .o(FE_OFN1535_n_10143) );
in01f04 FE_OFC1536_n_10143 ( .a(FE_OFN1533_n_10143), .o(FE_OFN1536_n_10143) );
in01f02 FE_OFC1537_n_10595 ( .a(n_10595), .o(FE_OFN1537_n_10595) );
in01f04 FE_OFC1538_n_10595 ( .a(FE_OFN1537_n_10595), .o(FE_OFN1538_n_10595) );
in01f04 FE_OFC1539_n_10595 ( .a(FE_OFN1537_n_10595), .o(FE_OFN1539_n_10595) );
in01f02 FE_OFC1540_n_10595 ( .a(n_10595), .o(FE_OFN1540_n_10595) );
in01f04 FE_OFC1541_n_10595 ( .a(n_10595), .o(FE_OFN1541_n_10595) );
in01f04 FE_OFC1542_n_10566 ( .a(n_10566), .o(FE_OFN1542_n_10566) );
in01f06 FE_OFC1543_n_10566 ( .a(n_10566), .o(FE_OFN1543_n_10566) );
in01f04 FE_OFC1544_n_10566 ( .a(n_10566), .o(FE_OFN1544_n_10566) );
in01f02 FE_OFC1545_n_10566 ( .a(FE_OFN1543_n_10566), .o(FE_OFN1545_n_10566) );
in01f08 FE_OFC1546_n_10566 ( .a(FE_OFN1543_n_10566), .o(FE_OFN1546_n_10566) );
in01f08 FE_OFC1547_n_10566 ( .a(FE_OFN1542_n_10566), .o(FE_OFN1547_n_10566) );
in01f08 FE_OFC1548_n_10566 ( .a(FE_OFN1544_n_10566), .o(FE_OFN1548_n_10566) );
in01f04 FE_OFC1549_n_12104 ( .a(n_12104), .o(FE_OFN1549_n_12104) );
in01f02 FE_OFC1550_n_12104 ( .a(n_12104), .o(FE_OFN1550_n_12104) );
in01f02 FE_OFC1551_n_12104 ( .a(FE_OFN1549_n_12104), .o(FE_OFN1551_n_12104) );
in01f06 FE_OFC1552_n_12104 ( .a(FE_OFN1549_n_12104), .o(FE_OFN1552_n_12104) );
in01f06 FE_OFC1553_n_12104 ( .a(FE_OFN1550_n_12104), .o(FE_OFN1553_n_12104) );
in01f06 FE_OFC1554_n_12104 ( .a(FE_OFN1549_n_12104), .o(FE_OFN1554_n_12104) );
in01f06 FE_OFC1556_n_12042 ( .a(FE_OCP_RBN2229_n_15969), .o(FE_OFN1556_n_12042) );
in01f04 FE_OFC1558_n_12042 ( .a(FE_OCP_RBN2229_n_15969), .o(FE_OFN1558_n_12042) );
in01f08 FE_OFC1559_n_12042 ( .a(FE_OFN2203_n_12042), .o(FE_OFN1559_n_12042) );
in01f04 FE_OFC1560_n_12502 ( .a(n_12502), .o(FE_OFN1560_n_12502) );
in01f02 FE_OFC1561_n_12502 ( .a(n_12502), .o(FE_OFN1561_n_12502) );
in01f04 FE_OFC1562_n_12502 ( .a(FE_OFN1561_n_12502), .o(FE_OFN1562_n_12502) );
in01f02 FE_OFC1563_n_12502 ( .a(FE_OFN1560_n_12502), .o(FE_OFN1563_n_12502) );
in01f04 FE_OFC1564_n_12502 ( .a(FE_OFN1561_n_12502), .o(FE_OFN1564_n_12502) );
in01f04 FE_OFC1565_n_12502 ( .a(FE_OFN1560_n_12502), .o(FE_OFN1565_n_12502) );
in01f06 FE_OFC1566_n_12502 ( .a(FE_OFN1560_n_12502), .o(FE_OFN1566_n_12502) );
in01f04 FE_OFC1568_n_11027 ( .a(FE_OCP_RBN2275_n_10268), .o(FE_OFN1568_n_11027) );
in01f04 FE_OFC1572_n_11027 ( .a(FE_OCP_RBN2274_n_10268), .o(FE_OFN1572_n_11027) );
in01f04 FE_OFC1573_n_12028 ( .a(n_12028), .o(FE_OFN1573_n_12028) );
in01f02 FE_OFC1574_n_12028 ( .a(FE_OFN1573_n_12028), .o(FE_OFN1574_n_12028) );
in01f08 FE_OFC1575_n_12028 ( .a(FE_OFN1573_n_12028), .o(FE_OFN1575_n_12028) );
in01f02 FE_OFC1576_n_12028 ( .a(n_12028), .o(FE_OFN1576_n_12028) );
in01f06 FE_OFC1577_n_12028 ( .a(FE_OFN1576_n_12028), .o(FE_OFN1577_n_12028) );
in01f06 FE_OFC1579_n_12306 ( .a(FE_OCP_RBN1928_n_10259), .o(FE_OFN1579_n_12306) );
in01f06 FE_OFC1581_n_12306 ( .a(FE_OCP_RBN1928_n_10259), .o(FE_OFN1581_n_12306) );
in01f06 FE_OFC1583_n_12306 ( .a(FE_OCP_RBN1927_n_10259), .o(FE_OFN1583_n_12306) );
in01f06 FE_OFC1584_n_12306 ( .a(FE_OCP_RBN1926_n_10259), .o(FE_OFN1584_n_12306) );
in01f06 FE_OFC1585_n_13736 ( .a(n_13736), .o(FE_OFN1585_n_13736) );
in01f06 FE_OFC1586_n_13736 ( .a(FE_OFN1585_n_13736), .o(FE_OFN1586_n_13736) );
in01f04 FE_OFC1587_n_13736 ( .a(FE_OFN1585_n_13736), .o(FE_OFN1587_n_13736) );
in01f06 FE_OFC1588_n_13736 ( .a(FE_OFN1585_n_13736), .o(FE_OFN1588_n_13736) );
in01f06 FE_OFC1589_n_13736 ( .a(FE_OFN1585_n_13736), .o(FE_OFN1589_n_13736) );
in01f02 FE_OFC1590_n_13741 ( .a(n_13741), .o(FE_OFN1590_n_13741) );
in01f02 FE_OFC1591_n_13741 ( .a(n_13741), .o(FE_OFN1591_n_13741) );
in01f02 FE_OFC1592_n_13741 ( .a(n_13741), .o(FE_OFN1592_n_13741) );
in01f06 FE_OFC1593_n_13741 ( .a(FE_OFN1590_n_13741), .o(FE_OFN1593_n_13741) );
in01f06 FE_OFC1596_n_13741 ( .a(FE_OFN1592_n_13741), .o(FE_OFN1596_n_13741) );
in01f08 FE_OFC1598_n_13995 ( .a(n_13995), .o(FE_OFN1598_n_13995) );
in01f06 FE_OFC1599_n_13995 ( .a(FE_OFN1598_n_13995), .o(FE_OFN1599_n_13995) );
in01f06 FE_OFC1600_n_13995 ( .a(FE_OFN1598_n_13995), .o(FE_OFN1600_n_13995) );
in01f06 FE_OFC1601_n_13995 ( .a(FE_OFN1598_n_13995), .o(FE_OFN1601_n_13995) );
in01f06 FE_OFC1602_n_13995 ( .a(FE_OFN1598_n_13995), .o(FE_OFN1602_n_13995) );
in01f04 FE_OFC1603_n_13997 ( .a(n_13997), .o(FE_OFN1603_n_13997) );
in01f04 FE_OFC1604_n_13997 ( .a(n_13997), .o(FE_OFN1604_n_13997) );
in01f08 FE_OFC1605_n_13997 ( .a(FE_OFN1603_n_13997), .o(FE_OFN1605_n_13997) );
in01f08 FE_OFC1606_n_13997 ( .a(FE_OFN1604_n_13997), .o(FE_OFN1606_n_13997) );
in01s06 FE_OFC1607_n_2122 ( .a(n_2122), .o(FE_OFN1607_n_2122) );
in01f06 FE_OFC1608_n_2122 ( .a(n_2122), .o(FE_OFN1608_n_2122) );
in01s06 FE_OFC1609_n_2122 ( .a(FE_OFN1607_n_2122), .o(FE_OFN1609_n_2122) );
in01s08 FE_OFC1610_n_2122 ( .a(FE_OFN1607_n_2122), .o(FE_OFN1610_n_2122) );
in01s08 FE_OFC1611_n_2122 ( .a(FE_OFN1608_n_2122), .o(FE_OFN1611_n_2122) );
in01m02 FE_OFC1612_n_2122 ( .a(FE_OFN1608_n_2122), .o(FE_OFN1612_n_2122) );
in01s02 FE_OFC1613_n_1787 ( .a(n_1787), .o(FE_OFN1613_n_1787) );
in01m02 FE_OFC1614_n_1787 ( .a(n_1787), .o(FE_OFN1614_n_1787) );
in01m04 FE_OFC1615_n_1787 ( .a(n_1787), .o(FE_OFN1615_n_1787) );
in01m02 FE_OFC1616_n_1787 ( .a(n_1787), .o(FE_OFN1616_n_1787) );
in01s06 FE_OFC1617_n_1787 ( .a(FE_OFN1613_n_1787), .o(FE_OFN1617_n_1787) );
in01s01 FE_OFC1618_n_1787 ( .a(FE_OFN1614_n_1787), .o(FE_OFN1618_n_1787) );
in01m04 FE_OFC1619_n_1787 ( .a(FE_OFN1614_n_1787), .o(FE_OFN1619_n_1787) );
in01m06 FE_OFC1620_n_1787 ( .a(FE_OFN1615_n_1787), .o(FE_OFN1620_n_1787) );
in01s06 FE_OFC1621_n_1787 ( .a(FE_OFN1616_n_1787), .o(FE_OFN1621_n_1787) );
in01s06 FE_OFC1622_n_4438 ( .a(n_4438), .o(FE_OFN1622_n_4438) );
in01s01 FE_OFC1623_n_4438 ( .a(FE_OFN1622_n_4438), .o(FE_OFN1623_n_4438) );
in01s03 FE_OFC1624_n_4438 ( .a(FE_OFN1622_n_4438), .o(FE_OFN1624_n_4438) );
in01s06 FE_OFC1625_n_4438 ( .a(FE_OFN1622_n_4438), .o(FE_OFN1625_n_4438) );
in01s06 FE_OFC1626_n_4438 ( .a(FE_OFN1622_n_4438), .o(FE_OFN1626_n_4438) );
in01s03 FE_OFC1627_n_4438 ( .a(FE_OFN1626_n_4438), .o(FE_OFN1627_n_4438) );
in01s06 FE_OFC1628_n_4438 ( .a(FE_OFN1627_n_4438), .o(FE_OFN1628_n_4438) );
in01s04 FE_OFC1629_n_9531 ( .a(n_9531), .o(FE_OFN1629_n_9531) );
in01m02 FE_OFC1630_n_9531 ( .a(n_9531), .o(FE_OFN1630_n_9531) );
in01m04 FE_OFC1631_n_9531 ( .a(FE_OFN1630_n_9531), .o(FE_OFN1631_n_9531) );
in01s01 FE_OFC1632_n_9531 ( .a(FE_OFN1630_n_9531), .o(FE_OFN1632_n_9531) );
in01m04 FE_OFC1633_n_9531 ( .a(FE_OFN1631_n_9531), .o(FE_OFN1633_n_9531) );
in01s04 FE_OFC1634_n_9531 ( .a(FE_OFN1633_n_9531), .o(FE_OFN1634_n_9531) );
in01s06 FE_OFC1635_n_9531 ( .a(FE_OFN1633_n_9531), .o(FE_OFN1635_n_9531) );
in01s08 FE_OFC1636_n_4460 ( .a(n_4460), .o(FE_OFN1636_n_4460) );
in01s02 FE_OFC1637_n_4671 ( .a(n_4671), .o(FE_OFN1637_n_4671) );
in01s04 FE_OFC1638_n_4671 ( .a(n_4671), .o(FE_OFN1638_n_4671) );
in01s01 FE_OFC1639_n_4671 ( .a(n_4671), .o(FE_OFN1639_n_4671) );
in01s06 FE_OFC1640_n_4671 ( .a(FE_OFN1638_n_4671), .o(FE_OFN1640_n_4671) );
in01s02 FE_OFC1641_n_4671 ( .a(n_4671), .o(FE_OFN1641_n_4671) );
in01s06 FE_OFC1642_n_4671 ( .a(FE_OFN1637_n_4671), .o(FE_OFN1642_n_4671) );
in01s04 FE_OFC1643_n_4671 ( .a(FE_OFN1639_n_4671), .o(FE_OFN1643_n_4671) );
in01s03 FE_OFC1644_n_4671 ( .a(FE_OFN1641_n_4671), .o(FE_OFN1644_n_4671) );
in01s01 FE_OFC1645_n_4671 ( .a(FE_OFN1641_n_4671), .o(FE_OFN1645_n_4671) );
in01s01 FE_OFC1646_n_9428 ( .a(n_9428), .o(FE_OFN1646_n_9428) );
in01s08 FE_OFC1647_n_9428 ( .a(n_9428), .o(FE_OFN1647_n_9428) );
in01s06 FE_OFC1648_n_9428 ( .a(FE_OFN1647_n_9428), .o(FE_OFN1648_n_9428) );
in01s06 FE_OFC1649_n_9428 ( .a(FE_OFN1647_n_9428), .o(FE_OFN1649_n_9428) );
in01s06 FE_OFC1650_n_9428 ( .a(FE_OFN1647_n_9428), .o(FE_OFN1650_n_9428) );
in01s03 FE_OFC1651_n_9428 ( .a(FE_OFN1647_n_9428), .o(FE_OFN1651_n_9428) );
in01s04 FE_OFC1652_n_9502 ( .a(n_9502), .o(FE_OFN1652_n_9502) );
in01m06 FE_OFC1653_n_9502 ( .a(n_9502), .o(FE_OFN1653_n_9502) );
in01s03 FE_OFC1654_n_9502 ( .a(FE_OFN1653_n_9502), .o(FE_OFN1654_n_9502) );
in01s02 FE_OFC1655_n_9502 ( .a(FE_OFN1653_n_9502), .o(FE_OFN1655_n_9502) );
in01s06 FE_OFC1656_n_9502 ( .a(FE_OFN1653_n_9502), .o(FE_OFN1656_n_9502) );
in01s06 FE_OFC1657_n_9502 ( .a(FE_OFN1653_n_9502), .o(FE_OFN1657_n_9502) );
in01s02 FE_OFC1658_n_4490 ( .a(n_4490), .o(FE_OFN1658_n_4490) );
in01s01 FE_OFC1659_n_4490 ( .a(FE_OFN1658_n_4490), .o(FE_OFN1659_n_4490) );
in01s03 FE_OFC1660_n_4490 ( .a(FE_OFN1658_n_4490), .o(FE_OFN1660_n_4490) );
in01s06 FE_OFC1661_n_4490 ( .a(n_4490), .o(FE_OFN1661_n_4490) );
in01s02 FE_OFC1662_n_4490 ( .a(n_4490), .o(FE_OFN1662_n_4490) );
in01s06 FE_OFC1663_n_4490 ( .a(FE_OFN1662_n_4490), .o(FE_OFN1663_n_4490) );
in01s01 FE_OFC1664_n_9477 ( .a(n_9477), .o(FE_OFN1664_n_9477) );
in01s06 FE_OFC1665_n_9477 ( .a(n_9477), .o(FE_OFN1665_n_9477) );
in01s06 FE_OFC1666_n_9477 ( .a(FE_OFN1665_n_9477), .o(FE_OFN1666_n_9477) );
in01s04 FE_OFC1667_n_9477 ( .a(FE_OFN1665_n_9477), .o(FE_OFN1667_n_9477) );
in01s03 FE_OFC1668_n_9477 ( .a(FE_OFN1665_n_9477), .o(FE_OFN1668_n_9477) );
in01s03 FE_OFC1669_n_9477 ( .a(FE_OFN1667_n_9477), .o(FE_OFN1669_n_9477) );
in01s03 FE_OFC1670_n_9477 ( .a(FE_OFN1669_n_9477), .o(FE_OFN1670_n_9477) );
in01s02 FE_OFC1671_n_9477 ( .a(FE_OFN1669_n_9477), .o(FE_OFN1671_n_9477) );
in01s02 FE_OFC1672_n_4655 ( .a(n_4655), .o(FE_OFN1672_n_4655) );
in01s02 FE_OFC1673_n_4655 ( .a(n_4655), .o(FE_OFN1673_n_4655) );
in01s02 FE_OFC1674_n_4655 ( .a(n_4655), .o(FE_OFN1674_n_4655) );
in01s02 FE_OFC1675_n_4655 ( .a(n_4655), .o(FE_OFN1675_n_4655) );
in01s06 FE_OFC1676_n_4655 ( .a(FE_OFN1673_n_4655), .o(FE_OFN1676_n_4655) );
in01s06 FE_OFC1677_n_4655 ( .a(FE_OFN1674_n_4655), .o(FE_OFN1677_n_4655) );
in01s06 FE_OFC1678_n_4655 ( .a(FE_OFN1675_n_4655), .o(FE_OFN1678_n_4655) );
in01s02 FE_OFC1679_n_4655 ( .a(FE_OFN1672_n_4655), .o(FE_OFN1679_n_4655) );
in01s03 FE_OFC1680_n_4655 ( .a(FE_OFN1672_n_4655), .o(FE_OFN1680_n_4655) );
in01s04 FE_OFC1681_n_4669 ( .a(n_4669), .o(FE_OFN1681_n_4669) );
in01s06 FE_OFC1682_n_4669 ( .a(n_4669), .o(FE_OFN1682_n_4669) );
in01s02 FE_OFC1683_n_9528 ( .a(n_9528), .o(FE_OFN1683_n_9528) );
in01s01 FE_OFC1684_n_9528 ( .a(n_9528), .o(FE_OFN1684_n_9528) );
in01s01 FE_OFC1685_n_9528 ( .a(n_9528), .o(FE_OFN1685_n_9528) );
in01s02 FE_OFC1686_n_9528 ( .a(n_9528), .o(FE_OFN1686_n_9528) );
in01s03 FE_OFC1687_n_9528 ( .a(FE_OFN1684_n_9528), .o(FE_OFN1687_n_9528) );
in01s01 FE_OFC1688_n_9528 ( .a(FE_OFN1686_n_9528), .o(FE_OFN1688_n_9528) );
in01s02 FE_OFC1689_n_9528 ( .a(FE_OFN1686_n_9528), .o(FE_OFN1689_n_9528) );
in01s03 FE_OFC1690_n_9528 ( .a(FE_OFN1685_n_9528), .o(FE_OFN1690_n_9528) );
in01s02 FE_OFC1691_n_9528 ( .a(FE_OFN1686_n_9528), .o(FE_OFN1691_n_9528) );
in01s01 FE_OFC1692_n_9528 ( .a(FE_OFN1686_n_9528), .o(FE_OFN1692_n_9528) );
in01f02 FE_OFC1693_n_3368 ( .a(n_3368), .o(FE_OFN1693_n_3368) );
in01f04 FE_OFC1694_n_3368 ( .a(FE_OFN1693_n_3368), .o(FE_OFN1694_n_3368) );
in01f04 FE_OFC1695_n_3368 ( .a(FE_OFN1693_n_3368), .o(FE_OFN1695_n_3368) );
in01f06 FE_OFC1696_n_5751 ( .a(n_5751), .o(FE_OFN1696_n_5751) );
in01m04 FE_OFC1697_n_5751 ( .a(FE_OFN1696_n_5751), .o(FE_OFN1697_n_5751) );
in01f04 FE_OFC1698_n_5751 ( .a(FE_OFN1696_n_5751), .o(FE_OFN1698_n_5751) );
in01f04 FE_OFC1699_n_5751 ( .a(FE_OFN1696_n_5751), .o(FE_OFN1699_n_5751) );
in01f08 FE_OFC1700_n_5751 ( .a(FE_OFN1696_n_5751), .o(FE_OFN1700_n_5751) );
in01f02 FE_OFC1701_n_4868 ( .a(n_4868), .o(FE_OFN1701_n_4868) );
in01f06 FE_OFC1702_n_4868 ( .a(n_4868), .o(FE_OFN1702_n_4868) );
in01f06 FE_OFC1703_n_4868 ( .a(n_4868), .o(FE_OFN1703_n_4868) );
in01m01 FE_OFC1704_n_4868 ( .a(n_4868), .o(FE_OFN1704_n_4868) );
in01f08 FE_OFC1705_n_4868 ( .a(FE_OFN1701_n_4868), .o(FE_OFN1705_n_4868) );
in01m08 FE_OFC1706_n_4868 ( .a(FE_OFN1703_n_4868), .o(FE_OFN1706_n_4868) );
in01f06 FE_OFC1707_n_4868 ( .a(FE_OFN1703_n_4868), .o(FE_OFN1707_n_4868) );
in01m06 FE_OFC1708_n_4868 ( .a(FE_OFN1704_n_4868), .o(FE_OFN1708_n_4868) );
in01m10 FE_OFC1709_n_4868 ( .a(FE_OFN1702_n_4868), .o(FE_OFN1709_n_4868) );
in01f06 FE_OFC1710_n_4868 ( .a(FE_OFN1702_n_4868), .o(FE_OFN1710_n_4868) );
in01f02 FE_OFC1711_n_13563 ( .a(n_13563), .o(FE_OFN1711_n_13563) );
in01f02 FE_OFC1712_n_13563 ( .a(FE_OFN1711_n_13563), .o(FE_OFN1712_n_13563) );
in01f02 FE_OFC1713_n_13650 ( .a(n_13650), .o(FE_OFN1713_n_13650) );
in01f02 FE_OFC1714_n_13650 ( .a(FE_OFN1713_n_13650), .o(FE_OFN1714_n_13650) );
in01f02 FE_OFC1716_n_16698 ( .a(FE_OCP_RBN2007_n_16698), .o(FE_OFN1716_n_16698) );
in01f04 FE_OFC1719_n_16891 ( .a(n_16891), .o(FE_OFN1719_n_16891) );
in01f08 FE_OFC1720_n_16891 ( .a(FE_OFN1719_n_16891), .o(FE_OFN1720_n_16891) );
in01m02 FE_OFC1721_n_16891 ( .a(n_16891), .o(FE_OFN1721_n_16891) );
in01f02 FE_OFC1722_n_16891 ( .a(n_16891), .o(FE_OFN1722_n_16891) );
in01f02 FE_OFC1723_n_16891 ( .a(FE_OFN1719_n_16891), .o(FE_OFN1723_n_16891) );
in01f06 FE_OFC1724_n_16891 ( .a(FE_OFN1722_n_16891), .o(FE_OFN1724_n_16891) );
in01f06 FE_OFC1725_n_16891 ( .a(FE_OFN1721_n_16891), .o(FE_OFN1725_n_16891) );
in01f04 FE_OFC1726_n_9975 ( .a(n_9975), .o(FE_OFN1726_n_9975) );
in01f08 FE_OFC1727_n_9975 ( .a(FE_OFN1726_n_9975), .o(FE_OFN1727_n_9975) );
in01f02 FE_OFC1728_n_9975 ( .a(FE_OFN1726_n_9975), .o(FE_OFN1728_n_9975) );
in01f04 FE_OFC1729_n_9975 ( .a(n_9975), .o(FE_OFN1729_n_9975) );
in01f06 FE_OFC1730_n_9975 ( .a(FE_OFN1729_n_9975), .o(FE_OFN1730_n_9975) );
in01f08 FE_OFC1731_n_9975 ( .a(FE_OFN1729_n_9975), .o(FE_OFN1731_n_9975) );
in01f06 FE_OFC1732_n_16317 ( .a(n_16317), .o(FE_OFN1732_n_16317) );
in01f02 FE_OFC1733_n_16317 ( .a(FE_OFN1732_n_16317), .o(FE_OFN1733_n_16317) );
in01f06 FE_OFC1734_n_16317 ( .a(FE_OFN1732_n_16317), .o(FE_OFN1734_n_16317) );
in01f06 FE_OFC1735_n_16317 ( .a(FE_OFN1732_n_16317), .o(FE_OFN1735_n_16317) );
in01f04 FE_OFC1736_n_16317 ( .a(FE_OFN1732_n_16317), .o(FE_OFN1736_n_16317) );
in01f06 FE_OFC1737_n_11019 ( .a(n_11019), .o(FE_OFN1737_n_11019) );
in01f02 FE_OFC1738_n_11019 ( .a(FE_OFN1737_n_11019), .o(FE_OFN1738_n_11019) );
in01f06 FE_OFC1739_n_11019 ( .a(FE_OFN1737_n_11019), .o(FE_OFN1739_n_11019) );
in01f01 FE_OFC1740_n_11019 ( .a(FE_OFN1737_n_11019), .o(FE_OFN1740_n_11019) );
in01f04 FE_OFC1741_n_11019 ( .a(FE_OFN1737_n_11019), .o(FE_OFN1741_n_11019) );
in01f04 FE_OFC1742_n_11019 ( .a(FE_OFN1737_n_11019), .o(FE_OFN1742_n_11019) );
in01f02 FE_OFC1743_n_12004 ( .a(n_12004), .o(FE_OFN1743_n_12004) );
in01f02 FE_OFC1744_n_12004 ( .a(n_12004), .o(FE_OFN1744_n_12004) );
in01f04 FE_OFC1745_n_12004 ( .a(n_12004), .o(FE_OFN1745_n_12004) );
in01f04 FE_OFC1746_n_12004 ( .a(FE_OFN1744_n_12004), .o(FE_OFN1746_n_12004) );
in01f04 FE_OFC1747_n_12004 ( .a(FE_OFN1743_n_12004), .o(FE_OFN1747_n_12004) );
in01f04 FE_OFC1748_n_12004 ( .a(FE_OFN1745_n_12004), .o(FE_OFN1748_n_12004) );
in01f08 FE_OFC1749_n_12004 ( .a(FE_OFN1745_n_12004), .o(FE_OFN1749_n_12004) );
in01f02 FE_OFC1751_n_12086 ( .a(FE_OCP_RBN1972_n_11767), .o(FE_OFN1751_n_12086) );
in01f04 FE_OFC1752_n_12086 ( .a(FE_OCP_RBN1972_n_11767), .o(FE_OFN1752_n_12086) );
in01f06 FE_OFC1753_n_12086 ( .a(FE_OCP_RBN1971_n_11767), .o(FE_OFN1753_n_12086) );
in01f04 FE_OFC1754_n_12681 ( .a(n_12681), .o(FE_OFN1754_n_12681) );
in01f02 FE_OFC1755_n_12681 ( .a(FE_OFN1754_n_12681), .o(FE_OFN1755_n_12681) );
in01f02 FE_OFC1756_n_12681 ( .a(FE_OFN1754_n_12681), .o(FE_OFN1756_n_12681) );
in01f08 FE_OFC1757_n_12681 ( .a(FE_OFN1754_n_12681), .o(FE_OFN1757_n_12681) );
in01f06 FE_OFC1758_n_10780 ( .a(n_10780), .o(FE_OFN1758_n_10780) );
in01f06 FE_OFC1759_n_10780 ( .a(FE_OFN1758_n_10780), .o(FE_OFN1759_n_10780) );
in01f06 FE_OFC1760_n_10780 ( .a(FE_OFN1758_n_10780), .o(FE_OFN1760_n_10780) );
in01f04 FE_OFC1761_n_10780 ( .a(FE_OFN1758_n_10780), .o(FE_OFN1761_n_10780) );
in01f06 FE_OFC1762_n_10780 ( .a(FE_OFN1758_n_10780), .o(FE_OFN1762_n_10780) );
in01f06 FE_OFC1767_n_14054 ( .a(n_14054), .o(FE_OFN1767_n_14054) );
in01f06 FE_OFC1768_n_14054 ( .a(FE_OFN1767_n_14054), .o(FE_OFN1768_n_14054) );
in01f06 FE_OFC1769_n_14054 ( .a(FE_OFN1767_n_14054), .o(FE_OFN1769_n_14054) );
in01f06 FE_OFC1770_n_14054 ( .a(FE_OFN1767_n_14054), .o(FE_OFN1770_n_14054) );
in01f06 FE_OFC1771_n_14054 ( .a(FE_OFN1767_n_14054), .o(FE_OFN1771_n_14054) );
in01f03 FE_OFC1773_n_13800 ( .a(FE_OFN1772_n_13800), .o(FE_OFN1773_n_13800) );
in01f06 FE_OFC1775_n_13800 ( .a(FE_OFN1772_n_13800), .o(FE_OFN1775_n_13800) );
in01f20 FE_OFC1776_parchk_pci_ad_reg_in_1222 ( .a(parchk_pci_ad_reg_in_1222), .o(FE_OFN1776_parchk_pci_ad_reg_in_1222) );
in01f08 FE_OFC1777_parchk_pci_ad_reg_in_1222 ( .a(FE_OFN1776_parchk_pci_ad_reg_in_1222), .o(FE_OFN1777_parchk_pci_ad_reg_in_1222) );
in01f03 FE_OFC1778_parchk_pci_ad_reg_in_1222 ( .a(FE_OFN1776_parchk_pci_ad_reg_in_1222), .o(FE_OFN1778_parchk_pci_ad_reg_in_1222) );
in01f20 FE_OFC1779_parchk_pci_ad_reg_in_1221 ( .a(parchk_pci_ad_reg_in_1221), .o(FE_OFN1779_parchk_pci_ad_reg_in_1221) );
in01m03 FE_OFC1780_parchk_pci_ad_reg_in_1221 ( .a(FE_OFN1779_parchk_pci_ad_reg_in_1221), .o(FE_OFN1780_parchk_pci_ad_reg_in_1221) );
in01f08 FE_OFC1781_parchk_pci_ad_reg_in_1221 ( .a(FE_OFN1779_parchk_pci_ad_reg_in_1221), .o(FE_OFN1781_parchk_pci_ad_reg_in_1221) );
in01s04 FE_OFC1782_n_1699 ( .a(n_1699), .o(FE_OFN1782_n_1699) );
in01s06 FE_OFC1783_n_1699 ( .a(FE_OFN1782_n_1699), .o(FE_OFN1783_n_1699) );
in01s02 FE_OFC1784_n_1699 ( .a(FE_OFN1782_n_1699), .o(FE_OFN1784_n_1699) );
in01s01 FE_OFC1785_n_1699 ( .a(FE_OFN1782_n_1699), .o(FE_OFN1785_n_1699) );
in01s02 FE_OFC1786_n_1699 ( .a(FE_OFN1782_n_1699), .o(FE_OFN1786_n_1699) );
in01s02 FE_OFC1789_n_9823 ( .a(FE_OFN530_n_9823), .o(FE_OFN1789_n_9823) );
in01f04 FE_OFC1790_n_2687 ( .a(n_2687), .o(FE_OFN1790_n_2687) );
in01s03 FE_OFC1791_n_9904 ( .a(FE_OFN607_n_9904), .o(FE_OFN1791_n_9904) );
in01s04 FE_OFC1792_n_9904 ( .a(FE_OFN607_n_9904), .o(FE_OFN1792_n_9904) );
in01s03 FE_OFC1793_n_9904 ( .a(FE_OFN1791_n_9904), .o(FE_OFN1793_n_9904) );
in01s03 FE_OFC1794_n_9904 ( .a(FE_OFN1791_n_9904), .o(FE_OFN1794_n_9904) );
in01s06 FE_OFC1795_n_9904 ( .a(FE_OFN1792_n_9904), .o(FE_OFN1795_n_9904) );
in01s03 FE_OFC1796_n_2299 ( .a(FE_OFN958_n_2299), .o(FE_OFN1796_n_2299) );
in01s06 FE_OFC1797_n_2299 ( .a(FE_OFN1796_n_2299), .o(FE_OFN1797_n_2299) );
in01s02 FE_OFC1798_n_9690 ( .a(FE_OFN541_n_9690), .o(FE_OFN1798_n_9690) );
in01s02 FE_OFC1799_n_9690 ( .a(FE_OFN541_n_9690), .o(FE_OFN1799_n_9690) );
in01s01 FE_OFC1800_n_9690 ( .a(FE_OFN1798_n_9690), .o(FE_OFN1800_n_9690) );
in01s03 FE_OFC1801_n_9690 ( .a(FE_OFN1798_n_9690), .o(FE_OFN1801_n_9690) );
in01s01 FE_OFC1802_n_9690 ( .a(FE_OFN1799_n_9690), .o(FE_OFN1802_n_9690) );
in01s03 FE_OFC1803_n_9690 ( .a(FE_OFN1799_n_9690), .o(FE_OFN1803_n_9690) );
in01s02 FE_OFC1804_n_4501 ( .a(FE_OFN613_n_4501), .o(FE_OFN1804_n_4501) );
in01s03 FE_OFC1805_n_4501 ( .a(FE_OFN613_n_4501), .o(FE_OFN1805_n_4501) );
in01s03 FE_OFC1806_n_4501 ( .a(FE_OFN1804_n_4501), .o(FE_OFN1806_n_4501) );
in01s06 FE_OFC1807_n_4501 ( .a(FE_OFN1805_n_4501), .o(FE_OFN1807_n_4501) );
in01s06 FE_OFC1808_n_4454 ( .a(FE_OFN632_n_4454), .o(FE_OFN1808_n_4454) );
in01s03 FE_OFC1809_n_4454 ( .a(FE_OFN1808_n_4454), .o(FE_OFN1809_n_4454) );
in01s06 FE_OFC1810_n_4454 ( .a(FE_OFN1808_n_4454), .o(FE_OFN1810_n_4454) );
in01m01 FE_OFC1811_n_7845 ( .a(FE_OFN700_n_7845), .o(FE_OFN1811_n_7845) );
in01s06 FE_OFC1812_n_7845 ( .a(FE_OFN1811_n_7845), .o(FE_OFN1812_n_7845) );
in01f02 FE_OFC1813_n_2919 ( .a(FE_OFN1819_n_2919), .o(FE_OFN1813_n_2919) );
in01m01 FE_OFC1814_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(FE_OFN1814_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid) );
in01s03 FE_OFC1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid ( .a(FE_OFN1814_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid) );
in01s03 FE_OFC1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid ( .a(FE_OFN1814_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid) );
in01f02 FE_OFC1819_n_2919 ( .a(n_2919), .o(FE_OFN1819_n_2919) );
in01f01 FE_OFC186_n_15768 ( .a(FE_OFN1503_n_15768), .o(FE_OFN186_n_15768) );
in01m02 FE_OFC190_n_1193 ( .a(n_1193), .o(FE_OFN190_n_1193) );
in01m04 FE_OFC191_n_1193 ( .a(FE_OFN190_n_1193), .o(FE_OFN191_n_1193) );
in01s02 FE_OFC1935_n_1781 ( .a(n_1781), .o(FE_OFN1935_n_1781) );
in01s02 FE_OFC1936_n_1781 ( .a(FE_OFN1935_n_1781), .o(FE_OFN1936_n_1781) );
in01s01 FE_OFC1937_g66085_p ( .a(g66085_p), .o(FE_OFN1937_g66085_p) );
in01s03 FE_OFC1938_g66085_p ( .a(FE_OFN1937_g66085_p), .o(FE_OFN1938_g66085_p) );
in01s01 FE_OFC1939_g66095_p ( .a(g66095_p), .o(FE_OFN1939_g66095_p) );
in01s03 FE_OFC1940_g66095_p ( .a(FE_OFN1939_g66095_p), .o(FE_OFN1940_g66095_p) );
in01f02 FE_OFC1941_n_3241 ( .a(n_3241), .o(FE_OFN1941_n_3241) );
in01f02 FE_OFC1942_n_3241 ( .a(FE_OFN1941_n_3241), .o(FE_OFN1942_n_3241) );
in01f02 FE_OFC1943_n_15813 ( .a(n_15813), .o(FE_OFN1943_n_15813) );
in01f02 FE_OFC1944_n_15813 ( .a(FE_OFN1943_n_15813), .o(FE_OFN1944_n_15813) );
in01m10 FE_OFC1945_n_13784 ( .a(n_13784), .o(FE_OFN1945_n_13784) );
in01f10 FE_OFC1946_n_13784 ( .a(FE_OFN1945_n_13784), .o(FE_OFN1946_n_13784) );
in01s01 FE_OFC196_n_2683 ( .a(n_2683), .o(FE_OFN196_n_2683) );
in01s02 FE_OFC197_n_2683 ( .a(FE_OFN196_n_2683), .o(FE_OFN197_n_2683) );
in01s02 FE_OFC198_n_3298 ( .a(n_3298), .o(FE_OFN198_n_3298) );
in01s02 FE_OFC199_n_3298 ( .a(FE_OFN198_n_3298), .o(FE_OFN199_n_3298) );
in01s04 FE_OFC1_n_4778 ( .a(FE_OFN1079_n_4778), .o(FE_OFN1_n_4778) );
in01s01 FE_OFC200_n_9230 ( .a(n_9230), .o(FE_OFN200_n_9230) );
in01s06 FE_OFC201_n_9230 ( .a(FE_OFN200_n_9230), .o(FE_OFN201_n_9230) );
in01s06 FE_OFC2020_n_4778 ( .a(FE_OFN1079_n_4778), .o(FE_OFN2020_n_4778) );
in01s08 FE_OFC2021_n_4778 ( .a(FE_OFN2020_n_4778), .o(FE_OFN2021_n_4778) );
in01s06 FE_OFC2022_n_4778 ( .a(FE_OFN2020_n_4778), .o(FE_OFN2022_n_4778) );
in01s02 FE_OFC202_n_9228 ( .a(n_9228), .o(FE_OFN202_n_9228) );
in01s06 FE_OFC203_n_9228 ( .a(FE_OFN202_n_9228), .o(FE_OFN203_n_9228) );
in01s02 FE_OFC204_n_9140 ( .a(n_9140), .o(FE_OFN204_n_9140) );
in01m02 FE_OFC2051_n_6965 ( .a(n_6965), .o(FE_OFN2051_n_6965) );
in01m02 FE_OFC2052_n_6965 ( .a(FE_OFN2051_n_6965), .o(FE_OFN2052_n_6965) );
in01s20 FE_OFC2053_n_8831 ( .a(n_8831), .o(FE_OFN2053_n_8831) );
in01s20 FE_OFC2054_n_8831 ( .a(FE_OFN2053_n_8831), .o(FE_OFN2054_n_8831) );
in01s08 FE_OFC2055_n_8831 ( .a(FE_OFN2053_n_8831), .o(FE_OFN2055_n_8831) );
in01s02 FE_OFC2056_n_2117 ( .a(n_2117), .o(FE_OFN2056_n_2117) );
in01s01 FE_OFC2057_n_2117 ( .a(FE_OFN2056_n_2117), .o(FE_OFN2057_n_2117) );
in01m08 FE_OFC2058_n_13447 ( .a(n_13447), .o(FE_OFN2058_n_13447) );
in01m08 FE_OFC2059_n_13447 ( .a(FE_OFN2058_n_13447), .o(FE_OFN2059_n_13447) );
in01s06 FE_OFC205_n_9140 ( .a(FE_OFN204_n_9140), .o(FE_OFN205_n_9140) );
in01s01 FE_OFC2060_g66087_p ( .a(g66087_p), .o(FE_OFN2060_g66087_p) );
in01s03 FE_OFC2061_g66087_p ( .a(FE_OFN2060_g66087_p), .o(FE_OFN2061_g66087_p) );
in01m08 FE_OFC2062_n_6391 ( .a(FE_OFN1223_n_6391), .o(FE_OFN2062_n_6391) );
in01s08 FE_OFC2063_n_6391 ( .a(FE_OFN2062_n_6391), .o(FE_OFN2063_n_6391) );
in01m08 FE_OFC2064_n_6391 ( .a(FE_OFN2062_n_6391), .o(FE_OFN2064_n_6391) );
in01s04 FE_OFC2069_n_15978 ( .a(FE_OFN1000_n_15978), .o(FE_OFN2069_n_15978) );
in01s02 FE_OFC206_n_9865 ( .a(n_9865), .o(FE_OFN206_n_9865) );
in01s02 FE_OFC2070_n_15978 ( .a(FE_OFN2069_n_15978), .o(FE_OFN2070_n_15978) );
in01s08 FE_OFC2071_n_15978 ( .a(FE_OFN1001_n_15978), .o(FE_OFN2071_n_15978) );
in01m03 FE_OFC2072_n_15978 ( .a(FE_OFN2071_n_15978), .o(FE_OFN2072_n_15978) );
in01m02 FE_OFC2073_n_2723 ( .a(n_2723), .o(FE_OFN2073_n_2723) );
in01m02 FE_OFC2074_n_2723 ( .a(FE_OFN2073_n_2723), .o(FE_OFN2074_n_2723) );
in01m06 FE_OFC2075_FE_OCPUNCON1952_FE_OFN697_n_16760 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(FE_OFN2075_FE_OCPUNCON1952_FE_OFN697_n_16760) );
in01m08 FE_OFC2076_FE_OCPUNCON1952_FE_OFN697_n_16760 ( .a(FE_OFN2075_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760) );
in01s08 FE_OFC2077_n_8069 ( .a(n_8069), .o(FE_OFN2077_n_8069) );
in01s08 FE_OFC2079_n_8069 ( .a(FE_OFN2077_n_8069), .o(FE_OFN2079_n_8069) );
in01s06 FE_OFC207_n_9865 ( .a(FE_OFN206_n_9865), .o(FE_OFN207_n_9865) );
in01s03 FE_OFC2080_n_8176 ( .a(n_8176), .o(FE_OFN2080_n_8176) );
in01s06 FE_OFC2081_n_8176 ( .a(FE_OFN2080_n_8176), .o(FE_OFN2081_n_8176) );
in01s06 FE_OFC2082_n_8407 ( .a(n_8407), .o(FE_OFN2082_n_8407) );
in01s04 FE_OFC2083_n_8407 ( .a(FE_OFN2082_n_8407), .o(FE_OFN2083_n_8407) );
in01s06 FE_OFC2084_n_8407 ( .a(FE_OFN2082_n_8407), .o(FE_OFN2084_n_8407) );
in01s01 FE_OFC2085_n_8448 ( .a(n_8448), .o(FE_OFN2085_n_8448) );
in01s02 FE_OFC2086_n_8448 ( .a(FE_OFN2085_n_8448), .o(FE_OFN2086_n_8448) );
in01s02 FE_OFC2088_n_13124 ( .a(FE_OFN2132_n_13124), .o(FE_OFN2088_n_13124) );
in01s01 FE_OFC208_n_9126 ( .a(n_9126), .o(FE_OFN208_n_9126) );
in01f10 FE_OFC2092_n_2301 ( .a(n_2301), .o(FE_OFN2092_n_2301) );
in01f10 FE_OFC2093_n_2301 ( .a(FE_OFN2092_n_2301), .o(FE_OFN2093_n_2301) );
in01s02 FE_OFC2094_n_2520 ( .a(n_2520), .o(FE_OFN2094_n_2520) );
in01s01 FE_OFC2095_n_2520 ( .a(FE_OFN2094_n_2520), .o(FE_OFN2095_n_2520) );
in01s01 FE_OFC2096_n_2520 ( .a(FE_OFN2094_n_2520), .o(FE_OFN2096_n_2520) );
in01m02 FE_OFC2099_n_3281 ( .a(n_3281), .o(FE_OFN2099_n_3281) );
in01s06 FE_OFC209_n_9126 ( .a(FE_OFN208_n_9126), .o(FE_OFN209_n_9126) );
in01m02 FE_OFC2100_n_3281 ( .a(FE_OFN2099_n_3281), .o(FE_OFN2100_n_3281) );
in01f02 FE_OFC2101_n_2834 ( .a(n_2834), .o(FE_OFN2101_n_2834) );
in01f02 FE_OFC2102_n_2834 ( .a(FE_OFN2101_n_2834), .o(FE_OFN2102_n_2834) );
in01m08 FE_OFC2103_g64577_p ( .a(FE_OFN1106_g64577_p), .o(FE_OFN2103_g64577_p) );
in01s06 FE_OFC2104_g64577_p ( .a(FE_OFN2103_g64577_p), .o(FE_OFN2104_g64577_p) );
in01s10 FE_OFC2105_g64577_p ( .a(FE_OFN2103_g64577_p), .o(FE_OFN2105_g64577_p) );
in01s06 FE_OFC2106_g64577_p ( .a(FE_OFN2103_g64577_p), .o(FE_OFN2106_g64577_p) );
in01m01 FE_OFC2107_n_2047 ( .a(FE_OFN1003_n_2047), .o(FE_OFN2107_n_2047) );
in01s06 FE_OFC2108_n_2047 ( .a(FE_OFN2107_n_2047), .o(FE_OFN2108_n_2047) );
in01s03 FE_OFC2109_n_2047 ( .a(FE_OFN2107_n_2047), .o(FE_OFN2109_n_2047) );
in01s02 FE_OFC210_n_9858 ( .a(n_9858), .o(FE_OFN210_n_9858) );
in01m01 FE_OFC2110_n_2248 ( .a(FE_OFN945_n_2248), .o(FE_OFN2110_n_2248) );
in01s06 FE_OFC2111_n_2248 ( .a(FE_OFN2110_n_2248), .o(FE_OFN2111_n_2248) );
in01s03 FE_OFC2112_n_2053 ( .a(FE_OFN1016_n_2053), .o(FE_OFN2112_n_2053) );
in01s06 FE_OFC2113_n_2053 ( .a(FE_OFN2112_n_2053), .o(FE_OFN2113_n_2053) );
in01s06 FE_OFC2114_wishbone_slave_unit_pci_initiator_if_data_source ( .a(wishbone_slave_unit_pci_initiator_if_data_source), .o(FE_OFN2114_wishbone_slave_unit_pci_initiator_if_data_source) );
in01m03 FE_OFC2115_wishbone_slave_unit_pci_initiator_if_data_source ( .a(wishbone_slave_unit_pci_initiator_if_data_source), .o(FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source) );
in01s06 FE_OFC2116_wishbone_slave_unit_pci_initiator_if_data_source ( .a(FE_OFN2114_wishbone_slave_unit_pci_initiator_if_data_source), .o(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source) );
in01s06 FE_OFC2118_wishbone_slave_unit_pci_initiator_if_data_source ( .a(FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source), .o(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source) );
in01s03 FE_OFC2119_wishbone_slave_unit_pci_initiator_if_data_source ( .a(FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source), .o(FE_OFN2119_wishbone_slave_unit_pci_initiator_if_data_source) );
in01s06 FE_OFC211_n_9858 ( .a(FE_OFN210_n_9858), .o(FE_OFN211_n_9858) );
in01f08 FE_OFC2121_n_2687 ( .a(FE_OFN1790_n_2687), .o(FE_OFN2121_n_2687) );
in01f08 FE_OFC2123_n_16497 ( .a(n_16497), .o(FE_OFN2123_n_16497) );
in01f06 FE_OFC2124_n_16497 ( .a(n_16497), .o(FE_OFN2124_n_16497) );
in01f04 FE_OFC2125_n_16497 ( .a(FE_OFN2124_n_16497), .o(FE_OFN2125_n_16497) );
in01f08 FE_OFC2126_n_16497 ( .a(FE_OFN2123_n_16497), .o(FE_OFN2126_n_16497) );
in01f08 FE_OFC2127_n_16497 ( .a(FE_OFN2124_n_16497), .o(FE_OFN2127_n_16497) );
in01f08 FE_OFC2128_n_16497 ( .a(FE_OFN2123_n_16497), .o(FE_OFN2128_n_16497) );
in01f04 FE_OFC2129_n_16720 ( .a(FE_OFN1060_n_16720), .o(FE_OFN2129_n_16720) );
in01m02 FE_OFC212_n_9124 ( .a(n_9124), .o(FE_OFN212_n_9124) );
in01f08 FE_OFC2130_n_10588 ( .a(FE_OFN1451_n_10588), .o(FE_OFN2130_n_10588) );
in01f06 FE_OFC2131_n_10588 ( .a(FE_OFN1451_n_10588), .o(FE_OFN2131_n_10588) );
in01m01 FE_OFC2132_n_13124 ( .a(FE_OFN1304_n_13124), .o(FE_OFN2132_n_13124) );
in01f08 FE_OFC2133_n_13124 ( .a(FE_OFN1304_n_13124), .o(FE_OFN2133_n_13124) );
in01f10 FE_OFC2134_n_13124 ( .a(FE_OFN2133_n_13124), .o(FE_OFN2134_n_13124) );
in01f06 FE_OFC2135_n_13124 ( .a(FE_OFN2133_n_13124), .o(FE_OFN2135_n_13124) );
in01f06 FE_OFC2136_n_13124 ( .a(FE_OFN2133_n_13124), .o(FE_OFN2136_n_13124) );
in01f08 FE_OFC2137_n_15534 ( .a(FE_OFN1481_n_15534), .o(FE_OFN2137_n_15534) );
in01f04 FE_OFC2139_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2139_n_16992) );
in01s06 FE_OFC213_n_9124 ( .a(FE_OFN212_n_9124), .o(FE_OFN213_n_9124) );
in01f01 FE_OFC2140_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2140_n_16992) );
in01f01 FE_OFC2141_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2141_n_16992) );
in01f08 FE_OFC2142_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2142_n_16992) );
in01f01 FE_OFC2143_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2143_n_16992) );
in01f01 FE_OFC2144_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2144_n_16992) );
in01f01 FE_OFC2145_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2145_n_16992) );
in01f06 FE_OFC2146_n_9320 ( .a(FE_OFN1488_n_9320), .o(FE_OFN2146_n_9320) );
in01f06 FE_OFC2147_n_10595 ( .a(FE_OFN1540_n_10595), .o(FE_OFN2147_n_10595) );
in01f01 FE_OFC2148_n_10595 ( .a(FE_OFN1540_n_10595), .o(FE_OFN2148_n_10595) );
in01f06 FE_OFC2149_n_10595 ( .a(FE_OFN1541_n_10595), .o(FE_OFN2149_n_10595) );
in01s02 FE_OFC214_n_9856 ( .a(n_9856), .o(FE_OFN214_n_9856) );
in01f06 FE_OFC2150_n_10595 ( .a(FE_OFN1541_n_10595), .o(FE_OFN2150_n_10595) );
in01f08 FE_OFC2151_n_16439 ( .a(FE_OFN1337_n_16439), .o(FE_OFN2151_n_16439) );
in01f02 FE_OFC2152_n_16439 ( .a(FE_OFN1337_n_16439), .o(FE_OFN2152_n_16439) );
in01f10 FE_OFC2153_n_16439 ( .a(FE_OFN2151_n_16439), .o(FE_OFN2153_n_16439) );
in01f06 FE_OFC2154_n_16439 ( .a(FE_OFN1337_n_16439), .o(FE_OFN2154_n_16439) );
in01f06 FE_OFC2155_n_16439 ( .a(FE_OFN2151_n_16439), .o(FE_OFN2155_n_16439) );
in01f06 FE_OFC2156_n_16439 ( .a(FE_OFN2152_n_16439), .o(FE_OFN2156_n_16439) );
in01f08 FE_OFC2157_n_16439 ( .a(FE_OFN2154_n_16439), .o(FE_OFN2157_n_16439) );
in01f06 FE_OFC2158_n_16439 ( .a(FE_OFN2154_n_16439), .o(FE_OFN2158_n_16439) );
in01f08 FE_OFC2159_n_16301 ( .a(n_16301), .o(FE_OFN2159_n_16301) );
in01s06 FE_OFC215_n_9856 ( .a(FE_OFN214_n_9856), .o(FE_OFN215_n_9856) );
in01f08 FE_OFC2160_n_16301 ( .a(n_16301), .o(FE_OFN2160_n_16301) );
in01f04 FE_OFC2161_n_16301 ( .a(n_16301), .o(FE_OFN2161_n_16301) );
in01f08 FE_OFC2162_n_16301 ( .a(FE_OFN2159_n_16301), .o(FE_OFN2162_n_16301) );
in01f08 FE_OFC2163_n_16301 ( .a(FE_OFN2161_n_16301), .o(FE_OFN2163_n_16301) );
in01f10 FE_OFC2164_n_16301 ( .a(FE_OFN2159_n_16301), .o(FE_OFN2164_n_16301) );
in01f10 FE_OFC2165_n_16301 ( .a(FE_OFN2160_n_16301), .o(FE_OFN2165_n_16301) );
in01f08 FE_OFC2166_n_8567 ( .a(FE_OFN1372_n_8567), .o(FE_OFN2166_n_8567) );
in01f08 FE_OFC2167_n_8567 ( .a(FE_OFN2166_n_8567), .o(FE_OFN2167_n_8567) );
in01f08 FE_OFC2168_n_8567 ( .a(FE_OFN2166_n_8567), .o(FE_OFN2168_n_8567) );
in01f08 FE_OFC2169_n_8567 ( .a(FE_OFN2166_n_8567), .o(FE_OFN2169_n_8567) );
in01s02 FE_OFC216_n_9889 ( .a(n_9889), .o(FE_OFN216_n_9889) );
in01f08 FE_OFC2170_n_8567 ( .a(FE_OFN2166_n_8567), .o(FE_OFN2170_n_8567) );
in01f08 FE_OFC2171_n_8567 ( .a(FE_OFN1373_n_8567), .o(FE_OFN2171_n_8567) );
in01f03 FE_OFC2172_n_8567 ( .a(FE_OFN1373_n_8567), .o(FE_OFN2172_n_8567) );
in01f08 FE_OFC2173_n_8567 ( .a(FE_OFN2171_n_8567), .o(FE_OFN2173_n_8567) );
in01f08 FE_OFC2174_n_8567 ( .a(FE_OFN2171_n_8567), .o(FE_OFN2174_n_8567) );
in01f06 FE_OFC2175_n_8567 ( .a(FE_OFN2172_n_8567), .o(FE_OFN2175_n_8567) );
in01f10 FE_OFC2176_n_8567 ( .a(FE_OFN1378_n_8567), .o(FE_OFN2176_n_8567) );
in01f10 FE_OFC2177_n_8567 ( .a(FE_OFN2176_n_8567), .o(FE_OFN2177_n_8567) );
in01f04 FE_OFC2178_n_8567 ( .a(FE_OFN2176_n_8567), .o(FE_OFN2178_n_8567) );
in01f08 FE_OFC2179_n_8567 ( .a(FE_OFN2176_n_8567), .o(FE_OFN2179_n_8567) );
in01s06 FE_OFC217_n_9889 ( .a(FE_OFN216_n_9889), .o(FE_OFN217_n_9889) );
in01f08 FE_OFC2180_n_8567 ( .a(FE_OFN2176_n_8567), .o(FE_OFN2180_n_8567) );
in01f10 FE_OFC2181_n_8567 ( .a(FE_OFN1394_n_8567), .o(FE_OFN2181_n_8567) );
in01f10 FE_OFC2182_n_8567 ( .a(FE_OFN2181_n_8567), .o(FE_OFN2182_n_8567) );
in01f08 FE_OFC2183_n_8567 ( .a(FE_OFN1394_n_8567), .o(FE_OFN2183_n_8567) );
in01f10 FE_OFC2184_n_8567 ( .a(FE_OFN2183_n_8567), .o(FE_OFN2184_n_8567) );
in01f10 FE_OFC2185_n_8567 ( .a(FE_OFN2181_n_8567), .o(FE_OFN2185_n_8567) );
in01f10 FE_OFC2186_n_8567 ( .a(FE_OFN1410_n_8567), .o(FE_OFN2186_n_8567) );
in01f08 FE_OFC2187_n_8567 ( .a(FE_OFN2186_n_8567), .o(FE_OFN2187_n_8567) );
in01f08 FE_OFC2188_n_8567 ( .a(FE_OFN2186_n_8567), .o(FE_OFN2188_n_8567) );
in01f04 FE_OFC2189_n_8567 ( .a(FE_OFN2186_n_8567), .o(FE_OFN2189_n_8567) );
in01s01 FE_OFC218_n_9853 ( .a(n_9853), .o(FE_OFN218_n_9853) );
in01f06 FE_OFC2190_n_8567 ( .a(FE_OFN2186_n_8567), .o(FE_OFN2190_n_8567) );
in01f08 FE_OFC2191_n_8567 ( .a(FE_OFN2186_n_8567), .o(FE_OFN2191_n_8567) );
in01f06 FE_OFC2192_n_16779 ( .a(FE_OFN1430_n_16779), .o(FE_OFN2192_n_16779) );
in01f06 FE_OFC2193_n_9163 ( .a(FE_OFN1447_n_9163), .o(FE_OFN2193_n_9163) );
in01f08 FE_OFC2194_n_9163 ( .a(FE_OFN1447_n_9163), .o(FE_OFN2194_n_9163) );
in01f02 FE_OFC2195_n_9163 ( .a(FE_OFN1447_n_9163), .o(FE_OFN2195_n_9163) );
in01f01 FE_OFC2196_n_9163 ( .a(FE_OFN1447_n_9163), .o(FE_OFN2196_n_9163) );
in01f10 FE_OFC2197_n_10256 ( .a(n_10256), .o(FE_OFN2197_n_10256) );
in01f10 FE_OFC2198_n_10256 ( .a(FE_OFN2197_n_10256), .o(FE_OFN2198_n_10256) );
in01f08 FE_OFC2199_n_10256 ( .a(n_10256), .o(FE_OFN2199_n_10256) );
in01s06 FE_OFC219_n_9853 ( .a(FE_OFN218_n_9853), .o(FE_OFN219_n_9853) );
in01m02 FE_OFC21_n_9372 ( .a(FE_OFN1434_n_9372), .o(FE_OFN21_n_9372) );
in01f10 FE_OFC2200_n_10256 ( .a(FE_OFN2199_n_10256), .o(FE_OFN2200_n_10256) );
in01f02 FE_OFC2201_n_12042 ( .a(n_15969), .o(FE_OFN2201_n_12042) );
in01f04 FE_OFC2202_n_12042 ( .a(n_15969), .o(FE_OFN2202_n_12042) );
in01f04 FE_OFC2203_n_12042 ( .a(FE_OFN2201_n_12042), .o(FE_OFN2203_n_12042) );
in01f01 FE_OFC2204_n_12028 ( .a(FE_OFN1576_n_12028), .o(FE_OFN2204_n_12028) );
in01f06 FE_OFC2205_n_10538 ( .a(FE_OFN1514_n_10538), .o(FE_OFN2205_n_10538) );
in01f02 FE_OFC2206_n_10892 ( .a(FE_OFN1520_n_10892), .o(FE_OFN2206_n_10892) );
in01f04 FE_OFC2207_n_10892 ( .a(FE_OFN1520_n_10892), .o(FE_OFN2207_n_10892) );
in01f06 FE_OFC2208_n_11795 ( .a(FE_OFN1459_n_11795), .o(FE_OFN2208_n_11795) );
in01f06 FE_OFC2209_n_11027 ( .a(FE_OCP_RBN2274_n_10268), .o(FE_OFN2209_n_11027) );
in01m02 FE_OFC220_n_9846 ( .a(n_9846), .o(FE_OFN220_n_9846) );
in01f04 FE_OFC2210_n_11027 ( .a(FE_OCP_RBN2274_n_10268), .o(FE_OFN2210_n_11027) );
in01s06 FE_OFC2211_n_8407 ( .a(FE_OFN2083_n_8407), .o(FE_OFN2211_n_8407) );
in01s08 FE_OFC2212_n_8407 ( .a(FE_OFN2211_n_8407), .o(FE_OFN2212_n_8407) );
in01s01 FE_OFC2213_n_15366 ( .a(FE_OFN995_n_15366), .o(FE_OFN2213_n_15366) );
in01f10 FE_OFC2214_n_15366 ( .a(FE_OFN995_n_15366), .o(FE_OFN2214_n_15366) );
in01s01 FE_OFC2215_n_15366 ( .a(FE_OFN2213_n_15366), .o(FE_OFN2215_n_15366) );
in01f06 FE_OFC2216_n_10143 ( .a(FE_OFN1531_n_10143), .o(FE_OFN2216_n_10143) );
in01s06 FE_OFC221_n_9846 ( .a(FE_OFN220_n_9846), .o(FE_OFN221_n_9846) );
in01s02 FE_OFC222_n_9844 ( .a(n_9844), .o(FE_OFN222_n_9844) );
in01s06 FE_OFC223_n_9844 ( .a(FE_OFN222_n_9844), .o(FE_OFN223_n_9844) );
in01f08 FE_OFC2240_g52675_p ( .a(FE_OFN1470_g52675_p), .o(FE_OFN2240_g52675_p) );
in01f03 FE_OFC2241_g52675_p ( .a(FE_OFN2240_g52675_p), .o(FE_OFN2241_g52675_p) );
in01f06 FE_OFC2242_g52675_p ( .a(FE_OFN2240_g52675_p), .o(FE_OFN2242_g52675_p) );
in01f10 FE_OFC2243_g52675_p ( .a(FE_OFN2240_g52675_p), .o(FE_OFN2243_g52675_p) );
in01m02 FE_OFC2244_n_4792 ( .a(n_4792), .o(FE_OFN2244_n_4792) );
in01s04 FE_OFC2245_n_4792 ( .a(FE_OFN2244_n_4792), .o(FE_OFN2245_n_4792) );
in01s01 FE_OFC2246_n_2113 ( .a(n_2113), .o(FE_OFN2246_n_2113) );
in01s01 FE_OFC2247_n_2113 ( .a(FE_OFN2246_n_2113), .o(FE_OFN2247_n_2113) );
in01s02 FE_OFC2248_n_1790 ( .a(n_1790), .o(FE_OFN2248_n_1790) );
in01s01 FE_OFC2249_n_1790 ( .a(FE_OFN2248_n_1790), .o(FE_OFN2249_n_1790) );
in01s02 FE_OFC224_n_9122 ( .a(n_9122), .o(FE_OFN224_n_9122) );
in01s02 FE_OFC2250_n_2101 ( .a(n_2101), .o(FE_OFN2250_n_2101) );
in01s02 FE_OFC2251_n_2101 ( .a(FE_OFN2250_n_2101), .o(FE_OFN2251_n_2101) );
in01s02 FE_OFC2252_n_9687 ( .a(FE_OFN602_n_9687), .o(FE_OFN2252_n_9687) );
in01s01 FE_OFC2253_n_9687 ( .a(FE_OFN2252_n_9687), .o(FE_OFN2253_n_9687) );
in01s01 FE_OFC2254_n_9687 ( .a(FE_OFN2252_n_9687), .o(FE_OFN2254_n_9687) );
in01s06 FE_OFC2255_n_8060 ( .a(n_8060), .o(FE_OFN2255_n_8060) );
in01s03 FE_OFC2256_n_8060 ( .a(FE_OFN2255_n_8060), .o(FE_OFN2256_n_8060) );
in01s04 FE_OFC2257_n_8060 ( .a(FE_OFN2255_n_8060), .o(FE_OFN2257_n_8060) );
in01s06 FE_OFC2258_n_8060 ( .a(FE_OFN2255_n_8060), .o(FE_OFN2258_n_8060) );
in01f02 FE_OFC2259_n_2775 ( .a(n_2775), .o(FE_OFN2259_n_2775) );
in01s06 FE_OFC225_n_9122 ( .a(FE_OFN224_n_9122), .o(FE_OFN225_n_9122) );
in01f02 FE_OFC2260_n_2775 ( .a(FE_OFN2259_n_2775), .o(FE_OFN2260_n_2775) );
in01m02 FE_OFC226_n_9841 ( .a(n_9841), .o(FE_OFN226_n_9841) );
in01s06 FE_OFC227_n_9841 ( .a(FE_OFN226_n_9841), .o(FE_OFN227_n_9841) );
in01s02 FE_OFC228_n_9120 ( .a(n_9120), .o(FE_OFN228_n_9120) );
in01s06 FE_OFC229_n_9120 ( .a(FE_OFN228_n_9120), .o(FE_OFN229_n_9120) );
in01s02 FE_OFC230_n_9839 ( .a(n_9839), .o(FE_OFN230_n_9839) );
in01s06 FE_OFC231_n_9839 ( .a(FE_OFN230_n_9839), .o(FE_OFN231_n_9839) );
in01m02 FE_OFC232_n_9876 ( .a(n_9876), .o(FE_OFN232_n_9876) );
in01s06 FE_OFC233_n_9876 ( .a(FE_OFN232_n_9876), .o(FE_OFN233_n_9876) );
in01m02 FE_OFC234_n_9834 ( .a(n_9834), .o(FE_OFN234_n_9834) );
in01s06 FE_OFC235_n_9834 ( .a(FE_OFN234_n_9834), .o(FE_OFN235_n_9834) );
in01s01 FE_OFC236_n_9118 ( .a(n_9118), .o(FE_OFN236_n_9118) );
in01s06 FE_OFC237_n_9118 ( .a(FE_OFN236_n_9118), .o(FE_OFN237_n_9118) );
in01m02 FE_OFC238_n_9832 ( .a(n_9832), .o(FE_OFN238_n_9832) );
in01s06 FE_OFC239_n_9832 ( .a(FE_OFN238_n_9832), .o(FE_OFN239_n_9832) );
in01s02 FE_OFC240_n_9830 ( .a(n_9830), .o(FE_OFN240_n_9830) );
in01s06 FE_OFC241_n_9830 ( .a(FE_OFN240_n_9830), .o(FE_OFN241_n_9830) );
in01m02 FE_OFC242_n_9116 ( .a(n_9116), .o(FE_OFN242_n_9116) );
in01s06 FE_OFC243_n_9116 ( .a(FE_OFN242_n_9116), .o(FE_OFN243_n_9116) );
in01s02 FE_OFC244_n_9114 ( .a(n_9114), .o(FE_OFN244_n_9114) );
in01s06 FE_OFC245_n_9114 ( .a(FE_OFN244_n_9114), .o(FE_OFN245_n_9114) );
in01s02 FE_OFC246_n_9112 ( .a(n_9112), .o(FE_OFN246_n_9112) );
in01s06 FE_OFC247_n_9112 ( .a(FE_OFN246_n_9112), .o(FE_OFN247_n_9112) );
in01s01 FE_OFC248_n_9789 ( .a(n_9789), .o(FE_OFN248_n_9789) );
in01s06 FE_OFC250_n_9789 ( .a(FE_OFN248_n_9789), .o(FE_OFN250_n_9789) );
in01s02 FE_OFC251_n_9868 ( .a(n_9868), .o(FE_OFN251_n_9868) );
in01s06 FE_OFC252_n_9868 ( .a(FE_OFN251_n_9868), .o(FE_OFN252_n_9868) );
in01s02 FE_OFC253_n_9825 ( .a(n_9825), .o(FE_OFN253_n_9825) );
in01s06 FE_OFC254_n_9825 ( .a(FE_OFN253_n_9825), .o(FE_OFN254_n_9825) );
in01s02 FE_OFC255_n_8969 ( .a(n_8969), .o(FE_OFN255_n_8969) );
in01s06 FE_OFC256_n_8969 ( .a(FE_OFN255_n_8969), .o(FE_OFN256_n_8969) );
in01m02 FE_OFC257_n_9862 ( .a(n_9862), .o(FE_OFN257_n_9862) );
in01s08 FE_OFC258_n_9862 ( .a(FE_OFN257_n_9862), .o(FE_OFN258_n_9862) );
in01s02 FE_OFC259_n_9860 ( .a(n_9860), .o(FE_OFN259_n_9860) );
in01s06 FE_OFC260_n_9860 ( .a(FE_OFN259_n_9860), .o(FE_OFN260_n_9860) );
in01m02 FE_OFC261_n_9851 ( .a(n_9851), .o(FE_OFN261_n_9851) );
in01s08 FE_OFC262_n_9851 ( .a(FE_OFN261_n_9851), .o(FE_OFN262_n_9851) );
in01m02 FE_OFC263_n_9849 ( .a(n_9849), .o(FE_OFN263_n_9849) );
in01s08 FE_OFC264_n_9849 ( .a(FE_OFN263_n_9849), .o(FE_OFN264_n_9849) );
in01s02 FE_OFC265_n_9884 ( .a(n_9884), .o(FE_OFN265_n_9884) );
in01s06 FE_OFC266_n_9884 ( .a(FE_OFN265_n_9884), .o(FE_OFN266_n_9884) );
in01m02 FE_OFC267_n_9880 ( .a(n_9880), .o(FE_OFN267_n_9880) );
in01s06 FE_OFC268_n_9880 ( .a(FE_OFN267_n_9880), .o(FE_OFN268_n_9880) );
in01s02 FE_OFC269_n_9836 ( .a(n_9836), .o(FE_OFN269_n_9836) );
in01s06 FE_OFC270_n_9836 ( .a(FE_OFN269_n_9836), .o(FE_OFN270_n_9836) );
in01s02 FE_OFC271_n_9828 ( .a(n_9828), .o(FE_OFN271_n_9828) );
in01s06 FE_OFC272_n_9828 ( .a(FE_OFN271_n_9828), .o(FE_OFN272_n_9828) );
in01m04 FE_OFC275_n_9941 ( .a(n_9941), .o(FE_OFN275_n_9941) );
in01m08 FE_OFC276_n_9941 ( .a(FE_OFN275_n_9941), .o(FE_OFN276_n_9941) );
in01s06 FE_OFC2_n_4778 ( .a(FE_OFN1_n_4778), .o(FE_OFN2_n_4778) );
in01s01 FE_OFC334_g66081_p ( .a(g66081_p), .o(FE_OFN334_g66081_p) );
in01s03 FE_OFC335_g66081_p ( .a(FE_OFN334_g66081_p), .o(FE_OFN335_g66081_p) );
in01s01 FE_OFC336_g66089_p ( .a(g66089_p), .o(FE_OFN336_g66089_p) );
in01s03 FE_OFC337_g66089_p ( .a(FE_OFN336_g66089_p), .o(FE_OFN337_g66089_p) );
in01s01 FE_OFC365_n_4093 ( .a(FE_OFN1245_n_4093), .o(FE_OFN365_n_4093) );
in01s01 FE_OFC369_n_4092 ( .a(FE_OFN1237_n_4092), .o(FE_OFN369_n_4092) );
in01s01 FE_OFC3_n_4778 ( .a(FE_OFN1_n_4778), .o(FE_OFN3_n_4778) );
in01s06 FE_OFC514_n_9697 ( .a(n_9697), .o(FE_OFN514_n_9697) );
in01s03 FE_OFC515_n_9697 ( .a(FE_OFN514_n_9697), .o(FE_OFN515_n_9697) );
in01s03 FE_OFC516_n_9697 ( .a(FE_OFN514_n_9697), .o(FE_OFN516_n_9697) );
in01s06 FE_OFC517_n_9697 ( .a(FE_OFN514_n_9697), .o(FE_OFN517_n_9697) );
in01s03 FE_OFC518_n_9697 ( .a(FE_OFN514_n_9697), .o(FE_OFN518_n_9697) );
in01s03 FE_OFC519_n_9697 ( .a(FE_OFN514_n_9697), .o(FE_OFN519_n_9697) );
in01s03 FE_OFC523_n_9428 ( .a(FE_OFN1646_n_9428), .o(FE_OFN523_n_9428) );
in01s06 FE_OFC524_n_9899 ( .a(n_9899), .o(FE_OFN524_n_9899) );
in01s02 FE_OFC525_n_9899 ( .a(FE_OFN524_n_9899), .o(FE_OFN525_n_9899) );
in01s02 FE_OFC526_n_9899 ( .a(FE_OFN524_n_9899), .o(FE_OFN526_n_9899) );
in01s10 FE_OFC527_n_9899 ( .a(FE_OFN524_n_9899), .o(FE_OFN527_n_9899) );
in01m02 FE_OFC528_n_9899 ( .a(FE_OFN524_n_9899), .o(FE_OFN528_n_9899) );
in01s03 FE_OFC529_n_9899 ( .a(FE_OFN524_n_9899), .o(FE_OFN529_n_9899) );
in01s06 FE_OFC530_n_9823 ( .a(n_9823), .o(FE_OFN530_n_9823) );
in01s02 FE_OFC531_n_9823 ( .a(FE_OFN530_n_9823), .o(FE_OFN531_n_9823) );
in01s02 FE_OFC532_n_9823 ( .a(FE_OFN530_n_9823), .o(FE_OFN532_n_9823) );
in01s06 FE_OFC533_n_9823 ( .a(FE_OFN530_n_9823), .o(FE_OFN533_n_9823) );
in01s02 FE_OFC534_n_9823 ( .a(FE_OFN530_n_9823), .o(FE_OFN534_n_9823) );
in01s08 FE_OFC535_n_9823 ( .a(FE_OFN530_n_9823), .o(FE_OFN535_n_9823) );
in01s04 FE_OFC537_n_9690 ( .a(n_9690), .o(FE_OFN537_n_9690) );
in01s02 FE_OFC539_n_9690 ( .a(FE_OFN537_n_9690), .o(FE_OFN539_n_9690) );
in01s02 FE_OFC540_n_9690 ( .a(FE_OFN537_n_9690), .o(FE_OFN540_n_9690) );
in01s04 FE_OFC541_n_9690 ( .a(FE_OFN537_n_9690), .o(FE_OFN541_n_9690) );
in01s02 FE_OFC542_n_9690 ( .a(FE_OFN537_n_9690), .o(FE_OFN542_n_9690) );
in01s02 FE_OFC543_n_9690 ( .a(FE_OFN537_n_9690), .o(FE_OFN543_n_9690) );
in01s02 FE_OFC548_n_9477 ( .a(FE_OFN1664_n_9477), .o(FE_OFN548_n_9477) );
in01s01 FE_OFC549_n_9864 ( .a(n_9864), .o(FE_OFN549_n_9864) );
in01m04 FE_OFC550_n_9864 ( .a(n_9864), .o(FE_OFN550_n_9864) );
in01s02 FE_OFC551_n_9864 ( .a(FE_OFN549_n_9864), .o(FE_OFN551_n_9864) );
in01s01 FE_OFC552_n_9864 ( .a(FE_OFN549_n_9864), .o(FE_OFN552_n_9864) );
in01s02 FE_OFC553_n_9864 ( .a(FE_OFN550_n_9864), .o(FE_OFN553_n_9864) );
in01s06 FE_OFC554_n_9864 ( .a(FE_OFN550_n_9864), .o(FE_OFN554_n_9864) );
in01s06 FE_OFC555_n_9864 ( .a(FE_OFN550_n_9864), .o(FE_OFN555_n_9864) );
in01s02 FE_OFC556_n_9864 ( .a(FE_OFN550_n_9864), .o(FE_OFN556_n_9864) );
in01s01 FE_OFC557_n_9895 ( .a(n_9895), .o(FE_OFN557_n_9895) );
in01s04 FE_OFC558_n_9895 ( .a(n_9895), .o(FE_OFN558_n_9895) );
in01s01 FE_OFC559_n_9895 ( .a(FE_OFN557_n_9895), .o(FE_OFN559_n_9895) );
in01s02 FE_OFC560_n_9895 ( .a(FE_OFN557_n_9895), .o(FE_OFN560_n_9895) );
in01s02 FE_OFC561_n_9895 ( .a(FE_OFN558_n_9895), .o(FE_OFN561_n_9895) );
in01s08 FE_OFC562_n_9895 ( .a(FE_OFN558_n_9895), .o(FE_OFN562_n_9895) );
in01s03 FE_OFC563_n_9895 ( .a(FE_OFN558_n_9895), .o(FE_OFN563_n_9895) );
in01s03 FE_OFC564_n_9895 ( .a(FE_OFN558_n_9895), .o(FE_OFN564_n_9895) );
in01s03 FE_OFC568_n_9528 ( .a(FE_OFN1683_n_9528), .o(FE_OFN568_n_9528) );
in01s03 FE_OFC569_n_9528 ( .a(FE_OFN1683_n_9528), .o(FE_OFN569_n_9528) );
in01s08 FE_OFC572_n_9502 ( .a(FE_OFN1652_n_9502), .o(FE_OFN572_n_9502) );
in01s06 FE_OFC573_n_9902 ( .a(n_9902), .o(FE_OFN573_n_9902) );
in01s04 FE_OFC574_n_9902 ( .a(FE_OFN573_n_9902), .o(FE_OFN574_n_9902) );
in01s03 FE_OFC575_n_9902 ( .a(FE_OFN573_n_9902), .o(FE_OFN575_n_9902) );
in01s04 FE_OFC576_n_9902 ( .a(FE_OFN573_n_9902), .o(FE_OFN576_n_9902) );
in01s08 FE_OFC577_n_9902 ( .a(FE_OFN573_n_9902), .o(FE_OFN577_n_9902) );
in01s03 FE_OFC579_n_9531 ( .a(FE_OFN1629_n_9531), .o(FE_OFN579_n_9531) );
in01s08 FE_OFC580_n_9531 ( .a(FE_OFN1629_n_9531), .o(FE_OFN580_n_9531) );
in01s04 FE_OFC582_n_9692 ( .a(n_9692), .o(FE_OFN582_n_9692) );
in01s01 FE_OFC583_n_9692 ( .a(n_9692), .o(FE_OFN583_n_9692) );
in01s04 FE_OFC584_n_9692 ( .a(FE_OFN582_n_9692), .o(FE_OFN584_n_9692) );
in01s03 FE_OFC585_n_9692 ( .a(FE_OFN583_n_9692), .o(FE_OFN585_n_9692) );
in01s06 FE_OFC587_n_9692 ( .a(FE_OFN582_n_9692), .o(FE_OFN587_n_9692) );
in01s04 FE_OFC588_n_9692 ( .a(FE_OFN582_n_9692), .o(FE_OFN588_n_9692) );
in01s02 FE_OFC589_n_9692 ( .a(FE_OFN582_n_9692), .o(FE_OFN589_n_9692) );
in01s06 FE_OFC590_n_9694 ( .a(n_9694), .o(FE_OFN590_n_9694) );
in01s01 FE_OFC591_n_9694 ( .a(n_9694), .o(FE_OFN591_n_9694) );
in01s02 FE_OFC592_n_9694 ( .a(FE_OFN590_n_9694), .o(FE_OFN592_n_9694) );
in01s02 FE_OFC593_n_9694 ( .a(FE_OFN591_n_9694), .o(FE_OFN593_n_9694) );
in01s08 FE_OFC595_n_9694 ( .a(FE_OFN590_n_9694), .o(FE_OFN595_n_9694) );
in01s03 FE_OFC596_n_9694 ( .a(FE_OFN590_n_9694), .o(FE_OFN596_n_9694) );
in01s02 FE_OFC597_n_9694 ( .a(FE_OFN590_n_9694), .o(FE_OFN597_n_9694) );
in01s04 FE_OFC598_n_9687 ( .a(n_9687), .o(FE_OFN598_n_9687) );
in01s01 FE_OFC599_n_9687 ( .a(n_9687), .o(FE_OFN599_n_9687) );
in01s03 FE_OFC600_n_9687 ( .a(FE_OFN598_n_9687), .o(FE_OFN600_n_9687) );
in01s06 FE_OFC601_n_9687 ( .a(FE_OFN598_n_9687), .o(FE_OFN601_n_9687) );
in01s06 FE_OFC602_n_9687 ( .a(FE_OFN598_n_9687), .o(FE_OFN602_n_9687) );
in01s02 FE_OFC603_n_9687 ( .a(FE_OFN599_n_9687), .o(FE_OFN603_n_9687) );
in01s06 FE_OFC605_n_9904 ( .a(n_9904), .o(FE_OFN605_n_9904) );
in01s08 FE_OFC606_n_9904 ( .a(FE_OFN605_n_9904), .o(FE_OFN606_n_9904) );
in01s06 FE_OFC607_n_9904 ( .a(FE_OFN605_n_9904), .o(FE_OFN607_n_9904) );
in01s01 FE_OFC608_n_9904 ( .a(FE_OFN605_n_9904), .o(FE_OFN608_n_9904) );
in01s06 FE_OFC611_n_4501 ( .a(n_4501), .o(FE_OFN611_n_4501) );
in01s06 FE_OFC612_n_4501 ( .a(FE_OFN611_n_4501), .o(FE_OFN612_n_4501) );
in01s03 FE_OFC613_n_4501 ( .a(FE_OFN611_n_4501), .o(FE_OFN613_n_4501) );
in01s03 FE_OFC614_n_4501 ( .a(FE_OFN611_n_4501), .o(FE_OFN614_n_4501) );
in01s06 FE_OFC615_n_4501 ( .a(FE_OFN611_n_4501), .o(FE_OFN615_n_4501) );
in01s06 FE_OFC618_n_4490 ( .a(FE_OFN1661_n_4490), .o(FE_OFN618_n_4490) );
in01s03 FE_OFC619_n_4490 ( .a(FE_OFN1661_n_4490), .o(FE_OFN619_n_4490) );
in01s03 FE_OFC620_n_4490 ( .a(FE_OFN1661_n_4490), .o(FE_OFN620_n_4490) );
in01s04 FE_OFC621_n_4409 ( .a(n_4409), .o(FE_OFN621_n_4409) );
in01s03 FE_OFC622_n_4409 ( .a(FE_OFN621_n_4409), .o(FE_OFN622_n_4409) );
in01s02 FE_OFC623_n_4409 ( .a(FE_OFN621_n_4409), .o(FE_OFN623_n_4409) );
in01s06 FE_OFC624_n_4409 ( .a(FE_OFN621_n_4409), .o(FE_OFN624_n_4409) );
in01s06 FE_OFC625_n_4409 ( .a(FE_OFN621_n_4409), .o(FE_OFN625_n_4409) );
in01m06 FE_OFC627_n_4454 ( .a(n_4454), .o(FE_OFN627_n_4454) );
in01s01 FE_OFC628_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN628_n_4454) );
in01s01 FE_OFC629_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN629_n_4454) );
in01s03 FE_OFC630_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN630_n_4454) );
in01s03 FE_OFC631_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN631_n_4454) );
in01s04 FE_OFC632_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN632_n_4454) );
in01s01 FE_OFC633_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN633_n_4454) );
in01s03 FE_OFC634_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN634_n_4454) );
in01s06 FE_OFC636_n_4669 ( .a(FE_OFN1682_n_4669), .o(FE_OFN636_n_4669) );
in01s01 FE_OFC638_n_4669 ( .a(FE_OFN1682_n_4669), .o(FE_OFN638_n_4669) );
in01s06 FE_OFC639_n_4669 ( .a(FE_OFN1682_n_4669), .o(FE_OFN639_n_4669) );
in01s08 FE_OFC640_n_4669 ( .a(FE_OFN1681_n_4669), .o(FE_OFN640_n_4669) );
in01s06 FE_OFC641_n_4677 ( .a(n_4677), .o(FE_OFN641_n_4677) );
in01s06 FE_OFC642_n_4677 ( .a(FE_OFN641_n_4677), .o(FE_OFN642_n_4677) );
in01s06 FE_OFC643_n_4677 ( .a(FE_OFN641_n_4677), .o(FE_OFN643_n_4677) );
in01s06 FE_OFC644_n_4677 ( .a(FE_OFN641_n_4677), .o(FE_OFN644_n_4677) );
in01s06 FE_OFC645_n_4497 ( .a(n_4497), .o(FE_OFN645_n_4497) );
in01s03 FE_OFC646_n_4497 ( .a(FE_OFN645_n_4497), .o(FE_OFN646_n_4497) );
in01s06 FE_OFC647_n_4497 ( .a(FE_OFN645_n_4497), .o(FE_OFN647_n_4497) );
in01s06 FE_OFC648_n_4497 ( .a(FE_OFN645_n_4497), .o(FE_OFN648_n_4497) );
in01s06 FE_OFC649_n_4497 ( .a(FE_OFN645_n_4497), .o(FE_OFN649_n_4497) );
in01s08 FE_OFC650_n_4508 ( .a(n_4508), .o(FE_OFN650_n_4508) );
in01s06 FE_OFC651_n_4508 ( .a(FE_OFN650_n_4508), .o(FE_OFN651_n_4508) );
in01s06 FE_OFC652_n_4508 ( .a(FE_OFN650_n_4508), .o(FE_OFN652_n_4508) );
in01s06 FE_OFC653_n_4508 ( .a(FE_OFN650_n_4508), .o(FE_OFN653_n_4508) );
in01s06 FE_OFC654_n_4508 ( .a(FE_OFN650_n_4508), .o(FE_OFN654_n_4508) );
in01s06 FE_OFC658_n_4392 ( .a(n_4392), .o(FE_OFN658_n_4392) );
in01s06 FE_OFC659_n_4392 ( .a(FE_OFN658_n_4392), .o(FE_OFN659_n_4392) );
in01s06 FE_OFC660_n_4392 ( .a(FE_OFN658_n_4392), .o(FE_OFN660_n_4392) );
in01s06 FE_OFC661_n_4392 ( .a(FE_OFN658_n_4392), .o(FE_OFN661_n_4392) );
in01s06 FE_OFC662_n_4392 ( .a(FE_OFN658_n_4392), .o(FE_OFN662_n_4392) );
in01s06 FE_OFC663_n_4495 ( .a(n_4495), .o(FE_OFN663_n_4495) );
in01s03 FE_OFC664_n_4495 ( .a(FE_OFN663_n_4495), .o(FE_OFN664_n_4495) );
in01s06 FE_OFC665_n_4495 ( .a(FE_OFN663_n_4495), .o(FE_OFN665_n_4495) );
in01s06 FE_OFC666_n_4495 ( .a(FE_OFN663_n_4495), .o(FE_OFN666_n_4495) );
in01s06 FE_OFC667_n_4495 ( .a(FE_OFN663_n_4495), .o(FE_OFN667_n_4495) );
in01m06 FE_OFC668_n_4505 ( .a(n_4505), .o(FE_OFN668_n_4505) );
in01s04 FE_OFC669_n_4505 ( .a(FE_OFN668_n_4505), .o(FE_OFN669_n_4505) );
in01s06 FE_OFC670_n_4505 ( .a(FE_OFN668_n_4505), .o(FE_OFN670_n_4505) );
in01s06 FE_OFC671_n_4505 ( .a(FE_OFN668_n_4505), .o(FE_OFN671_n_4505) );
in01s03 FE_OFC672_n_4505 ( .a(FE_OFN668_n_4505), .o(FE_OFN672_n_4505) );
in01s01 FE_OFC678_n_4460 ( .a(FE_OFN1636_n_4460), .o(FE_OFN678_n_4460) );
in01s06 FE_OFC679_n_4460 ( .a(FE_OFN1636_n_4460), .o(FE_OFN679_n_4460) );
in01s06 FE_OFC681_n_4460 ( .a(FE_OFN1636_n_4460), .o(FE_OFN681_n_4460) );
in01s06 FE_OFC682_n_4460 ( .a(FE_OFN1636_n_4460), .o(FE_OFN682_n_4460) );
in01s08 FE_OFC683_n_4417 ( .a(n_4417), .o(FE_OFN683_n_4417) );
in01s02 FE_OFC684_n_4417 ( .a(FE_OFN683_n_4417), .o(FE_OFN684_n_4417) );
in01s06 FE_OFC685_n_4417 ( .a(FE_OFN683_n_4417), .o(FE_OFN685_n_4417) );
in01s06 FE_OFC686_n_4417 ( .a(FE_OFN683_n_4417), .o(FE_OFN686_n_4417) );
in01s06 FE_OFC687_n_4417 ( .a(FE_OFN683_n_4417), .o(FE_OFN687_n_4417) );
in01s02 FE_OFC689_n_4438 ( .a(FE_OFN1622_n_4438), .o(FE_OFN689_n_4438) );
in01f01 FE_OFC697_n_16760 ( .a(FE_OFN1026_n_16760), .o(FE_OFN697_n_16760) );
in01s08 FE_OFC698_n_7845 ( .a(n_7845), .o(FE_OFN698_n_7845) );
in01s06 FE_OFC699_n_7845 ( .a(FE_OFN698_n_7845), .o(FE_OFN699_n_7845) );
in01s04 FE_OFC700_n_7845 ( .a(FE_OFN698_n_7845), .o(FE_OFN700_n_7845) );
in01s03 FE_OFC701_n_7845 ( .a(FE_OFN698_n_7845), .o(FE_OFN701_n_7845) );
in01s06 FE_OFC702_n_7845 ( .a(FE_OFN698_n_7845), .o(FE_OFN702_n_7845) );
in01s03 FE_OFC703_n_8069 ( .a(n_8069), .o(FE_OFN703_n_8069) );
in01s06 FE_OFC704_n_8069 ( .a(FE_OFN703_n_8069), .o(FE_OFN704_n_8069) );
in01s06 FE_OFC705_n_8119 ( .a(n_8119), .o(FE_OFN705_n_8119) );
in01s06 FE_OFC706_n_8119 ( .a(FE_OFN705_n_8119), .o(FE_OFN706_n_8119) );
in01s06 FE_OFC707_n_8119 ( .a(FE_OFN705_n_8119), .o(FE_OFN707_n_8119) );
in01s06 FE_OFC708_n_8232 ( .a(n_8232), .o(FE_OFN708_n_8232) );
in01s06 FE_OFC709_n_8232 ( .a(FE_OFN708_n_8232), .o(FE_OFN709_n_8232) );
in01s06 FE_OFC710_n_8232 ( .a(FE_OFN708_n_8232), .o(FE_OFN710_n_8232) );
in01s08 FE_OFC711_n_8140 ( .a(n_8140), .o(FE_OFN711_n_8140) );
in01s06 FE_OFC712_n_8140 ( .a(FE_OFN711_n_8140), .o(FE_OFN712_n_8140) );
in01s06 FE_OFC713_n_8140 ( .a(FE_OFN711_n_8140), .o(FE_OFN713_n_8140) );
in01s06 FE_OFC714_n_8140 ( .a(FE_OFN711_n_8140), .o(FE_OFN714_n_8140) );
in01s06 FE_OFC715_n_8176 ( .a(n_8176), .o(FE_OFN715_n_8176) );
in01s06 FE_OFC716_n_8176 ( .a(FE_OFN715_n_8176), .o(FE_OFN716_n_8176) );
in01s06 FE_OFC717_n_8176 ( .a(FE_OFN715_n_8176), .o(FE_OFN717_n_8176) );
in01s08 FE_OFC718_n_8060 ( .a(FE_OFN2258_n_8060), .o(FE_OFN718_n_8060) );
in01s06 FE_OFC719_n_8060 ( .a(FE_OFN718_n_8060), .o(FE_OFN719_n_8060) );
in01s06 FE_OFC720_n_8060 ( .a(FE_OFN718_n_8060), .o(FE_OFN720_n_8060) );
in01m06 FE_OFC732_n_7498 ( .a(FE_OFN1156_n_7498), .o(FE_OFN732_n_7498) );
in01s03 FE_OFC775_n_15366 ( .a(FE_OFN2215_n_15366), .o(FE_OFN775_n_15366) );
in01s03 FE_OFC776_n_15366 ( .a(FE_OFN2215_n_15366), .o(FE_OFN776_n_15366) );
in01s02 FE_OFC777_n_4152 ( .a(n_4152), .o(FE_OFN777_n_4152) );
in01s06 FE_OFC778_n_4152 ( .a(FE_OFN777_n_4152), .o(FE_OFN778_n_4152) );
in01s01 FE_OFC779_n_2746 ( .a(n_2746), .o(FE_OFN779_n_2746) );
in01s02 FE_OFC780_n_2746 ( .a(FE_OFN779_n_2746), .o(FE_OFN780_n_2746) );
in01s01 FE_OFC781_n_2746 ( .a(FE_OFN779_n_2746), .o(FE_OFN781_n_2746) );
in01m04 FE_OFC782_n_2678 ( .a(n_2678), .o(FE_OFN782_n_2678) );
in01m01 FE_OFC783_n_2678 ( .a(n_2678), .o(FE_OFN783_n_2678) );
in01s04 FE_OFC784_n_2678 ( .a(FE_OFN782_n_2678), .o(FE_OFN784_n_2678) );
in01s08 FE_OFC785_n_2678 ( .a(FE_OFN782_n_2678), .o(FE_OFN785_n_2678) );
in01s04 FE_OFC786_n_2678 ( .a(FE_OFN782_n_2678), .o(FE_OFN786_n_2678) );
in01s02 FE_OFC787_n_2678 ( .a(FE_OFN783_n_2678), .o(FE_OFN787_n_2678) );
in01s04 FE_OFC789_n_2678 ( .a(FE_OFN782_n_2678), .o(FE_OFN789_n_2678) );
in01s01 FE_OFC792_n_2547 ( .a(n_2547), .o(FE_OFN792_n_2547) );
in01s01 FE_OFC793_n_2547 ( .a(FE_OFN792_n_2547), .o(FE_OFN793_n_2547) );
in01s01 FE_OFC794_n_2520 ( .a(n_2520), .o(FE_OFN794_n_2520) );
in01s02 FE_OFC795_n_2520 ( .a(FE_OFN794_n_2520), .o(FE_OFN795_n_2520) );
in01s06 FE_OFC877_g64577_p ( .a(FE_OFN1099_g64577_p), .o(FE_OFN877_g64577_p) );
in01s03 FE_OFC881_g64577_p ( .a(FE_OFN1086_g64577_p), .o(FE_OFN881_g64577_p) );
in01s06 FE_OFC882_g64577_p ( .a(FE_OFN1098_g64577_p), .o(FE_OFN882_g64577_p) );
in01m04 FE_OFC8_n_11877 ( .a(FE_OFN1020_n_11877), .o(FE_OFN8_n_11877) );
in01s01 FE_OFC900_n_4736 ( .a(n_4736), .o(FE_OFN900_n_4736) );
in01s06 FE_OFC901_n_4736 ( .a(n_4736), .o(FE_OFN901_n_4736) );
in01s01 FE_OFC902_n_4736 ( .a(FE_OFN900_n_4736), .o(FE_OFN902_n_4736) );
in01s02 FE_OFC903_n_4736 ( .a(FE_OFN900_n_4736), .o(FE_OFN903_n_4736) );
in01s03 FE_OFC904_n_4736 ( .a(FE_OFN901_n_4736), .o(FE_OFN904_n_4736) );
in01s06 FE_OFC905_n_4736 ( .a(FE_OFN901_n_4736), .o(FE_OFN905_n_4736) );
in01s06 FE_OFC906_n_4736 ( .a(FE_OFN901_n_4736), .o(FE_OFN906_n_4736) );
in01s03 FE_OFC908_n_4734 ( .a(FE_OFN1007_n_4734), .o(FE_OFN908_n_4734) );
in01s04 FE_OFC912_n_4727 ( .a(FE_OFN1052_n_4727), .o(FE_OFN912_n_4727) );
in01s08 FE_OFC915_n_4725 ( .a(n_4725), .o(FE_OFN915_n_4725) );
in01s04 FE_OFC916_n_4725 ( .a(FE_OFN915_n_4725), .o(FE_OFN916_n_4725) );
in01s06 FE_OFC917_n_4725 ( .a(FE_OFN915_n_4725), .o(FE_OFN917_n_4725) );
in01s06 FE_OFC918_n_4725 ( .a(FE_OFN915_n_4725), .o(FE_OFN918_n_4725) );
in01s04 FE_OFC923_n_4740 ( .a(FE_OFN1072_n_4740), .o(FE_OFN923_n_4740) );
in01s06 FE_OFC926_n_4730 ( .a(n_4730), .o(FE_OFN926_n_4730) );
in01s03 FE_OFC927_n_4730 ( .a(FE_OFN926_n_4730), .o(FE_OFN927_n_4730) );
in01s06 FE_OFC928_n_4730 ( .a(FE_OFN926_n_4730), .o(FE_OFN928_n_4730) );
in01s04 FE_OFC929_n_4730 ( .a(FE_OFN926_n_4730), .o(FE_OFN929_n_4730) );
in01s04 FE_OFC930_n_4730 ( .a(FE_OFN926_n_4730), .o(FE_OFN930_n_4730) );
in01s06 FE_OFC934_n_2292 ( .a(n_2292), .o(FE_OFN934_n_2292) );
in01s03 FE_OFC935_n_2292 ( .a(FE_OFN934_n_2292), .o(FE_OFN935_n_2292) );
in01s06 FE_OFC936_n_2292 ( .a(FE_OFN934_n_2292), .o(FE_OFN936_n_2292) );
in01s03 FE_OFC937_n_2292 ( .a(FE_OFN934_n_2292), .o(FE_OFN937_n_2292) );
in01s03 FE_OFC938_n_2292 ( .a(FE_OFN934_n_2292), .o(FE_OFN938_n_2292) );
in01s03 FE_OFC941_n_2047 ( .a(FE_OFN1002_n_2047), .o(FE_OFN941_n_2047) );
in01s06 FE_OFC944_n_2248 ( .a(n_2248), .o(FE_OFN944_n_2248) );
in01s06 FE_OFC945_n_2248 ( .a(FE_OFN944_n_2248), .o(FE_OFN945_n_2248) );
in01s03 FE_OFC946_n_2248 ( .a(FE_OFN944_n_2248), .o(FE_OFN946_n_2248) );
in01s06 FE_OFC947_n_2248 ( .a(FE_OFN2111_n_2248), .o(FE_OFN947_n_2248) );
in01s06 FE_OFC948_n_2248 ( .a(FE_OFN947_n_2248), .o(FE_OFN948_n_2248) );
in01s06 FE_OFC949_n_2055 ( .a(n_2055), .o(FE_OFN949_n_2055) );
in01s06 FE_OFC950_n_2055 ( .a(FE_OFN949_n_2055), .o(FE_OFN950_n_2055) );
in01s06 FE_OFC951_n_2055 ( .a(FE_OFN949_n_2055), .o(FE_OFN951_n_2055) );
in01s03 FE_OFC952_n_2055 ( .a(FE_OFN949_n_2055), .o(FE_OFN952_n_2055) );
in01s06 FE_OFC953_n_2055 ( .a(FE_OFN949_n_2055), .o(FE_OFN953_n_2055) );
in01s06 FE_OFC954_n_1699 ( .a(FE_OFN1783_n_1699), .o(FE_OFN954_n_1699) );
in01s06 FE_OFC955_n_1699 ( .a(FE_OFN954_n_1699), .o(FE_OFN955_n_1699) );
in01s06 FE_OFC956_n_1699 ( .a(FE_OFN954_n_1699), .o(FE_OFN956_n_1699) );
in01s06 FE_OFC957_n_2299 ( .a(n_2299), .o(FE_OFN957_n_2299) );
in01s01 FE_OFC958_n_2299 ( .a(FE_OFN957_n_2299), .o(FE_OFN958_n_2299) );
in01s06 FE_OFC959_n_2299 ( .a(FE_OFN957_n_2299), .o(FE_OFN959_n_2299) );
in01m02 FE_OFC966_n_2233 ( .a(n_2233), .o(FE_OFN966_n_2233) );
in01s02 FE_OFC967_n_2233 ( .a(FE_OFN966_n_2233), .o(FE_OFN967_n_2233) );
in01f08 FE_OFC968_n_13784 ( .a(FE_OFN1946_n_13784), .o(FE_OFN968_n_13784) );
in01f10 FE_OFC969_n_13784 ( .a(FE_OFN968_n_13784), .o(FE_OFN969_n_13784) );
in01m02 FE_OFC982_n_2700 ( .a(n_2700), .o(FE_OFN982_n_2700) );
in01s02 FE_OFC983_n_2700 ( .a(FE_OFN982_n_2700), .o(FE_OFN983_n_2700) );
in01s02 FE_OFC984_n_2697 ( .a(n_2697), .o(FE_OFN984_n_2697) );
in01s03 FE_OFC985_n_2697 ( .a(FE_OFN984_n_2697), .o(FE_OFN985_n_2697) );
in01s02 FE_OFC986_n_2696 ( .a(n_2696), .o(FE_OFN986_n_2696) );
in01s02 FE_OFC987_n_2696 ( .a(FE_OFN986_n_2696), .o(FE_OFN987_n_2696) );
in01s04 FE_OFC988_n_574 ( .a(n_574), .o(FE_OFN988_n_574) );
in01s06 FE_OFC989_n_574 ( .a(FE_OFN988_n_574), .o(FE_OFN989_n_574) );
in01s02 FE_OFC991_n_2373 ( .a(n_2373), .o(FE_OFN991_n_2373) );
in01s02 FE_OFC992_n_2373 ( .a(FE_OFN991_n_2373), .o(FE_OFN992_n_2373) );
in01f06 FE_OFC994_n_15366 ( .a(FE_OFN993_n_15366), .o(FE_OFN994_n_15366) );
in01f08 FE_OFC995_n_15366 ( .a(FE_OFN994_n_15366), .o(FE_OFN995_n_15366) );
in01f08 FE_OFC996_n_15366 ( .a(FE_OFN993_n_15366), .o(FE_OFN996_n_15366) );
in01m03 FE_OFC999_n_15978 ( .a(FE_OFN997_n_15978), .o(FE_OFN999_n_15978) );
in01m02 FE_OFC9_n_11877 ( .a(FE_OFN1020_n_11877), .o(FE_OFN9_n_11877) );
in01f20 FE_RC_0_0 ( .a(pci_target_unit_wishbone_master_first_data_is_burst_reg), .o(FE_RN_0_0) );
in01f06 FE_RC_1000_0 ( .a(n_3078), .o(FE_RN_695_0) );
oa12f02 FE_RC_1002_0 ( .a(FE_RN_694_0), .b(FE_RN_695_0), .c(FE_RN_693_0), .o(FE_RN_697_0) );
na02f04 FE_RC_1003_0 ( .a(n_2835), .b(n_419), .o(FE_RN_698_0) );
oa12f02 FE_RC_1004_0 ( .a(FE_RN_698_0), .b(n_2835), .c(n_419), .o(FE_RN_699_0) );
no02f02 FE_RC_1005_0 ( .a(FE_RN_697_0), .b(FE_RN_699_0), .o(FE_RN_700_0) );
na02f02 FE_RC_1006_0 ( .a(FE_RN_691_0), .b(FE_RN_700_0), .o(FE_RN_701_0) );
no02f02 FE_RC_1007_0 ( .a(FE_RN_684_0), .b(FE_RN_701_0), .o(FE_RN_702_0) );
na02s02 TIMEBOOST_cell_43007 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__Q), .b(g58301_sb), .o(TIMEBOOST_net_13742) );
na02s01 TIMEBOOST_cell_39534 ( .a(TIMEBOOST_net_12005), .b(g61933_sb), .o(n_7957) );
na02f02 TIMEBOOST_cell_22580 ( .a(FE_OFN1749_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__Q), .o(TIMEBOOST_net_6547) );
na02m02 TIMEBOOST_cell_32520 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__Q), .o(TIMEBOOST_net_10171) );
na02f02 TIMEBOOST_cell_37126 ( .a(FE_OFN1601_n_13995), .b(TIMEBOOST_net_10801), .o(g53302_p) );
na02s02 TIMEBOOST_cell_36728 ( .a(TIMEBOOST_net_10602), .b(g63600_sb), .o(n_4768) );
na02f06 FE_RC_1013_0 ( .a(n_16330), .b(FE_RN_707_0), .o(n_16331) );
in01f08 FE_RC_1014_0 ( .a(n_15998), .o(n_15746) );
in01f04 FE_RC_1015_0 ( .a(n_15998), .o(FE_RN_708_0) );
na02f04 FE_RC_1016_0 ( .a(FE_RN_708_0), .b(n_15924), .o(n_15754) );
in01f04 FE_RC_1017_0 ( .a(n_15924), .o(FE_RN_709_0) );
na02s01 TIMEBOOST_cell_37273 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__Q), .b(FE_OFN671_n_4505), .o(TIMEBOOST_net_10875) );
na04f04 FE_RC_1019_0 ( .a(n_11097), .b(n_11788), .c(n_11095), .d(n_11096), .o(n_12545) );
in01f10 FE_RC_101_0 ( .a(wishbone_slave_unit_fifos_outGreyCount_2_), .o(FE_RN_57_0) );
in01s01 FE_RC_1020_0 ( .a(n_7822), .o(FE_RN_710_0) );
in01f02 FE_RC_1021_0 ( .a(n_12981), .o(FE_RN_711_0) );
na02s02 TIMEBOOST_cell_42036 ( .a(TIMEBOOST_net_13256), .b(g62582_sb), .o(n_6388) );
na02f02 TIMEBOOST_cell_40910 ( .a(TIMEBOOST_net_12693), .b(g57533_sb), .o(n_10312) );
na04f04 FE_RC_1025_0 ( .a(n_10154), .b(n_10151), .c(n_9307), .d(n_9306), .o(n_12158) );
in01f02 FE_RC_1026_0 ( .a(n_9274), .o(FE_RN_713_0) );
in01f02 FE_RC_1027_0 ( .a(n_17043), .o(FE_RN_714_0) );
no02f02 FE_RC_1028_0 ( .a(FE_RN_714_0), .b(FE_RN_713_0), .o(FE_RN_715_0) );
na02s02 TIMEBOOST_cell_42978 ( .a(TIMEBOOST_net_13727), .b(TIMEBOOST_net_9856), .o(n_5543) );
in01f08 FE_RC_102_0 ( .a(wishbone_slave_unit_fifos_pci_clk_inGreyCount_2_), .o(FE_RN_58_0) );
ao22f02 FE_RC_1031_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__Q), .b(FE_OCP_RBN1968_FE_OFN1532_n_10143), .c(n_10185), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__Q), .o(n_10599) );
ao22f02 FE_RC_1032_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__Q), .b(FE_OFN2149_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__Q), .d(FE_OFN1522_n_10892), .o(n_10728) );
in01f02 FE_RC_1033_0 ( .a(FE_RN_716_0), .o(n_16317) );
na02f02 FE_RC_1034_0 ( .a(n_16313), .b(n_16445), .o(FE_RN_716_0) );
na04f04 FE_RC_1035_0 ( .a(n_12036), .b(n_12310), .c(n_12037), .d(n_12038), .o(n_12818) );
na04f04 FE_RC_1036_0 ( .a(n_12195), .b(n_12196), .c(n_12112), .d(n_12341), .o(n_12868) );
in01m01 FE_RC_1037_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q), .o(FE_RN_717_0) );
na02s02 TIMEBOOST_cell_43514 ( .a(TIMEBOOST_net_13995), .b(FE_OFN1230_n_6391), .o(TIMEBOOST_net_12633) );
na02s01 TIMEBOOST_cell_45574 ( .a(TIMEBOOST_net_15025), .b(g64997_db), .o(n_4354) );
na02s02 TIMEBOOST_cell_42668 ( .a(TIMEBOOST_net_13572), .b(g64096_da), .o(TIMEBOOST_net_11305) );
in01s01 FE_RC_1041_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__531), .o(FE_RN_720_0) );
ao22f02 FE_RC_1043_0 ( .a(FE_RN_720_0), .b(FE_OFN1581_n_12306), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__Q), .d(FE_OFN1759_n_10780), .o(n_12721) );
in01m01 FE_RC_1044_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__Q), .o(FE_RN_722_0) );
in01f02 FE_RC_1045_0 ( .a(FE_OFN1559_n_12042), .o(FE_RN_723_0) );
na02s02 TIMEBOOST_cell_45226 ( .a(TIMEBOOST_net_14851), .b(FE_OFN1270_n_4095), .o(TIMEBOOST_net_12593) );
na02s01 TIMEBOOST_cell_43149 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q), .b(n_4308), .o(TIMEBOOST_net_13813) );
in01m01 FE_RC_1048_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__Q), .o(FE_RN_725_0) );
in01f02 FE_RC_1049_0 ( .a(FE_OFN1556_n_12042), .o(FE_RN_726_0) );
na02s01 TIMEBOOST_cell_37272 ( .a(TIMEBOOST_net_10874), .b(g64771_sb), .o(TIMEBOOST_net_221) );
na02f02 TIMEBOOST_cell_44560 ( .a(TIMEBOOST_net_14518), .b(FE_OFN2180_n_8567), .o(TIMEBOOST_net_12997) );
na02f02 TIMEBOOST_cell_22483 ( .a(TIMEBOOST_net_6498), .b(FE_OFN1551_n_12104), .o(n_12508) );
in01m01 FE_RC_1052_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__Q), .o(FE_RN_728_0) );
in01f02 FE_RC_1053_0 ( .a(FE_OFN1556_n_12042), .o(FE_RN_729_0) );
na02f02 TIMEBOOST_cell_43770 ( .a(TIMEBOOST_net_14123), .b(FE_OFN1422_n_8567), .o(TIMEBOOST_net_12900) );
na02f02 TIMEBOOST_cell_22485 ( .a(TIMEBOOST_net_6499), .b(FE_OCP_RBN1977_n_10273), .o(n_12520) );
na03f02 FE_RC_1056_0 ( .a(n_14535), .b(n_14497), .c(n_14407), .o(n_14579) );
na02s01 TIMEBOOST_cell_41939 ( .a(g65414_da), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__Q), .o(TIMEBOOST_net_13208) );
in01f10 FE_RC_105_0 ( .a(wishbone_slave_unit_fifos_pci_clk_inGreyCount_1_), .o(FE_RN_60_0) );
ao22f02 FE_RC_1060_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__Q), .b(FE_OFN1511_n_15587), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__Q), .d(FE_OFN1725_n_16891), .o(n_16845) );
ao22f02 FE_RC_1061_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__Q), .b(FE_OCP_RBN1969_FE_OFN1532_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__Q), .d(n_10195), .o(n_10078) );
in01m10 FE_RC_1062_0 ( .a(parchk_pci_ad_out_in_1174), .o(FE_RN_731_0) );
in01m10 FE_RC_1063_0 ( .a(parchk_pci_ad_out_in_1173), .o(FE_RN_732_0) );
na02s01 TIMEBOOST_cell_43150 ( .a(TIMEBOOST_net_13813), .b(FE_OFN1212_n_4151), .o(TIMEBOOST_net_12065) );
na03f02 TIMEBOOST_cell_34083 ( .a(TIMEBOOST_net_9676), .b(g54332_sb), .c(FE_OFN2128_n_16497), .o(n_12984) );
in01s02 FE_RC_1066_0 ( .a(n_13415), .o(FE_RN_734_0) );
in01f02 FE_RC_1067_0 ( .a(n_7312), .o(FE_RN_735_0) );
no02f03 FE_RC_1068_0 ( .a(FE_RN_735_0), .b(FE_RN_734_0), .o(FE_RN_736_0) );
no02f04 FE_RC_1069_0 ( .a(FE_RN_736_0), .b(n_13725), .o(n_13787) );
in01f10 FE_RC_106_0 ( .a(wishbone_slave_unit_fifos_outGreyCount_1_), .o(FE_RN_61_0) );
in01f02 FE_RC_1070_0 ( .a(n_3070), .o(FE_RN_737_0) );
in01f02 FE_RC_1071_0 ( .a(n_3292), .o(FE_RN_738_0) );
no02f02 FE_RC_1072_0 ( .a(FE_RN_737_0), .b(FE_RN_738_0), .o(FE_RN_739_0) );
na02m02 TIMEBOOST_cell_44259 ( .a(n_9808), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__Q), .o(TIMEBOOST_net_14368) );
in01s01 FE_RC_1074_0 ( .a(n_2284), .o(FE_RN_740_0) );
in01s01 FE_RC_1075_0 ( .a(n_2137), .o(FE_RN_741_0) );
no02s01 FE_RC_1076_0 ( .a(FE_RN_741_0), .b(FE_RN_740_0), .o(FE_RN_742_0) );
no02f02 FE_RC_1077_0 ( .a(FE_RN_742_0), .b(n_14532), .o(n_14622) );
na02s02 TIMEBOOST_cell_43646 ( .a(TIMEBOOST_net_14061), .b(FE_OFN2063_n_6391), .o(TIMEBOOST_net_12154) );
na04f04 FE_RC_1079_0 ( .a(n_11056), .b(n_11053), .c(n_11055), .d(n_11054), .o(n_12533) );
na02f02 TIMEBOOST_cell_37033 ( .a(FE_OFN1771_n_14054), .b(TIMEBOOST_net_10140), .o(TIMEBOOST_net_10755) );
na02s01 TIMEBOOST_cell_45227 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__Q), .b(n_4435), .o(TIMEBOOST_net_14852) );
na02f02 TIMEBOOST_cell_41024 ( .a(TIMEBOOST_net_12750), .b(g57418_sb), .o(n_11322) );
in01f02 FE_RC_1083_0 ( .a(n_10688), .o(FE_RN_743_0) );
in01f02 FE_RC_1084_0 ( .a(FE_RN_179_0), .o(FE_RN_744_0) );
no02f02 FE_RC_1085_0 ( .a(FE_RN_743_0), .b(FE_RN_744_0), .o(FE_RN_745_0) );
na02f02 FE_RC_1086_0 ( .a(FE_RN_745_0), .b(n_12579), .o(n_12841) );
ao22f02 FE_RC_1087_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__Q), .b(FE_OFN1511_n_15587), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__Q), .d(FE_OFN1725_n_16891), .o(n_16985) );
in01f02 FE_RC_1088_0 ( .a(n_10851), .o(FE_RN_746_0) );
in01f02 FE_RC_1089_0 ( .a(FE_RN_465_0), .o(FE_RN_747_0) );
na02s01 TIMEBOOST_cell_42979 ( .a(FE_OFN237_n_9118), .b(g58189_sb), .o(TIMEBOOST_net_13728) );
no02f02 FE_RC_1090_0 ( .a(FE_RN_746_0), .b(FE_RN_747_0), .o(FE_RN_748_0) );
na02f02 FE_RC_1091_0 ( .a(n_12559), .b(FE_RN_748_0), .o(n_12821) );
na02s01 TIMEBOOST_cell_40373 ( .a(TIMEBOOST_net_986), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__Q), .o(TIMEBOOST_net_12425) );
in01s01 FE_RC_1093_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__Q), .o(FE_RN_749_0) );
in01f02 FE_RC_1094_0 ( .a(FE_OFN1720_n_16891), .o(FE_RN_750_0) );
no02f02 FE_RC_1095_0 ( .a(FE_RN_749_0), .b(FE_RN_750_0), .o(FE_RN_751_0) );
no02f02 FE_RC_1096_0 ( .a(n_15592), .b(FE_RN_751_0), .o(n_15593) );
ao22f02 FE_RC_1097_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__Q), .b(FE_OFN2147_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__Q), .d(FE_OFN1523_n_10892), .o(n_10596) );
na02s02 TIMEBOOST_cell_41943 ( .a(TIMEBOOST_net_1824), .b(FE_OFN1083_n_13221), .o(TIMEBOOST_net_13210) );
ao22f02 FE_RC_1099_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__Q), .b(FE_OCP_RBN1968_FE_OFN1532_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__Q), .d(n_10185), .o(n_10188) );
in01f10 FE_RC_109_0 ( .a(wishbone_slave_unit_fifos_pci_clk_inGreyCount_0_), .o(FE_RN_63_0) );
in01f04 FE_RC_10_0 ( .a(n_16021), .o(FE_RN_6_0) );
ao22f02 FE_RC_1100_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__Q), .b(FE_OFN1511_n_15587), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__Q), .d(FE_OFN1725_n_16891), .o(n_9982) );
ao22f02 FE_RC_1101_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__Q), .b(FE_OCP_RBN1968_FE_OFN1532_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__Q), .d(n_10185), .o(n_10026) );
na02s02 TIMEBOOST_cell_16831 ( .a(TIMEBOOST_net_3672), .b(g65318_db), .o(n_3564) );
ao22f02 FE_RC_1103_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__Q), .b(FE_OFN2147_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__Q), .d(FE_OFN1523_n_10892), .o(n_10173) );
ao22f02 FE_RC_1104_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__Q), .b(FE_OFN2147_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__Q), .d(FE_OFN1523_n_10892), .o(n_10877) );
ao22f02 FE_RC_1105_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__Q), .b(FE_OFN2146_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__Q), .d(FE_OFN1547_n_10566), .o(n_9979) );
in01f02 FE_RC_1106_0 ( .a(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(FE_RN_752_0) );
in01m06 FE_RC_1107_0 ( .a(n_15859), .o(FE_RN_753_0) );
na02f06 FE_RC_1108_0 ( .a(FE_RN_752_0), .b(FE_RN_753_0), .o(FE_OFN997_n_15978) );
no02m06 FE_RC_1109_0 ( .a(wishbone_slave_unit_pci_initiator_if_del_read_req), .b(n_15859), .o(FE_OFN1000_n_15978) );
in01f10 FE_RC_110_0 ( .a(wishbone_slave_unit_fifos_outGreyCount_0_), .o(FE_RN_64_0) );
in01f10 FE_RC_1110_0 ( .a(wishbone_slave_unit_pci_initiator_if_err_recovery), .o(FE_RN_754_0) );
na02s01 TIMEBOOST_cell_45228 ( .a(TIMEBOOST_net_14852), .b(FE_OFN1249_n_4093), .o(TIMEBOOST_net_12561) );
no02f20 FE_RC_1112_0 ( .a(wbu_pciif_devsel_reg_in), .b(n_16763), .o(n_15798) );
na02f06 FE_RC_1114_0 ( .a(g75418_da), .b(g75418_db), .o(n_16974) );
in01f02 FE_RC_1115_0 ( .a(g75418_db), .o(FE_RN_755_0) );
in01f02 FE_RC_1116_0 ( .a(g75418_da), .o(FE_RN_756_0) );
no02f08 FE_RC_1117_0 ( .a(FE_RN_756_0), .b(FE_RN_755_0), .o(n_16205) );
in01f06 FE_RC_1118_0 ( .a(n_16966), .o(n_16967) );
na02s02 TIMEBOOST_cell_41705 ( .a(g58786_sb), .b(wbu_addr_in_276), .o(TIMEBOOST_net_13091) );
na03s02 TIMEBOOST_cell_6343 ( .a(n_4450), .b(FE_OFN1680_n_4655), .c(g65350_da), .o(n_4258) );
na03s02 TIMEBOOST_cell_42987 ( .a(g64100_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__Q), .c(FE_OFN882_g64577_p), .o(TIMEBOOST_net_13732) );
in01f02 FE_RC_1123_0 ( .a(n_16974), .o(FE_RN_758_0) );
na02f04 FE_RC_1124_0 ( .a(FE_OCP_RBN2016_n_16970), .b(n_16967), .o(FE_RN_759_0) );
no02f08 FE_RC_1125_0 ( .a(FE_RN_758_0), .b(FE_RN_759_0), .o(n_13901) );
na02f02 TIMEBOOST_cell_44681 ( .a(TIMEBOOST_net_10051), .b(FE_OFN1376_n_8567), .o(TIMEBOOST_net_14579) );
in01f10 FE_RC_1130_0 ( .a(n_16516), .o(FE_RN_764_0) );
na04f04 FE_RC_1135_0 ( .a(n_14536), .b(n_13930), .c(n_14499), .d(n_13849), .o(n_14580) );
na02f02 TIMEBOOST_cell_40912 ( .a(TIMEBOOST_net_12694), .b(g57106_sb), .o(n_11639) );
in01f02 FE_RC_1138_0 ( .a(n_13854), .o(FE_RN_767_0) );
in01s01 FE_RC_1139_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__Q), .o(FE_RN_768_0) );
in01f04 FE_RC_113_0 ( .a(n_15401), .o(FE_RN_66_0) );
in01f02 FE_RC_1140_0 ( .a(FE_OCP_RBN1996_n_13971), .o(FE_RN_769_0) );
na02s02 TIMEBOOST_cell_42362 ( .a(TIMEBOOST_net_13419), .b(g54353_sb), .o(n_13088) );
na02s02 TIMEBOOST_cell_45575 ( .a(n_4498), .b(g64937_sb), .o(TIMEBOOST_net_15026) );
na02s01 TIMEBOOST_cell_45016 ( .a(TIMEBOOST_net_14746), .b(g65304_db), .o(n_3573) );
ao22f02 FE_RC_1144_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__Q), .b(FE_OFN1462_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__Q), .d(FE_OFN1457_n_11138), .o(n_17017) );
ao22f02 FE_RC_1145_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__Q), .b(FE_OCP_RBN2010_n_16698), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__Q), .d(FE_OFN1465_n_10789), .o(n_11093) );
na02f02 TIMEBOOST_cell_44348 ( .a(TIMEBOOST_net_14412), .b(FE_OFN1422_n_8567), .o(TIMEBOOST_net_12733) );
na02f02 TIMEBOOST_cell_44275 ( .a(n_9615), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__Q), .o(TIMEBOOST_net_14376) );
in01f03 FE_RC_114_0 ( .a(n_16798), .o(FE_RN_67_0) );
in01f06 FE_RC_1153_0 ( .a(n_16264), .o(n_15823) );
no02f20 FE_RC_1155_0 ( .a(FE_OCP_RBN2270_g75061_p), .b(n_16264), .o(FE_RN_772_0) );
na02f20 FE_RC_1156_0 ( .a(n_16599), .b(FE_RN_772_0), .o(n_16980) );
in01f02 FE_RC_1157_0 ( .a(n_16154), .o(FE_RN_773_0) );
in01f02 FE_RC_1158_0 ( .a(n_16153), .o(FE_RN_774_0) );
no02f04 FE_RC_1159_0 ( .a(FE_RN_774_0), .b(FE_RN_773_0), .o(FE_RN_775_0) );
na03s01 TIMEBOOST_cell_34039 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(g64083_sb), .c(g64083_db), .o(n_4072) );
na02f06 FE_RC_1160_0 ( .a(FE_RN_775_0), .b(n_16980), .o(n_16156) );
in01f02 FE_RC_1161_0 ( .a(FE_RN_776_0), .o(n_3421) );
na02f04 FE_RC_1162_0 ( .a(FE_OCP_RBN2238_g74749_p), .b(n_3310), .o(FE_RN_776_0) );
in01f01 FE_RC_1166_0 ( .a(n_16966), .o(FE_RN_778_0) );
no02f03 FE_RC_1167_0 ( .a(FE_OCP_RBN2279_n_16974), .b(FE_RN_778_0), .o(FE_RN_779_0) );
na02f06 FE_RC_1168_0 ( .a(FE_RN_779_0), .b(FE_OCP_RBN2017_n_16970), .o(FE_OFN1772_n_13800) );
na02f04 FE_RC_1169_0 ( .a(FE_OCP_RBN2019_n_16970), .b(n_16966), .o(FE_RN_780_0) );
na02s02 TIMEBOOST_cell_37788 ( .a(TIMEBOOST_net_11132), .b(FE_OFN2256_n_8060), .o(TIMEBOOST_net_4354) );
no02f10 FE_RC_1170_0 ( .a(FE_RN_780_0), .b(FE_OCP_RBN2278_n_16974), .o(FE_OFN1774_n_13800) );
in01f10 FE_RC_117_0 ( .a(pci_target_unit_pci_target_sm_rd_from_fifo), .o(FE_RN_69_0) );
in01f10 FE_RC_118_0 ( .a(pci_target_unit_pci_target_sm_same_read_reg), .o(FE_RN_70_0) );
in01f02 FE_RC_1194_0 ( .a(FE_RN_8_0), .o(FE_RN_795_0) );
no02f02 FE_RC_1195_0 ( .a(n_15919), .b(FE_RN_795_0), .o(n_15917) );
in01f02 FE_RC_1196_0 ( .a(n_16075), .o(n_16076) );
in01f02 FE_RC_1197_0 ( .a(n_16075), .o(FE_RN_796_0) );
na02f02 FE_RC_1198_0 ( .a(n_16444), .b(FE_RN_796_0), .o(n_15581) );
in01m10 FE_RC_1199_0 ( .a(parchk_pci_ad_out_in), .o(FE_RN_797_0) );
no02f08 FE_RC_119_0 ( .a(FE_RN_69_0), .b(FE_RN_70_0), .o(FE_RN_71_0) );
in01f04 FE_RC_11_0 ( .a(n_16914), .o(FE_RN_7_0) );
in01m10 FE_RC_1200_0 ( .a(parchk_pci_ad_out_in_1168), .o(FE_RN_798_0) );
na02s01 TIMEBOOST_cell_37451 ( .a(pci_target_unit_del_sync_addr_in_232), .b(parchk_pci_ad_reg_in_1233), .o(TIMEBOOST_net_10964) );
na02s02 TIMEBOOST_cell_38104 ( .a(TIMEBOOST_net_11290), .b(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_4618) );
in01s01 FE_RC_1203_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__Q), .o(FE_RN_800_0) );
no02f04 FE_RC_1204_0 ( .a(FE_OCPN1856_FE_OFN1774_n_13800), .b(FE_RN_800_0), .o(FE_RN_801_0) );
in01f02 FE_RC_1205_0 ( .a(FE_RN_802_0), .o(g53187_p) );
ao12f02 FE_RC_1206_0 ( .a(FE_RN_801_0), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__Q), .c(FE_OFN1771_n_14054), .o(FE_RN_802_0) );
na02s01 TIMEBOOST_cell_38646 ( .a(TIMEBOOST_net_11561), .b(g59111_sb), .o(n_8707) );
na02f02 TIMEBOOST_cell_44682 ( .a(TIMEBOOST_net_14579), .b(g57256_sb), .o(n_11497) );
na02s01 TIMEBOOST_cell_39536 ( .a(TIMEBOOST_net_12006), .b(g61726_sb), .o(n_8368) );
in01s01 TIMEBOOST_cell_45874 ( .a(TIMEBOOST_net_15180), .o(TIMEBOOST_net_15181) );
in01f02 FE_RC_1211_0 ( .a(n_14963), .o(FE_RN_805_0) );
in01s01 FE_RC_1212_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__Q), .o(FE_RN_806_0) );
in01f02 FE_RC_1213_0 ( .a(FE_OCP_RBN1985_FE_OFN1591_n_13741), .o(FE_RN_807_0) );
na02s01 TIMEBOOST_cell_42918 ( .a(TIMEBOOST_net_13697), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_11181) );
na02s02 TIMEBOOST_cell_45229 ( .a(n_4913), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__Q), .o(TIMEBOOST_net_14853) );
na02s02 TIMEBOOST_cell_45230 ( .a(TIMEBOOST_net_14853), .b(FE_OFN1274_n_4096), .o(TIMEBOOST_net_12563) );
na03s02 TIMEBOOST_cell_42037 ( .a(n_3640), .b(FE_OFN1276_n_4096), .c(n_84), .o(TIMEBOOST_net_13257) );
na02s01 TIMEBOOST_cell_45017 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__30__Q), .b(g65382_sb), .o(TIMEBOOST_net_14747) );
in01s02 FE_RC_121_0 ( .a(n_2629), .o(FE_RN_72_0) );
ao22f02 FE_RC_1220_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__Q), .b(FE_OFN1727_n_9975), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__Q), .d(FE_OCP_RBN2005_FE_RN_459_0), .o(n_9303) );
ao22f02 FE_RC_1221_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__Q), .b(FE_OFN2149_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__Q), .d(FE_OFN1522_n_10892), .o(n_17046) );
ao22f02 FE_RC_1222_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q), .b(FE_OFN2147_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__Q), .d(FE_OFN1523_n_10892), .o(n_10054) );
ao22f02 FE_RC_1223_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__Q), .b(FE_OFN2149_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__Q), .d(FE_OFN1522_n_10892), .o(n_10930) );
ao22f02 FE_RC_1224_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__Q), .b(FE_OFN1536_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__Q), .d(n_10141), .o(n_17045) );
na02m02 TIMEBOOST_cell_41583 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_22__Q), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_13030) );
ao22f06 FE_RC_1226_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_1_), .c(n_16175), .d(FE_OCP_RBN2290_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .o(n_16433) );
na02f06 FE_RC_1227_0 ( .a(FE_OCP_RBN1955_n_16981), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q), .o(FE_RN_809_0) );
in01f02 FE_RC_1229_0 ( .a(n_13856), .o(FE_RN_810_0) );
in01m02 FE_RC_122_0 ( .a(n_2623), .o(FE_RN_73_0) );
in01s01 FE_RC_1230_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__Q), .o(FE_RN_811_0) );
in01f02 FE_RC_1231_0 ( .a(FE_OCP_RBN1995_n_13971), .o(FE_RN_812_0) );
na02f02 TIMEBOOST_cell_22581 ( .a(n_12273), .b(TIMEBOOST_net_6547), .o(n_12707) );
na02f02 TIMEBOOST_cell_38910 ( .a(TIMEBOOST_net_11693), .b(FE_OFN2200_n_10256), .o(TIMEBOOST_net_10698) );
in01f02 FE_RC_1234_0 ( .a(n_13990), .o(FE_RN_814_0) );
in01f02 FE_RC_1235_0 ( .a(n_13991), .o(FE_RN_815_0) );
no02f02 FE_RC_1236_0 ( .a(FE_RN_814_0), .b(FE_RN_815_0), .o(n_14283) );
in01f02 FE_RC_1237_0 ( .a(n_14197), .o(FE_RN_816_0) );
in01s01 FE_RC_1238_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__Q), .o(FE_RN_817_0) );
in01f02 FE_RC_1239_0 ( .a(FE_OFN1769_n_14054), .o(FE_RN_818_0) );
na02s01 TIMEBOOST_cell_37275 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__Q), .b(FE_OFN670_n_4505), .o(TIMEBOOST_net_10876) );
na02s02 TIMEBOOST_cell_40878 ( .a(TIMEBOOST_net_12677), .b(g62501_sb), .o(n_6580) );
na02m02 TIMEBOOST_cell_32374 ( .a(wbs_wbb3_2_wbb2_dat_o_i_119), .b(wbs_dat_o_20_), .o(TIMEBOOST_net_10098) );
na02f02 TIMEBOOST_cell_40914 ( .a(TIMEBOOST_net_12695), .b(g57052_sb), .o(n_11684) );
na02f10 FE_RC_1243_0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_control_in_86), .b(n_16501), .o(FE_RN_820_0) );
in01f10 FE_RC_1244_0 ( .a(pci_target_unit_wishbone_master_burst_chopped_delayed), .o(FE_RN_821_0) );
na02s01 TIMEBOOST_cell_45748 ( .a(TIMEBOOST_net_15112), .b(FE_OFN2081_n_8176), .o(TIMEBOOST_net_11037) );
na02f06 FE_RC_1246_0 ( .a(n_16499), .b(FE_RN_822_0), .o(n_16513) );
na02s02 TIMEBOOST_cell_37888 ( .a(TIMEBOOST_net_11182), .b(g58334_sb), .o(n_9483) );
in01f02 FE_RC_1250_0 ( .a(FE_RN_824_0), .o(n_14054) );
na03f02 FE_RC_1251_0 ( .a(n_16974), .b(n_16966), .c(n_16970), .o(FE_RN_824_0) );
na02s02 TIMEBOOST_cell_43342 ( .a(TIMEBOOST_net_13909), .b(g62634_sb), .o(n_6284) );
na02s02 TIMEBOOST_cell_40880 ( .a(TIMEBOOST_net_12678), .b(g62442_sb), .o(n_6712) );
na02s01 TIMEBOOST_cell_42038 ( .a(TIMEBOOST_net_13257), .b(g62641_sb), .o(n_6266) );
in01f02 FE_RC_1256_0 ( .a(n_13847), .o(FE_RN_827_0) );
in01s01 FE_RC_1257_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__Q), .o(FE_RN_828_0) );
in01f02 FE_RC_1258_0 ( .a(FE_OCP_RBN1996_n_13971), .o(FE_RN_829_0) );
na02s01 TIMEBOOST_cell_39216 ( .a(TIMEBOOST_net_11846), .b(n_1565), .o(TIMEBOOST_net_11475) );
na02s02 TIMEBOOST_cell_17467 ( .a(TIMEBOOST_net_3990), .b(g65292_da), .o(n_4283) );
in01f02 FE_RC_1261_0 ( .a(n_14099), .o(FE_RN_831_0) );
in01s01 FE_RC_1262_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__Q), .o(FE_RN_832_0) );
in01f02 FE_RC_1263_0 ( .a(FE_OCPN2218_n_13997), .o(FE_RN_833_0) );
na02f04 TIMEBOOST_cell_36295 ( .a(FE_RN_597_0), .b(FE_RN_598_0), .o(TIMEBOOST_net_10386) );
na02f10 TIMEBOOST_cell_36284 ( .a(TIMEBOOST_net_10380), .b(n_3030), .o(n_2380) );
in01f02 FE_RC_1266_0 ( .a(n_14507), .o(FE_RN_835_0) );
na02f02 TIMEBOOST_cell_40916 ( .a(TIMEBOOST_net_12696), .b(g57274_sb), .o(n_11480) );
na02s01 TIMEBOOST_cell_39287 ( .a(TIMEBOOST_net_9344), .b(FE_OFN956_n_1699), .o(TIMEBOOST_net_11882) );
na02f02 TIMEBOOST_cell_42388 ( .a(TIMEBOOST_net_13432), .b(g57050_sb), .o(n_11685) );
na04f04 FE_RC_1270_0 ( .a(n_11101), .b(n_11099), .c(n_11102), .d(n_11100), .o(n_12546) );
na04f04 FE_RC_1271_0 ( .a(n_12248), .b(n_11960), .c(n_12246), .d(n_11819), .o(n_12814) );
ao22f02 FE_RC_1273_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q), .b(FE_OFN2137_n_15534), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q), .d(FE_OFN2144_n_16992), .o(n_16984) );
ao22f02 FE_RC_1274_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__Q), .b(FE_OFN2149_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__Q), .d(FE_OFN1522_n_10892), .o(n_10524) );
ao22f02 FE_RC_1275_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__Q), .b(FE_OFN2216_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__Q), .d(n_11728), .o(n_11733) );
ao22f02 FE_RC_1276_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__Q), .b(FE_OFN2146_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__Q), .d(FE_OFN1547_n_10566), .o(n_9311) );
ao22f02 FE_RC_1277_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__Q), .b(FE_OFN1535_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__Q), .d(n_11728), .o(n_10947) );
ao22f02 FE_RC_1278_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__Q), .b(FE_OFN1493_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__Q), .d(FE_OFN1546_n_10566), .o(n_10903) );
ao22f02 FE_RC_1279_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__Q), .b(FE_OFN1478_n_16637), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__Q), .d(FE_OFN2193_n_9163), .o(n_11118) );
na03f02 FE_RC_1280_0 ( .a(FE_RN_113_0), .b(n_13051), .c(n_12787), .o(n_13134) );
ao22f02 FE_RC_1281_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__8__Q), .b(FE_OFN2131_n_10588), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__8__Q), .d(FE_OFN1528_n_10853), .o(n_10533) );
ao22f02 FE_RC_1282_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__Q), .b(FE_OFN1508_n_15587), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__Q), .d(FE_OFN1720_n_16891), .o(n_9988) );
ao22f02 FE_RC_1283_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__Q), .b(FE_OFN2216_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__Q), .d(n_11728), .o(n_11726) );
ao22f02 FE_RC_1284_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__Q), .b(FE_OFN1727_n_9975), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__Q), .d(FE_OCP_RBN1932_FE_OFN1515_n_10538), .o(n_17044) );
ao22f02 FE_RC_1285_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__Q), .b(FE_OFN1493_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__Q), .d(FE_OFN1546_n_10566), .o(n_10702) );
ao22f02 FE_RC_1286_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__Q), .b(n_16637), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__Q), .d(FE_OFN2194_n_9163), .o(n_11091) );
ao22f02 FE_RC_1287_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__Q), .b(FE_OCP_RBN2010_n_16698), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__Q), .d(FE_OFN1465_n_10789), .o(n_11059) );
ao22f02 FE_RC_1288_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__Q), .b(FE_OFN1479_n_16637), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__Q), .d(FE_OFN2194_n_9163), .o(n_11073) );
in01f04 FE_RC_1289_0 ( .a(n_16358), .o(FE_RN_836_0) );
in01f08 FE_RC_1291_0 ( .a(FE_RN_0_0), .o(FE_RN_837_0) );
in01f02 FE_RC_1293_0 ( .a(n_16513), .o(FE_RN_839_0) );
no02f04 FE_RC_1294_0 ( .a(FE_RN_839_0), .b(FE_RN_462_0), .o(FE_RN_840_0) );
na02s02 TIMEBOOST_cell_19082 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q), .b(g58361_sb), .o(TIMEBOOST_net_4798) );
na02m02 TIMEBOOST_cell_36364 ( .a(TIMEBOOST_net_1091), .b(TIMEBOOST_net_10420), .o(n_9122) );
na03s02 TIMEBOOST_cell_5529 ( .a(n_4470), .b(g65049_sb), .c(g65049_db), .o(n_4322) );
na02s02 TIMEBOOST_cell_43518 ( .a(TIMEBOOST_net_13997), .b(FE_OFN1225_n_6391), .o(TIMEBOOST_net_12537) );
in01f02 FE_RC_1299_0 ( .a(n_14111), .o(FE_RN_843_0) );
no02f04 FE_RC_12_0 ( .a(FE_RN_7_0), .b(FE_RN_6_0), .o(FE_RN_8_0) );
in01s01 FE_RC_1300_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__Q), .o(FE_RN_844_0) );
in01f02 FE_RC_1301_0 ( .a(FE_OFN1602_n_13995), .o(FE_RN_845_0) );
na02s01 TIMEBOOST_cell_36285 ( .a(parchk_pci_ad_reg_in_1233), .b(g67094_db), .o(TIMEBOOST_net_10381) );
na02s01 TIMEBOOST_cell_41938 ( .a(TIMEBOOST_net_13207), .b(g58439_db), .o(n_9200) );
ao22f02 FE_RC_1305_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__Q), .b(FE_OFN2146_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__Q), .d(FE_OFN1547_n_10566), .o(n_10023) );
ao22f02 FE_RC_1306_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__Q), .b(FE_OFN1489_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__Q), .d(FE_OFN1548_n_10566), .o(n_9287) );
ao22f02 FE_RC_1307_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__Q), .b(FE_OFN2146_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__Q), .d(FE_OFN1547_n_10566), .o(n_9297) );
ao22f02 FE_RC_1308_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__Q), .b(FE_OCP_RBN2011_n_16698), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__Q), .d(FE_OFN1467_n_10789), .o(n_10791) );
na03f08 FE_RC_1309_0 ( .a(FE_OFN996_n_15366), .b(n_16049), .c(n_16046), .o(n_16310) );
na03s02 TIMEBOOST_cell_41963 ( .a(n_3660), .b(FE_OFN1250_n_4093), .c(n_119), .o(TIMEBOOST_net_13220) );
ao22f02 FE_RC_1310_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__Q), .b(FE_OFN2146_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__Q), .d(FE_OFN1547_n_10566), .o(n_9319) );
ao22f02 FE_RC_1311_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__Q), .b(FE_OCP_RBN2009_n_16698), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__Q), .d(FE_OFN1466_n_10789), .o(n_11137) );
na04f04 FE_RC_1312_0 ( .a(n_12052), .b(n_12053), .c(n_12054), .d(n_12055), .o(n_12819) );
in01f02 FE_RC_1335_0 ( .a(n_16403), .o(FE_RN_862_0) );
in01f02 FE_RC_1336_0 ( .a(n_16406), .o(FE_RN_863_0) );
na03f02 FE_RC_1338_0 ( .a(FE_RN_107_0), .b(n_13059), .c(n_12799), .o(n_13141) );
in01f02 FE_RC_1364_0 ( .a(n_16547), .o(FE_RN_880_0) );
in01f02 FE_RC_1365_0 ( .a(n_16550), .o(FE_RN_881_0) );
no02f06 FE_RC_1366_0 ( .a(FE_RN_881_0), .b(FE_RN_880_0), .o(n_16552) );
na02s01 TIMEBOOST_cell_43151 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__Q), .b(n_3703), .o(TIMEBOOST_net_13814) );
na02s01 TIMEBOOST_cell_45018 ( .a(TIMEBOOST_net_14747), .b(g65382_db), .o(n_3526) );
na03f02 FE_RC_1369_0 ( .a(n_12928), .b(FE_RN_236_0), .c(n_13120), .o(n_13323) );
na02s02 TIMEBOOST_cell_45231 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__Q), .b(n_3693), .o(TIMEBOOST_net_14854) );
na02s01 TIMEBOOST_cell_39538 ( .a(TIMEBOOST_net_12007), .b(g61717_sb), .o(n_8391) );
no02f04 FE_RC_1372_0 ( .a(n_3448), .b(n_3320), .o(FE_RN_882_0) );
na02f04 FE_RC_1373_0 ( .a(FE_RN_882_0), .b(n_16507), .o(FE_RN_883_0) );
na02s02 TIMEBOOST_cell_45711 ( .a(n_4418), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__14__Q), .o(TIMEBOOST_net_15094) );
no02f04 FE_RC_1375_0 ( .a(FE_RN_430_0), .b(FE_RN_428_0), .o(FE_OFN1026_n_16760) );
na02f02 TIMEBOOST_cell_43814 ( .a(TIMEBOOST_net_14145), .b(FE_OFN1416_n_8567), .o(TIMEBOOST_net_12843) );
ao22f02 FE_RC_1377_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__Q), .b(FE_OFN1493_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__Q), .d(FE_OFN1546_n_10566), .o(n_10741) );
ao22f02 FE_RC_1378_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__Q), .b(FE_OFN2130_n_10588), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q), .d(FE_OFN1530_n_10853), .o(n_10951) );
na02f02 TIMEBOOST_cell_39540 ( .a(TIMEBOOST_net_12008), .b(n_5230), .o(TIMEBOOST_net_531) );
in01s10 FE_RC_137_0 ( .a(configuration_sync_command_bit1), .o(FE_RN_81_0) );
no02f06 FE_RC_1383_0 ( .a(FE_OCP_RBN2271_g75061_p), .b(n_16433), .o(n_16434) );
na02f08 FE_RC_1384_0 ( .a(FE_RN_809_0), .b(g75413_db), .o(n_16966) );
na02f02 FE_RC_1385_0 ( .a(g75413_db), .b(FE_RN_809_0), .o(n_14939) );
na02m02 TIMEBOOST_cell_32372 ( .a(wbs_wbb3_2_wbb2_dat_o_i_102), .b(wbs_dat_o_3_), .o(TIMEBOOST_net_10097) );
na02f02 TIMEBOOST_cell_40882 ( .a(TIMEBOOST_net_12679), .b(n_7685), .o(TIMEBOOST_net_6441) );
na02f02 FE_RC_1388_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__Q), .b(n_13891), .o(FE_RN_887_0) );
in01s01 FE_RC_1389_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q), .o(FE_RN_888_0) );
in01s10 FE_RC_138_0 ( .a(conf_pci_init_complete_out), .o(FE_RN_82_0) );
oa12f02 FE_RC_1390_0 ( .a(FE_RN_887_0), .b(FE_RN_888_0), .c(FE_OCP_RBN1964_FE_OFN1591_n_13741), .o(g53206_p) );
na02m02 TIMEBOOST_cell_32370 ( .a(wbs_wbb3_2_wbb2_dat_o_i_114), .b(wbs_dat_o_15_), .o(TIMEBOOST_net_10096) );
na02m02 TIMEBOOST_cell_40884 ( .a(TIMEBOOST_net_12680), .b(n_3356), .o(n_14838) );
no02f02 FE_RC_1393_0 ( .a(n_14268), .b(FE_RN_890_0), .o(n_14556) );
ao22f02 FE_RC_1394_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__Q), .b(FE_OFN1478_n_16637), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__Q), .d(FE_OFN2193_n_9163), .o(n_11104) );
ao22f01 FE_RC_1395_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__Q), .b(n_15566), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__Q), .d(n_15558), .o(n_9328) );
ao22f02 FE_RC_1396_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__Q), .b(n_15566), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__Q), .d(FE_OFN1499_n_15558), .o(n_10002) );
ao22f02 FE_RC_1397_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__Q), .b(FE_OFN2137_n_15534), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__Q), .d(FE_OCPN1873_FE_OFN474_n_16992), .o(n_10755) );
ao22f02 FE_RC_1398_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__Q), .b(FE_OFN1485_n_15534), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__Q), .d(FE_OCPN1888_FE_OFN473_n_16992), .o(n_10758) );
ao22f02 FE_RC_1399_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__Q), .b(FE_OFN1433_n_16779), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__Q), .d(FE_OFN1445_n_11125), .o(n_11051) );
no02m06 FE_RC_139_0 ( .a(FE_RN_81_0), .b(FE_RN_82_0), .o(FE_RN_83_0) );
ao22f02 FE_RC_1400_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__Q), .b(FE_OFN1432_n_16779), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__Q), .d(FE_OFN1445_n_11125), .o(n_11113) );
ao22f02 FE_RC_1401_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__Q), .b(FE_OFN2208_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__Q), .d(FE_OFN1455_n_11138), .o(n_11777) );
ao22f02 FE_RC_1402_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__Q), .b(FE_OFN1462_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__Q), .d(FE_OFN1457_n_11138), .o(n_11107) );
na02m02 TIMEBOOST_cell_32368 ( .a(wbs_wbb3_2_wbb2_dat_o_i_104), .b(wbs_dat_o_5_), .o(TIMEBOOST_net_10095) );
na03m02 TIMEBOOST_cell_33985 ( .a(pci_target_unit_pcit_if_strd_addr_in_692), .b(g52651_sb), .c(g52651_db), .o(n_14671) );
na02f02 TIMEBOOST_cell_40886 ( .a(TIMEBOOST_net_12681), .b(g57115_db), .o(n_11631) );
na02m02 TIMEBOOST_cell_32366 ( .a(wbs_wbb3_2_wbb2_dat_o_i_101), .b(wbs_dat_o_2_), .o(TIMEBOOST_net_10094) );
no02f02 FE_RC_1407_0 ( .a(FE_RN_893_0), .b(n_14505), .o(n_14539) );
na02m06 TIMEBOOST_cell_45019 ( .a(TIMEBOOST_net_4221), .b(TIMEBOOST_net_870), .o(TIMEBOOST_net_14748) );
na02s01 TIMEBOOST_cell_16805 ( .a(TIMEBOOST_net_3659), .b(g64970_db), .o(n_3653) );
in01s01 TIMEBOOST_cell_45942 ( .a(TIMEBOOST_net_15248), .o(TIMEBOOST_net_15249) );
ao22f02 FE_RC_1410_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__Q), .b(FE_OFN1460_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__Q), .d(FE_OFN1456_n_11138), .o(n_11058) );
na03f02 FE_RC_1411_0 ( .a(FE_RN_863_0), .b(FE_RN_862_0), .c(n_13067), .o(n_13408) );
ao22f02 FE_RC_1412_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__Q), .b(FE_OFN1731_n_9975), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__Q), .d(FE_OCP_RBN2006_FE_RN_459_0), .o(n_10530) );
ao22f02 FE_RC_1413_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__Q), .b(n_15566), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__Q), .d(FE_OFN1501_n_15558), .o(n_9265) );
ao22f02 FE_RC_1414_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q), .b(FE_OCPN1884_n_15566), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__Q), .d(FE_OFN1498_n_15558), .o(n_10179) );
ao22f02 FE_RC_1415_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__Q), .b(FE_OFN2208_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__Q), .d(FE_OFN1455_n_11138), .o(n_11048) );
ao22f02 FE_RC_1416_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__Q), .b(FE_OCP_RBN2009_n_16698), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__Q), .d(FE_OFN1466_n_10789), .o(n_11106) );
ao22f02 FE_RC_1417_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__Q), .b(FE_OFN1484_n_15534), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__Q), .d(n_16992), .o(n_16834) );
ao22f02 FE_RC_1418_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__Q), .b(FE_OFN1462_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__Q), .d(FE_OFN1457_n_11138), .o(n_11139) );
ao22f02 FE_RC_1419_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__Q), .b(FE_OFN2208_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__Q), .d(FE_OFN1455_n_11138), .o(n_11796) );
in01f02 FE_RC_1420_0 ( .a(n_15917), .o(FE_RN_894_0) );
no02f04 FE_RC_1421_0 ( .a(FE_RN_894_0), .b(FE_RN_390_0), .o(FE_RN_895_0) );
in01f03 FE_RC_1423_0 ( .a(n_16523), .o(FE_RN_896_0) );
oa22f04 FE_RC_1424_0 ( .a(n_16523), .b(FE_RN_493_0), .c(FE_RN_896_0), .d(FE_RN_491_0), .o(n_16075) );
in01m01 FE_RC_1425_0 ( .a(FE_RN_15_0), .o(FE_RN_897_0) );
in01f01 FE_RC_1426_0 ( .a(FE_RN_899_0), .o(FE_RN_898_0) );
no02f06 FE_RC_1427_0 ( .a(FE_RN_897_0), .b(FE_RN_898_0), .o(n_14971) );
na02f03 FE_RC_1428_0 ( .a(n_15915), .b(n_16524), .o(FE_RN_899_0) );
in01f02 FE_RC_1429_0 ( .a(FE_RN_15_0), .o(FE_RN_900_0) );
in01f04 FE_RC_1430_0 ( .a(n_135), .o(FE_RN_901_0) );
no02f02 FE_RC_1431_0 ( .a(FE_RN_900_0), .b(FE_RN_901_0), .o(FE_RN_902_0) );
na02f04 FE_RC_1432_0 ( .a(FE_RN_899_0), .b(FE_RN_902_0), .o(n_16564) );
ao22f02 FE_RC_1433_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__Q), .b(n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__Q), .d(n_11728), .o(n_10931) );
na02f03 FE_RC_1436_0 ( .a(wbm_dat_o_22_), .b(n_14800), .o(FE_RN_904_0) );
in01s01 FE_RC_1437_0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_71), .o(FE_RN_905_0) );
oa12f02 FE_RC_1438_0 ( .a(FE_RN_904_0), .b(FE_RN_905_0), .c(n_14725), .o(FE_RN_906_0) );
in01f02 FE_RC_1439_0 ( .a(FE_RN_907_0), .o(n_16304) );
ao22f02 FE_RC_1440_0 ( .a(n_16300), .b(FE_RN_906_0), .c(wbm_dat_o_22_), .d(FE_OFN2164_n_16301), .o(FE_RN_907_0) );
na03s02 TIMEBOOST_cell_37803 ( .a(n_1896), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__Q), .c(FE_OFN706_n_8119), .o(TIMEBOOST_net_11140) );
in01f02 FE_RC_1443_0 ( .a(n_12753), .o(FE_RN_909_0) );
in01f02 FE_RC_1444_0 ( .a(FE_RN_908_0), .o(FE_RN_910_0) );
na02s01 TIMEBOOST_cell_45744 ( .a(TIMEBOOST_net_15110), .b(FE_OFN706_n_8119), .o(TIMEBOOST_net_11038) );
na02s02 TIMEBOOST_cell_44892 ( .a(TIMEBOOST_net_14684), .b(g65747_db), .o(n_1925) );
in01f02 FE_RC_1447_0 ( .a(n_16022), .o(FE_RN_911_0) );
no02f04 FE_RC_1448_0 ( .a(n_15919), .b(FE_RN_911_0), .o(n_15914) );
in01f02 FE_RC_1449_0 ( .a(FE_RN_912_0), .o(n_16313) );
na02f02 FE_RC_1450_0 ( .a(n_16554), .b(n_16547), .o(FE_RN_912_0) );
in01f02 FE_RC_1451_0 ( .a(n_12257), .o(FE_RN_913_0) );
in01f02 FE_RC_1452_0 ( .a(n_11975), .o(FE_RN_914_0) );
no02f02 FE_RC_1453_0 ( .a(FE_RN_913_0), .b(FE_RN_914_0), .o(n_16411) );
in01f02 FE_RC_1454_0 ( .a(n_12031), .o(FE_RN_915_0) );
no02f02 FE_RC_1455_0 ( .a(FE_RN_25_0), .b(FE_RN_915_0), .o(FE_RN_26_0) );
in01f02 FE_RC_1456_0 ( .a(n_15935), .o(FE_RN_916_0) );
in01f02 FE_RC_1457_0 ( .a(n_15937), .o(FE_RN_917_0) );
ao22f02 FE_RC_1459_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__Q), .b(FE_OFN1479_n_16637), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__Q), .d(FE_OFN2195_n_9163), .o(n_11077) );
na02s01 TIMEBOOST_cell_16854 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__Q), .b(g64287_sb), .o(TIMEBOOST_net_3684) );
na04f04 FE_RC_1461_0 ( .a(FE_RN_917_0), .b(n_15940), .c(FE_RN_916_0), .d(n_15941), .o(n_15942) );
na03f02 FE_RC_148_0 ( .a(n_14269), .b(n_14456), .c(n_14557), .o(n_14602) );
in01f02 FE_RC_149_0 ( .a(n_10650), .o(FE_RN_87_0) );
in01f02 FE_RC_150_0 ( .a(n_10647), .o(FE_RN_88_0) );
no02f02 FE_RC_151_0 ( .a(FE_RN_87_0), .b(FE_RN_88_0), .o(FE_RN_89_0) );
in01f02 FE_RC_153_0 ( .a(n_10179), .o(FE_RN_90_0) );
in01f02 FE_RC_154_0 ( .a(n_10754), .o(FE_RN_91_0) );
no02f02 FE_RC_155_0 ( .a(FE_RN_90_0), .b(FE_RN_91_0), .o(FE_RN_92_0) );
na02s02 TIMEBOOST_cell_45232 ( .a(TIMEBOOST_net_14854), .b(FE_OFN1213_n_4151), .o(TIMEBOOST_net_12564) );
in01f02 FE_RC_157_0 ( .a(n_10750), .o(FE_RN_93_0) );
in01f02 FE_RC_158_0 ( .a(n_10747), .o(FE_RN_94_0) );
no02f02 FE_RC_159_0 ( .a(FE_RN_93_0), .b(FE_RN_94_0), .o(FE_RN_95_0) );
in01f06 FE_RC_15_0 ( .a(n_16159), .o(FE_RN_9_0) );
na02s02 TIMEBOOST_cell_22279 ( .a(n_10277), .b(TIMEBOOST_net_6396), .o(n_11875) );
in01f02 FE_RC_161_0 ( .a(n_10774), .o(FE_RN_96_0) );
in01f02 FE_RC_162_0 ( .a(n_10771), .o(FE_RN_97_0) );
no02f02 FE_RC_163_0 ( .a(FE_RN_96_0), .b(FE_RN_97_0), .o(FE_RN_98_0) );
na02m02 TIMEBOOST_cell_44657 ( .a(n_9205), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__Q), .o(TIMEBOOST_net_14567) );
in01f02 FE_RC_165_0 ( .a(n_10544), .o(FE_RN_99_0) );
in01f02 FE_RC_166_0 ( .a(n_10541), .o(FE_RN_100_0) );
no02f02 FE_RC_167_0 ( .a(FE_RN_99_0), .b(FE_RN_100_0), .o(FE_RN_101_0) );
na02m02 TIMEBOOST_cell_39542 ( .a(TIMEBOOST_net_2018), .b(TIMEBOOST_net_12009), .o(n_13426) );
in01f08 FE_RC_169_0 ( .a(parchk_pci_cbe_reg_in_1236), .o(FE_RN_102_0) );
in01f06 FE_RC_170_0 ( .a(n_2071), .o(FE_RN_103_0) );
na02m02 TIMEBOOST_cell_42157 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__Q), .b(n_9667), .o(TIMEBOOST_net_13317) );
na02f02 TIMEBOOST_cell_42158 ( .a(TIMEBOOST_net_13317), .b(FE_OFN1384_n_8567), .o(TIMEBOOST_net_12281) );
in01f02 FE_RC_173_0 ( .a(n_12922), .o(FE_RN_105_0) );
in01f02 FE_RC_174_0 ( .a(n_12923), .o(FE_RN_106_0) );
no02f02 FE_RC_175_0 ( .a(FE_RN_105_0), .b(FE_RN_106_0), .o(FE_RN_107_0) );
in01f02 FE_RC_178_0 ( .a(n_12949), .o(FE_RN_108_0) );
in01f02 FE_RC_179_0 ( .a(n_12950), .o(FE_RN_109_0) );
na02s01 TIMEBOOST_cell_42902 ( .a(TIMEBOOST_net_13689), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_11166) );
no02f02 FE_RC_180_0 ( .a(FE_RN_108_0), .b(FE_RN_109_0), .o(FE_RN_110_0) );
na02s02 TIMEBOOST_cell_45233 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__14__Q), .b(n_4436), .o(TIMEBOOST_net_14855) );
in01f02 FE_RC_182_0 ( .a(n_12889), .o(FE_RN_111_0) );
in01f02 FE_RC_183_0 ( .a(n_12890), .o(FE_RN_112_0) );
no02f02 FE_RC_184_0 ( .a(FE_RN_112_0), .b(FE_RN_111_0), .o(FE_RN_113_0) );
in01f02 FE_RC_186_0 ( .a(n_12913), .o(FE_RN_114_0) );
in01f02 FE_RC_187_0 ( .a(n_12912), .o(FE_RN_115_0) );
no02f02 FE_RC_188_0 ( .a(FE_RN_115_0), .b(FE_RN_114_0), .o(FE_RN_116_0) );
na03f02 FE_RC_189_0 ( .a(n_13118), .b(FE_RN_116_0), .c(n_12795), .o(n_13320) );
na02f02 TIMEBOOST_cell_38912 ( .a(TIMEBOOST_net_11694), .b(FE_OFN2200_n_10256), .o(TIMEBOOST_net_10700) );
in01s01 FE_RC_196_0 ( .a(n_16635), .o(FE_RN_120_0) );
in01s02 FE_RC_197_0 ( .a(n_1963), .o(FE_RN_121_0) );
no02s02 FE_RC_198_0 ( .a(FE_RN_120_0), .b(FE_RN_121_0), .o(FE_RN_122_0) );
na02s01 TIMEBOOST_cell_43033 ( .a(FE_OFN201_n_9230), .b(g58410_sb), .o(TIMEBOOST_net_13755) );
in01f02 FE_RC_201_0 ( .a(n_13672), .o(FE_RN_124_0) );
na03s02 TIMEBOOST_cell_38409 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__Q), .b(FE_OFN1112_g64577_p), .c(n_4006), .o(TIMEBOOST_net_11443) );
na02m02 TIMEBOOST_cell_43815 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__Q), .b(n_9090), .o(TIMEBOOST_net_14146) );
in01f02 FE_RC_205_0 ( .a(n_13651), .o(FE_RN_127_0) );
na02s01 TIMEBOOST_cell_36309 ( .a(parchk_pci_ad_reg_in_1213), .b(g67059_db), .o(TIMEBOOST_net_10393) );
na02f02 TIMEBOOST_cell_40918 ( .a(TIMEBOOST_net_12697), .b(g57237_sb), .o(n_11519) );
in01f02 FE_RC_209_0 ( .a(n_13661), .o(FE_RN_130_0) );
na02s01 TIMEBOOST_cell_44789 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__Q), .b(FE_OFN527_n_9899), .o(TIMEBOOST_net_14633) );
na02s01 TIMEBOOST_cell_30916 ( .a(pci_target_unit_pcit_if_strd_addr_in_695), .b(pci_target_unit_del_sync_addr_in_213), .o(TIMEBOOST_net_9369) );
na02f02 TIMEBOOST_cell_22064 ( .a(n_13997), .b(TIMEBOOST_net_2873), .o(TIMEBOOST_net_6289) );
na04f04 FE_RC_217_0 ( .a(n_14960), .b(n_14142), .c(n_14961), .d(n_14144), .o(n_16222) );
in01f02 FE_RC_218_0 ( .a(n_11733), .o(FE_RN_135_0) );
in01f02 FE_RC_219_0 ( .a(n_10908), .o(FE_RN_136_0) );
no02f02 FE_RC_220_0 ( .a(FE_RN_135_0), .b(FE_RN_136_0), .o(FE_RN_137_0) );
na02s01 TIMEBOOST_cell_16874 ( .a(pci_target_unit_fifos_pcir_data_in_172), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__Q), .o(TIMEBOOST_net_3694) );
in01f02 FE_RC_222_0 ( .a(n_10699), .o(FE_RN_138_0) );
in01f02 FE_RC_223_0 ( .a(n_10702), .o(FE_RN_139_0) );
no02f02 FE_RC_224_0 ( .a(FE_RN_138_0), .b(FE_RN_139_0), .o(FE_RN_140_0) );
na02s01 TIMEBOOST_cell_41841 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__Q), .b(FE_OFN553_n_9864), .o(TIMEBOOST_net_13159) );
in01f02 FE_RC_227_0 ( .a(n_11719), .o(FE_RN_141_0) );
in01f02 FE_RC_228_0 ( .a(n_10866), .o(FE_RN_142_0) );
no02f02 FE_RC_229_0 ( .a(FE_RN_141_0), .b(FE_RN_142_0), .o(FE_RN_143_0) );
na02s01 TIMEBOOST_cell_45134 ( .a(TIMEBOOST_net_14805), .b(FE_OFN1125_g64577_p), .o(TIMEBOOST_net_11434) );
in01f02 FE_RC_231_0 ( .a(n_10608), .o(FE_RN_144_0) );
in01f02 FE_RC_232_0 ( .a(n_11735), .o(FE_RN_145_0) );
no02f02 FE_RC_233_0 ( .a(FE_RN_144_0), .b(FE_RN_145_0), .o(FE_RN_146_0) );
na02m02 TIMEBOOST_cell_43566 ( .a(TIMEBOOST_net_14021), .b(FE_OFN1315_n_6624), .o(TIMEBOOST_net_12254) );
in01f06 FE_RC_238_0 ( .a(FE_OCPN1850_n_15998), .o(FE_RN_147_0) );
in01f06 FE_RC_239_0 ( .a(FE_OCPN1852_n_16538), .o(FE_RN_148_0) );
na02f10 FE_RC_240_0 ( .a(FE_RN_148_0), .b(FE_RN_147_0), .o(FE_RN_149_0) );
in01f02 FE_RC_242_0 ( .a(n_1399), .o(FE_RN_150_0) );
in01f02 FE_RC_243_0 ( .a(n_2227), .o(FE_RN_151_0) );
na02s02 TIMEBOOST_cell_45234 ( .a(TIMEBOOST_net_14855), .b(FE_OFN1241_n_4092), .o(TIMEBOOST_net_12566) );
na02s02 TIMEBOOST_cell_45235 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__Q), .b(n_3579), .o(TIMEBOOST_net_14856) );
in01f02 FE_RC_246_0 ( .a(n_2250), .o(FE_RN_153_0) );
in01f02 FE_RC_247_0 ( .a(n_3466), .o(FE_RN_154_0) );
na02s01 TIMEBOOST_cell_36319 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__Q), .b(g65964_sb), .o(TIMEBOOST_net_10398) );
na02s01 TIMEBOOST_cell_15834 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_94), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3174) );
na02s01 TIMEBOOST_cell_36488 ( .a(TIMEBOOST_net_10482), .b(g66398_sb), .o(n_2545) );
in01m01 FE_RC_251_0 ( .a(n_16160), .o(FE_RN_156_0) );
no02m02 FE_RC_253_0 ( .a(FE_RN_156_0), .b(FE_RN_9_0), .o(FE_RN_158_0) );
na02s01 TIMEBOOST_cell_30870 ( .a(FE_OFN219_n_9853), .b(g57986_sb), .o(TIMEBOOST_net_9346) );
in01m02 FE_RC_255_0 ( .a(n_4874), .o(FE_RN_159_0) );
in01f02 FE_RC_256_0 ( .a(n_3432), .o(FE_RN_160_0) );
na02s02 TIMEBOOST_cell_39544 ( .a(TIMEBOOST_net_12010), .b(g59089_sb), .o(n_8589) );
na02s01 TIMEBOOST_cell_39261 ( .a(pci_target_unit_fifos_pciw_addr_data_in_136), .b(g64150_sb), .o(TIMEBOOST_net_11869) );
na02s01 TIMEBOOST_cell_42732 ( .a(TIMEBOOST_net_13604), .b(FE_OFN707_n_8119), .o(TIMEBOOST_net_11105) );
na02s02 TIMEBOOST_cell_43008 ( .a(TIMEBOOST_net_13742), .b(g58301_db), .o(n_9029) );
na03s02 TIMEBOOST_cell_38157 ( .a(TIMEBOOST_net_3548), .b(g64357_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__Q), .o(TIMEBOOST_net_11317) );
in01f02 FE_RC_282_0 ( .a(FE_RN_176_0), .o(n_13577) );
na02s02 TIMEBOOST_cell_38106 ( .a(TIMEBOOST_net_11291), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_4700) );
na03f02 FE_RC_285_0 ( .a(n_14292), .b(n_14473), .c(n_14565), .o(n_14610) );
na03f02 FE_RC_286_0 ( .a(n_14273), .b(n_14460), .c(n_14559), .o(n_14604) );
in01f02 FE_RC_287_0 ( .a(n_10951), .o(FE_RN_177_0) );
in01f02 FE_RC_288_0 ( .a(n_10691), .o(FE_RN_178_0) );
no02f04 FE_RC_289_0 ( .a(FE_RN_177_0), .b(FE_RN_178_0), .o(FE_RN_179_0) );
in01f02 FE_RC_291_0 ( .a(n_10875), .o(FE_RN_180_0) );
in01f02 FE_RC_292_0 ( .a(n_10873), .o(FE_RN_181_0) );
no02f02 FE_RC_293_0 ( .a(FE_RN_180_0), .b(FE_RN_181_0), .o(FE_RN_182_0) );
in01f02 FE_RC_295_0 ( .a(n_10579), .o(FE_RN_183_0) );
in01f02 FE_RC_296_0 ( .a(n_11726), .o(FE_RN_184_0) );
no02f02 FE_RC_297_0 ( .a(FE_RN_183_0), .b(FE_RN_184_0), .o(FE_RN_185_0) );
na02s02 TIMEBOOST_cell_16838 ( .a(n_3770), .b(g64872_sb), .o(TIMEBOOST_net_3676) );
in01f02 FE_RC_299_0 ( .a(n_10891), .o(FE_RN_186_0) );
in01f02 FE_RC_300_0 ( .a(n_10576), .o(FE_RN_187_0) );
no02f02 FE_RC_301_0 ( .a(FE_RN_186_0), .b(FE_RN_187_0), .o(FE_RN_188_0) );
na02s01 TIMEBOOST_cell_16826 ( .a(n_3749), .b(g65062_sb), .o(TIMEBOOST_net_3670) );
in01f02 FE_RC_303_0 ( .a(n_10109), .o(FE_RN_189_0) );
in01f02 FE_RC_304_0 ( .a(n_10685), .o(FE_RN_190_0) );
no02f02 FE_RC_305_0 ( .a(FE_RN_189_0), .b(FE_RN_190_0), .o(FE_RN_191_0) );
na02s01 TIMEBOOST_cell_16837 ( .a(TIMEBOOST_net_3675), .b(g65342_db), .o(n_3546) );
in01f02 FE_RC_307_0 ( .a(n_10147), .o(FE_RN_192_0) );
in01f02 FE_RC_308_0 ( .a(n_10970), .o(FE_RN_193_0) );
no02f02 FE_RC_309_0 ( .a(FE_RN_192_0), .b(FE_RN_193_0), .o(FE_RN_194_0) );
na02s01 TIMEBOOST_cell_45085 ( .a(g58040_sb), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_14781) );
in01f02 FE_RC_311_0 ( .a(n_10041), .o(FE_RN_195_0) );
in01f02 FE_RC_312_0 ( .a(n_10038), .o(FE_RN_196_0) );
no02f02 FE_RC_313_0 ( .a(FE_RN_195_0), .b(FE_RN_196_0), .o(FE_RN_197_0) );
na02s02 TIMEBOOST_cell_45196 ( .a(TIMEBOOST_net_14836), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_12649) );
in01s01 FE_RC_315_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__Q), .o(FE_RN_198_0) );
in01f02 FE_RC_316_0 ( .a(FE_OFN1453_n_10588), .o(FE_RN_199_0) );
no02f02 FE_RC_317_0 ( .a(FE_RN_198_0), .b(FE_RN_199_0), .o(FE_RN_200_0) );
no02f02 FE_RC_318_0 ( .a(FE_RN_200_0), .b(n_15590), .o(n_15591) );
in01f02 FE_RC_319_0 ( .a(n_12914), .o(FE_RN_201_0) );
na02f02 TIMEBOOST_cell_41116 ( .a(TIMEBOOST_net_12796), .b(g57380_sb), .o(n_11367) );
in01f02 FE_RC_320_0 ( .a(n_12915), .o(FE_RN_202_0) );
no02f02 FE_RC_321_0 ( .a(FE_RN_201_0), .b(FE_RN_202_0), .o(FE_RN_203_0) );
na04f04 FE_RC_324_0 ( .a(n_12122), .b(n_11992), .c(n_12276), .d(n_12393), .o(n_12920) );
na02s02 TIMEBOOST_cell_43053 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__Q), .b(n_3776), .o(TIMEBOOST_net_13765) );
na02s02 TIMEBOOST_cell_43009 ( .a(n_1094), .b(wishbone_slave_unit_fifos_outGreyCount_1_), .o(TIMEBOOST_net_13743) );
na02f02 TIMEBOOST_cell_44683 ( .a(TIMEBOOST_net_10052), .b(FE_OFN1376_n_8567), .o(TIMEBOOST_net_14580) );
na02f02 TIMEBOOST_cell_44684 ( .a(TIMEBOOST_net_14580), .b(g57315_sb), .o(n_11436) );
ao22f02 FE_RC_329_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__Q), .b(FE_OFN1731_n_9975), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__Q), .d(FE_OCP_RBN2005_FE_RN_459_0), .o(n_9332) );
na03f40 FE_RC_32_0 ( .a(n_326), .b(n_15204), .c(n_16910), .o(n_15317) );
na02s01 TIMEBOOST_cell_30776 ( .a(parchk_pci_ad_reg_in_1231), .b(pci_target_unit_del_sync_addr_in_230), .o(TIMEBOOST_net_9299) );
in01m08 FE_RC_335_0 ( .a(pci_target_unit_wishbone_master_read_bound), .o(FE_RN_207_0) );
in01f02 FE_RC_336_0 ( .a(n_16275), .o(FE_RN_208_0) );
no02f04 FE_RC_337_0 ( .a(FE_RN_207_0), .b(FE_RN_208_0), .o(FE_RN_209_0) );
na02s01 TIMEBOOST_cell_38461 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__Q), .b(g58266_sb), .o(TIMEBOOST_net_11469) );
na02f02 TIMEBOOST_cell_22074 ( .a(n_13873), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__Q), .o(TIMEBOOST_net_6294) );
in01s01 TIMEBOOST_cell_45864 ( .a(TIMEBOOST_net_15171), .o(TIMEBOOST_net_15170) );
in01m02 FE_RC_341_0 ( .a(n_13667), .o(FE_RN_211_0) );
na02f02 TIMEBOOST_cell_42500 ( .a(TIMEBOOST_net_13488), .b(g57137_sb), .o(n_11613) );
na02s02 TIMEBOOST_cell_42068 ( .a(TIMEBOOST_net_13272), .b(g62557_sb), .o(n_6448) );
na02s01 TIMEBOOST_cell_36289 ( .a(n_2509), .b(g67056_db), .o(TIMEBOOST_net_10383) );
in01f02 FE_RC_345_0 ( .a(n_13571), .o(FE_RN_214_0) );
in01f02 FE_RC_346_0 ( .a(FE_RN_215_0), .o(n_13768) );
na02f04 FE_RC_347_0 ( .a(FE_RN_214_0), .b(FE_RN_213_0), .o(FE_RN_215_0) );
na02f06 FE_RC_348_0 ( .a(n_16492), .b(n_16494), .o(FE_RN_216_0) );
in01f04 FE_RC_349_0 ( .a(n_16490), .o(FE_RN_217_0) );
in01f02 FE_RC_34_0 ( .a(n_15645), .o(FE_RN_15_0) );
in01f08 FE_RC_350_0 ( .a(FE_RN_218_0), .o(n_16495) );
no02f08 FE_RC_351_0 ( .a(FE_RN_216_0), .b(FE_RN_217_0), .o(FE_RN_218_0) );
na02s01 TIMEBOOST_cell_45086 ( .a(TIMEBOOST_net_14781), .b(g58040_db), .o(n_9748) );
in01f02 FE_RC_353_0 ( .a(n_10075), .o(FE_RN_219_0) );
in01f02 FE_RC_354_0 ( .a(n_10659), .o(FE_RN_220_0) );
no02f02 FE_RC_355_0 ( .a(FE_RN_219_0), .b(FE_RN_220_0), .o(FE_RN_221_0) );
na02s01 TIMEBOOST_cell_16833 ( .a(TIMEBOOST_net_3673), .b(g64796_db), .o(n_3759) );
in01f06 FE_RC_358_0 ( .a(pci_target_unit_pcit_if_strd_bc_in_717), .o(FE_RN_222_0) );
in01m10 FE_RC_359_0 ( .a(pci_target_unit_pcit_if_strd_bc_in_718), .o(FE_RN_223_0) );
no02f08 FE_RC_360_0 ( .a(FE_RN_222_0), .b(FE_RN_223_0), .o(FE_RN_224_0) );
na02f06 FE_RC_361_0 ( .a(FE_RN_224_0), .b(n_1219), .o(n_1507) );
na02s02 TIMEBOOST_cell_43529 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__Q), .b(n_3644), .o(TIMEBOOST_net_14003) );
in01f02 FE_RC_364_0 ( .a(n_10901), .o(FE_RN_225_0) );
in01f02 FE_RC_365_0 ( .a(n_10902), .o(FE_RN_226_0) );
no02f02 FE_RC_366_0 ( .a(FE_RN_225_0), .b(FE_RN_226_0), .o(FE_RN_227_0) );
na02s02 TIMEBOOST_cell_39546 ( .a(TIMEBOOST_net_12011), .b(g58290_db), .o(n_9514) );
in01f02 FE_RC_368_0 ( .a(n_10569), .o(FE_RN_228_0) );
in01f02 FE_RC_369_0 ( .a(n_11723), .o(FE_RN_229_0) );
no02f02 FE_RC_370_0 ( .a(FE_RN_228_0), .b(FE_RN_229_0), .o(FE_RN_230_0) );
na02s01 TIMEBOOST_cell_16825 ( .a(TIMEBOOST_net_3669), .b(g65311_db), .o(n_3569) );
na02s01 TIMEBOOST_cell_16850 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__Q), .b(g64279_sb), .o(TIMEBOOST_net_3682) );
na02f04 TIMEBOOST_cell_44872 ( .a(TIMEBOOST_net_14674), .b(n_4674), .o(TIMEBOOST_net_1424) );
na02s02 TIMEBOOST_cell_39548 ( .a(TIMEBOOST_net_12012), .b(g58283_db), .o(n_9519) );
in01f02 FE_RC_375_0 ( .a(n_9979), .o(FE_RN_231_0) );
in01f02 FE_RC_376_0 ( .a(n_10877), .o(FE_RN_232_0) );
no02f02 FE_RC_377_0 ( .a(FE_RN_231_0), .b(FE_RN_232_0), .o(FE_RN_233_0) );
na03f02 FE_RC_379_0 ( .a(n_16228), .b(n_16230), .c(n_16227), .o(n_16231) );
na03f02 FE_RC_380_0 ( .a(n_16625), .b(n_16624), .c(n_14446), .o(n_14597) );
na02m06 TIMEBOOST_cell_45020 ( .a(TIMEBOOST_net_14748), .b(FE_OFN1147_n_13249), .o(TIMEBOOST_net_13205) );
na03f02 FE_RC_382_0 ( .a(n_14402), .b(n_14534), .c(n_14494), .o(n_14578) );
na03f02 FE_RC_383_0 ( .a(n_14435), .b(n_14250), .c(n_14547), .o(n_14592) );
na03f02 FE_RC_384_0 ( .a(n_14541), .b(n_14420), .c(n_14421), .o(n_14585) );
na03f02 FE_RC_385_0 ( .a(n_14286), .b(n_14563), .c(n_14468), .o(n_14608) );
na02s02 TIMEBOOST_cell_43647 ( .a(n_3612), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__Q), .o(TIMEBOOST_net_14062) );
na02f02 TIMEBOOST_cell_41935 ( .a(TIMEBOOST_net_9851), .b(FE_OCPN1911_FE_OFN1152_n_13249), .o(TIMEBOOST_net_13206) );
na03f02 FE_RC_389_0 ( .a(n_16622), .b(n_16623), .c(n_14261), .o(n_14598) );
na02m02 TIMEBOOST_cell_41944 ( .a(TIMEBOOST_net_13210), .b(TIMEBOOST_net_9874), .o(n_13502) );
na03f02 FE_RC_391_0 ( .a(n_12960), .b(n_13034), .c(n_12677), .o(n_13319) );
in01f02 FE_RC_392_0 ( .a(n_12721), .o(FE_RN_234_0) );
in01f02 FE_RC_393_0 ( .a(n_12929), .o(FE_RN_235_0) );
no02f02 FE_RC_394_0 ( .a(FE_RN_235_0), .b(FE_RN_234_0), .o(FE_RN_236_0) );
na04f04 FE_RC_396_0 ( .a(n_13054), .b(n_12902), .c(n_12791), .d(n_12903), .o(n_13137) );
na02s02 TIMEBOOST_cell_43648 ( .a(TIMEBOOST_net_14062), .b(FE_OFN1231_n_6391), .o(TIMEBOOST_net_12630) );
in01s01 FE_RC_401_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__Q), .o(FE_RN_237_0) );
in01f02 FE_RC_402_0 ( .a(FE_OFN1565_n_12502), .o(FE_RN_238_0) );
no02f02 FE_RC_403_0 ( .a(FE_RN_237_0), .b(FE_RN_238_0), .o(FE_RN_239_0) );
no02f02 FE_RC_404_0 ( .a(FE_RN_239_0), .b(n_12460), .o(n_12799) );
in01s01 FE_RC_405_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__Q), .o(FE_RN_240_0) );
in01f02 FE_RC_406_0 ( .a(FE_OFN1563_n_12502), .o(FE_RN_241_0) );
no02f02 FE_RC_407_0 ( .a(FE_RN_240_0), .b(FE_RN_241_0), .o(FE_RN_242_0) );
no02f02 FE_RC_408_0 ( .a(n_12446), .b(FE_RN_242_0), .o(n_12778) );
in01s01 FE_RC_409_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__Q), .o(FE_RN_243_0) );
in01m01 FE_RC_410_0 ( .a(FE_OFN1563_n_12502), .o(FE_RN_244_0) );
no02f02 FE_RC_411_0 ( .a(FE_RN_243_0), .b(FE_RN_244_0), .o(FE_RN_245_0) );
no02f02 FE_RC_412_0 ( .a(n_12457), .b(FE_RN_245_0), .o(n_12795) );
in01s01 FE_RC_413_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__Q), .o(FE_RN_246_0) );
in01f01 FE_RC_414_0 ( .a(FE_OFN1563_n_12502), .o(FE_RN_247_0) );
no02f02 FE_RC_415_0 ( .a(FE_RN_246_0), .b(FE_RN_247_0), .o(FE_RN_248_0) );
no02f02 FE_RC_416_0 ( .a(FE_RN_248_0), .b(n_12454), .o(n_12790) );
na02m02 TIMEBOOST_cell_41584 ( .a(FE_OFN1439_n_9372), .b(TIMEBOOST_net_13030), .o(TIMEBOOST_net_11668) );
na04f04 FE_RC_418_0 ( .a(n_11961), .b(n_12379), .c(n_12117), .d(n_11962), .o(n_12904) );
na02s02 TIMEBOOST_cell_45598 ( .a(TIMEBOOST_net_15037), .b(g65232_sb), .o(n_2655) );
in01f02 FE_RC_41_0 ( .a(n_12881), .o(FE_RN_18_0) );
in01f02 FE_RC_422_0 ( .a(n_11991), .o(FE_RN_249_0) );
in01f02 FE_RC_423_0 ( .a(n_11990), .o(FE_RN_250_0) );
no02f02 FE_RC_424_0 ( .a(FE_RN_250_0), .b(FE_RN_249_0), .o(FE_RN_251_0) );
na02f02 FE_RC_425_0 ( .a(FE_RN_29_0), .b(FE_RN_251_0), .o(n_12816) );
in01f02 FE_RC_42_0 ( .a(n_12880), .o(FE_RN_19_0) );
in01f02 FE_RC_437_0 ( .a(FE_RN_259_0), .o(n_13410) );
na02f02 FE_RC_438_0 ( .a(n_13122), .b(n_16299), .o(FE_RN_259_0) );
in01s10 FE_RC_439_0 ( .a(pci_target_unit_pci_target_sm_wr_to_fifo), .o(FE_RN_260_0) );
no02f02 FE_RC_43_0 ( .a(FE_RN_18_0), .b(FE_RN_19_0), .o(FE_RN_20_0) );
in01f04 FE_RC_440_0 ( .a(n_978), .o(FE_RN_261_0) );
no02f06 FE_RC_441_0 ( .a(FE_RN_261_0), .b(FE_RN_260_0), .o(FE_RN_262_0) );
in01f02 FE_RC_442_0 ( .a(n_653), .o(FE_RN_263_0) );
no02f04 FE_RC_443_0 ( .a(pci_target_unit_pci_target_sm_state_transfere_reg), .b(FE_RN_263_0), .o(FE_RN_264_0) );
na02s02 TIMEBOOST_cell_45599 ( .a(TIMEBOOST_net_9368), .b(FE_OFN789_n_2678), .o(TIMEBOOST_net_15038) );
na02s01 TIMEBOOST_cell_38552 ( .a(TIMEBOOST_net_11514), .b(g62046_sb), .o(n_7766) );
na03s01 TIMEBOOST_cell_6271 ( .a(FE_OFN254_n_9825), .b(g58010_sb), .c(g58038_db), .o(n_9751) );
na02s01 TIMEBOOST_cell_37274 ( .a(TIMEBOOST_net_10875), .b(g64797_sb), .o(TIMEBOOST_net_225) );
no02f02 FE_RC_448_0 ( .a(n_1724), .b(pci_target_unit_pci_target_sm_cnf_progress), .o(FE_RN_269_0) );
in01f02 FE_RC_449_0 ( .a(n_2031), .o(FE_RN_270_0) );
na02f02 TIMEBOOST_cell_40920 ( .a(TIMEBOOST_net_12698), .b(g57042_sb), .o(n_11692) );
in01s08 FE_RC_450_0 ( .a(pci_target_unit_pci_target_sm_state_backoff_reg_reg_Q), .o(FE_RN_271_0) );
na02s02 TIMEBOOST_cell_42066 ( .a(TIMEBOOST_net_13271), .b(g62934_sb), .o(n_6013) );
na02s01 TIMEBOOST_cell_31073 ( .a(TIMEBOOST_net_9447), .b(g65006_db), .o(n_4350) );
oa12f04 FE_RC_453_0 ( .a(FE_RN_267_0), .b(FE_RN_268_0), .c(FE_RN_273_0), .o(n_8566) );
in01f20 FE_RC_454_0 ( .a(n_2078), .o(FE_RN_274_0) );
na02f20 FE_RC_455_0 ( .a(FE_RN_274_0), .b(n_525), .o(n_16287) );
in01s01 FE_RC_456_0 ( .a(parchk_pci_cbe_out_in_1204), .o(FE_RN_275_0) );
in01f02 FE_RC_457_0 ( .a(n_4702), .o(FE_RN_276_0) );
ao22f02 FE_RC_458_0 ( .a(FE_RN_275_0), .b(FE_RN_276_0), .c(parchk_pci_cbe_out_in_1204), .d(n_4702), .o(n_4703) );
in01s01 FE_RC_460_0 ( .a(n_532), .o(FE_RN_278_0) );
na02s02 FE_RC_461_0 ( .a(n_1196), .b(FE_RN_278_0), .o(FE_RN_279_0) );
na02f02 FE_RC_462_0 ( .a(FE_RN_279_0), .b(n_15292), .o(FE_RN_280_0) );
in01m02 FE_RC_463_0 ( .a(n_15607), .o(FE_RN_281_0) );
na02s01 TIMEBOOST_cell_42695 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__Q), .b(FE_OFN1651_n_9428), .o(TIMEBOOST_net_13586) );
na02s01 TIMEBOOST_cell_15961 ( .a(TIMEBOOST_net_3237), .b(g65957_db), .o(n_2165) );
no02f04 FE_RC_466_0 ( .a(FE_RN_283_0), .b(FE_RN_280_0), .o(n_15611) );
in01s06 FE_RC_467_0 ( .a(parchk_pci_cbe_out_in), .o(FE_RN_284_0) );
in01f02 FE_RC_468_0 ( .a(n_4703), .o(FE_RN_285_0) );
na02f02 TIMEBOOST_cell_43816 ( .a(TIMEBOOST_net_14146), .b(FE_OFN1394_n_8567), .o(TIMEBOOST_net_12950) );
na02s02 TIMEBOOST_cell_45236 ( .a(TIMEBOOST_net_14856), .b(FE_OFN1288_n_4098), .o(TIMEBOOST_net_12568) );
na04f20 FE_RC_481_0 ( .a(pci_target_unit_pci_target_sm_rd_from_fifo), .b(pci_target_unit_pci_target_sm_same_read_reg), .c(n_1724), .d(n_653), .o(FE_RN_294_0) );
no02f08 FE_RC_482_0 ( .a(FE_RN_294_0), .b(n_1435), .o(n_15401) );
no02f20 FE_RC_483_0 ( .a(wbm_ack_i), .b(FE_RN_295_0), .o(n_1445) );
na02f40 FE_RC_484_0 ( .a(n_705), .b(wbm_err_i), .o(FE_RN_295_0) );
na04f04 FE_RC_490_0 ( .a(n_11092), .b(n_11093), .c(n_11094), .d(n_11091), .o(n_12544) );
na02m02 TIMEBOOST_cell_43817 ( .a(n_9776), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__Q), .o(TIMEBOOST_net_14147) );
in01f10 FE_RC_493_0 ( .a(FE_RN_299_0), .o(n_15981) );
na02s02 TIMEBOOST_cell_41741 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__Q), .b(g58264_sb), .o(TIMEBOOST_net_13109) );
na02f02 FE_RC_497_0 ( .a(n_16268), .b(n_16511), .o(n_14967) );
na02s02 TIMEBOOST_cell_45215 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__15__Q), .b(n_3686), .o(TIMEBOOST_net_14846) );
na02f02 TIMEBOOST_cell_40888 ( .a(TIMEBOOST_net_12682), .b(g57489_db), .o(n_11247) );
na02f02 FE_RC_49_0 ( .a(FE_RN_23_0), .b(n_13061), .o(n_13321) );
na02f02 TIMEBOOST_cell_4173 ( .a(TIMEBOOST_net_666), .b(n_9325), .o(n_12163) );
in01m10 FE_RC_501_0 ( .a(pciu_bar0_in_378), .o(FE_RN_303_0) );
in01f06 FE_RC_502_0 ( .a(n_396), .o(FE_RN_304_0) );
ao22f06 FE_RC_503_0 ( .a(FE_RN_303_0), .b(FE_RN_304_0), .c(pciu_bar0_in_378), .d(n_396), .o(FE_RN_305_0) );
na02s02 TIMEBOOST_cell_37985 ( .a(g62848_sb), .b(g62848_db), .o(TIMEBOOST_net_11231) );
no02m06 FE_RC_505_0 ( .a(pciu_bar0_in_379), .b(parchk_pci_ad_reg_in_1235), .o(FE_RN_307_0) );
ao12f02 FE_RC_506_0 ( .a(FE_RN_307_0), .b(pciu_bar0_in_379), .c(parchk_pci_ad_reg_in_1235), .o(FE_RN_308_0) );
no02m10 FE_RC_507_0 ( .a(pciu_bar0_in_376), .b(parchk_pci_ad_reg_in_1232), .o(FE_RN_309_0) );
ao12f04 FE_RC_508_0 ( .a(FE_RN_309_0), .b(pciu_bar0_in_376), .c(parchk_pci_ad_reg_in_1232), .o(FE_RN_310_0) );
no02m10 FE_RC_509_0 ( .a(pciu_bar0_in_377), .b(parchk_pci_ad_reg_in_1233), .o(FE_RN_311_0) );
ao12f04 FE_RC_510_0 ( .a(FE_RN_311_0), .b(pciu_bar0_in_377), .c(parchk_pci_ad_reg_in_1233), .o(FE_RN_312_0) );
no02f04 FE_RC_511_0 ( .a(FE_RN_310_0), .b(FE_RN_312_0), .o(FE_RN_313_0) );
no02m10 FE_RC_512_0 ( .a(pciu_bar0_in), .b(parchk_pci_ad_reg_in_1216), .o(FE_RN_314_0) );
ao12f06 FE_RC_513_0 ( .a(FE_RN_314_0), .b(pciu_bar0_in), .c(parchk_pci_ad_reg_in_1216), .o(FE_RN_315_0) );
no02m10 FE_RC_514_0 ( .a(pciu_bar0_in_362), .b(parchk_pci_ad_reg_in_1218), .o(FE_RN_316_0) );
ao12f06 FE_RC_515_0 ( .a(FE_RN_316_0), .b(pciu_bar0_in_362), .c(parchk_pci_ad_reg_in_1218), .o(FE_RN_317_0) );
na02m10 FE_RC_516_0 ( .a(pciu_bar0_in_363), .b(parchk_pci_ad_reg_in_1219), .o(FE_RN_318_0) );
oa12f04 FE_RC_517_0 ( .a(FE_RN_318_0), .b(pciu_bar0_in_363), .c(parchk_pci_ad_reg_in_1219), .o(FE_RN_319_0) );
na02m10 FE_RC_518_0 ( .a(pciu_bar0_in_361), .b(parchk_pci_ad_reg_in_1217), .o(FE_RN_320_0) );
oa12f04 FE_RC_519_0 ( .a(FE_RN_320_0), .b(pciu_bar0_in_361), .c(parchk_pci_ad_reg_in_1217), .o(FE_RN_321_0) );
in01f02 FE_RC_51_0 ( .a(n_12032), .o(FE_RN_25_0) );
na02f04 FE_RC_520_0 ( .a(FE_RN_319_0), .b(FE_RN_321_0), .o(FE_RN_322_0) );
na02s01 TIMEBOOST_cell_43034 ( .a(TIMEBOOST_net_13755), .b(g58410_db), .o(n_9207) );
na02m10 FE_RC_522_0 ( .a(pciu_bar0_in_367), .b(parchk_pci_ad_reg_in_1223), .o(FE_RN_324_0) );
oa12f04 FE_RC_523_0 ( .a(FE_RN_324_0), .b(pciu_bar0_in_367), .c(parchk_pci_ad_reg_in_1223), .o(FE_RN_325_0) );
na02m10 FE_RC_524_0 ( .a(pciu_bar0_in_364), .b(parchk_pci_ad_reg_in_1220), .o(FE_RN_326_0) );
oa12f04 FE_RC_525_0 ( .a(FE_RN_326_0), .b(pciu_bar0_in_364), .c(parchk_pci_ad_reg_in_1220), .o(FE_RN_327_0) );
na02f04 FE_RC_526_0 ( .a(FE_RN_325_0), .b(FE_RN_327_0), .o(FE_RN_328_0) );
no02f02 FE_RC_527_0 ( .a(pciu_bar0_in_365), .b(FE_OFN1780_parchk_pci_ad_reg_in_1221), .o(FE_RN_329_0) );
ao12f02 FE_RC_528_0 ( .a(FE_RN_329_0), .b(pciu_bar0_in_365), .c(FE_OFN1780_parchk_pci_ad_reg_in_1221), .o(FE_RN_330_0) );
no02f04 FE_RC_529_0 ( .a(pciu_bar0_in_366), .b(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(FE_RN_331_0) );
ao12f02 FE_RC_530_0 ( .a(FE_RN_331_0), .b(pciu_bar0_in_366), .c(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(FE_RN_332_0) );
na02s01 TIMEBOOST_cell_40404 ( .a(g63603_da), .b(TIMEBOOST_net_12440), .o(n_7207) );
na02m08 FE_RC_532_0 ( .a(pciu_bar0_in_368), .b(parchk_pci_ad_reg_in_1224), .o(FE_RN_334_0) );
oa12f04 FE_RC_533_0 ( .a(FE_RN_334_0), .b(pciu_bar0_in_368), .c(parchk_pci_ad_reg_in_1224), .o(FE_RN_335_0) );
na02m08 FE_RC_534_0 ( .a(pciu_bar0_in_369), .b(parchk_pci_ad_reg_in_1225), .o(FE_RN_336_0) );
oa12f04 FE_RC_535_0 ( .a(FE_RN_336_0), .b(pciu_bar0_in_369), .c(parchk_pci_ad_reg_in_1225), .o(FE_RN_337_0) );
na02f02 FE_RC_536_0 ( .a(FE_RN_335_0), .b(FE_RN_337_0), .o(FE_RN_338_0) );
na02m10 FE_RC_537_0 ( .a(pciu_bar0_in_373), .b(parchk_pci_ad_reg_in_1229), .o(FE_RN_339_0) );
oa12f04 FE_RC_538_0 ( .a(FE_RN_339_0), .b(pciu_bar0_in_373), .c(parchk_pci_ad_reg_in_1229), .o(FE_RN_340_0) );
na02m10 FE_RC_539_0 ( .a(pciu_bar0_in_374), .b(parchk_pci_ad_reg_in_1230), .o(FE_RN_341_0) );
na02s02 TIMEBOOST_cell_43519 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__Q), .b(n_3621), .o(TIMEBOOST_net_13998) );
oa12f04 FE_RC_540_0 ( .a(FE_RN_341_0), .b(pciu_bar0_in_374), .c(parchk_pci_ad_reg_in_1230), .o(FE_RN_342_0) );
na02f02 FE_RC_541_0 ( .a(FE_RN_340_0), .b(FE_RN_342_0), .o(FE_RN_343_0) );
na02m08 FE_RC_542_0 ( .a(pciu_bar0_in_370), .b(parchk_pci_ad_reg_in_1226), .o(FE_RN_344_0) );
oa12f04 FE_RC_543_0 ( .a(FE_RN_344_0), .b(pciu_bar0_in_370), .c(parchk_pci_ad_reg_in_1226), .o(FE_RN_345_0) );
na02m08 FE_RC_544_0 ( .a(pciu_bar0_in_371), .b(parchk_pci_ad_reg_in_1227), .o(FE_RN_346_0) );
oa12f04 FE_RC_545_0 ( .a(FE_RN_346_0), .b(pciu_bar0_in_371), .c(parchk_pci_ad_reg_in_1227), .o(FE_RN_347_0) );
na02f02 FE_RC_546_0 ( .a(FE_RN_345_0), .b(FE_RN_347_0), .o(FE_RN_348_0) );
na02m08 FE_RC_547_0 ( .a(pciu_bar0_in_372), .b(parchk_pci_ad_reg_in_1228), .o(FE_RN_349_0) );
oa12f04 FE_RC_548_0 ( .a(FE_RN_349_0), .b(pciu_bar0_in_372), .c(parchk_pci_ad_reg_in_1228), .o(FE_RN_350_0) );
na02m08 FE_RC_549_0 ( .a(pciu_bar0_in_375), .b(parchk_pci_ad_reg_in_1231), .o(FE_RN_351_0) );
in01f02 FE_RC_54_0 ( .a(n_12275), .o(FE_RN_27_0) );
oa12f04 FE_RC_550_0 ( .a(FE_RN_351_0), .b(pciu_bar0_in_375), .c(parchk_pci_ad_reg_in_1231), .o(FE_RN_352_0) );
na02f02 FE_RC_551_0 ( .a(FE_RN_350_0), .b(FE_RN_352_0), .o(FE_RN_353_0) );
na02f02 TIMEBOOST_cell_41420 ( .a(TIMEBOOST_net_12948), .b(g57152_sb), .o(n_11598) );
na03f06 TIMEBOOST_cell_33631 ( .a(n_15908), .b(n_319), .c(FE_OCP_RBN2221_n_15347), .o(g74563_p) );
no02f02 FE_RC_554_0 ( .a(FE_RN_308_0), .b(FE_RN_355_0), .o(FE_RN_356_0) );
na02m02 TIMEBOOST_cell_41659 ( .a(TIMEBOOST_net_6243), .b(n_16070), .o(TIMEBOOST_net_13068) );
in01f10 FE_RC_557_0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_control_in), .o(FE_RN_357_0) );
na02f10 FE_RC_558_0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_control_in_85), .b(FE_RN_357_0), .o(FE_RN_358_0) );
in01f02 FE_RC_559_0 ( .a(n_16980), .o(FE_RN_359_0) );
in01f02 FE_RC_55_0 ( .a(n_12274), .o(FE_RN_28_0) );
no02f04 FE_RC_560_0 ( .a(FE_RN_359_0), .b(FE_RN_358_0), .o(FE_RN_360_0) );
in01s01 FE_RC_562_0 ( .a(n_13763), .o(FE_RN_361_0) );
in01m02 FE_RC_563_0 ( .a(n_13666), .o(FE_RN_362_0) );
na03s02 TIMEBOOST_cell_36753 ( .a(g64340_da), .b(g64340_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__Q), .o(TIMEBOOST_net_10615) );
na02f02 TIMEBOOST_cell_42390 ( .a(TIMEBOOST_net_13433), .b(g57402_sb), .o(n_11340) );
na02f04 FE_RC_566_0 ( .a(n_13784), .b(FE_OFN1714_n_13650), .o(FE_RN_364_0) );
in01f02 FE_RC_567_0 ( .a(n_13566), .o(FE_RN_365_0) );
in01f02 FE_RC_568_0 ( .a(FE_RN_366_0), .o(n_13761) );
na02f04 FE_RC_569_0 ( .a(FE_RN_365_0), .b(FE_RN_364_0), .o(FE_RN_366_0) );
no02f02 FE_RC_56_0 ( .a(FE_RN_28_0), .b(FE_RN_27_0), .o(FE_RN_29_0) );
na02m02 TIMEBOOST_cell_11487 ( .a(n_14392), .b(TIMEBOOST_net_2310), .o(n_14397) );
in01f02 FE_RC_571_0 ( .a(n_13568), .o(FE_RN_368_0) );
in01f02 FE_RC_572_0 ( .a(FE_RN_369_0), .o(n_13764) );
na02f04 FE_RC_573_0 ( .a(FE_RN_367_0), .b(FE_RN_368_0), .o(FE_RN_369_0) );
in01s01 FE_RC_574_0 ( .a(n_7822), .o(FE_RN_370_0) );
in01f02 FE_RC_575_0 ( .a(n_13028), .o(FE_RN_371_0) );
in01s01 TIMEBOOST_cell_45886 ( .a(TIMEBOOST_net_15192), .o(TIMEBOOST_net_15193) );
na02m02 TIMEBOOST_cell_45237 ( .a(TIMEBOOST_net_570), .b(g53897_sb), .o(TIMEBOOST_net_14857) );
in01s01 FE_RC_578_0 ( .a(n_13354), .o(FE_RN_373_0) );
in01f02 FE_RC_579_0 ( .a(n_12982), .o(FE_RN_374_0) );
in01s01 TIMEBOOST_cell_45887 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_), .o(TIMEBOOST_net_15194) );
na03s02 TIMEBOOST_cell_33786 ( .a(FE_OFN254_n_9825), .b(g58197_sb), .c(g58197_db), .o(n_9589) );
in01s02 FE_RC_582_0 ( .a(n_13354), .o(FE_RN_376_0) );
in01f02 FE_RC_583_0 ( .a(n_12984), .o(FE_RN_377_0) );
in01s01 TIMEBOOST_cell_45888 ( .a(TIMEBOOST_net_15194), .o(TIMEBOOST_net_15195) );
na02s02 TIMEBOOST_cell_43649 ( .a(n_3614), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__Q), .o(TIMEBOOST_net_14063) );
na02s01 TIMEBOOST_cell_31063 ( .a(TIMEBOOST_net_9442), .b(g64995_db), .o(n_4356) );
na02s01 TIMEBOOST_cell_31062 ( .a(n_4488), .b(g64995_sb), .o(TIMEBOOST_net_9442) );
na02s01 TIMEBOOST_cell_40374 ( .a(TIMEBOOST_net_12425), .b(FE_OFN2079_n_8069), .o(TIMEBOOST_net_11076) );
in01f08 FE_RC_589_0 ( .a(FE_RN_381_0), .o(n_16791) );
na02f06 FE_RC_590_0 ( .a(n_15755), .b(n_16002), .o(FE_RN_381_0) );
in01f02 FE_RC_591_0 ( .a(n_16578), .o(FE_RN_382_0) );
no02f02 FE_RC_592_0 ( .a(FE_RN_382_0), .b(n_16573), .o(n_15453) );
na02s01 FE_RC_593_0 ( .a(parchk_pci_ad_out_in_1191), .b(FE_OFN1709_n_4868), .o(FE_RN_383_0) );
na02f02 FE_RC_594_0 ( .a(FE_RN_383_0), .b(n_14345), .o(n_14376) );
na02s02 TIMEBOOST_cell_17749 ( .a(TIMEBOOST_net_4131), .b(g61757_sb), .o(n_8299) );
na02s02 TIMEBOOST_cell_43456 ( .a(TIMEBOOST_net_13966), .b(FE_OFN1234_n_6391), .o(TIMEBOOST_net_12164) );
in01s01 TIMEBOOST_cell_45943 ( .a(wbm_dat_i_2_), .o(TIMEBOOST_net_15250) );
in01f08 FE_RC_599_0 ( .a(FE_RN_384_0), .o(n_15919) );
na02f08 FE_RC_600_0 ( .a(n_16015), .b(n_16016), .o(FE_RN_384_0) );
in01f03 FE_RC_601_0 ( .a(FE_RN_385_0), .o(n_8800) );
no02f04 FE_RC_602_0 ( .a(n_9175), .b(n_16331), .o(FE_RN_385_0) );
no02f20 FE_RC_604_0 ( .a(n_16275), .b(configuration_sync_cache_lsize_to_wb_bits_reg_3__Q), .o(FE_RN_387_0) );
na02f10 FE_RC_605_0 ( .a(FE_RN_387_0), .b(FE_RN_386_0), .o(n_16280) );
in01s08 FE_RC_606_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_), .o(FE_RN_388_0) );
na02f04 FE_RC_607_0 ( .a(n_16576), .b(FE_RN_388_0), .o(FE_RN_389_0) );
oa12f04 FE_RC_608_0 ( .a(FE_RN_389_0), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_), .c(n_16576), .o(n_16577) );
in01f02 FE_RC_60_0 ( .a(n_10202), .o(FE_RN_30_0) );
na02f06 FE_RC_610_0 ( .a(n_15014), .b(n_15055), .o(FE_RN_390_0) );
no02s02 FE_RC_612_0 ( .a(n_12179), .b(n_15762), .o(FE_RN_392_0) );
in01m02 FE_RC_613_0 ( .a(n_15760), .o(FE_RN_393_0) );
in01f02 FE_RC_614_0 ( .a(n_15759), .o(FE_RN_394_0) );
no02f06 FE_RC_615_0 ( .a(FE_RN_393_0), .b(FE_RN_394_0), .o(FE_RN_395_0) );
ao12f08 FE_RC_616_0 ( .a(FE_RN_392_0), .b(FE_RN_395_0), .c(n_15758), .o(FE_OFN1503_n_15768) );
in01m08 FE_RC_617_0 ( .a(n_13784), .o(FE_RN_396_0) );
na02f02 FE_RC_618_0 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_8__Q), .b(FE_OFN2126_n_16497), .o(FE_RN_397_0) );
in01s01 FE_RC_619_0 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_773), .o(FE_RN_398_0) );
in01f02 FE_RC_61_0 ( .a(n_10205), .o(FE_RN_31_0) );
oa12f02 FE_RC_620_0 ( .a(FE_RN_397_0), .b(FE_RN_398_0), .c(FE_OFN2126_n_16497), .o(FE_RN_399_0) );
na02f02 FE_RC_621_0 ( .a(n_12595), .b(FE_RN_399_0), .o(FE_RN_400_0) );
in01m01 FE_RC_622_0 ( .a(n_3295), .o(FE_RN_401_0) );
ao22m02 FE_RC_623_0 ( .a(configuration_pci_err_cs_bit8), .b(n_3252), .c(configuration_sync_command_bit8), .d(n_3248), .o(FE_RN_402_0) );
ao22f02 FE_RC_624_0 ( .a(configuration_wb_err_addr_540), .b(n_15444), .c(n_2844), .d(n_16000), .o(FE_RN_403_0) );
na02f02 TIMEBOOST_cell_44265 ( .a(n_9115), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__Q), .o(TIMEBOOST_net_14371) );
ao22f02 FE_RC_626_0 ( .a(configuration_pci_err_addr_478), .b(FE_OFN1006_n_16288), .c(wbu_latency_tim_val_in), .d(FE_OFN1694_n_3368), .o(FE_RN_405_0) );
in01s03 FE_RC_627_0 ( .a(configuration_wb_err_data_578), .o(FE_RN_406_0) );
in01f02 FE_RC_628_0 ( .a(FE_OFN1068_n_15729), .o(FE_RN_407_0) );
no02f02 FE_RC_62_0 ( .a(FE_RN_30_0), .b(FE_RN_31_0), .o(FE_RN_32_0) );
in01f02 FE_RC_630_0 ( .a(FE_OCPN1845_n_16427), .o(FE_RN_409_0) );
oa22f02 FE_RC_631_0 ( .a(FE_RN_406_0), .b(FE_RN_407_0), .c(FE_RN_678_0), .d(FE_RN_409_0), .o(FE_RN_410_0) );
na02f02 FE_RC_632_0 ( .a(FE_OCPN1901_n_16810), .b(n_14911), .o(FE_RN_411_0) );
na02s01 TIMEBOOST_cell_45083 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__Q), .b(FE_OFN528_n_9899), .o(TIMEBOOST_net_14780) );
na02f02 FE_RC_634_0 ( .a(n_16543), .b(configuration_wb_err_cs_bit8), .o(FE_RN_413_0) );
na02s01 TIMEBOOST_cell_37989 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__Q), .b(FE_OFN881_g64577_p), .o(TIMEBOOST_net_11233) );
no02f02 FE_RC_637_0 ( .a(FE_RN_415_0), .b(FE_RN_410_0), .o(FE_RN_416_0) );
na02f02 FE_RC_638_0 ( .a(FE_RN_416_0), .b(FE_RN_405_0), .o(FE_RN_417_0) );
no02f02 FE_RC_639_0 ( .a(FE_RN_417_0), .b(FE_RN_404_0), .o(FE_RN_418_0) );
na02s02 TIMEBOOST_cell_16839 ( .a(TIMEBOOST_net_3676), .b(g64872_db), .o(n_3711) );
oa12f02 FE_RC_640_0 ( .a(FE_RN_400_0), .b(n_12595), .c(FE_RN_418_0), .o(FE_RN_419_0) );
ao22s02 FE_RC_641_0 ( .a(conf_wb_err_addr_in_949), .b(n_2115), .c(wishbone_slave_unit_pcim_sm_data_in_642), .d(FE_OFN1610_n_2122), .o(FE_RN_420_0) );
na02f02 FE_RC_642_0 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__Q), .b(FE_OCPN1913_FE_OFN1150_n_13249), .o(FE_RN_421_0) );
in01s01 FE_RC_643_0 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_391), .o(FE_RN_422_0) );
oa12f02 FE_RC_644_0 ( .a(FE_RN_421_0), .b(FE_RN_422_0), .c(FE_OCPN1913_FE_OFN1150_n_13249), .o(FE_RN_423_0) );
na03s01 TIMEBOOST_cell_33540 ( .a(TIMEBOOST_net_271), .b(g61777_sb), .c(g61777_db), .o(n_8253) );
na03s01 TIMEBOOST_cell_33539 ( .a(TIMEBOOST_net_273), .b(g61783_sb), .c(g61783_db), .o(n_8239) );
ao22f02 FE_RC_647_0 ( .a(FE_RN_396_0), .b(FE_RN_419_0), .c(n_13784), .d(FE_RN_425_0), .o(FE_RN_426_0) );
in01f02 FE_RC_648_0 ( .a(FE_RN_427_0), .o(n_14323) );
no02f02 FE_RC_649_0 ( .a(FE_RN_426_0), .b(FE_OFN1708_n_4868), .o(FE_RN_427_0) );
in01f02 FE_RC_64_0 ( .a(n_10738), .o(FE_RN_33_0) );
na02f06 FE_RC_650_0 ( .a(n_16462), .b(n_15823), .o(FE_RN_428_0) );
no02f06 FE_RC_651_0 ( .a(FE_OCP_RBN2270_g75061_p), .b(n_16262), .o(FE_RN_429_0) );
na02f08 FE_RC_652_0 ( .a(FE_RN_429_0), .b(n_15824), .o(FE_RN_430_0) );
in01s01 FE_RC_654_0 ( .a(n_7822), .o(FE_RN_431_0) );
ao22f02 FE_RC_655_0 ( .a(configuration_pci_err_data_520), .b(FE_OFN1063_n_15808), .c(n_14922), .d(FE_OCPN1900_n_16810), .o(FE_RN_432_0) );
ao22f02 FE_RC_656_0 ( .a(configuration_wb_err_data_589), .b(FE_OFN1069_n_15729), .c(n_15598), .d(FE_OCPN1845_n_16427), .o(FE_RN_433_0) );
na02f02 FE_RC_657_0 ( .a(FE_RN_432_0), .b(FE_RN_433_0), .o(FE_RN_434_0) );
na02f02 FE_RC_658_0 ( .a(n_16791), .b(pciu_bar0_in_367), .o(FE_RN_435_0) );
na02f02 TIMEBOOST_cell_39127 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_10184), .o(TIMEBOOST_net_11802) );
in01f02 FE_RC_65_0 ( .a(n_10160), .o(FE_RN_34_0) );
ao22f02 FE_RC_660_0 ( .a(configuration_wb_err_addr_551), .b(n_15445), .c(configuration_pci_err_addr_489), .d(FE_OFN1006_n_16288), .o(FE_RN_437_0) );
ao22f02 FE_RC_661_0 ( .a(pciu_am1_in_528), .b(FE_OCPN1903_FE_OFN1061_n_16720), .c(pciu_bar0_in_367), .d(FE_OCPN1898_n_3231), .o(FE_RN_438_0) );
na02s01 TIMEBOOST_cell_41898 ( .a(TIMEBOOST_net_13187), .b(g62122_sb), .o(TIMEBOOST_net_11978) );
no02f02 FE_RC_663_0 ( .a(FE_RN_434_0), .b(FE_RN_439_0), .o(FE_RN_440_0) );
na02f02 FE_RC_664_0 ( .a(FE_RN_440_0), .b(n_4880), .o(FE_RN_441_0) );
na02f02 FE_RC_665_0 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_19__Q), .b(FE_OFN2126_n_16497), .o(FE_RN_442_0) );
in01s01 FE_RC_666_0 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_784), .o(FE_RN_443_0) );
oa12f02 FE_RC_667_0 ( .a(FE_RN_442_0), .b(FE_RN_443_0), .c(FE_OFN2126_n_16497), .o(FE_RN_444_0) );
ao22f02 FE_RC_668_0 ( .a(FE_RN_431_0), .b(FE_RN_441_0), .c(n_7822), .d(FE_RN_444_0), .o(FE_RN_445_0) );
no02f02 FE_RC_669_0 ( .a(FE_RN_445_0), .b(n_13784), .o(FE_RN_446_0) );
no02f02 FE_RC_66_0 ( .a(FE_RN_33_0), .b(FE_RN_34_0), .o(FE_RN_35_0) );
ao22s02 FE_RC_670_0 ( .a(conf_wb_err_addr_in_960), .b(FE_OFN1620_n_1787), .c(wishbone_slave_unit_pcim_sm_data_in_653), .d(FE_OFN1611_n_2122), .o(FE_RN_447_0) );
na02f02 FE_RC_671_0 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__Q), .b(FE_OCPN1911_FE_OFN1152_n_13249), .o(FE_RN_448_0) );
in01s01 FE_RC_672_0 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_402), .o(FE_RN_449_0) );
oa12f02 FE_RC_673_0 ( .a(FE_RN_448_0), .b(FE_RN_449_0), .c(FE_OCPN1911_FE_OFN1152_n_13249), .o(FE_RN_450_0) );
na02s02 TIMEBOOST_cell_43010 ( .a(TIMEBOOST_net_13743), .b(n_8590), .o(TIMEBOOST_net_12010) );
na02s01 TIMEBOOST_cell_9339 ( .a(TIMEBOOST_net_1236), .b(g64135_db), .o(n_4027) );
ao12f02 FE_RC_676_0 ( .a(FE_RN_446_0), .b(n_13781), .c(FE_RN_452_0), .o(FE_RN_453_0) );
in01f02 FE_RC_677_0 ( .a(FE_RN_454_0), .o(n_14351) );
no02f02 FE_RC_678_0 ( .a(FE_RN_453_0), .b(FE_OFN1706_n_4868), .o(FE_RN_454_0) );
na02f02 FE_RC_679_0 ( .a(n_13781), .b(n_13649), .o(FE_RN_455_0) );
na02s01 TIMEBOOST_cell_16836 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__Q), .b(g65342_sb), .o(TIMEBOOST_net_3675) );
in01f02 FE_RC_680_0 ( .a(n_13565), .o(FE_RN_456_0) );
in01f02 FE_RC_681_0 ( .a(FE_RN_457_0), .o(n_13760) );
na02f04 FE_RC_682_0 ( .a(FE_RN_456_0), .b(FE_RN_455_0), .o(FE_RN_457_0) );
in01f02 FE_RC_683_0 ( .a(FE_RN_458_0), .o(n_10595) );
na02f02 FE_RC_684_0 ( .a(n_8867), .b(n_15453), .o(FE_RN_458_0) );
na02f02 FE_RC_686_0 ( .a(n_8863), .b(n_16579), .o(FE_RN_459_0) );
no02f06 FE_RC_688_0 ( .a(n_15371), .b(n_4853), .o(FE_RN_460_0) );
na02f06 FE_RC_689_0 ( .a(FE_RN_460_0), .b(n_4815), .o(n_16435) );
in01f04 FE_RC_68_0 ( .a(n_16307), .o(FE_RN_36_0) );
in01f02 FE_RC_693_0 ( .a(n_10855), .o(FE_RN_463_0) );
in01f02 FE_RC_694_0 ( .a(n_11715), .o(FE_RN_464_0) );
no02f04 FE_RC_695_0 ( .a(FE_RN_463_0), .b(FE_RN_464_0), .o(FE_RN_465_0) );
in01f02 FE_RC_697_0 ( .a(n_10230), .o(FE_RN_466_0) );
in01f02 FE_RC_698_0 ( .a(n_10768), .o(FE_RN_467_0) );
no02f02 FE_RC_699_0 ( .a(FE_RN_466_0), .b(FE_RN_467_0), .o(FE_RN_468_0) );
in01f04 FE_RC_69_0 ( .a(n_16309), .o(FE_RN_37_0) );
na02f02 TIMEBOOST_cell_40922 ( .a(TIMEBOOST_net_12699), .b(g57066_sb), .o(n_11676) );
in01f02 FE_RC_701_0 ( .a(n_10679), .o(FE_RN_469_0) );
in01f02 FE_RC_702_0 ( .a(n_10681), .o(FE_RN_470_0) );
no02f02 FE_RC_703_0 ( .a(FE_RN_469_0), .b(FE_RN_470_0), .o(FE_RN_471_0) );
na02f02 TIMEBOOST_cell_45238 ( .a(TIMEBOOST_net_14857), .b(g54202_da), .o(TIMEBOOST_net_4813) );
in01f02 FE_RC_705_0 ( .a(n_10637), .o(FE_RN_472_0) );
in01f02 FE_RC_706_0 ( .a(n_10060), .o(FE_RN_473_0) );
no02f02 FE_RC_707_0 ( .a(FE_RN_472_0), .b(FE_RN_473_0), .o(FE_RN_474_0) );
in01f02 FE_RC_709_0 ( .a(n_10905), .o(FE_RN_475_0) );
na02s02 TIMEBOOST_cell_18422 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_18__Q), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_4468) );
in01f02 FE_RC_710_0 ( .a(n_11732), .o(FE_RN_476_0) );
no02f02 FE_RC_711_0 ( .a(FE_RN_475_0), .b(FE_RN_476_0), .o(FE_RN_477_0) );
na02s02 TIMEBOOST_cell_22277 ( .a(n_10190), .b(TIMEBOOST_net_6395), .o(n_11860) );
in01f02 FE_RC_713_0 ( .a(n_10981), .o(FE_RN_478_0) );
in01f02 FE_RC_714_0 ( .a(n_10758), .o(FE_RN_479_0) );
no02f02 FE_RC_715_0 ( .a(FE_RN_478_0), .b(FE_RN_479_0), .o(FE_RN_480_0) );
na02s02 TIMEBOOST_cell_39550 ( .a(TIMEBOOST_net_12013), .b(g58363_db), .o(n_9461) );
na02s01 TIMEBOOST_cell_36490 ( .a(TIMEBOOST_net_10483), .b(g66398_sb), .o(n_2542) );
in01m02 FE_RC_718_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_0_), .o(FE_RN_481_0) );
na02s02 TIMEBOOST_cell_37391 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_20__Q), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_403), .o(TIMEBOOST_net_10934) );
in01s06 FE_RC_720_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_), .o(FE_RN_483_0) );
oa22f04 FE_RC_721_0 ( .a(FE_OCP_RBN2225_n_16322), .b(FE_RN_481_0), .c(FE_RN_483_0), .d(n_16322), .o(n_16368) );
in01s01 FE_RC_722_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_4__213), .o(FE_RN_484_0) );
na02f02 FE_RC_724_0 ( .a(n_10680), .b(FE_RN_484_0), .o(FE_RN_486_0) );
na02f02 FE_RC_725_0 ( .a(n_9303), .b(FE_RN_486_0), .o(n_15590) );
na03f02 FE_RC_726_0 ( .a(n_16595), .b(n_14478), .c(n_16594), .o(n_14614) );
na03f02 FE_RC_728_0 ( .a(n_14257), .b(n_14551), .c(n_14258), .o(n_14596) );
na03f02 FE_RC_729_0 ( .a(n_14543), .b(n_14426), .c(n_14427), .o(n_14588) );
na03f02 FE_RC_731_0 ( .a(n_14272), .b(n_14558), .c(n_14271), .o(n_14603) );
na02s02 TIMEBOOST_cell_41941 ( .a(TIMEBOOST_net_1823), .b(FE_OFN1083_n_13221), .o(TIMEBOOST_net_13209) );
na03f02 FE_RC_733_0 ( .a(n_14564), .b(n_14290), .c(n_14471), .o(n_14609) );
na03f02 FE_RC_736_0 ( .a(n_14301), .b(n_14480), .c(n_14569), .o(n_14613) );
na02s01 TIMEBOOST_cell_41940 ( .a(TIMEBOOST_net_13208), .b(g65414_db), .o(TIMEBOOST_net_10658) );
na03f02 FE_RC_738_0 ( .a(n_14251), .b(n_14438), .c(n_14548), .o(n_14593) );
in01f06 FE_RC_73_0 ( .a(conf_w_addr_in_931), .o(FE_RN_39_0) );
no02f02 FE_RC_742_0 ( .a(g53222_p), .b(g53223_p), .o(FE_RN_489_0) );
na02f02 FE_RC_743_0 ( .a(FE_RN_489_0), .b(n_14554), .o(n_14599) );
in01f10 FE_RC_744_0 ( .a(wishbone_slave_unit_wishbone_slave_img_wallow), .o(FE_RN_490_0) );
na02f08 FE_RC_745_0 ( .a(n_15919), .b(FE_RN_490_0), .o(n_15908) );
in01m02 FE_RC_746_0 ( .a(n_16071), .o(FE_RN_491_0) );
in01s06 FE_RC_748_0 ( .a(n_16070), .o(FE_RN_493_0) );
in01f04 FE_RC_74_0 ( .a(parchk_pci_cbe_reg_in_1236), .o(FE_RN_40_0) );
na02f06 FE_RC_751_0 ( .a(FE_OCP_RBN2280_g74996_p), .b(n_16364), .o(FE_RN_494_0) );
na03f02 FE_RC_752_0 ( .a(n_13058), .b(FE_RN_203_0), .c(n_12695), .o(n_13139) );
na04f04 FE_RC_753_0 ( .a(n_12790), .b(n_13053), .c(n_12900), .d(n_12899), .o(n_13136) );
na02f02 TIMEBOOST_cell_40890 ( .a(TIMEBOOST_net_12683), .b(FE_OFN1403_n_8567), .o(TIMEBOOST_net_6161) );
na02s02 TIMEBOOST_cell_43152 ( .a(TIMEBOOST_net_13814), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_12138) );
na02s01 TIMEBOOST_cell_42669 ( .a(g64189_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__Q), .o(TIMEBOOST_net_13573) );
na04f04 FE_RC_759_0 ( .a(n_13045), .b(n_12780), .c(n_12869), .d(n_12870), .o(n_13129) );
no02f06 FE_RC_75_0 ( .a(FE_RN_40_0), .b(FE_RN_39_0), .o(FE_RN_41_0) );
na02s02 TIMEBOOST_cell_43650 ( .a(TIMEBOOST_net_14063), .b(FE_OFN1231_n_6391), .o(TIMEBOOST_net_12614) );
na02s02 TIMEBOOST_cell_44431 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_788), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_23__Q), .o(TIMEBOOST_net_14454) );
na02s02 TIMEBOOST_cell_43651 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__Q), .b(n_3604), .o(TIMEBOOST_net_14064) );
na02s01 TIMEBOOST_cell_42657 ( .a(TIMEBOOST_net_3407), .b(FE_OFN917_n_4725), .o(TIMEBOOST_net_13567) );
ao22f02 FE_RC_764_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__Q), .b(FE_OFN1734_n_16317), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__Q), .d(FE_OFN1739_n_11019), .o(FE_RN_496_0) );
na02s02 TIMEBOOST_cell_31999 ( .a(TIMEBOOST_net_9910), .b(FE_OFN1181_n_3476), .o(TIMEBOOST_net_4892) );
in01f02 FE_RC_766_0 ( .a(FE_RN_498_0), .o(n_12912) );
na02m02 TIMEBOOST_cell_41585 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_25__Q), .b(FE_OFN229_n_9120), .o(TIMEBOOST_net_13031) );
na03f08 FE_RC_76_0 ( .a(n_15959), .b(FE_RN_41_0), .c(conf_w_addr_in), .o(n_16046) );
in01f02 FE_RC_770_0 ( .a(n_8452), .o(FE_RN_500_0) );
na03s01 TIMEBOOST_cell_34006 ( .a(conf_wb_err_addr_in_956), .b(g62116_sb), .c(g62116_db), .o(n_5580) );
na02f02 FE_RC_772_0 ( .a(n_4699), .b(n_2963), .o(FE_RN_501_0) );
in01f02 FE_RC_773_0 ( .a(FE_RN_502_0), .o(n_7093) );
oa12f02 FE_RC_774_0 ( .a(FE_RN_501_0), .b(n_4699), .c(n_2963), .o(FE_RN_502_0) );
in01f02 FE_RC_775_0 ( .a(n_1397), .o(FE_RN_503_0) );
no02f04 FE_RC_777_0 ( .a(FE_RN_503_0), .b(FE_OCP_RBN2000_n_1403), .o(FE_RN_505_0) );
na03s02 TIMEBOOST_cell_39467 ( .a(TIMEBOOST_net_3958), .b(g64341_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__Q), .o(TIMEBOOST_net_11972) );
in01m10 FE_RC_779_0 ( .a(FE_RN_506_0), .o(n_1679) );
na02s02 TIMEBOOST_cell_43652 ( .a(TIMEBOOST_net_14064), .b(n_6645), .o(TIMEBOOST_net_12198) );
na02m20 FE_RC_780_0 ( .a(wbu_addr_in_252), .b(wbu_addr_in_251), .o(FE_RN_506_0) );
no02f20 FE_RC_781_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_0_), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_0_), .o(FE_RN_507_0) );
ao12f10 FE_RC_782_0 ( .a(FE_RN_507_0), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_0_), .c(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_0_), .o(FE_RN_508_0) );
no02f20 FE_RC_783_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_2_), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_2_), .o(FE_RN_509_0) );
ao12f10 FE_RC_784_0 ( .a(FE_RN_509_0), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_2_), .c(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_2_), .o(FE_RN_510_0) );
no02f20 FE_RC_785_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_1_), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_1_), .o(FE_RN_511_0) );
ao12f10 FE_RC_786_0 ( .a(FE_RN_511_0), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_1_), .c(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_1_), .o(FE_RN_512_0) );
no02f20 FE_RC_787_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_3_), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_3_), .o(FE_RN_513_0) );
ao12f10 FE_RC_788_0 ( .a(FE_RN_513_0), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_3_), .c(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_3_), .o(FE_RN_514_0) );
na02s01 TIMEBOOST_cell_45600 ( .a(TIMEBOOST_net_15038), .b(g65245_sb), .o(n_2637) );
in01f02 FE_RC_78_0 ( .a(n_551), .o(FE_RN_42_0) );
na02f08 FE_RC_790_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .o(FE_RN_515_0) );
oa12f06 FE_RC_791_0 ( .a(FE_RN_515_0), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .o(FE_RN_516_0) );
na02f08 FE_RC_792_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .o(FE_RN_517_0) );
oa12f04 FE_RC_793_0 ( .a(FE_RN_517_0), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .o(FE_RN_518_0) );
in01m10 FE_RC_794_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_), .o(FE_RN_519_0) );
in01m08 FE_RC_795_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .o(FE_RN_520_0) );
oa22f04 FE_RC_796_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .c(FE_RN_519_0), .d(FE_RN_520_0), .o(FE_RN_521_0) );
na02s02 TIMEBOOST_cell_45239 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__Q), .b(n_4499), .o(TIMEBOOST_net_14858) );
in01f08 FE_RC_798_0 ( .a(FE_RN_522_0), .o(n_2809) );
na02m20 FE_RC_799_0 ( .a(pciu_bar1_in_385), .b(pciu_am1_in_523), .o(FE_RN_522_0) );
in01f02 FE_RC_79_0 ( .a(n_16690), .o(FE_RN_43_0) );
na02m02 TIMEBOOST_cell_44341 ( .a(n_9791), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__Q), .o(TIMEBOOST_net_14409) );
in01f02 FE_RC_801_0 ( .a(n_2961), .o(FE_RN_523_0) );
in01f02 FE_RC_802_0 ( .a(n_2962), .o(FE_RN_524_0) );
ao22f04 FE_RC_803_0 ( .a(FE_RN_523_0), .b(FE_RN_524_0), .c(n_2961), .d(n_2962), .o(n_4702) );
in01m03 FE_RC_804_0 ( .a(FE_OCPN1852_n_16538), .o(FE_RN_525_0) );
in01f02 FE_RC_805_0 ( .a(FE_OCPN1843_n_16033), .o(FE_RN_526_0) );
na02f04 FE_RC_806_0 ( .a(FE_RN_525_0), .b(FE_RN_526_0), .o(n_16034) );
in01f04 FE_RC_807_0 ( .a(n_15744), .o(FE_RN_527_0) );
in01f03 FE_RC_808_0 ( .a(n_15748), .o(FE_RN_528_0) );
no02f06 FE_RC_809_0 ( .a(FE_OCPN1843_n_16033), .b(FE_OCPN1852_n_16538), .o(FE_RN_529_0) );
no02f04 FE_RC_80_0 ( .a(FE_RN_43_0), .b(FE_RN_42_0), .o(FE_RN_44_0) );
na02s02 TIMEBOOST_cell_45594 ( .a(TIMEBOOST_net_15035), .b(g65244_sb), .o(n_2638) );
na02s01 TIMEBOOST_cell_39552 ( .a(TIMEBOOST_net_12014), .b(g58295_db), .o(n_9510) );
na02s01 FE_RC_812_0 ( .a(n_565), .b(parchk_pci_trdy_en_in), .o(n_1088) );
na02f20 FE_RC_813_0 ( .a(parchk_pci_trdy_en_in), .b(n_565), .o(FE_RN_530_0) );
no02f08 FE_RC_814_0 ( .a(FE_OCP_RBN1930_parchk_pci_trdy_reg_in), .b(FE_RN_530_0), .o(n_1616) );
in01f02 FE_RC_815_0 ( .a(FE_RN_71_0), .o(FE_RN_531_0) );
in01f02 FE_RC_816_0 ( .a(n_1616), .o(FE_RN_532_0) );
no02f04 FE_RC_817_0 ( .a(FE_RN_531_0), .b(FE_RN_532_0), .o(FE_RN_533_0) );
na02f04 TIMEBOOST_cell_44774 ( .a(TIMEBOOST_net_14625), .b(n_3123), .o(TIMEBOOST_net_1530) );
na02s02 TIMEBOOST_cell_43530 ( .a(TIMEBOOST_net_14003), .b(FE_OFN1234_n_6391), .o(TIMEBOOST_net_12187) );
na02f08 FE_RC_81_0 ( .a(n_1072), .b(FE_RN_44_0), .o(n_2552) );
na02f10 FE_RC_820_0 ( .a(n_16284), .b(n_16285), .o(n_16289) );
na02f06 FE_RC_821_0 ( .a(n_16284), .b(n_16285), .o(FE_OCPN1868_n_16289) );
na02f02 FE_RC_822_0 ( .a(FE_RN_535_0), .b(n_16474), .o(n_16475) );
na02f04 FE_RC_823_0 ( .a(FE_OCP_RBN1954_FE_RN_462_0), .b(n_16513), .o(FE_RN_535_0) );
na02s01 TIMEBOOST_cell_17864 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__Q), .b(g65321_sb), .o(TIMEBOOST_net_4189) );
na02s02 TIMEBOOST_cell_17865 ( .a(TIMEBOOST_net_4189), .b(g65321_db), .o(n_3561) );
in01m01 FE_RC_828_0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_), .o(FE_RN_538_0) );
in01f02 FE_RC_829_0 ( .a(n_15512), .o(FE_RN_539_0) );
in01f06 FE_RC_82_0 ( .a(n_8728), .o(FE_RN_45_0) );
na02s02 TIMEBOOST_cell_43637 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__Q), .b(n_3714), .o(TIMEBOOST_net_14057) );
na02s01 TIMEBOOST_cell_36286 ( .a(TIMEBOOST_net_10381), .b(g67057_sb), .o(n_1677) );
na02s03 TIMEBOOST_cell_45769 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__Q), .b(n_13172), .o(TIMEBOOST_net_15123) );
in01s01 FE_RC_833_0 ( .a(n_7822), .o(FE_RN_541_0) );
in01f02 FE_RC_834_0 ( .a(n_12983), .o(FE_RN_542_0) );
na02s01 TIMEBOOST_cell_44790 ( .a(TIMEBOOST_net_14633), .b(g57911_sb), .o(TIMEBOOST_net_12448) );
na02f02 TIMEBOOST_cell_42392 ( .a(TIMEBOOST_net_13434), .b(g57442_sb), .o(n_11293) );
in01s02 FE_RC_837_0 ( .a(n_13354), .o(FE_RN_544_0) );
in01f02 FE_RC_838_0 ( .a(n_12988), .o(FE_RN_545_0) );
in01s01 TIMEBOOST_cell_45889 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_), .o(TIMEBOOST_net_15196) );
in01f02 FE_RC_83_0 ( .a(n_3334), .o(FE_RN_46_0) );
na02s01 TIMEBOOST_cell_42032 ( .a(TIMEBOOST_net_13254), .b(g62580_sb), .o(n_6393) );
in01s01 FE_RC_841_0 ( .a(n_3404), .o(FE_RN_547_0) );
in01m01 FE_RC_842_0 ( .a(n_16000), .o(FE_RN_548_0) );
no02m02 FE_RC_843_0 ( .a(FE_RN_548_0), .b(FE_RN_547_0), .o(FE_RN_549_0) );
no02f02 FE_RC_844_0 ( .a(n_5724), .b(FE_RN_549_0), .o(n_7308) );
na02s02 TIMEBOOST_cell_41742 ( .a(TIMEBOOST_net_13109), .b(g58264_db), .o(n_9535) );
in01f20 FE_RC_846_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_), .o(FE_RN_551_0) );
na02m02 TIMEBOOST_cell_42118 ( .a(TIMEBOOST_net_13297), .b(FE_OFN1323_n_6436), .o(TIMEBOOST_net_11587) );
na02s01 TIMEBOOST_cell_41743 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__Q), .b(g65426_sb), .o(TIMEBOOST_net_13110) );
in01f10 FE_RC_849_0 ( .a(configuration_sync_cache_lsize_to_wb_bits_reg_2__Q), .o(FE_RN_553_0) );
no02f04 FE_RC_84_0 ( .a(FE_RN_45_0), .b(FE_RN_46_0), .o(FE_RN_47_0) );
no02f10 FE_RC_850_0 ( .a(FE_RN_553_0), .b(n_3319), .o(n_3320) );
in01f10 FE_RC_851_0 ( .a(n_681), .o(FE_RN_554_0) );
no02f20 FE_RC_852_0 ( .a(n_1200), .b(FE_RN_554_0), .o(n_16474) );
in01f08 FE_RC_854_0 ( .a(FE_RN_555_0), .o(FE_OFN993_n_15366) );
na02f10 FE_RC_855_0 ( .a(n_15365), .b(pci_target_unit_pci_target_sm_previous_frame), .o(FE_RN_555_0) );
in01f06 FE_RC_856_0 ( .a(FE_RN_556_0), .o(n_16351) );
no02f10 FE_RC_857_0 ( .a(n_16350), .b(parchk_pci_cbe_reg_in_1236), .o(FE_RN_556_0) );
in01f08 FE_RC_858_0 ( .a(FE_RN_557_0), .o(n_16307) );
na02f10 FE_RC_859_0 ( .a(n_16390), .b(n_16027), .o(FE_RN_557_0) );
in01f08 FE_RC_860_0 ( .a(n_15958), .o(FE_RN_558_0) );
na02f08 FE_RC_861_0 ( .a(FE_RN_558_0), .b(n_15959), .o(n_16388) );
no04f40 FE_RC_862_0 ( .a(pciu_cache_line_size_in_776), .b(configuration_sync_cache_lsize_to_wb_bits_reg_4__Q), .c(pciu_cache_line_size_in_777), .d(pciu_cache_line_size_in_775), .o(FE_RN_386_0) );
in01s01 FE_RC_863_0 ( .a(n_12595), .o(FE_RN_559_0) );
in01s01 FE_RC_864_0 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_789), .o(FE_RN_560_0) );
no02f02 FE_RC_865_0 ( .a(FE_RN_560_0), .b(FE_OCPN1909_n_16497), .o(FE_RN_561_0) );
ao12f02 FE_RC_866_0 ( .a(FE_RN_561_0), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_24__Q), .c(FE_OCPN1909_n_16497), .o(FE_RN_562_0) );
na02s02 TIMEBOOST_cell_36737 ( .a(n_2795), .b(n_2995), .o(TIMEBOOST_net_10607) );
ao22f01 FE_RC_868_0 ( .a(configuration_pci_err_data_525), .b(FE_OFN1066_n_15808), .c(configuration_wb_err_cs_bit31_24), .d(n_16543), .o(FE_RN_564_0) );
na02f02 FE_RC_869_0 ( .a(FE_RN_564_0), .b(n_2768), .o(FE_RN_565_0) );
ao22f01 FE_RC_870_0 ( .a(configuration_status_bit8), .b(n_3248), .c(n_2815), .d(n_16000), .o(FE_RN_566_0) );
ao22f01 FE_RC_871_0 ( .a(configuration_pci_err_addr_494), .b(FE_OFN1005_n_16288), .c(configuration_pci_err_cs_bit31_24), .d(n_3252), .o(FE_RN_567_0) );
na02f01 FE_RC_872_0 ( .a(n_15444), .b(configuration_wb_err_addr_556), .o(FE_RN_568_0) );
na03s01 TIMEBOOST_cell_34286 ( .a(n_3908), .b(g63052_sb), .c(g63052_db), .o(n_5146) );
ao22f01 FE_RC_874_0 ( .a(n_14927), .b(n_16810), .c(pciu_am1_in_533), .d(FE_OFN2129_n_16720), .o(FE_RN_570_0) );
ao22f01 FE_RC_875_0 ( .a(configuration_wb_err_data_594), .b(FE_OFN1070_n_15729), .c(n_2815), .d(FE_OCPN1845_n_16427), .o(FE_RN_571_0) );
na02f01 FE_RC_876_0 ( .a(n_3290), .b(pciu_bar0_in_372), .o(FE_RN_572_0) );
na02s02 TIMEBOOST_cell_41817 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__Q), .b(g58371_sb), .o(TIMEBOOST_net_13147) );
na02f02 TIMEBOOST_cell_44741 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__Q), .b(FE_OFN1584_n_12306), .o(TIMEBOOST_net_14609) );
na02f02 TIMEBOOST_cell_40924 ( .a(TIMEBOOST_net_12700), .b(g57102_sb), .o(n_11644) );
in01f02 TIMEBOOST_cell_15782 ( .a(TIMEBOOST_net_3147), .o(n_7608) );
in01m04 FE_RC_882_0 ( .a(FE_OFN969_n_13784), .o(FE_RN_578_0) );
na02s01 TIMEBOOST_cell_42733 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__Q), .b(n_2059), .o(TIMEBOOST_net_13605) );
na02m02 TIMEBOOST_cell_40481 ( .a(g54186_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_405), .o(TIMEBOOST_net_12479) );
na02s01 TIMEBOOST_cell_40434 ( .a(TIMEBOOST_net_12455), .b(n_3914), .o(n_5163) );
in01s02 FE_RC_886_0 ( .a(n_504), .o(FE_RN_582_0) );
in01m02 FE_RC_887_0 ( .a(FE_OFN1151_n_13249), .o(FE_RN_583_0) );
ao22f02 FE_RC_888_0 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__Q), .b(FE_OCPN1911_FE_OFN1152_n_13249), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_407), .d(FE_RN_583_0), .o(FE_RN_584_0) );
na02f02 TIMEBOOST_cell_22383 ( .a(n_8896), .b(TIMEBOOST_net_6448), .o(n_9931) );
in01f04 FE_RC_88_0 ( .a(n_13754), .o(FE_RN_48_0) );
na02s01 TIMEBOOST_cell_43653 ( .a(n_4518), .b(g61877_sb), .o(TIMEBOOST_net_14065) );
na02s01 TIMEBOOST_cell_37990 ( .a(TIMEBOOST_net_11233), .b(TIMEBOOST_net_9746), .o(n_5448) );
no02m02 TIMEBOOST_cell_36366 ( .a(TIMEBOOST_net_1154), .b(TIMEBOOST_net_10421), .o(g63943_p) );
in01f02 FE_RC_893_0 ( .a(FE_RN_589_0), .o(n_14345) );
na02f02 TIMEBOOST_cell_22587 ( .a(TIMEBOOST_net_6550), .b(n_14072), .o(n_14532) );
in01f02 FE_RC_895_0 ( .a(n_2440), .o(FE_RN_590_0) );
in01f06 FE_RC_896_0 ( .a(FE_OFN2093_n_2301), .o(FE_RN_591_0) );
no02f06 FE_RC_897_0 ( .a(FE_RN_590_0), .b(FE_RN_591_0), .o(FE_RN_592_0) );
no02m02 FE_RC_898_0 ( .a(n_8511), .b(n_16326), .o(FE_RN_593_0) );
in01f04 FE_RC_899_0 ( .a(n_2833), .o(FE_RN_594_0) );
in01f02 FE_RC_89_0 ( .a(n_13654), .o(FE_RN_49_0) );
in01f02 FE_RC_900_0 ( .a(n_307), .o(FE_RN_595_0) );
oa22f02 FE_RC_901_0 ( .a(n_2833), .b(n_307), .c(FE_RN_594_0), .d(FE_RN_595_0), .o(FE_RN_596_0) );
in01f02 FE_RC_902_0 ( .a(n_2841), .o(FE_RN_597_0) );
in01f02 FE_RC_903_0 ( .a(n_385), .o(FE_RN_598_0) );
na02s01 TIMEBOOST_cell_31061 ( .a(TIMEBOOST_net_9441), .b(g64989_db), .o(n_4359) );
na02f04 FE_RC_905_0 ( .a(n_2841), .b(n_385), .o(FE_RN_600_0) );
na02s02 TIMEBOOST_cell_31060 ( .a(n_4498), .b(g64989_sb), .o(TIMEBOOST_net_9441) );
no02f02 FE_RC_907_0 ( .a(FE_RN_596_0), .b(FE_RN_601_0), .o(FE_RN_602_0) );
na02s10 FE_RC_908_0 ( .a(pciu_am1_in_540), .b(conf_pci_init_complete_out), .o(FE_RN_603_0) );
in01s10 FE_RC_909_0 ( .a(configuration_sync_command_bit0), .o(FE_RN_604_0) );
na02s01 TIMEBOOST_cell_44873 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__Q), .b(g64276_sb), .o(TIMEBOOST_net_14675) );
in01f02 FE_RC_910_0 ( .a(n_2380), .o(FE_RN_605_0) );
na02s01 TIMEBOOST_cell_41744 ( .a(TIMEBOOST_net_13110), .b(g65426_db), .o(n_3509) );
in01f04 FE_RC_912_0 ( .a(n_2815), .o(FE_RN_607_0) );
in01f02 FE_RC_913_0 ( .a(n_227), .o(FE_RN_608_0) );
ao22f02 FE_RC_914_0 ( .a(FE_RN_607_0), .b(FE_RN_608_0), .c(n_2815), .d(n_227), .o(FE_RN_609_0) );
na02f04 FE_RC_915_0 ( .a(n_2851), .b(n_233), .o(FE_RN_610_0) );
oa12f02 FE_RC_916_0 ( .a(FE_RN_610_0), .b(n_2851), .c(n_233), .o(FE_RN_611_0) );
na02f04 FE_RC_917_0 ( .a(n_2854), .b(n_277), .o(FE_RN_612_0) );
oa12f02 FE_RC_918_0 ( .a(FE_RN_612_0), .b(n_2854), .c(n_277), .o(FE_RN_613_0) );
na02f04 FE_RC_919_0 ( .a(n_2825), .b(n_302), .o(FE_RN_614_0) );
na02s01 TIMEBOOST_cell_31998 ( .a(configuration_pci_err_addr_498), .b(wbm_adr_o_28_), .o(TIMEBOOST_net_9910) );
oa12f02 FE_RC_920_0 ( .a(FE_RN_614_0), .b(n_2825), .c(n_302), .o(FE_RN_615_0) );
in01f04 FE_RC_921_0 ( .a(n_3592), .o(FE_RN_616_0) );
in01f02 FE_RC_922_0 ( .a(n_372), .o(FE_RN_617_0) );
oa22f02 FE_RC_923_0 ( .a(n_3592), .b(n_372), .c(FE_RN_616_0), .d(FE_RN_617_0), .o(FE_RN_618_0) );
na02m02 TIMEBOOST_cell_32556 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__Q), .o(TIMEBOOST_net_10189) );
na02f04 FE_RC_925_0 ( .a(n_2856), .b(n_336), .o(FE_RN_620_0) );
oa12f02 FE_RC_926_0 ( .a(FE_RN_620_0), .b(n_2856), .c(n_336), .o(FE_RN_621_0) );
in01f02 FE_RC_927_0 ( .a(n_3404), .o(FE_RN_622_0) );
in01f02 FE_RC_928_0 ( .a(n_290), .o(FE_RN_623_0) );
na02s01 TIMEBOOST_cell_31059 ( .a(TIMEBOOST_net_9440), .b(g64987_db), .o(n_4361) );
na02m02 TIMEBOOST_cell_44249 ( .a(n_9666), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__Q), .o(TIMEBOOST_net_14363) );
in01s01 TIMEBOOST_cell_45944 ( .a(TIMEBOOST_net_15250), .o(TIMEBOOST_net_15251) );
na02s01 TIMEBOOST_cell_31058 ( .a(n_4498), .b(g64987_sb), .o(TIMEBOOST_net_9440) );
in01f02 FE_RC_932_0 ( .a(n_2869), .o(FE_RN_627_0) );
in01f02 FE_RC_933_0 ( .a(n_287), .o(FE_RN_628_0) );
na02s02 TIMEBOOST_cell_22303 ( .a(n_10275), .b(TIMEBOOST_net_6408), .o(n_11872) );
in01s01 TIMEBOOST_cell_32828 ( .a(TIMEBOOST_net_10329), .o(wbs_dat_i_22_) );
na02f02 TIMEBOOST_cell_43818 ( .a(TIMEBOOST_net_14147), .b(FE_OFN1409_n_8567), .o(TIMEBOOST_net_12888) );
in01f02 FE_RC_937_0 ( .a(n_15598), .o(FE_RN_632_0) );
in01f02 FE_RC_938_0 ( .a(n_360), .o(FE_RN_633_0) );
na02s02 TIMEBOOST_cell_41707 ( .a(g58779_sb), .b(wbu_addr_in_269), .o(TIMEBOOST_net_13092) );
in01m02 FE_RC_93_0 ( .a(n_3365), .o(FE_RN_51_0) );
na02s01 TIMEBOOST_cell_44893 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__Q), .b(FE_OFN1793_n_9904), .o(TIMEBOOST_net_14685) );
na02s02 TIMEBOOST_cell_32013 ( .a(TIMEBOOST_net_9917), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4899) );
in01f02 FE_RC_942_0 ( .a(n_2866), .o(FE_RN_637_0) );
in01f02 FE_RC_943_0 ( .a(n_300), .o(FE_RN_638_0) );
na02f02 TIMEBOOST_cell_41660 ( .a(TIMEBOOST_net_13068), .b(n_14971), .o(TIMEBOOST_net_11704) );
in01s01 TIMEBOOST_cell_32827 ( .a(TIMEBOOST_net_10328), .o(TIMEBOOST_net_10327) );
na02s01 TIMEBOOST_cell_30898 ( .a(pci_target_unit_pcit_if_strd_addr_in_687), .b(n_2515), .o(TIMEBOOST_net_9360) );
in01f02 FE_RC_947_0 ( .a(n_2809), .o(FE_RN_642_0) );
in01f02 FE_RC_948_0 ( .a(n_413), .o(FE_RN_643_0) );
na02f04 FE_RC_949_0 ( .a(FE_RN_642_0), .b(FE_RN_643_0), .o(FE_RN_644_0) );
in01m02 FE_RC_94_0 ( .a(n_3046), .o(FE_RN_52_0) );
in01f02 FE_RC_950_0 ( .a(n_2809), .o(FE_RN_645_0) );
in01f02 FE_RC_951_0 ( .a(n_413), .o(FE_RN_646_0) );
oa12f02 FE_RC_952_0 ( .a(FE_RN_644_0), .b(FE_RN_645_0), .c(FE_RN_646_0), .o(FE_RN_647_0) );
in01f04 FE_RC_953_0 ( .a(n_2831), .o(FE_RN_648_0) );
in01m06 FE_RC_954_0 ( .a(n_303), .o(FE_RN_649_0) );
na02f04 FE_RC_955_0 ( .a(FE_RN_648_0), .b(FE_RN_649_0), .o(FE_RN_650_0) );
in01f02 FE_RC_956_0 ( .a(n_2831), .o(FE_RN_651_0) );
oa12f02 FE_RC_958_0 ( .a(FE_RN_650_0), .b(FE_RN_651_0), .c(FE_RN_649_0), .o(FE_RN_653_0) );
in01f02 FE_RC_959_0 ( .a(n_2812), .o(FE_RN_654_0) );
no02f02 FE_RC_95_0 ( .a(FE_RN_51_0), .b(FE_RN_52_0), .o(FE_RN_53_0) );
in01f04 FE_RC_960_0 ( .a(n_389), .o(FE_RN_655_0) );
na02f04 FE_RC_961_0 ( .a(FE_RN_654_0), .b(FE_RN_655_0), .o(FE_RN_656_0) );
in01f02 FE_RC_962_0 ( .a(n_2812), .o(FE_RN_657_0) );
oa12f02 FE_RC_964_0 ( .a(FE_RN_656_0), .b(FE_RN_657_0), .c(FE_RN_655_0), .o(FE_RN_659_0) );
in01f02 FE_RC_965_0 ( .a(n_16428), .o(FE_RN_660_0) );
in01f04 FE_RC_966_0 ( .a(n_297), .o(FE_RN_661_0) );
na02f04 FE_RC_967_0 ( .a(FE_RN_660_0), .b(FE_RN_661_0), .o(FE_RN_662_0) );
in01f02 FE_RC_968_0 ( .a(n_16428), .o(FE_RN_663_0) );
na02f02 FE_RC_96_0 ( .a(n_7697), .b(FE_RN_53_0), .o(n_8488) );
oa12f02 FE_RC_970_0 ( .a(FE_RN_662_0), .b(FE_RN_663_0), .c(FE_RN_661_0), .o(FE_RN_665_0) );
na02s02 TIMEBOOST_cell_45601 ( .a(TIMEBOOST_net_9345), .b(FE_OFN787_n_2678), .o(TIMEBOOST_net_15039) );
in01f02 FE_RC_972_0 ( .a(n_231), .o(FE_RN_667_0) );
in01f02 FE_RC_973_0 ( .a(n_2818), .o(FE_RN_668_0) );
no02f02 FE_RC_974_0 ( .a(FE_RN_667_0), .b(FE_RN_668_0), .o(FE_RN_669_0) );
no02f04 FE_RC_975_0 ( .a(n_2822), .b(n_439), .o(FE_RN_670_0) );
no02f04 FE_RC_976_0 ( .a(n_2818), .b(n_231), .o(FE_RN_671_0) );
in01f02 FE_RC_977_0 ( .a(n_439), .o(FE_RN_672_0) );
in01f02 FE_RC_978_0 ( .a(n_2822), .o(FE_RN_673_0) );
no02f02 FE_RC_979_0 ( .a(FE_RN_672_0), .b(FE_RN_673_0), .o(FE_RN_674_0) );
in01s01 TIMEBOOST_cell_45940 ( .a(TIMEBOOST_net_15246), .o(TIMEBOOST_net_15247) );
na02f02 TIMEBOOST_cell_22075 ( .a(n_14024), .b(TIMEBOOST_net_6294), .o(n_14416) );
in01f02 FE_RC_982_0 ( .a(n_376), .o(FE_RN_677_0) );
in01f04 FE_RC_983_0 ( .a(n_2844), .o(FE_RN_678_0) );
na02f02 TIMEBOOST_cell_44128 ( .a(TIMEBOOST_net_14302), .b(FE_OFN1407_n_8567), .o(TIMEBOOST_net_13386) );
in01f02 FE_RC_985_0 ( .a(n_298), .o(FE_RN_680_0) );
in01f02 FE_RC_986_0 ( .a(n_2838), .o(FE_RN_681_0) );
oa22f02 FE_RC_987_0 ( .a(n_298), .b(n_2838), .c(FE_RN_680_0), .d(FE_RN_681_0), .o(FE_RN_682_0) );
na02s01 TIMEBOOST_cell_43654 ( .a(TIMEBOOST_net_14065), .b(g61877_db), .o(n_8076) );
na02f02 FE_RC_989_0 ( .a(FE_RN_675_0), .b(FE_RN_683_0), .o(FE_RN_684_0) );
in01f08 FE_RC_98_0 ( .a(n_15798), .o(FE_RN_55_0) );
in01f02 FE_RC_990_0 ( .a(n_2864), .o(FE_RN_685_0) );
in01f02 FE_RC_991_0 ( .a(n_436), .o(FE_RN_686_0) );
na02f04 FE_RC_993_0 ( .a(n_2828), .b(n_204), .o(FE_RN_688_0) );
oa12f02 FE_RC_994_0 ( .a(FE_RN_688_0), .b(n_2828), .c(n_204), .o(FE_RN_689_0) );
na02s01 TIMEBOOST_cell_41915 ( .a(TIMEBOOST_net_4251), .b(g64084_db), .o(TIMEBOOST_net_13196) );
na02s01 TIMEBOOST_cell_41916 ( .a(TIMEBOOST_net_13196), .b(TIMEBOOST_net_4398), .o(n_5521) );
in01f06 FE_RC_998_0 ( .a(n_357), .o(FE_RN_693_0) );
na02f04 FE_RC_999_0 ( .a(FE_RN_695_0), .b(FE_RN_693_0), .o(FE_RN_694_0) );
no02f08 FE_RC_99_0 ( .a(FE_RN_55_0), .b(parchk_pci_trdy_reg_in), .o(FE_RN_56_0) );
ms00f80 configuration_cache_line_size_reg_reg_0__u0 ( .ck(ispd_clk), .d(n_7598), .o(configuration_cache_line_size_reg) );
ms00f80 configuration_cache_line_size_reg_reg_1__u0 ( .ck(ispd_clk), .d(n_7596), .o(configuration_cache_line_size_reg_2996) );
ms00f80 configuration_cache_line_size_reg_reg_2__u0 ( .ck(ispd_clk), .d(n_7595), .o(wbu_cache_line_size_in_206) );
ms00f80 configuration_cache_line_size_reg_reg_3__u0 ( .ck(ispd_clk), .d(n_8437), .o(wbu_cache_line_size_in_207) );
ms00f80 configuration_cache_line_size_reg_reg_4__u0 ( .ck(ispd_clk), .d(n_8436), .o(wbu_cache_line_size_in_208) );
ms00f80 configuration_cache_line_size_reg_reg_5__u0 ( .ck(ispd_clk), .d(n_8434), .o(wbu_cache_line_size_in_209) );
ms00f80 configuration_cache_line_size_reg_reg_6__u0 ( .ck(ispd_clk), .d(n_7590), .o(wbu_cache_line_size_in_210) );
ms00f80 configuration_cache_line_size_reg_reg_7__u0 ( .ck(ispd_clk), .d(n_8433), .o(wbu_cache_line_size_in_211) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wbu_cache_line_size_in_206), .o(configuration_meta_cache_lsize_to_wb_bits) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(wbu_cache_line_size_in_207), .o(configuration_meta_cache_lsize_to_wb_bits_926) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(wbu_cache_line_size_in_208), .o(configuration_meta_cache_lsize_to_wb_bits_927) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_3__u0 ( .ck(ispd_clk), .d(wbu_cache_line_size_in_209), .o(configuration_meta_cache_lsize_to_wb_bits_928) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_4__u0 ( .ck(ispd_clk), .d(wbu_cache_line_size_in_210), .o(configuration_meta_cache_lsize_to_wb_bits_929) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_5__u0 ( .ck(ispd_clk), .d(wbu_cache_line_size_in_211), .o(configuration_meta_cache_lsize_to_wb_bits_930) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_6__u0 ( .ck(ispd_clk), .d(n_1625), .o(configuration_meta_cache_lsize_to_wb_bits_931) );
ms00f80 configuration_command_bit2_0_reg_0__u0 ( .ck(ispd_clk), .d(n_8456), .o(configuration_sync_command_bit0) );
ms00f80 configuration_command_bit2_0_reg_1__u0 ( .ck(ispd_clk), .d(n_8455), .o(configuration_sync_command_bit1) );
ms00f80 configuration_command_bit2_0_reg_2__u0 ( .ck(ispd_clk), .d(n_8454), .o(configuration_command_bit) );
ms00f80 configuration_command_bit6_reg_u0 ( .ck(ispd_clk), .d(n_8453), .o(configuration_sync_command_bit6) );
ms00f80 configuration_command_bit8_reg_u0 ( .ck(ispd_clk), .d(n_8464), .o(configuration_sync_command_bit8) );
ms00f80 configuration_command_bit_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(configuration_command_bit), .o(configuration_meta_command_bit) );
ms00f80 configuration_i_wb_init_complete_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(FE_OFN992_n_2373), .o(configuration_sync_init_complete) );
ms00f80 configuration_icr_bit2_0_reg_0__u0 ( .ck(ispd_clk), .d(n_7820), .o(configuration_icr_bit2_0) );
ms00f80 configuration_icr_bit2_0_reg_1__u0 ( .ck(ispd_clk), .d(n_7819), .o(configuration_icr_bit_2961) );
ms00f80 configuration_icr_bit2_0_reg_2__u0 ( .ck(ispd_clk), .d(n_7817), .o(configuration_icr_bit_2967) );
ms00f80 configuration_icr_bit31_reg_u0 ( .ck(ispd_clk), .d(n_7627), .o(pci_resi_conf_soft_res_in) );
ms00f80 configuration_init_complete_reg_u0 ( .ck(ispd_clk), .d(n_1385), .o(conf_pci_init_complete_out) );
ms00f80 configuration_int_pin_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_1545), .o(configuration_int_meta) );
ms00f80 configuration_interrupt_line_reg_0__u0 ( .ck(ispd_clk), .d(n_8463), .o(configuration_interrupt_line) );
ms00f80 configuration_interrupt_line_reg_1__u0 ( .ck(ispd_clk), .d(n_8462), .o(configuration_interrupt_line_37) );
ms00f80 configuration_interrupt_line_reg_2__u0 ( .ck(ispd_clk), .d(n_8461), .o(configuration_interrupt_line_38) );
ms00f80 configuration_interrupt_line_reg_3__u0 ( .ck(ispd_clk), .d(n_8442), .o(configuration_interrupt_line_39) );
ms00f80 configuration_interrupt_line_reg_4__u0 ( .ck(ispd_clk), .d(n_8441), .o(configuration_interrupt_line_40) );
ms00f80 configuration_interrupt_line_reg_5__u0 ( .ck(ispd_clk), .d(n_8439), .o(configuration_interrupt_line_41) );
ms00f80 configuration_interrupt_line_reg_6__u0 ( .ck(ispd_clk), .d(n_8457), .o(configuration_interrupt_line_42) );
ms00f80 configuration_interrupt_line_reg_7__u0 ( .ck(ispd_clk), .d(n_8438), .o(configuration_interrupt_line_43) );
ms00f80 configuration_interrupt_out_reg_u0 ( .ck(ispd_clk), .d(configuration_int_meta), .o(configuration_interrupt_out_reg_Q) );
in01s01 configuration_interrupt_out_reg_u1 ( .a(configuration_interrupt_out_reg_Q), .o(pci_inti_conf_int_in) );
ms00f80 configuration_isr_bit0_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_536), .o(configuration_isr_bit_1461) );
ms00f80 configuration_isr_bit2_0_reg_0__u0 ( .ck(ispd_clk), .d(configuration_isr_bit_1461), .o(configuration_isr_bit_631) );
ms00f80 configuration_isr_bit2_0_reg_1__u0 ( .ck(ispd_clk), .d(n_8508), .o(configuration_isr_bit_2975) );
ms00f80 configuration_isr_bit2_0_reg_2__u0 ( .ck(ispd_clk), .d(configuration_isr_bit_1457), .o(configuration_isr_bit_618) );
ms00f80 configuration_isr_bit2_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_1084), .o(configuration_isr_bit_1457) );
ms00f80 configuration_latency_timer_reg_0__u0 ( .ck(ispd_clk), .d(n_7607), .o(wbu_latency_tim_val_in) );
ms00f80 configuration_latency_timer_reg_1__u0 ( .ck(ispd_clk), .d(n_7606), .o(wbu_latency_tim_val_in_243) );
ms00f80 configuration_latency_timer_reg_2__u0 ( .ck(ispd_clk), .d(n_7605), .o(wbu_latency_tim_val_in_244) );
ms00f80 configuration_latency_timer_reg_3__u0 ( .ck(ispd_clk), .d(n_7604), .o(wbu_latency_tim_val_in_245) );
ms00f80 configuration_latency_timer_reg_4__u0 ( .ck(ispd_clk), .d(n_7602), .o(wbu_latency_tim_val_in_246) );
ms00f80 configuration_latency_timer_reg_5__u0 ( .ck(ispd_clk), .d(n_7601), .o(wbu_latency_tim_val_in_247) );
ms00f80 configuration_latency_timer_reg_6__u0 ( .ck(ispd_clk), .d(n_7600), .o(wbu_latency_tim_val_in_248) );
ms00f80 configuration_latency_timer_reg_7__u0 ( .ck(ispd_clk), .d(n_7599), .o(wbu_latency_tim_val_in_249) );
ms00f80 configuration_pci_am1_reg_10__u0 ( .ck(ispd_clk), .d(n_7453), .o(pciu_am1_in_519) );
ms00f80 configuration_pci_am1_reg_11__u0 ( .ck(ispd_clk), .d(n_7452), .o(pciu_am1_in_520) );
ms00f80 configuration_pci_am1_reg_12__u0 ( .ck(ispd_clk), .d(n_7451), .o(pciu_am1_in_521) );
ms00f80 configuration_pci_am1_reg_13__u0 ( .ck(ispd_clk), .d(n_7450), .o(pciu_am1_in_522) );
ms00f80 configuration_pci_am1_reg_14__u0 ( .ck(ispd_clk), .d(n_7449), .o(pciu_am1_in_523) );
ms00f80 configuration_pci_am1_reg_15__u0 ( .ck(ispd_clk), .d(n_7448), .o(pciu_am1_in_524) );
ms00f80 configuration_pci_am1_reg_16__u0 ( .ck(ispd_clk), .d(n_7447), .o(pciu_am1_in_525) );
ms00f80 configuration_pci_am1_reg_17__u0 ( .ck(ispd_clk), .d(n_7446), .o(pciu_am1_in_526) );
ms00f80 configuration_pci_am1_reg_18__u0 ( .ck(ispd_clk), .d(n_7445), .o(pciu_am1_in_527) );
ms00f80 configuration_pci_am1_reg_19__u0 ( .ck(ispd_clk), .d(n_7433), .o(pciu_am1_in_528) );
ms00f80 configuration_pci_am1_reg_20__u0 ( .ck(ispd_clk), .d(n_7444), .o(pciu_am1_in_529) );
ms00f80 configuration_pci_am1_reg_21__u0 ( .ck(ispd_clk), .d(n_7443), .o(pciu_am1_in_530) );
ms00f80 configuration_pci_am1_reg_22__u0 ( .ck(ispd_clk), .d(n_7458), .o(pciu_am1_in_531) );
ms00f80 configuration_pci_am1_reg_23__u0 ( .ck(ispd_clk), .d(n_7439), .o(pciu_am1_in_532) );
ms00f80 configuration_pci_am1_reg_24__u0 ( .ck(ispd_clk), .d(n_7436), .o(pciu_am1_in_533) );
ms00f80 configuration_pci_am1_reg_25__u0 ( .ck(ispd_clk), .d(n_7435), .o(pciu_am1_in_534) );
ms00f80 configuration_pci_am1_reg_26__u0 ( .ck(ispd_clk), .d(n_7456), .o(pciu_am1_in_535) );
ms00f80 configuration_pci_am1_reg_27__u0 ( .ck(ispd_clk), .d(n_7432), .o(pciu_am1_in_536) );
ms00f80 configuration_pci_am1_reg_28__u0 ( .ck(ispd_clk), .d(n_7431), .o(pciu_am1_in_537) );
ms00f80 configuration_pci_am1_reg_29__u0 ( .ck(ispd_clk), .d(n_7470), .o(pciu_am1_in_538) );
ms00f80 configuration_pci_am1_reg_30__u0 ( .ck(ispd_clk), .d(n_7464), .o(pciu_am1_in_539) );
ms00f80 configuration_pci_am1_reg_31__u0 ( .ck(ispd_clk), .d(n_7430), .o(pciu_am1_in_540) );
ms00f80 configuration_pci_am1_reg_8__u0 ( .ck(ispd_clk), .d(n_7460), .o(pciu_am1_in) );
ms00f80 configuration_pci_am1_reg_9__u0 ( .ck(ispd_clk), .d(n_7429), .o(pciu_am1_in_518) );
ms00f80 configuration_pci_ba0_bit31_8_reg_12__u0 ( .ck(ispd_clk), .d(n_7594), .o(pciu_bar0_in) );
ms00f80 configuration_pci_ba0_bit31_8_reg_13__u0 ( .ck(ispd_clk), .d(n_7593), .o(pciu_bar0_in_361) );
ms00f80 configuration_pci_ba0_bit31_8_reg_14__u0 ( .ck(ispd_clk), .d(n_7592), .o(pciu_bar0_in_362) );
ms00f80 configuration_pci_ba0_bit31_8_reg_15__u0 ( .ck(ispd_clk), .d(n_7597), .o(pciu_bar0_in_363) );
ms00f80 configuration_pci_ba0_bit31_8_reg_16__u0 ( .ck(ispd_clk), .d(n_7603), .o(pciu_bar0_in_364) );
ms00f80 configuration_pci_ba0_bit31_8_reg_17__u0 ( .ck(ispd_clk), .d(n_7589), .o(pciu_bar0_in_365) );
ms00f80 configuration_pci_ba0_bit31_8_reg_18__u0 ( .ck(ispd_clk), .d(n_7591), .o(pciu_bar0_in_366) );
ms00f80 configuration_pci_ba0_bit31_8_reg_19__u0 ( .ck(ispd_clk), .d(n_7588), .o(pciu_bar0_in_367) );
ms00f80 configuration_pci_ba0_bit31_8_reg_20__u0 ( .ck(ispd_clk), .d(n_7587), .o(pciu_bar0_in_368) );
ms00f80 configuration_pci_ba0_bit31_8_reg_21__u0 ( .ck(ispd_clk), .d(n_7586), .o(pciu_bar0_in_369) );
ms00f80 configuration_pci_ba0_bit31_8_reg_22__u0 ( .ck(ispd_clk), .d(n_7585), .o(pciu_bar0_in_370) );
ms00f80 configuration_pci_ba0_bit31_8_reg_23__u0 ( .ck(ispd_clk), .d(n_7584), .o(pciu_bar0_in_371) );
ms00f80 configuration_pci_ba0_bit31_8_reg_24__u0 ( .ck(ispd_clk), .d(n_7583), .o(pciu_bar0_in_372) );
ms00f80 configuration_pci_ba0_bit31_8_reg_25__u0 ( .ck(ispd_clk), .d(n_7582), .o(pciu_bar0_in_373) );
ms00f80 configuration_pci_ba0_bit31_8_reg_26__u0 ( .ck(ispd_clk), .d(n_7581), .o(pciu_bar0_in_374) );
ms00f80 configuration_pci_ba0_bit31_8_reg_27__u0 ( .ck(ispd_clk), .d(n_7580), .o(pciu_bar0_in_375) );
ms00f80 configuration_pci_ba0_bit31_8_reg_28__u0 ( .ck(ispd_clk), .d(n_7579), .o(pciu_bar0_in_376) );
ms00f80 configuration_pci_ba0_bit31_8_reg_29__u0 ( .ck(ispd_clk), .d(n_7578), .o(pciu_bar0_in_377) );
ms00f80 configuration_pci_ba0_bit31_8_reg_30__u0 ( .ck(ispd_clk), .d(n_7577), .o(pciu_bar0_in_378) );
ms00f80 configuration_pci_ba0_bit31_8_reg_31__u0 ( .ck(ispd_clk), .d(n_7576), .o(pciu_bar0_in_379) );
ms00f80 configuration_pci_ba1_bit31_8_reg_10__u0 ( .ck(ispd_clk), .d(n_7483), .o(pciu_bar1_in_381) );
ms00f80 configuration_pci_ba1_bit31_8_reg_11__u0 ( .ck(ispd_clk), .d(n_7482), .o(pciu_bar1_in_382) );
ms00f80 configuration_pci_ba1_bit31_8_reg_12__u0 ( .ck(ispd_clk), .d(n_7481), .o(pciu_bar1_in_383) );
ms00f80 configuration_pci_ba1_bit31_8_reg_13__u0 ( .ck(ispd_clk), .d(n_7480), .o(pciu_bar1_in_384) );
ms00f80 configuration_pci_ba1_bit31_8_reg_14__u0 ( .ck(ispd_clk), .d(n_7479), .o(pciu_bar1_in_385) );
ms00f80 configuration_pci_ba1_bit31_8_reg_15__u0 ( .ck(ispd_clk), .d(n_7478), .o(pciu_bar1_in_386) );
ms00f80 configuration_pci_ba1_bit31_8_reg_16__u0 ( .ck(ispd_clk), .d(n_7477), .o(pciu_bar1_in_387) );
ms00f80 configuration_pci_ba1_bit31_8_reg_17__u0 ( .ck(ispd_clk), .d(n_7476), .o(pciu_bar1_in_388) );
ms00f80 configuration_pci_ba1_bit31_8_reg_18__u0 ( .ck(ispd_clk), .d(n_7500), .o(pciu_bar1_in_389) );
ms00f80 configuration_pci_ba1_bit31_8_reg_19__u0 ( .ck(ispd_clk), .d(n_7499), .o(pciu_bar1_in_390) );
ms00f80 configuration_pci_ba1_bit31_8_reg_20__u0 ( .ck(ispd_clk), .d(n_7497), .o(pciu_bar1_in_391) );
ms00f80 configuration_pci_ba1_bit31_8_reg_21__u0 ( .ck(ispd_clk), .d(n_7495), .o(pciu_bar1_in_392) );
ms00f80 configuration_pci_ba1_bit31_8_reg_22__u0 ( .ck(ispd_clk), .d(n_7496), .o(pciu_bar1_in_393) );
ms00f80 configuration_pci_ba1_bit31_8_reg_23__u0 ( .ck(ispd_clk), .d(n_7494), .o(pciu_bar1_in_394) );
ms00f80 configuration_pci_ba1_bit31_8_reg_24__u0 ( .ck(ispd_clk), .d(n_7493), .o(pciu_bar1_in_395) );
ms00f80 configuration_pci_ba1_bit31_8_reg_25__u0 ( .ck(ispd_clk), .d(n_7492), .o(pciu_bar1_in_396) );
ms00f80 configuration_pci_ba1_bit31_8_reg_26__u0 ( .ck(ispd_clk), .d(n_7491), .o(pciu_bar1_in_397) );
ms00f80 configuration_pci_ba1_bit31_8_reg_27__u0 ( .ck(ispd_clk), .d(n_7490), .o(pciu_bar1_in_398) );
ms00f80 configuration_pci_ba1_bit31_8_reg_28__u0 ( .ck(ispd_clk), .d(n_7489), .o(pciu_bar1_in_399) );
ms00f80 configuration_pci_ba1_bit31_8_reg_29__u0 ( .ck(ispd_clk), .d(n_7488), .o(pciu_bar1_in_400) );
ms00f80 configuration_pci_ba1_bit31_8_reg_30__u0 ( .ck(ispd_clk), .d(n_7487), .o(pciu_bar1_in_401) );
ms00f80 configuration_pci_ba1_bit31_8_reg_31__u0 ( .ck(ispd_clk), .d(n_7486), .o(pciu_bar1_in_402) );
ms00f80 configuration_pci_ba1_bit31_8_reg_8__u0 ( .ck(ispd_clk), .d(n_7484), .o(pciu_bar1_in) );
ms00f80 configuration_pci_ba1_bit31_8_reg_9__u0 ( .ck(ispd_clk), .d(n_7485), .o(pciu_bar1_in_380) );
ms00f80 configuration_pci_err_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_4851), .o(configuration_pci_err_addr) );
ms00f80 configuration_pci_err_addr_reg_10__u0 ( .ck(ispd_clk), .d(n_4849), .o(configuration_pci_err_addr_480) );
ms00f80 configuration_pci_err_addr_reg_11__u0 ( .ck(ispd_clk), .d(n_4848), .o(configuration_pci_err_addr_481) );
ms00f80 configuration_pci_err_addr_reg_12__u0 ( .ck(ispd_clk), .d(n_4847), .o(configuration_pci_err_addr_482) );
ms00f80 configuration_pci_err_addr_reg_13__u0 ( .ck(ispd_clk), .d(n_4846), .o(configuration_pci_err_addr_483) );
ms00f80 configuration_pci_err_addr_reg_14__u0 ( .ck(ispd_clk), .d(n_4845), .o(configuration_pci_err_addr_484) );
ms00f80 configuration_pci_err_addr_reg_15__u0 ( .ck(ispd_clk), .d(n_4844), .o(configuration_pci_err_addr_485) );
ms00f80 configuration_pci_err_addr_reg_16__u0 ( .ck(ispd_clk), .d(n_4843), .o(configuration_pci_err_addr_486) );
ms00f80 configuration_pci_err_addr_reg_17__u0 ( .ck(ispd_clk), .d(n_4842), .o(configuration_pci_err_addr_487) );
ms00f80 configuration_pci_err_addr_reg_18__u0 ( .ck(ispd_clk), .d(n_4841), .o(configuration_pci_err_addr_488) );
ms00f80 configuration_pci_err_addr_reg_19__u0 ( .ck(ispd_clk), .d(n_4840), .o(configuration_pci_err_addr_489) );
ms00f80 configuration_pci_err_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_4839), .o(configuration_pci_err_addr_471) );
ms00f80 configuration_pci_err_addr_reg_20__u0 ( .ck(ispd_clk), .d(n_4838), .o(configuration_pci_err_addr_490) );
ms00f80 configuration_pci_err_addr_reg_21__u0 ( .ck(ispd_clk), .d(n_4837), .o(configuration_pci_err_addr_491) );
ms00f80 configuration_pci_err_addr_reg_22__u0 ( .ck(ispd_clk), .d(n_4836), .o(configuration_pci_err_addr_492) );
ms00f80 configuration_pci_err_addr_reg_23__u0 ( .ck(ispd_clk), .d(n_4835), .o(configuration_pci_err_addr_493) );
ms00f80 configuration_pci_err_addr_reg_24__u0 ( .ck(ispd_clk), .d(n_4834), .o(configuration_pci_err_addr_494) );
ms00f80 configuration_pci_err_addr_reg_25__u0 ( .ck(ispd_clk), .d(n_4833), .o(configuration_pci_err_addr_495) );
ms00f80 configuration_pci_err_addr_reg_26__u0 ( .ck(ispd_clk), .d(n_4831), .o(configuration_pci_err_addr_496) );
ms00f80 configuration_pci_err_addr_reg_27__u0 ( .ck(ispd_clk), .d(n_4832), .o(configuration_pci_err_addr_497) );
ms00f80 configuration_pci_err_addr_reg_28__u0 ( .ck(ispd_clk), .d(n_4830), .o(configuration_pci_err_addr_498) );
ms00f80 configuration_pci_err_addr_reg_29__u0 ( .ck(ispd_clk), .d(n_4828), .o(configuration_pci_err_addr_499) );
ms00f80 configuration_pci_err_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_5712), .o(configuration_pci_err_addr_472) );
ms00f80 configuration_pci_err_addr_reg_30__u0 ( .ck(ispd_clk), .d(n_5710), .o(configuration_pci_err_addr_500) );
ms00f80 configuration_pci_err_addr_reg_31__u0 ( .ck(ispd_clk), .d(n_5709), .o(configuration_pci_err_addr_501) );
ms00f80 configuration_pci_err_addr_reg_3__u0 ( .ck(ispd_clk), .d(n_5708), .o(configuration_pci_err_addr_473) );
ms00f80 configuration_pci_err_addr_reg_4__u0 ( .ck(ispd_clk), .d(n_5707), .o(configuration_pci_err_addr_474) );
ms00f80 configuration_pci_err_addr_reg_5__u0 ( .ck(ispd_clk), .d(n_5705), .o(configuration_pci_err_addr_475) );
ms00f80 configuration_pci_err_addr_reg_6__u0 ( .ck(ispd_clk), .d(n_5704), .o(configuration_pci_err_addr_476) );
ms00f80 configuration_pci_err_addr_reg_7__u0 ( .ck(ispd_clk), .d(n_5703), .o(configuration_pci_err_addr_477) );
ms00f80 configuration_pci_err_addr_reg_8__u0 ( .ck(ispd_clk), .d(n_5702), .o(configuration_pci_err_addr_478) );
ms00f80 configuration_pci_err_addr_reg_9__u0 ( .ck(ispd_clk), .d(n_5701), .o(configuration_pci_err_addr_479) );
ms00f80 configuration_pci_err_cs_bit0_reg_u0 ( .ck(ispd_clk), .d(n_8519), .o(configuration_pci_err_cs_bit0) );
ms00f80 configuration_pci_err_cs_bit10_reg_u0 ( .ck(ispd_clk), .d(n_4873), .o(configuration_pci_err_cs_bit10) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_24__u0 ( .ck(ispd_clk), .d(n_5699), .o(configuration_pci_err_cs_bit31_24) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_25__u0 ( .ck(ispd_clk), .d(n_5696), .o(configuration_pci_err_cs_bit_464) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_26__u0 ( .ck(ispd_clk), .d(n_5694), .o(configuration_pci_err_cs_bit_465) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_27__u0 ( .ck(ispd_clk), .d(n_5691), .o(configuration_pci_err_cs_bit_466) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_28__u0 ( .ck(ispd_clk), .d(n_4867), .o(configuration_pci_err_cs_bit_467) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_29__u0 ( .ck(ispd_clk), .d(n_4866), .o(configuration_pci_err_cs_bit_468) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_30__u0 ( .ck(ispd_clk), .d(n_4864), .o(configuration_pci_err_cs_bit_469) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_31__u0 ( .ck(ispd_clk), .d(n_4863), .o(configuration_pci_err_cs_bit_470) );
ms00f80 configuration_pci_err_cs_bit8_reg_u0 ( .ck(ispd_clk), .d(configuration_meta_pci_err_cs_bits), .o(configuration_pci_err_cs_bit8) );
ms00f80 configuration_pci_err_cs_bit9_reg_u0 ( .ck(ispd_clk), .d(n_4872), .o(configuration_pci_err_cs_bit9) );
ms00f80 configuration_pci_err_cs_bits_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_736), .o(configuration_meta_pci_err_cs_bits) );
ms00f80 configuration_pci_err_data_reg_0__u0 ( .ck(ispd_clk), .d(n_5689), .o(configuration_pci_err_data) );
ms00f80 configuration_pci_err_data_reg_10__u0 ( .ck(ispd_clk), .d(n_5688), .o(configuration_pci_err_data_511) );
ms00f80 configuration_pci_err_data_reg_11__u0 ( .ck(ispd_clk), .d(n_5687), .o(configuration_pci_err_data_512) );
ms00f80 configuration_pci_err_data_reg_12__u0 ( .ck(ispd_clk), .d(n_5686), .o(configuration_pci_err_data_513) );
ms00f80 configuration_pci_err_data_reg_13__u0 ( .ck(ispd_clk), .d(n_5684), .o(configuration_pci_err_data_514) );
ms00f80 configuration_pci_err_data_reg_14__u0 ( .ck(ispd_clk), .d(n_5682), .o(configuration_pci_err_data_515) );
ms00f80 configuration_pci_err_data_reg_15__u0 ( .ck(ispd_clk), .d(n_5681), .o(configuration_pci_err_data_516) );
ms00f80 configuration_pci_err_data_reg_16__u0 ( .ck(ispd_clk), .d(n_5679), .o(configuration_pci_err_data_517) );
ms00f80 configuration_pci_err_data_reg_17__u0 ( .ck(ispd_clk), .d(n_5678), .o(configuration_pci_err_data_518) );
ms00f80 configuration_pci_err_data_reg_18__u0 ( .ck(ispd_clk), .d(n_5676), .o(configuration_pci_err_data_519) );
ms00f80 configuration_pci_err_data_reg_19__u0 ( .ck(ispd_clk), .d(n_5675), .o(configuration_pci_err_data_520) );
ms00f80 configuration_pci_err_data_reg_1__u0 ( .ck(ispd_clk), .d(n_5673), .o(configuration_pci_err_data_502) );
ms00f80 configuration_pci_err_data_reg_20__u0 ( .ck(ispd_clk), .d(n_5672), .o(configuration_pci_err_data_521) );
ms00f80 configuration_pci_err_data_reg_21__u0 ( .ck(ispd_clk), .d(n_5670), .o(configuration_pci_err_data_522) );
ms00f80 configuration_pci_err_data_reg_22__u0 ( .ck(ispd_clk), .d(n_5669), .o(configuration_pci_err_data_523) );
ms00f80 configuration_pci_err_data_reg_23__u0 ( .ck(ispd_clk), .d(n_5668), .o(configuration_pci_err_data_524) );
ms00f80 configuration_pci_err_data_reg_24__u0 ( .ck(ispd_clk), .d(n_5666), .o(configuration_pci_err_data_525) );
ms00f80 configuration_pci_err_data_reg_25__u0 ( .ck(ispd_clk), .d(n_5664), .o(configuration_pci_err_data_526) );
ms00f80 configuration_pci_err_data_reg_26__u0 ( .ck(ispd_clk), .d(n_5663), .o(configuration_pci_err_data_527) );
ms00f80 configuration_pci_err_data_reg_27__u0 ( .ck(ispd_clk), .d(n_5662), .o(configuration_pci_err_data_528) );
ms00f80 configuration_pci_err_data_reg_28__u0 ( .ck(ispd_clk), .d(n_5660), .o(configuration_pci_err_data_529) );
ms00f80 configuration_pci_err_data_reg_29__u0 ( .ck(ispd_clk), .d(n_5658), .o(configuration_pci_err_data_530) );
ms00f80 configuration_pci_err_data_reg_2__u0 ( .ck(ispd_clk), .d(n_5648), .o(configuration_pci_err_data_503) );
ms00f80 configuration_pci_err_data_reg_30__u0 ( .ck(ispd_clk), .d(n_5657), .o(configuration_pci_err_data_531) );
ms00f80 configuration_pci_err_data_reg_31__u0 ( .ck(ispd_clk), .d(n_5656), .o(configuration_pci_err_data_532) );
ms00f80 configuration_pci_err_data_reg_3__u0 ( .ck(ispd_clk), .d(n_5655), .o(configuration_pci_err_data_504) );
ms00f80 configuration_pci_err_data_reg_4__u0 ( .ck(ispd_clk), .d(n_5654), .o(configuration_pci_err_data_505) );
ms00f80 configuration_pci_err_data_reg_5__u0 ( .ck(ispd_clk), .d(n_5652), .o(configuration_pci_err_data_506) );
ms00f80 configuration_pci_err_data_reg_6__u0 ( .ck(ispd_clk), .d(n_5646), .o(configuration_pci_err_data_507) );
ms00f80 configuration_pci_err_data_reg_7__u0 ( .ck(ispd_clk), .d(n_5651), .o(configuration_pci_err_data_508) );
ms00f80 configuration_pci_err_data_reg_8__u0 ( .ck(ispd_clk), .d(n_5650), .o(configuration_pci_err_data_509) );
ms00f80 configuration_pci_err_data_reg_9__u0 ( .ck(ispd_clk), .d(n_5649), .o(configuration_pci_err_data_510) );
ms00f80 configuration_pci_img_ctrl1_bit2_1_reg_1__u0 ( .ck(ispd_clk), .d(n_8523), .o(pciu_pref_en_in_320) );
ms00f80 configuration_pci_img_ctrl1_bit2_1_reg_2__u0 ( .ck(ispd_clk), .d(n_8522), .o(n_14910) );
ms00f80 configuration_pci_ta1_reg_10__u0 ( .ck(ispd_clk), .d(n_7271), .o(n_14913) );
ms00f80 configuration_pci_ta1_reg_11__u0 ( .ck(ispd_clk), .d(n_7264), .o(n_14914) );
ms00f80 configuration_pci_ta1_reg_12__u0 ( .ck(ispd_clk), .d(n_7263), .o(n_14915) );
ms00f80 configuration_pci_ta1_reg_13__u0 ( .ck(ispd_clk), .d(n_7262), .o(n_14916) );
ms00f80 configuration_pci_ta1_reg_14__u0 ( .ck(ispd_clk), .d(n_7261), .o(n_14917) );
ms00f80 configuration_pci_ta1_reg_15__u0 ( .ck(ispd_clk), .d(n_7228), .o(n_14918) );
ms00f80 configuration_pci_ta1_reg_16__u0 ( .ck(ispd_clk), .d(n_7258), .o(n_14919) );
ms00f80 configuration_pci_ta1_reg_17__u0 ( .ck(ispd_clk), .d(n_7257), .o(n_14920) );
ms00f80 configuration_pci_ta1_reg_18__u0 ( .ck(ispd_clk), .d(n_7256), .o(n_14921) );
ms00f80 configuration_pci_ta1_reg_19__u0 ( .ck(ispd_clk), .d(n_7298), .o(n_14922) );
ms00f80 configuration_pci_ta1_reg_20__u0 ( .ck(ispd_clk), .d(n_7253), .o(n_14923) );
ms00f80 configuration_pci_ta1_reg_21__u0 ( .ck(ispd_clk), .d(n_7252), .o(n_14924) );
ms00f80 configuration_pci_ta1_reg_22__u0 ( .ck(ispd_clk), .d(n_7251), .o(n_14925) );
ms00f80 configuration_pci_ta1_reg_23__u0 ( .ck(ispd_clk), .d(n_7248), .o(n_14926) );
ms00f80 configuration_pci_ta1_reg_24__u0 ( .ck(ispd_clk), .d(n_7247), .o(n_14927) );
ms00f80 configuration_pci_ta1_reg_25__u0 ( .ck(ispd_clk), .d(n_7246), .o(n_14928) );
ms00f80 configuration_pci_ta1_reg_26__u0 ( .ck(ispd_clk), .d(n_7243), .o(n_14929) );
ms00f80 configuration_pci_ta1_reg_27__u0 ( .ck(ispd_clk), .d(n_7281), .o(n_14930) );
ms00f80 configuration_pci_ta1_reg_28__u0 ( .ck(ispd_clk), .d(n_7229), .o(n_14931) );
ms00f80 configuration_pci_ta1_reg_29__u0 ( .ck(ispd_clk), .d(n_7297), .o(n_14932) );
ms00f80 configuration_pci_ta1_reg_30__u0 ( .ck(ispd_clk), .d(n_7227), .o(n_14933) );
ms00f80 configuration_pci_ta1_reg_31__u0 ( .ck(ispd_clk), .d(n_7238), .o(n_14934) );
ms00f80 configuration_pci_ta1_reg_8__u0 ( .ck(ispd_clk), .d(n_7237), .o(n_14911) );
ms00f80 configuration_pci_ta1_reg_9__u0 ( .ck(ispd_clk), .d(n_7236), .o(n_14912) );
ms00f80 configuration_rst_inactive_reg_u0 ( .ck(ispd_clk), .d(configuration_rst_inactive_sync), .o(configuration_rst_inactive) );
ms00f80 configuration_rst_inactive_sync_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15175), .o(configuration_rst_inactive_sync) );
ms00f80 configuration_set_isr_bit2_reg_u0 ( .ck(ispd_clk), .d(n_5730), .o(configuration_set_isr_bit2_reg_Q) );
in01s01 configuration_set_isr_bit2_reg_u1 ( .a(configuration_set_isr_bit2_reg_Q), .o(configuration_set_isr_bit2) );
ms00f80 configuration_set_pci_err_cs_bit8_reg_u0 ( .ck(ispd_clk), .d(n_4695), .o(configuration_set_pci_err_cs_bit8_reg_Q) );
in01s01 configuration_set_pci_err_cs_bit8_reg_u1 ( .a(configuration_set_pci_err_cs_bit8_reg_Q), .o(configuration_set_pci_err_cs_bit8) );
ms00f80 configuration_status_bit15_11_reg_11__u0 ( .ck(ispd_clk), .d(n_8472), .o(configuration_status_bit_435) );
ms00f80 configuration_status_bit15_11_reg_12__u0 ( .ck(ispd_clk), .d(n_8509), .o(configuration_status_bit_407) );
ms00f80 configuration_status_bit15_11_reg_13__u0 ( .ck(ispd_clk), .d(n_8506), .o(configuration_status_bit_379) );
ms00f80 configuration_status_bit15_11_reg_14__u0 ( .ck(ispd_clk), .d(n_14080), .o(configuration_status_bit_351) );
ms00f80 configuration_status_bit15_11_reg_15__u0 ( .ck(ispd_clk), .d(n_14491), .o(configuration_status_bit_322) );
ms00f80 configuration_status_bit8_reg_u0 ( .ck(ispd_clk), .d(n_14901), .o(configuration_status_bit8) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_2__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits), .o(configuration_sync_cache_lsize_to_wb_bits_reg_2__Q) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_3__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits_926), .o(configuration_sync_cache_lsize_to_wb_bits_reg_3__Q) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_4__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits_927), .o(configuration_sync_cache_lsize_to_wb_bits_reg_4__Q) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_5__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits_928), .o(pciu_cache_line_size_in_775) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_6__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits_929), .o(pciu_cache_line_size_in_776) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_7__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits_930), .o(pciu_cache_line_size_in_777) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_8__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits_931), .o(pciu_cache_lsize_not_zero_in) );
ms00f80 configuration_sync_command_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_meta_command_bit), .o(configuration_sync_command_bit2) );
ms00f80 configuration_sync_isr_2_clear_delete_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(configuration_sync_isr_2_sync_del_bit), .o(configuration_sync_isr_2_meta_bckp_bit) );
ms00f80 configuration_sync_isr_2_del_bit_reg_u0 ( .ck(ispd_clk), .d(n_8432), .o(configuration_sync_isr_2_del_bit_reg_Q) );
ms00f80 configuration_sync_isr_2_delayed_bckp_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_isr_2_sync_bckp_bit), .o(configuration_sync_isr_2_delayed_bckp_bit_reg_Q) );
in01s01 configuration_sync_isr_2_delayed_bckp_bit_reg_u1 ( .a(configuration_sync_isr_2_delayed_bckp_bit_reg_Q), .o(configuration_sync_isr_2_delayed_bckp_bit) );
ms00f80 configuration_sync_isr_2_delayed_del_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_isr_2_sync_del_bit), .o(configuration_sync_isr_2_delayed_del_bit_reg_Q) );
in01s01 configuration_sync_isr_2_delayed_del_bit_reg_u1 ( .a(configuration_sync_isr_2_delayed_del_bit_reg_Q), .o(configuration_sync_isr_2_delayed_del_bit) );
ms00f80 configuration_sync_isr_2_delete_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(configuration_sync_isr_2_del_bit_reg_Q), .o(configuration_sync_isr_2_meta_del_bit) );
ms00f80 configuration_sync_isr_2_sync_bckp_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_isr_2_meta_bckp_bit), .o(configuration_sync_isr_2_sync_bckp_bit) );
ms00f80 configuration_sync_isr_2_sync_del_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_isr_2_meta_del_bit), .o(configuration_sync_isr_2_sync_del_bit) );
ms00f80 configuration_sync_pci_err_cs_8_clear_delete_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(configuration_sync_pci_err_cs_8_sync_del_bit), .o(configuration_sync_pci_err_cs_8_meta_bckp_bit) );
ms00f80 configuration_sync_pci_err_cs_8_del_bit_reg_u0 ( .ck(ispd_clk), .d(n_8431), .o(configuration_sync_pci_err_cs_8_del_bit_reg_Q) );
ms00f80 configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_pci_err_cs_8_sync_bckp_bit), .o(configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg_Q) );
in01s01 configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg_u1 ( .a(configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg_Q), .o(configuration_sync_pci_err_cs_8_delayed_bckp_bit) );
ms00f80 configuration_sync_pci_err_cs_8_delayed_del_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_pci_err_cs_8_sync_del_bit), .o(configuration_sync_pci_err_cs_8_delayed_del_bit_reg_Q) );
in01s01 configuration_sync_pci_err_cs_8_delayed_del_bit_reg_u1 ( .a(configuration_sync_pci_err_cs_8_delayed_del_bit_reg_Q), .o(configuration_sync_pci_err_cs_8_delayed_del_bit) );
ms00f80 configuration_sync_pci_err_cs_8_delete_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(configuration_sync_pci_err_cs_8_del_bit_reg_Q), .o(configuration_sync_pci_err_cs_8_meta_del_bit) );
ms00f80 configuration_sync_pci_err_cs_8_sync_bckp_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_pci_err_cs_8_meta_bckp_bit), .o(configuration_sync_pci_err_cs_8_sync_bckp_bit) );
ms00f80 configuration_sync_pci_err_cs_8_sync_del_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_pci_err_cs_8_meta_del_bit), .o(configuration_sync_pci_err_cs_8_sync_del_bit) );
ms00f80 configuration_wb_am1_reg_31__u0 ( .ck(ispd_clk), .d(n_8542), .o(wbu_am1_in) );
ms00f80 configuration_wb_am2_reg_31__u0 ( .ck(ispd_clk), .d(n_8541), .o(wbu_am2_in) );
ms00f80 configuration_wb_ba1_bit0_reg_u0 ( .ck(ispd_clk), .d(n_8470), .o(wbu_map_in_131) );
ms00f80 configuration_wb_ba1_bit31_12_reg_31__u0 ( .ck(ispd_clk), .d(n_8469), .o(wbu_bar1_in) );
ms00f80 configuration_wb_ba2_bit0_reg_u0 ( .ck(ispd_clk), .d(n_8467), .o(wbu_map_in_132) );
ms00f80 configuration_wb_ba2_bit31_12_reg_31__u0 ( .ck(ispd_clk), .d(n_8466), .o(wbu_bar2_in) );
ms00f80 configuration_wb_err_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_5718), .o(configuration_wb_err_addr) );
ms00f80 configuration_wb_err_addr_reg_10__u0 ( .ck(ispd_clk), .d(n_5587), .o(configuration_wb_err_addr_542) );
ms00f80 configuration_wb_err_addr_reg_11__u0 ( .ck(ispd_clk), .d(n_5585), .o(configuration_wb_err_addr_543) );
ms00f80 configuration_wb_err_addr_reg_12__u0 ( .ck(ispd_clk), .d(n_5583), .o(configuration_wb_err_addr_544) );
ms00f80 configuration_wb_err_addr_reg_13__u0 ( .ck(ispd_clk), .d(n_5582), .o(configuration_wb_err_addr_545) );
ms00f80 configuration_wb_err_addr_reg_14__u0 ( .ck(ispd_clk), .d(n_5581), .o(configuration_wb_err_addr_546) );
ms00f80 configuration_wb_err_addr_reg_15__u0 ( .ck(ispd_clk), .d(n_5580), .o(configuration_wb_err_addr_547) );
ms00f80 configuration_wb_err_addr_reg_16__u0 ( .ck(ispd_clk), .d(n_5579), .o(configuration_wb_err_addr_548) );
ms00f80 configuration_wb_err_addr_reg_17__u0 ( .ck(ispd_clk), .d(n_5578), .o(configuration_wb_err_addr_549) );
ms00f80 configuration_wb_err_addr_reg_18__u0 ( .ck(ispd_clk), .d(n_5577), .o(configuration_wb_err_addr_550) );
ms00f80 configuration_wb_err_addr_reg_19__u0 ( .ck(ispd_clk), .d(n_5576), .o(configuration_wb_err_addr_551) );
ms00f80 configuration_wb_err_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_4891), .o(configuration_wb_err_addr_533) );
ms00f80 configuration_wb_err_addr_reg_20__u0 ( .ck(ispd_clk), .d(n_5575), .o(configuration_wb_err_addr_552) );
ms00f80 configuration_wb_err_addr_reg_21__u0 ( .ck(ispd_clk), .d(n_5574), .o(configuration_wb_err_addr_553) );
ms00f80 configuration_wb_err_addr_reg_22__u0 ( .ck(ispd_clk), .d(n_5573), .o(configuration_wb_err_addr_554) );
ms00f80 configuration_wb_err_addr_reg_23__u0 ( .ck(ispd_clk), .d(n_5572), .o(configuration_wb_err_addr_555) );
ms00f80 configuration_wb_err_addr_reg_24__u0 ( .ck(ispd_clk), .d(n_5571), .o(configuration_wb_err_addr_556) );
ms00f80 configuration_wb_err_addr_reg_25__u0 ( .ck(ispd_clk), .d(n_5570), .o(configuration_wb_err_addr_557) );
ms00f80 configuration_wb_err_addr_reg_26__u0 ( .ck(ispd_clk), .d(n_5569), .o(configuration_wb_err_addr_558) );
ms00f80 configuration_wb_err_addr_reg_27__u0 ( .ck(ispd_clk), .d(n_5568), .o(configuration_wb_err_addr_559) );
ms00f80 configuration_wb_err_addr_reg_28__u0 ( .ck(ispd_clk), .d(n_5567), .o(configuration_wb_err_addr_560) );
ms00f80 configuration_wb_err_addr_reg_29__u0 ( .ck(ispd_clk), .d(n_5566), .o(configuration_wb_err_addr_561) );
ms00f80 configuration_wb_err_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_5565), .o(configuration_wb_err_addr_534) );
ms00f80 configuration_wb_err_addr_reg_30__u0 ( .ck(ispd_clk), .d(n_5563), .o(configuration_wb_err_addr_562) );
ms00f80 configuration_wb_err_addr_reg_31__u0 ( .ck(ispd_clk), .d(n_5561), .o(configuration_wb_err_addr_563) );
ms00f80 configuration_wb_err_addr_reg_3__u0 ( .ck(ispd_clk), .d(n_5559), .o(configuration_wb_err_addr_535) );
ms00f80 configuration_wb_err_addr_reg_4__u0 ( .ck(ispd_clk), .d(n_5558), .o(configuration_wb_err_addr_536) );
ms00f80 configuration_wb_err_addr_reg_5__u0 ( .ck(ispd_clk), .d(n_5557), .o(configuration_wb_err_addr_537) );
ms00f80 configuration_wb_err_addr_reg_6__u0 ( .ck(ispd_clk), .d(n_5556), .o(configuration_wb_err_addr_538) );
ms00f80 configuration_wb_err_addr_reg_7__u0 ( .ck(ispd_clk), .d(n_5555), .o(configuration_wb_err_addr_539) );
ms00f80 configuration_wb_err_addr_reg_8__u0 ( .ck(ispd_clk), .d(n_5554), .o(configuration_wb_err_addr_540) );
ms00f80 configuration_wb_err_addr_reg_9__u0 ( .ck(ispd_clk), .d(n_5553), .o(configuration_wb_err_addr_541) );
ms00f80 configuration_wb_err_cs_bit0_reg_u0 ( .ck(ispd_clk), .d(n_8518), .o(configuration_wb_err_cs_bit0) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_24__u0 ( .ck(ispd_clk), .d(n_5552), .o(configuration_wb_err_cs_bit31_24) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_25__u0 ( .ck(ispd_clk), .d(n_5639), .o(configuration_wb_err_cs_bit_564) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_26__u0 ( .ck(ispd_clk), .d(n_5638), .o(configuration_wb_err_cs_bit_565) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_27__u0 ( .ck(ispd_clk), .d(n_5637), .o(configuration_wb_err_cs_bit_566) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_28__u0 ( .ck(ispd_clk), .d(n_5636), .o(configuration_wb_err_cs_bit_567) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_29__u0 ( .ck(ispd_clk), .d(n_5635), .o(configuration_wb_err_cs_bit_568) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_30__u0 ( .ck(ispd_clk), .d(n_5634), .o(configuration_wb_err_cs_bit_569) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_31__u0 ( .ck(ispd_clk), .d(n_5632), .o(configuration_wb_err_cs_bit_570) );
ms00f80 configuration_wb_err_cs_bit8_reg_u0 ( .ck(ispd_clk), .d(n_8510), .o(configuration_wb_err_cs_bit8) );
ms00f80 configuration_wb_err_cs_bit9_reg_u0 ( .ck(ispd_clk), .d(n_6218), .o(configuration_wb_err_cs_bit9) );
ms00f80 configuration_wb_err_data_reg_0__u0 ( .ck(ispd_clk), .d(n_5631), .o(configuration_wb_err_data) );
ms00f80 configuration_wb_err_data_reg_10__u0 ( .ck(ispd_clk), .d(n_5630), .o(configuration_wb_err_data_580) );
ms00f80 configuration_wb_err_data_reg_11__u0 ( .ck(ispd_clk), .d(n_5628), .o(configuration_wb_err_data_581) );
ms00f80 configuration_wb_err_data_reg_12__u0 ( .ck(ispd_clk), .d(n_5627), .o(configuration_wb_err_data_582) );
ms00f80 configuration_wb_err_data_reg_13__u0 ( .ck(ispd_clk), .d(n_5626), .o(configuration_wb_err_data_583) );
ms00f80 configuration_wb_err_data_reg_14__u0 ( .ck(ispd_clk), .d(n_5625), .o(configuration_wb_err_data_584) );
ms00f80 configuration_wb_err_data_reg_15__u0 ( .ck(ispd_clk), .d(n_5623), .o(configuration_wb_err_data_585) );
ms00f80 configuration_wb_err_data_reg_16__u0 ( .ck(ispd_clk), .d(n_5622), .o(configuration_wb_err_data_586) );
ms00f80 configuration_wb_err_data_reg_17__u0 ( .ck(ispd_clk), .d(n_5620), .o(configuration_wb_err_data_587) );
ms00f80 configuration_wb_err_data_reg_18__u0 ( .ck(ispd_clk), .d(n_5619), .o(configuration_wb_err_data_588) );
ms00f80 configuration_wb_err_data_reg_19__u0 ( .ck(ispd_clk), .d(n_5618), .o(configuration_wb_err_data_589) );
ms00f80 configuration_wb_err_data_reg_1__u0 ( .ck(ispd_clk), .d(n_5617), .o(configuration_wb_err_data_571) );
ms00f80 configuration_wb_err_data_reg_20__u0 ( .ck(ispd_clk), .d(n_5616), .o(configuration_wb_err_data_590) );
ms00f80 configuration_wb_err_data_reg_21__u0 ( .ck(ispd_clk), .d(n_5614), .o(configuration_wb_err_data_591) );
ms00f80 configuration_wb_err_data_reg_22__u0 ( .ck(ispd_clk), .d(n_5612), .o(configuration_wb_err_data_592) );
ms00f80 configuration_wb_err_data_reg_23__u0 ( .ck(ispd_clk), .d(n_5611), .o(configuration_wb_err_data_593) );
ms00f80 configuration_wb_err_data_reg_24__u0 ( .ck(ispd_clk), .d(n_5609), .o(configuration_wb_err_data_594) );
ms00f80 configuration_wb_err_data_reg_25__u0 ( .ck(ispd_clk), .d(n_5608), .o(configuration_wb_err_data_595) );
ms00f80 configuration_wb_err_data_reg_26__u0 ( .ck(ispd_clk), .d(n_5607), .o(configuration_wb_err_data_596) );
ms00f80 configuration_wb_err_data_reg_27__u0 ( .ck(ispd_clk), .d(n_5606), .o(configuration_wb_err_data_597) );
ms00f80 configuration_wb_err_data_reg_28__u0 ( .ck(ispd_clk), .d(n_5604), .o(configuration_wb_err_data_598) );
ms00f80 configuration_wb_err_data_reg_29__u0 ( .ck(ispd_clk), .d(n_5603), .o(configuration_wb_err_data_599) );
ms00f80 configuration_wb_err_data_reg_2__u0 ( .ck(ispd_clk), .d(n_5601), .o(configuration_wb_err_data_572) );
ms00f80 configuration_wb_err_data_reg_30__u0 ( .ck(ispd_clk), .d(n_5600), .o(configuration_wb_err_data_600) );
ms00f80 configuration_wb_err_data_reg_31__u0 ( .ck(ispd_clk), .d(n_5598), .o(configuration_wb_err_data_601) );
ms00f80 configuration_wb_err_data_reg_3__u0 ( .ck(ispd_clk), .d(n_5597), .o(configuration_wb_err_data_573) );
ms00f80 configuration_wb_err_data_reg_4__u0 ( .ck(ispd_clk), .d(n_5595), .o(configuration_wb_err_data_574) );
ms00f80 configuration_wb_err_data_reg_5__u0 ( .ck(ispd_clk), .d(n_5594), .o(configuration_wb_err_data_575) );
ms00f80 configuration_wb_err_data_reg_6__u0 ( .ck(ispd_clk), .d(n_5593), .o(configuration_wb_err_data_576) );
ms00f80 configuration_wb_err_data_reg_7__u0 ( .ck(ispd_clk), .d(n_5591), .o(configuration_wb_err_data_577) );
ms00f80 configuration_wb_err_data_reg_8__u0 ( .ck(ispd_clk), .d(n_5589), .o(configuration_wb_err_data_578) );
ms00f80 configuration_wb_err_data_reg_9__u0 ( .ck(ispd_clk), .d(n_5588), .o(configuration_wb_err_data_579) );
ms00f80 configuration_wb_img_ctrl1_bit2_0_reg_0__u0 ( .ck(ispd_clk), .d(n_8478), .o(wbu_mrl_en_in_141) );
ms00f80 configuration_wb_img_ctrl1_bit2_0_reg_1__u0 ( .ck(ispd_clk), .d(n_8474), .o(wbu_pref_en_in_136) );
ms00f80 configuration_wb_img_ctrl1_bit2_0_reg_2__u0 ( .ck(ispd_clk), .d(n_8477), .o(n_14907) );
ms00f80 configuration_wb_img_ctrl2_bit2_0_reg_0__u0 ( .ck(ispd_clk), .d(n_8460), .o(wbu_mrl_en_in_142) );
ms00f80 configuration_wb_img_ctrl2_bit2_0_reg_1__u0 ( .ck(ispd_clk), .d(n_8459), .o(wbu_pref_en_in_137) );
ms00f80 configuration_wb_img_ctrl2_bit2_0_reg_2__u0 ( .ck(ispd_clk), .d(n_8458), .o(n_14906) );
ms00f80 configuration_wb_init_complete_out_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_init_complete), .o(wbu_wb_init_complete_in) );
ms00f80 configuration_wb_ta1_reg_31__u0 ( .ck(ispd_clk), .d(n_8520), .o(n_14909) );
ms00f80 configuration_wb_ta2_reg_31__u0 ( .ck(ispd_clk), .d(n_8516), .o(n_14908) );
na02f80 g10_u0 ( .a(wbs_cti_i_0_), .b(wbs_cti_i_2_), .o(n_16963) );
na02f20 g13_u0 ( .a(parchk_pci_cbe_reg_in_1238), .b(parchk_pci_cbe_reg_in_1236), .o(n_15958) );
in01f06 g14_u0 ( .a(n_15959), .o(n_15960) );
na02f40 g15_u0 ( .a(parchk_pci_cbe_reg_in), .b(parchk_pci_cbe_reg_in_1237), .o(g15_p) );
in01f10 g15_u1 ( .a(g15_p), .o(n_15959) );
in01f40 g16_u0 ( .a(parchk_pci_cbe_reg_in_1238), .o(n_1061) );
na02f02 g17_u0 ( .a(wishbone_slave_unit_pcim_sm_rdy_in), .b(n_15262), .o(g17_p) );
in01f02 g17_u1 ( .a(g17_p), .o(n_15054) );
na02s01 TIMEBOOST_cell_42696 ( .a(TIMEBOOST_net_13586), .b(g58440_sb), .o(TIMEBOOST_net_10971) );
no02f10 g20_u0 ( .a(n_15999), .b(n_15998), .o(n_16001) );
na02s01 TIMEBOOST_cell_31689 ( .a(TIMEBOOST_net_9755), .b(FE_OFN262_n_9851), .o(n_9852) );
in01f02 g21_u0 ( .a(n_16577), .o(n_16578) );
no02f10 g22_u0 ( .a(n_1323), .b(n_15371), .o(g22_p) );
in01f08 g22_u1 ( .a(g22_p), .o(n_15055) );
na02f04 g23_dup_u0 ( .a(n_16487), .b(n_16089), .o(n_16576) );
in01s08 g23_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_1_), .o(n_16071) );
no02f08 g25_u0 ( .a(FE_OCPN1852_n_16538), .b(n_15210), .o(n_15065) );
no02f08 g27_u0 ( .a(n_15924), .b(n_15998), .o(n_15231) );
na02f06 g28_dup74417_u0 ( .a(n_15746), .b(n_15924), .o(n_15748) );
no02f02 g28_dup_u0 ( .a(n_15403), .b(n_15397), .o(n_15512) );
ao22f06 g31_u0 ( .a(configuration_pci_err_data_510), .b(FE_OFN1063_n_15808), .c(n_16810), .d(n_14912), .o(n_15813) );
na03s02 TIMEBOOST_cell_33535 ( .a(pci_target_unit_del_sync_bc_in), .b(g65215_sb), .c(g65239_db), .o(n_2644) );
no02f20 g33_u0 ( .a(n_16460), .b(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(n_16914) );
na02f10 g34_u0 ( .a(n_370), .b(n_931), .o(n_16021) );
na02m02 TIMEBOOST_cell_32364 ( .a(wbs_wbb3_2_wbb2_dat_o_i_120), .b(wbs_dat_o_21_), .o(TIMEBOOST_net_10093) );
na02m02 TIMEBOOST_cell_32474 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__Q), .o(TIMEBOOST_net_10148) );
na02m04 TIMEBOOST_cell_45822 ( .a(TIMEBOOST_net_15149), .b(FE_OFN2134_n_13124), .o(TIMEBOOST_net_14991) );
na02s03 TIMEBOOST_cell_44771 ( .a(FE_OFN2055_n_8831), .b(g58771_sb), .o(TIMEBOOST_net_14624) );
no02f08 g46_u0 ( .a(n_1177), .b(n_906), .o(n_16154) );
in01f10 g47_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_control_in_86), .o(n_16157) );
oa12s02 g52241_u0 ( .a(n_7740), .b(n_14888), .c(parity_checker_master_perr_report), .o(n_14901) );
na03f02 g52244_u0 ( .a(n_14900), .b(n_14306), .c(n_14902), .o(n_14904) );
na03f02 g52245_u0 ( .a(n_14899), .b(n_14304), .c(n_14902), .o(n_14903) );
ao12s01 g52246_u0 ( .a(parity_checker_pci_perr_en_reg), .b(parity_checker_perr_sampled), .c(n_13766), .o(n_14888) );
no02f02 g52252_u0 ( .a(n_14892), .b(n_14898), .o(g52252_p) );
in01f02 g52252_u1 ( .a(g52252_p), .o(n_14900) );
no02f02 g52253_u0 ( .a(n_14891), .b(n_14898), .o(g52253_p) );
in01f02 g52253_u1 ( .a(g52253_p), .o(n_14899) );
na02m02 TIMEBOOST_cell_43819 ( .a(n_8994), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__Q), .o(TIMEBOOST_net_14148) );
na02s01 TIMEBOOST_cell_16827 ( .a(TIMEBOOST_net_3670), .b(g65062_db), .o(n_3611) );
na02s01 TIMEBOOST_cell_16828 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__Q), .b(g65327_sb), .o(TIMEBOOST_net_3671) );
in01s01 TIMEBOOST_cell_45945 ( .a(wbm_dat_i_30_), .o(TIMEBOOST_net_15252) );
na02s01 TIMEBOOST_cell_16830 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__Q), .b(g65318_sb), .o(TIMEBOOST_net_3672) );
ao12f02 g52353_u0 ( .a(n_14889), .b(n_14890), .c(wbm_cti_o_0_), .o(n_14892) );
ao12f02 g52354_u0 ( .a(n_14889), .b(n_14890), .c(wbm_cti_o_2_), .o(n_14891) );
oa12f02 g52390_u0 ( .a(n_14308), .b(n_14586), .c(n_9178), .o(n_14630) );
no02s01 g52391_u0 ( .a(n_14662), .b(parity_checker_check_perr), .o(n_14765) );
ao12f02 g52392_u0 ( .a(n_14806), .b(n_14764), .c(n_14967), .o(n_14889) );
in01s02 g52393_u0 ( .a(n_8757), .o(g52393_sb) );
na02f06 TIMEBOOST_cell_3855 ( .a(n_15915), .b(TIMEBOOST_net_507), .o(n_16273) );
na02s02 TIMEBOOST_cell_42988 ( .a(TIMEBOOST_net_13732), .b(TIMEBOOST_net_4267), .o(TIMEBOOST_net_4511) );
na02f02 TIMEBOOST_cell_42394 ( .a(TIMEBOOST_net_13435), .b(g57058_sb), .o(n_11679) );
in01s02 g52394_u0 ( .a(n_8757), .o(g52394_sb) );
na02s01 TIMEBOOST_cell_42734 ( .a(TIMEBOOST_net_13605), .b(FE_OFN717_n_8176), .o(TIMEBOOST_net_11103) );
na03s02 TIMEBOOST_cell_6301 ( .a(FE_OFN231_n_9839), .b(g58215_sb), .c(g58215_db), .o(n_9571) );
in01s01 TIMEBOOST_cell_45915 ( .a(wbm_dat_i_17_), .o(TIMEBOOST_net_15222) );
in01s02 g52395_u0 ( .a(n_14839), .o(g52395_sb) );
na02s02 TIMEBOOST_cell_37942 ( .a(TIMEBOOST_net_11209), .b(g58179_sb), .o(n_9608) );
na02s02 TIMEBOOST_cell_38441 ( .a(FE_OFN201_n_9230), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__Q), .o(TIMEBOOST_net_11459) );
na02s02 TIMEBOOST_cell_19297 ( .a(TIMEBOOST_net_4905), .b(g60655_sb), .o(n_5668) );
in01s02 g52396_u0 ( .a(n_8757), .o(g52396_sb) );
na02s01 TIMEBOOST_cell_16064 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__Q), .b(g65860_sb), .o(TIMEBOOST_net_3289) );
na02m02 TIMEBOOST_cell_43343 ( .a(TIMEBOOST_net_9971), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_13910) );
na02s01 TIMEBOOST_cell_15835 ( .a(TIMEBOOST_net_3174), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_407), .o(TIMEBOOST_net_69) );
in01s02 g52397_u0 ( .a(n_14839), .o(g52397_sb) );
na02f06 TIMEBOOST_cell_36888 ( .a(TIMEBOOST_net_10682), .b(n_8489), .o(n_8567) );
na02s02 g52397_u2 ( .a(n_14755), .b(n_14839), .o(g52397_db) );
na02s01 TIMEBOOST_cell_40436 ( .a(TIMEBOOST_net_12456), .b(g62123_sb), .o(n_5573) );
in01m01 g52398_u0 ( .a(n_14839), .o(g52398_sb) );
na02f02 TIMEBOOST_cell_3861 ( .a(TIMEBOOST_net_510), .b(n_3438), .o(n_4877) );
na02s02 g52398_u2 ( .a(n_14753), .b(n_14839), .o(g52398_db) );
na02s02 TIMEBOOST_cell_38108 ( .a(TIMEBOOST_net_11292), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_4516) );
in01s02 g52399_u0 ( .a(n_8757), .o(g52399_sb) );
na02s01 TIMEBOOST_cell_39218 ( .a(TIMEBOOST_net_11847), .b(n_1655), .o(TIMEBOOST_net_11476) );
na02s02 g52399_u2 ( .a(n_14751), .b(n_8757), .o(g52399_db) );
na02s01 TIMEBOOST_cell_45602 ( .a(TIMEBOOST_net_15039), .b(g65215_sb), .o(n_2653) );
in01m02 g52400_u0 ( .a(n_14839), .o(g52400_sb) );
na02f02 TIMEBOOST_cell_41560 ( .a(TIMEBOOST_net_13018), .b(g57406_sb), .o(n_10828) );
na02s06 g52400_u2 ( .a(n_14749), .b(n_14839), .o(g52400_db) );
na02f02 TIMEBOOST_cell_43781 ( .a(TIMEBOOST_net_10046), .b(g57290_sb), .o(TIMEBOOST_net_14129) );
in01s02 g52401_u0 ( .a(n_8757), .o(g52401_sb) );
na02m02 TIMEBOOST_cell_4001 ( .a(TIMEBOOST_net_580), .b(n_8596), .o(n_8680) );
na02f02 TIMEBOOST_cell_41671 ( .a(TIMEBOOST_net_10134), .b(FE_OFN1769_n_14054), .o(TIMEBOOST_net_13074) );
na02s01 TIMEBOOST_cell_18463 ( .a(TIMEBOOST_net_4488), .b(g62863_sb), .o(n_5240) );
in01m01 g52402_u0 ( .a(n_14837), .o(g52402_sb) );
na02m02 TIMEBOOST_cell_36739 ( .a(g52402_sb), .b(g52643_da), .o(TIMEBOOST_net_10608) );
na02s01 TIMEBOOST_cell_36492 ( .a(TIMEBOOST_net_10484), .b(g66398_sb), .o(n_2527) );
na02s01 TIMEBOOST_cell_38648 ( .a(TIMEBOOST_net_11562), .b(g62777_db), .o(n_5438) );
in01m02 g52403_u0 ( .a(n_8757), .o(g52403_sb) );
na02f02 TIMEBOOST_cell_4111 ( .a(TIMEBOOST_net_635), .b(n_16167), .o(n_12956) );
na02m02 g52403_u2 ( .a(n_14744), .b(n_8757), .o(g52403_db) );
na02f01 TIMEBOOST_cell_4112 ( .a(n_14967), .b(pci_target_unit_wbm_sm_pciw_fifo_control_in_84), .o(TIMEBOOST_net_636) );
in01s02 g52404_u0 ( .a(n_14839), .o(g52404_sb) );
na02s02 TIMEBOOST_cell_37924 ( .a(TIMEBOOST_net_11200), .b(g58421_sb), .o(n_9426) );
na02s02 TIMEBOOST_cell_38110 ( .a(TIMEBOOST_net_11293), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_4587) );
na02s01 TIMEBOOST_cell_44894 ( .a(TIMEBOOST_net_14685), .b(g58055_sb), .o(TIMEBOOST_net_12428) );
in01m02 g52405_u0 ( .a(n_14839), .o(g52405_sb) );
na02f08 TIMEBOOST_cell_3987 ( .a(TIMEBOOST_net_573), .b(g54131_da), .o(n_13679) );
na02s01 TIMEBOOST_cell_37790 ( .a(TIMEBOOST_net_11133), .b(g64078_sb), .o(TIMEBOOST_net_469) );
na02s01 TIMEBOOST_cell_39169 ( .a(TIMEBOOST_net_1102), .b(FE_OFN945_n_2248), .o(TIMEBOOST_net_11823) );
oa12m02 g52406_u0 ( .a(n_13398), .b(n_14802), .c(FE_OFN2163_n_16301), .o(n_14887) );
oa12m02 g52408_u0 ( .a(n_13395), .b(n_14799), .c(FE_OFN2165_n_16301), .o(n_14885) );
oa12m02 g52409_u0 ( .a(n_13394), .b(n_14798), .c(FE_OFN2165_n_16301), .o(n_14884) );
oa12m02 g52410_u0 ( .a(n_13393), .b(n_14797), .c(FE_OFN2165_n_16301), .o(n_14883) );
oa12m02 g52411_u0 ( .a(n_13392), .b(n_14796), .c(FE_OFN2165_n_16301), .o(n_14881) );
oa12m02 g52412_u0 ( .a(n_13391), .b(n_14763), .c(n_16305), .o(n_14851) );
oa12m02 g52413_u0 ( .a(n_13389), .b(n_14793), .c(FE_OFN2165_n_16301), .o(n_14880) );
oa12m02 g52414_u0 ( .a(n_13390), .b(n_14794), .c(FE_OFN2165_n_16301), .o(n_14879) );
oa12m02 g52415_u0 ( .a(n_13388), .b(n_14762), .c(FE_OFN2165_n_16301), .o(n_14850) );
oa12m02 g52416_u0 ( .a(n_13387), .b(n_14792), .c(FE_OFN2165_n_16301), .o(n_14877) );
oa12m02 g52417_u0 ( .a(n_13386), .b(n_14791), .c(FE_OFN2163_n_16301), .o(n_14875) );
oa12m02 g52418_u0 ( .a(n_13384), .b(n_14790), .c(FE_OFN2165_n_16301), .o(n_14873) );
oa12m02 g52419_u0 ( .a(n_13383), .b(n_14789), .c(FE_OFN2165_n_16301), .o(n_14871) );
oa12m02 g52421_u0 ( .a(n_13381), .b(n_14786), .c(FE_OFN2165_n_16301), .o(n_14869) );
oa12m02 g52422_u0 ( .a(n_13380), .b(n_14784), .c(FE_OFN2162_n_16301), .o(n_14867) );
oa12m02 g52423_u0 ( .a(n_13379), .b(n_14783), .c(FE_OFN2162_n_16301), .o(n_14866) );
oa12m02 g52424_u0 ( .a(n_13378), .b(n_14781), .c(FE_OFN2164_n_16301), .o(n_14865) );
oa12m02 g52425_u0 ( .a(n_13376), .b(n_14778), .c(FE_OFN2162_n_16301), .o(n_14864) );
oa12m02 g52426_u0 ( .a(n_13377), .b(n_14780), .c(FE_OFN2164_n_16301), .o(n_14863) );
oa12m02 g52427_u0 ( .a(n_13375), .b(n_14777), .c(FE_OFN2162_n_16301), .o(n_14862) );
oa12m02 g52428_u0 ( .a(n_13374), .b(n_14776), .c(FE_OFN2162_n_16301), .o(n_14861) );
oa12m02 g52429_u0 ( .a(n_13373), .b(n_14775), .c(FE_OFN2162_n_16301), .o(n_14860) );
oa12m02 g52430_u0 ( .a(n_13371), .b(n_14772), .c(FE_OFN2163_n_16301), .o(n_14859) );
oa12m02 g52431_u0 ( .a(n_13370), .b(n_14770), .c(n_16305), .o(n_14858) );
oa12m02 g52432_u0 ( .a(n_13372), .b(n_14773), .c(n_16305), .o(n_14856) );
oa12m02 g52433_u0 ( .a(n_13369), .b(n_14769), .c(n_16305), .o(n_14855) );
oa12m02 g52434_u0 ( .a(n_13368), .b(n_14768), .c(FE_OFN2163_n_16301), .o(n_14854) );
oa12m02 g52435_u0 ( .a(n_13367), .b(n_14761), .c(FE_OFN2164_n_16301), .o(n_14849) );
oa12m02 g52436_u0 ( .a(n_13366), .b(n_14767), .c(FE_OFN2164_n_16301), .o(n_14853) );
oa12m02 g52437_u0 ( .a(n_13365), .b(n_14766), .c(FE_OFN2164_n_16301), .o(n_14852) );
na02m04 TIMEBOOST_cell_3853 ( .a(TIMEBOOST_net_506), .b(n_3130), .o(n_3141) );
na02f02 TIMEBOOST_cell_44236 ( .a(TIMEBOOST_net_14356), .b(FE_OFN1382_n_8567), .o(TIMEBOOST_net_12740) );
na02f04 TIMEBOOST_cell_3854 ( .a(n_16524), .b(FE_OCPN1823_n_16560), .o(TIMEBOOST_net_507) );
in01m01 g52440_u0 ( .a(n_14839), .o(g52440_sb) );
na02s02 TIMEBOOST_cell_38112 ( .a(TIMEBOOST_net_11294), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_4488) );
na02m02 g52440_u2 ( .a(n_14681), .b(n_14839), .o(g52440_db) );
na02s02 TIMEBOOST_cell_38114 ( .a(TIMEBOOST_net_11295), .b(FE_OFN1135_g64577_p), .o(TIMEBOOST_net_4586) );
in01s01 g52441_u0 ( .a(n_14839), .o(g52441_sb) );
na02s02 TIMEBOOST_cell_37944 ( .a(TIMEBOOST_net_11210), .b(g58019_sb), .o(n_9771) );
na03s02 TIMEBOOST_cell_38219 ( .a(g64196_da), .b(g64196_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__Q), .o(TIMEBOOST_net_11348) );
na02s02 TIMEBOOST_cell_37890 ( .a(TIMEBOOST_net_11183), .b(g58041_sb), .o(n_9747) );
in01s02 g52442_u0 ( .a(n_8757), .o(g52442_sb) );
na02s01 TIMEBOOST_cell_18629 ( .a(TIMEBOOST_net_4571), .b(g63106_sb), .o(n_5042) );
na02s02 TIMEBOOST_cell_37858 ( .a(TIMEBOOST_net_11167), .b(g58018_sb), .o(n_9773) );
na02s02 TIMEBOOST_cell_18657 ( .a(TIMEBOOST_net_4585), .b(g63074_sb), .o(n_5102) );
in01s02 g52443_u0 ( .a(n_8757), .o(g52443_sb) );
na02m02 TIMEBOOST_cell_19126 ( .a(wbm_adr_o_14_), .b(FE_OFN1700_n_5751), .o(TIMEBOOST_net_4820) );
na02s01 TIMEBOOST_cell_37577 ( .a(parchk_pci_ad_reg_in_1232), .b(g65893_sb), .o(TIMEBOOST_net_11027) );
na02s02 TIMEBOOST_cell_19291 ( .a(TIMEBOOST_net_4902), .b(g60651_sb), .o(n_5673) );
in01m01 g52444_u0 ( .a(n_14839), .o(g52444_sb) );
na02s02 TIMEBOOST_cell_19124 ( .a(wbm_adr_o_15_), .b(FE_OFN1700_n_5751), .o(TIMEBOOST_net_4819) );
na03s02 TIMEBOOST_cell_38331 ( .a(n_3874), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q), .c(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_11404) );
na02s02 TIMEBOOST_cell_19293 ( .a(TIMEBOOST_net_4903), .b(g60653_sb), .o(n_5670) );
na02f02 TIMEBOOST_cell_42240 ( .a(TIMEBOOST_net_13358), .b(FE_OFN1394_n_8567), .o(TIMEBOOST_net_12315) );
na02f01 g52445_u2 ( .a(n_14678), .b(n_14837), .o(g52445_db) );
na02s01 TIMEBOOST_cell_37688 ( .a(TIMEBOOST_net_11082), .b(g61908_sb), .o(n_8005) );
in01s02 g52446_u0 ( .a(n_8757), .o(g52446_sb) );
na02s01 TIMEBOOST_cell_43397 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__Q), .b(n_4315), .o(TIMEBOOST_net_13937) );
na02s01 TIMEBOOST_cell_38000 ( .a(TIMEBOOST_net_11238), .b(g61873_sb), .o(n_8087) );
na02s02 TIMEBOOST_cell_40876 ( .a(TIMEBOOST_net_12676), .b(g62427_sb), .o(n_7386) );
in01m02 g52447_u0 ( .a(n_14839), .o(g52447_sb) );
na02s01 TIMEBOOST_cell_18294 ( .a(g61923_sb), .b(g61987_db), .o(TIMEBOOST_net_4404) );
na02s01 TIMEBOOST_cell_39370 ( .a(TIMEBOOST_net_11923), .b(g65884_sb), .o(n_1863) );
na02s01 TIMEBOOST_cell_37690 ( .a(TIMEBOOST_net_11083), .b(g61919_sb), .o(n_7983) );
in01s01 g52448_u0 ( .a(n_14839), .o(g52448_sb) );
na02m04 TIMEBOOST_cell_2901 ( .a(n_521), .b(TIMEBOOST_net_30), .o(n_1639) );
na02m02 g52448_u2 ( .a(n_14746), .b(n_14839), .o(g52448_db) );
na02s02 TIMEBOOST_cell_43153 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__14__Q), .b(n_4486), .o(TIMEBOOST_net_13815) );
in01s01 g52449_u0 ( .a(n_14839), .o(g52449_sb) );
na02f02 TIMEBOOST_cell_43820 ( .a(TIMEBOOST_net_14148), .b(FE_OFN1412_n_8567), .o(TIMEBOOST_net_12844) );
na02m02 g52449_u2 ( .a(n_14741), .b(n_14839), .o(g52449_db) );
in01f02 TIMEBOOST_cell_15783 ( .a(TIMEBOOST_net_3148), .o(TIMEBOOST_net_3147) );
in01s01 g52450_u0 ( .a(n_14839), .o(g52450_sb) );
na02m02 TIMEBOOST_cell_44503 ( .a(n_9419), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__Q), .o(TIMEBOOST_net_14490) );
na02m02 g52450_u2 ( .a(n_14740), .b(n_14839), .o(g52450_db) );
na02m02 TIMEBOOST_cell_43655 ( .a(n_4678), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__Q), .o(TIMEBOOST_net_14066) );
in01s01 g52451_u0 ( .a(n_14839), .o(g52451_sb) );
na02s02 TIMEBOOST_cell_37866 ( .a(TIMEBOOST_net_11171), .b(g57910_sb), .o(n_9903) );
na02s02 g52451_u2 ( .a(n_14738), .b(n_14839), .o(g52451_db) );
na03s02 TIMEBOOST_cell_38139 ( .a(TIMEBOOST_net_4027), .b(g64326_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__Q), .o(TIMEBOOST_net_11308) );
in01s01 g52452_u0 ( .a(n_14839), .o(g52452_sb) );
na02s02 TIMEBOOST_cell_43154 ( .a(TIMEBOOST_net_13815), .b(FE_OFN1295_n_4098), .o(TIMEBOOST_net_12558) );
na02s02 TIMEBOOST_cell_37798 ( .a(TIMEBOOST_net_11137), .b(g61942_sb), .o(n_7939) );
na02s02 TIMEBOOST_cell_45135 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__Q), .b(n_3981), .o(TIMEBOOST_net_14806) );
na02m04 TIMEBOOST_cell_3859 ( .a(TIMEBOOST_net_509), .b(n_3221), .o(n_7818) );
na02s01 TIMEBOOST_cell_36494 ( .a(TIMEBOOST_net_10485), .b(g66398_sb), .o(n_2508) );
in01s01 TIMEBOOST_cell_32832 ( .a(TIMEBOOST_net_10333), .o(wbs_dat_i_13_) );
in01s01 g52454_u0 ( .a(n_14839), .o(g52454_sb) );
na02s02 TIMEBOOST_cell_37946 ( .a(TIMEBOOST_net_11211), .b(g58321_sb), .o(n_9492) );
na02m02 g52454_u2 ( .a(n_14734), .b(n_14839), .o(g52454_db) );
na02s02 TIMEBOOST_cell_37892 ( .a(TIMEBOOST_net_11184), .b(g58170_sb), .o(n_9621) );
in01m01 g52455_u0 ( .a(n_8757), .o(g52455_sb) );
in01s01 TIMEBOOST_cell_45890 ( .a(TIMEBOOST_net_15196), .o(TIMEBOOST_net_15197) );
na02m02 g52455_u2 ( .a(n_14733), .b(n_8757), .o(g52455_db) );
na02s02 TIMEBOOST_cell_19285 ( .a(TIMEBOOST_net_4899), .b(g60644_sb), .o(n_5684) );
in01s02 g52456_u0 ( .a(FE_OFN1021_n_11877), .o(g52456_sb) );
na02s01 g52456_u1 ( .a(wbs_adr_i_10_), .b(g52456_sb), .o(g52456_da) );
in01s01 TIMEBOOST_cell_45865 ( .a(TIMEBOOST_net_15172), .o(wishbone_slave_unit_del_sync_sync_req_comp_pending) );
na02f02 TIMEBOOST_cell_44504 ( .a(TIMEBOOST_net_14490), .b(FE_OFN2180_n_8567), .o(TIMEBOOST_net_13451) );
in01m02 g52457_u0 ( .a(FE_OFN1022_n_11877), .o(g52457_sb) );
na02s01 g52457_u1 ( .a(wbs_adr_i_11_), .b(g52457_sb), .o(g52457_da) );
na02m02 TIMEBOOST_cell_43821 ( .a(n_9896), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__Q), .o(TIMEBOOST_net_14149) );
na02f02 TIMEBOOST_cell_43822 ( .a(TIMEBOOST_net_14149), .b(FE_OFN1420_n_8567), .o(TIMEBOOST_net_12931) );
in01m02 g52458_u0 ( .a(FE_OFN1022_n_11877), .o(g52458_sb) );
na02s01 g52458_u1 ( .a(wbs_adr_i_12_), .b(g52458_sb), .o(g52458_da) );
na02s01 TIMEBOOST_cell_30971 ( .a(TIMEBOOST_net_9396), .b(g64938_db), .o(n_3676) );
na02m02 TIMEBOOST_cell_43823 ( .a(n_9139), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__Q), .o(TIMEBOOST_net_14150) );
in01m02 g52459_u0 ( .a(FE_OFN1022_n_11877), .o(g52459_sb) );
na02s01 TIMEBOOST_cell_18002 ( .a(pci_target_unit_fifos_pciw_cbe_in), .b(g64111_sb), .o(TIMEBOOST_net_4258) );
na02f02 TIMEBOOST_cell_42396 ( .a(TIMEBOOST_net_13436), .b(g57468_sb), .o(n_11264) );
na02s02 TIMEBOOST_cell_45603 ( .a(TIMEBOOST_net_9362), .b(FE_OFN789_n_2678), .o(TIMEBOOST_net_15040) );
in01s02 g52460_u0 ( .a(FE_OFN1021_n_11877), .o(g52460_sb) );
na02s01 g52460_u1 ( .a(wbs_adr_i_15_), .b(g52460_sb), .o(g52460_da) );
na02f02 TIMEBOOST_cell_42398 ( .a(TIMEBOOST_net_13437), .b(g57055_sb), .o(n_11681) );
na02s01 TIMEBOOST_cell_43531 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__Q), .b(n_4349), .o(TIMEBOOST_net_14004) );
in01m02 g52461_u0 ( .a(FE_OFN1022_n_11877), .o(g52461_sb) );
na02s01 g52461_u1 ( .a(wbs_adr_i_14_), .b(g52461_sb), .o(g52461_da) );
na02s01 TIMEBOOST_cell_30969 ( .a(TIMEBOOST_net_9395), .b(g64936_sb), .o(n_3677) );
na02s02 TIMEBOOST_cell_30970 ( .a(n_3780), .b(g64938_sb), .o(TIMEBOOST_net_9396) );
in01m02 g52462_u0 ( .a(FE_OFN1022_n_11877), .o(g52462_sb) );
na02s01 TIMEBOOST_cell_44895 ( .a(g65721_db), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__Q), .o(TIMEBOOST_net_14686) );
na02f02 TIMEBOOST_cell_41380 ( .a(TIMEBOOST_net_12928), .b(g57476_sb), .o(n_10336) );
na02f02 TIMEBOOST_cell_44129 ( .a(n_9824), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__Q), .o(TIMEBOOST_net_14303) );
in01m02 g52463_u0 ( .a(FE_OFN1022_n_11877), .o(g52463_sb) );
na02s01 g52463_u1 ( .a(wbs_adr_i_17_), .b(g52463_sb), .o(g52463_da) );
na02s01 TIMEBOOST_cell_30978 ( .a(pci_target_unit_fifos_pcir_data_in_164), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__Q), .o(TIMEBOOST_net_9400) );
na02s02 TIMEBOOST_cell_42121 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__Q), .b(n_3623), .o(TIMEBOOST_net_13299) );
in01s02 g52464_u0 ( .a(FE_OFN1021_n_11877), .o(g52464_sb) );
na02s01 g52464_u1 ( .a(wbs_adr_i_18_), .b(g52464_sb), .o(g52464_da) );
na02s02 TIMEBOOST_cell_42122 ( .a(TIMEBOOST_net_13299), .b(FE_OFN1314_n_6624), .o(TIMEBOOST_net_11592) );
na02s01 TIMEBOOST_cell_30920 ( .a(pci_target_unit_pcit_if_strd_addr_in_703), .b(pci_target_unit_del_sync_addr_in_221), .o(TIMEBOOST_net_9371) );
na02s01 g52465_u1 ( .a(wbs_adr_i_19_), .b(g52461_sb), .o(g52465_da) );
na02s02 TIMEBOOST_cell_45240 ( .a(TIMEBOOST_net_14858), .b(FE_OFN1268_n_4095), .o(TIMEBOOST_net_12116) );
na02s01 TIMEBOOST_cell_45241 ( .a(n_75), .b(n_3727), .o(TIMEBOOST_net_14859) );
in01s02 g52466_u0 ( .a(FE_OFN1021_n_11877), .o(g52466_sb) );
na02s01 g52466_u1 ( .a(wbs_adr_i_20_), .b(g52466_sb), .o(g52466_da) );
na02f04 TIMEBOOST_cell_44707 ( .a(wbu_addr_in_267), .b(g52602_sb), .o(TIMEBOOST_net_14592) );
na02f02 TIMEBOOST_cell_36992 ( .a(TIMEBOOST_net_10734), .b(g58830_sb), .o(n_8607) );
na02s01 g52467_u1 ( .a(wbs_adr_i_21_), .b(g52457_sb), .o(g52467_da) );
na02f02 TIMEBOOST_cell_22599 ( .a(TIMEBOOST_net_6556), .b(FE_OFN1577_n_12028), .o(n_12599) );
na02m02 TIMEBOOST_cell_43656 ( .a(TIMEBOOST_net_14066), .b(FE_OFN1316_n_6624), .o(TIMEBOOST_net_12256) );
na02s01 TIMEBOOST_cell_44896 ( .a(TIMEBOOST_net_14686), .b(g65721_da), .o(TIMEBOOST_net_10974) );
na02f02 TIMEBOOST_cell_44272 ( .a(TIMEBOOST_net_14374), .b(FE_OFN1416_n_8567), .o(TIMEBOOST_net_12837) );
na02s01 TIMEBOOST_cell_39220 ( .a(TIMEBOOST_net_11848), .b(n_1934), .o(TIMEBOOST_net_10938) );
na02s01 g52469_u1 ( .a(wbs_adr_i_23_), .b(g52458_sb), .o(g52469_da) );
na03f04 TIMEBOOST_cell_22362 ( .a(n_10931), .b(n_10661), .c(n_10660), .o(TIMEBOOST_net_6438) );
na02s01 TIMEBOOST_cell_31018 ( .a(n_4444), .b(g64836_sb), .o(TIMEBOOST_net_9420) );
in01m04 g52470_u0 ( .a(FE_OFN1023_n_11877), .o(g52470_sb) );
na02s01 g52470_u1 ( .a(wbs_adr_i_24_), .b(g52470_sb), .o(g52470_da) );
na02s01 TIMEBOOST_cell_31017 ( .a(TIMEBOOST_net_9419), .b(g64828_db), .o(n_4453) );
na02s02 TIMEBOOST_cell_31016 ( .a(n_4452), .b(g64828_sb), .o(TIMEBOOST_net_9419) );
na02s01 g52471_u1 ( .a(wbs_adr_i_25_), .b(g52459_sb), .o(g52471_da) );
na02f02 TIMEBOOST_cell_22601 ( .a(TIMEBOOST_net_6557), .b(FE_OFN1566_n_12502), .o(n_12488) );
na02s02 TIMEBOOST_cell_42670 ( .a(TIMEBOOST_net_13573), .b(g64189_da), .o(TIMEBOOST_net_11303) );
na02s01 g52472_u1 ( .a(wbs_adr_i_26_), .b(g52458_sb), .o(g52472_da) );
na02s01 TIMEBOOST_cell_45604 ( .a(TIMEBOOST_net_15040), .b(g65238_sb), .o(n_2645) );
na02f02 TIMEBOOST_cell_42400 ( .a(TIMEBOOST_net_13438), .b(g57588_sb), .o(n_11164) );
na02s01 g52473_u1 ( .a(wbs_adr_i_27_), .b(g52457_sb), .o(g52473_da) );
na02f02 TIMEBOOST_cell_22603 ( .a(TIMEBOOST_net_6558), .b(FE_OFN1565_n_12502), .o(n_12620) );
na03s02 TIMEBOOST_cell_43339 ( .a(n_3526), .b(FE_OFN1193_n_6935), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__30__Q), .o(TIMEBOOST_net_13908) );
na02s01 g52474_u1 ( .a(wbs_adr_i_28_), .b(g52462_sb), .o(g52474_da) );
na02f02 TIMEBOOST_cell_22605 ( .a(TIMEBOOST_net_6559), .b(FE_OFN1564_n_12502), .o(n_12643) );
na02s02 TIMEBOOST_cell_43155 ( .a(n_3596), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__Q), .o(TIMEBOOST_net_13816) );
na03f02 TIMEBOOST_cell_36198 ( .a(FE_OCP_RBN1973_n_12381), .b(TIMEBOOST_net_10297), .c(n_11831), .o(n_12703) );
na02f02 TIMEBOOST_cell_22487 ( .a(TIMEBOOST_net_6500), .b(FE_OFN1581_n_12306), .o(n_12498) );
na02s02 TIMEBOOST_cell_43657 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__Q), .b(n_3700), .o(TIMEBOOST_net_14067) );
in01s02 g52476_u0 ( .a(FE_OFN1021_n_11877), .o(g52476_sb) );
na02s01 g52476_u1 ( .a(wbs_adr_i_30_), .b(g52476_sb), .o(g52476_da) );
na02s02 TIMEBOOST_cell_42123 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__Q), .b(n_3737), .o(TIMEBOOST_net_13300) );
na02s01 TIMEBOOST_cell_43035 ( .a(FE_OFN201_n_9230), .b(g57906_sb), .o(TIMEBOOST_net_13756) );
in01m02 g52477_u0 ( .a(FE_OFN1025_n_11877), .o(g52477_sb) );
na02s01 g52477_u1 ( .a(wbs_adr_i_29_), .b(g52477_sb), .o(g52477_da) );
na03s02 TIMEBOOST_cell_5685 ( .a(n_4442), .b(g64925_sb), .c(g64925_db), .o(n_4390) );
na02f02 TIMEBOOST_cell_22607 ( .a(TIMEBOOST_net_6560), .b(FE_OFN1564_n_12502), .o(n_12648) );
in01s02 g52478_u0 ( .a(FE_OFN8_n_11877), .o(g52478_sb) );
na02s01 g52478_u1 ( .a(wbs_adr_i_31_), .b(g52478_sb), .o(g52478_da) );
na02s02 TIMEBOOST_cell_43156 ( .a(TIMEBOOST_net_13816), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_12560) );
na03s02 TIMEBOOST_cell_5676 ( .a(n_4447), .b(g64861_sb), .c(g64861_db), .o(n_4428) );
in01m02 g52479_u0 ( .a(FE_OFN1024_n_11877), .o(g52479_sb) );
na02s01 g52479_u1 ( .a(wbs_adr_i_3_), .b(g52479_sb), .o(g52479_da) );
na03s01 TIMEBOOST_cell_33787 ( .a(FE_OFN254_n_9825), .b(g58006_sb), .c(g58006_db), .o(n_9788) );
na02m02 TIMEBOOST_cell_44255 ( .a(n_9095), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__Q), .o(TIMEBOOST_net_14366) );
na02s01 g52480_u1 ( .a(wbs_adr_i_4_), .b(g52479_sb), .o(g52480_da) );
na02s02 TIMEBOOST_cell_43060 ( .a(TIMEBOOST_net_13768), .b(FE_OFN1293_n_4098), .o(TIMEBOOST_net_12021) );
na03s02 TIMEBOOST_cell_5456 ( .a(n_4447), .b(g64792_sb), .c(g64792_db), .o(n_4472) );
na02m01 g52481_u1 ( .a(wbs_adr_i_5_), .b(g52479_sb), .o(g52481_da) );
na02m02 TIMEBOOST_cell_44273 ( .a(n_9835), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__Q), .o(TIMEBOOST_net_14375) );
na02s01 TIMEBOOST_cell_17857 ( .a(TIMEBOOST_net_4185), .b(g65356_db), .o(n_3538) );
in01s02 g52482_u0 ( .a(FE_OFN8_n_11877), .o(g52482_sb) );
na02m01 g52482_u1 ( .a(wbs_adr_i_6_), .b(g52482_sb), .o(g52482_da) );
na02s02 TIMEBOOST_cell_31015 ( .a(TIMEBOOST_net_9418), .b(g64818_db), .o(n_4457) );
na02s02 TIMEBOOST_cell_31014 ( .a(n_4482), .b(g64818_sb), .o(TIMEBOOST_net_9418) );
na02s01 g52483_u1 ( .a(wbs_adr_i_7_), .b(g52470_sb), .o(g52483_da) );
na02f02 TIMEBOOST_cell_40892 ( .a(TIMEBOOST_net_12684), .b(FE_OFN1391_n_8567), .o(TIMEBOOST_net_11644) );
na02s01 TIMEBOOST_cell_45242 ( .a(TIMEBOOST_net_14859), .b(FE_OFN1293_n_4098), .o(TIMEBOOST_net_12605) );
na02m01 g52484_u1 ( .a(wbs_adr_i_8_), .b(g52477_sb), .o(g52484_da) );
na02s01 TIMEBOOST_cell_42615 ( .a(FE_OFN245_n_9114), .b(g58003_sb), .o(TIMEBOOST_net_13546) );
na02s02 TIMEBOOST_cell_45605 ( .a(TIMEBOOST_net_9373), .b(FE_OFN789_n_2678), .o(TIMEBOOST_net_15041) );
na02s01 g52485_u1 ( .a(wbs_adr_i_9_), .b(g52470_sb), .o(g52485_da) );
na02s02 TIMEBOOST_cell_31013 ( .a(TIMEBOOST_net_9417), .b(g64812_db), .o(n_4461) );
na02s02 TIMEBOOST_cell_45243 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__Q), .b(n_4350), .o(TIMEBOOST_net_14860) );
na02f02 g52494_u0 ( .a(n_14693), .b(n_14482), .o(n_14806) );
no02f02 g52495_u0 ( .a(n_14760), .b(FE_OFN2163_n_16301), .o(g52495_p) );
in01f02 g52495_u1 ( .a(g52495_p), .o(n_14833) );
no02f02 g52496_u0 ( .a(n_14759), .b(FE_OFN2163_n_16301), .o(g52496_p) );
in01f02 g52496_u1 ( .a(g52496_p), .o(n_14832) );
no02f02 g52497_u0 ( .a(n_14757), .b(FE_OFN2163_n_16301), .o(g52497_p) );
in01f02 g52497_u1 ( .a(g52497_p), .o(n_14830) );
no02f02 g52498_u0 ( .a(n_14756), .b(FE_OFN2163_n_16301), .o(g52498_p) );
in01f02 g52498_u1 ( .a(g52498_p), .o(n_14829) );
oa12f01 g52499_u0 ( .a(n_10793), .b(FE_OFN3_n_4778), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(n_11844) );
na02m02 g52500_u0 ( .a(n_8880), .b(n_14691), .o(n_14804) );
na02m02 g52501_u0 ( .a(n_8879), .b(n_14690), .o(n_14805) );
ao12s01 g52502_u0 ( .a(n_14624), .b(parchk_pci_perr_out_in), .c(out_bckp_perr_en_out), .o(n_14662) );
in01f02 g52503_u0 ( .a(FE_OFN2243_g52675_p), .o(g52503_sb) );
na02s02 TIMEBOOST_cell_31997 ( .a(TIMEBOOST_net_9909), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_4891) );
na02m02 TIMEBOOST_cell_41665 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_8__Q), .o(TIMEBOOST_net_13071) );
na02s02 TIMEBOOST_cell_31012 ( .a(n_4476), .b(g64812_sb), .o(TIMEBOOST_net_9417) );
in01f01 g52504_u0 ( .a(FE_OFN1471_g52675_p), .o(g52504_sb) );
na02s01 TIMEBOOST_cell_31996 ( .a(configuration_pci_err_addr_495), .b(wbm_adr_o_25_), .o(TIMEBOOST_net_9909) );
na02f02 TIMEBOOST_cell_42142 ( .a(TIMEBOOST_net_13309), .b(g57079_sb), .o(n_11663) );
na03s02 TIMEBOOST_cell_5534 ( .a(n_4493), .b(g65072_sb), .c(g65072_db), .o(n_4310) );
in01f02 g52505_u0 ( .a(FE_OFN2243_g52675_p), .o(g52505_sb) );
na02s02 TIMEBOOST_cell_31995 ( .a(TIMEBOOST_net_9908), .b(FE_OFN1179_n_3476), .o(TIMEBOOST_net_4890) );
na02s01 TIMEBOOST_cell_31011 ( .a(TIMEBOOST_net_9416), .b(g64801_db), .o(n_4467) );
na02s02 TIMEBOOST_cell_31010 ( .a(n_4479), .b(g64801_sb), .o(TIMEBOOST_net_9416) );
in01f01 g52506_u0 ( .a(FE_OFN1471_g52675_p), .o(g52506_sb) );
na02s01 TIMEBOOST_cell_31994 ( .a(configuration_pci_err_addr_493), .b(wbm_adr_o_23_), .o(TIMEBOOST_net_9908) );
na02f02 TIMEBOOST_cell_42402 ( .a(TIMEBOOST_net_13439), .b(g57356_sb), .o(n_11391) );
na03s02 TIMEBOOST_cell_5536 ( .a(n_4442), .b(g65078_sb), .c(g65078_db), .o(n_4308) );
in01f02 g52507_u0 ( .a(FE_OFN2243_g52675_p), .o(g52507_sb) );
na02s02 TIMEBOOST_cell_38078 ( .a(TIMEBOOST_net_11277), .b(FE_OFN1135_g64577_p), .o(TIMEBOOST_net_4689) );
na04f04 TIMEBOOST_cell_35714 ( .a(n_9441), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__Q), .c(FE_OFN2187_n_8567), .d(g57532_sb), .o(n_11209) );
in01f02 g52508_u0 ( .a(FE_OFN2242_g52675_p), .o(g52508_sb) );
na02s01 TIMEBOOST_cell_31992 ( .a(configuration_pci_err_addr_497), .b(wbm_adr_o_27_), .o(TIMEBOOST_net_9907) );
na02s02 TIMEBOOST_cell_31007 ( .a(TIMEBOOST_net_9414), .b(n_4447), .o(n_4377) );
na02s02 TIMEBOOST_cell_43658 ( .a(TIMEBOOST_net_14067), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_12257) );
in01f01 g52509_u0 ( .a(FE_OFN1472_g52675_p), .o(g52509_sb) );
na02f02 TIMEBOOST_cell_44124 ( .a(TIMEBOOST_net_14300), .b(FE_OFN1413_n_8567), .o(TIMEBOOST_net_12706) );
na02f02 TIMEBOOST_cell_32361 ( .a(TIMEBOOST_net_10091), .b(g58653_sb), .o(TIMEBOOST_net_6264) );
na02m02 TIMEBOOST_cell_44561 ( .a(n_9203), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__Q), .o(TIMEBOOST_net_14519) );
in01f02 g52510_u0 ( .a(FE_OFN2243_g52675_p), .o(g52510_sb) );
na02s02 TIMEBOOST_cell_31991 ( .a(TIMEBOOST_net_9906), .b(FE_OFN1183_n_3476), .o(TIMEBOOST_net_4888) );
na02s01 TIMEBOOST_cell_31006 ( .a(g64953_sb), .b(g64953_db), .o(TIMEBOOST_net_9414) );
na02s01 TIMEBOOST_cell_31005 ( .a(TIMEBOOST_net_9413), .b(g65073_db), .o(n_4309) );
in01f02 g52511_u0 ( .a(FE_OFN2243_g52675_p), .o(g52511_sb) );
na02s01 TIMEBOOST_cell_31990 ( .a(configuration_pci_err_data_503), .b(wbm_dat_o_2_), .o(TIMEBOOST_net_9906) );
na02s01 TIMEBOOST_cell_31004 ( .a(n_4476), .b(g65073_sb), .o(TIMEBOOST_net_9413) );
na02s01 TIMEBOOST_cell_43121 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__Q), .b(n_3571), .o(TIMEBOOST_net_13799) );
in01f02 g52512_u0 ( .a(FE_OFN2243_g52675_p), .o(g52512_sb) );
na02s02 TIMEBOOST_cell_31989 ( .a(TIMEBOOST_net_9905), .b(FE_OFN1185_n_3476), .o(TIMEBOOST_net_4887) );
na02f02 TIMEBOOST_cell_22611 ( .a(TIMEBOOST_net_6562), .b(FE_OFN1566_n_12502), .o(n_12525) );
no02f08 TIMEBOOST_cell_15784 ( .a(conf_wb_err_bc_in), .b(conf_wb_err_bc_in_846), .o(TIMEBOOST_net_3149) );
in01f02 g52513_u0 ( .a(FE_OFN2243_g52675_p), .o(g52513_sb) );
na02s01 TIMEBOOST_cell_31988 ( .a(configuration_pci_err_addr_485), .b(wbm_adr_o_15_), .o(TIMEBOOST_net_9905) );
na02s01 TIMEBOOST_cell_31003 ( .a(TIMEBOOST_net_9412), .b(g65071_db), .o(n_4311) );
na02s02 TIMEBOOST_cell_31002 ( .a(n_4476), .b(g65071_sb), .o(TIMEBOOST_net_9412) );
in01f02 g52514_u0 ( .a(FE_OFN2243_g52675_p), .o(g52514_sb) );
na02s02 TIMEBOOST_cell_31987 ( .a(TIMEBOOST_net_9904), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_4885) );
na02f02 TIMEBOOST_cell_40887 ( .a(n_9471), .b(g57489_sb), .o(TIMEBOOST_net_12682) );
na02s01 TIMEBOOST_cell_31001 ( .a(TIMEBOOST_net_9411), .b(g64790_db), .o(n_4475) );
in01f01 g52515_u0 ( .a(FE_OFN1472_g52675_p), .o(g52515_sb) );
na02s02 TIMEBOOST_cell_42671 ( .a(n_4488), .b(n_4677), .o(TIMEBOOST_net_13574) );
na02s02 TIMEBOOST_cell_43157 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__Q), .b(n_3599), .o(TIMEBOOST_net_13817) );
na02s01 TIMEBOOST_cell_15786 ( .a(parchk_pci_ad_reg_in_1212), .b(g67043_db), .o(TIMEBOOST_net_3150) );
in01f02 g52516_u0 ( .a(FE_OFN2243_g52675_p), .o(g52516_sb) );
na02s02 TIMEBOOST_cell_45244 ( .a(TIMEBOOST_net_14860), .b(FE_OFN1293_n_4098), .o(TIMEBOOST_net_12120) );
na02f02 TIMEBOOST_cell_32359 ( .a(TIMEBOOST_net_10090), .b(g58652_sb), .o(TIMEBOOST_net_6262) );
na02s02 TIMEBOOST_cell_43158 ( .a(TIMEBOOST_net_13817), .b(FE_OFN1288_n_4098), .o(TIMEBOOST_net_12562) );
in01f01 g52517_u0 ( .a(FE_OFN1472_g52675_p), .o(g52517_sb) );
na02s02 TIMEBOOST_cell_43159 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__Q), .b(n_3789), .o(TIMEBOOST_net_13818) );
na02s02 TIMEBOOST_cell_43659 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__Q), .b(n_3706), .o(TIMEBOOST_net_14068) );
na02s02 TIMEBOOST_cell_31000 ( .a(n_4498), .b(g64790_sb), .o(TIMEBOOST_net_9411) );
in01f02 g52518_u0 ( .a(FE_OFN2241_g52675_p), .o(g52518_sb) );
na02s01 TIMEBOOST_cell_31986 ( .a(configuration_pci_err_data_532), .b(wbm_dat_o_31_), .o(TIMEBOOST_net_9904) );
na02s01 TIMEBOOST_cell_30999 ( .a(TIMEBOOST_net_9410), .b(g64758_db), .o(n_4496) );
na02s01 TIMEBOOST_cell_30998 ( .a(n_4482), .b(g64758_sb), .o(TIMEBOOST_net_9410) );
in01f01 g52519_u0 ( .a(FE_OFN1471_g52675_p), .o(g52519_sb) );
na02s02 TIMEBOOST_cell_31985 ( .a(TIMEBOOST_net_9903), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4884) );
na03s02 TIMEBOOST_cell_5537 ( .a(n_4645), .b(g65080_sb), .c(g65080_db), .o(n_4307) );
na03s02 TIMEBOOST_cell_5538 ( .a(n_4488), .b(g65082_sb), .c(g65082_db), .o(n_4305) );
in01f02 g52520_u0 ( .a(FE_OFN2242_g52675_p), .o(g52520_sb) );
na02s01 TIMEBOOST_cell_31984 ( .a(configuration_pci_err_addr_483), .b(wbm_adr_o_13_), .o(TIMEBOOST_net_9903) );
na02s01 TIMEBOOST_cell_30997 ( .a(TIMEBOOST_net_9409), .b(g61776_db), .o(TIMEBOOST_net_3509) );
na02s02 TIMEBOOST_cell_45245 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__Q), .b(n_4329), .o(TIMEBOOST_net_14861) );
in01f02 g52521_u0 ( .a(FE_OFN2242_g52675_p), .o(g52521_sb) );
na02s02 TIMEBOOST_cell_31983 ( .a(TIMEBOOST_net_9902), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_4883) );
na02s01 TIMEBOOST_cell_30996 ( .a(g65781_sb), .b(pci_target_unit_fifos_pcir_data_in_158), .o(TIMEBOOST_net_9409) );
na02s01 TIMEBOOST_cell_30995 ( .a(TIMEBOOST_net_9408), .b(g64843_sb), .o(n_3726) );
in01f02 g52522_u0 ( .a(FE_OFN2243_g52675_p), .o(g52522_sb) );
na02s01 TIMEBOOST_cell_31982 ( .a(configuration_pci_err_data_530), .b(wbm_dat_o_29_), .o(TIMEBOOST_net_9902) );
na02f02 TIMEBOOST_cell_43824 ( .a(TIMEBOOST_net_14150), .b(FE_OFN1377_n_8567), .o(TIMEBOOST_net_12889) );
na02s01 TIMEBOOST_cell_45006 ( .a(TIMEBOOST_net_14741), .b(g64204_db), .o(n_3965) );
in01f02 g52523_u0 ( .a(FE_OFN2241_g52675_p), .o(g52523_sb) );
na02s02 TIMEBOOST_cell_31981 ( .a(TIMEBOOST_net_9901), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_4882) );
na02s02 TIMEBOOST_cell_43660 ( .a(TIMEBOOST_net_14068), .b(FE_OFN1268_n_4095), .o(TIMEBOOST_net_11549) );
na02s01 TIMEBOOST_cell_30993 ( .a(TIMEBOOST_net_9407), .b(g64824_db), .o(n_3734) );
in01f02 g52524_u0 ( .a(FE_OFN2242_g52675_p), .o(g52524_sb) );
na02s01 TIMEBOOST_cell_31980 ( .a(configuration_pci_err_data_528), .b(wbm_dat_o_27_), .o(TIMEBOOST_net_9901) );
na02s02 TIMEBOOST_cell_45246 ( .a(TIMEBOOST_net_14861), .b(FE_OFN1253_n_4143), .o(TIMEBOOST_net_12036) );
na02s02 TIMEBOOST_cell_30992 ( .a(n_3764), .b(g64824_sb), .o(TIMEBOOST_net_9407) );
in01f01 g52525_u0 ( .a(FE_OFN1472_g52675_p), .o(g52525_sb) );
na02s01 TIMEBOOST_cell_30991 ( .a(TIMEBOOST_net_9406), .b(g64817_db), .o(n_3742) );
na02f02 TIMEBOOST_cell_32357 ( .a(TIMEBOOST_net_10089), .b(g58654_sb), .o(TIMEBOOST_net_6265) );
na02s01 TIMEBOOST_cell_15844 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_78), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3179) );
in01f02 g52526_u0 ( .a(FE_OFN2243_g52675_p), .o(g52526_sb) );
na02s02 TIMEBOOST_cell_31979 ( .a(TIMEBOOST_net_9900), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_4881) );
na02s01 TIMEBOOST_cell_30990 ( .a(n_3741), .b(g64817_sb), .o(TIMEBOOST_net_9406) );
na02f02 TIMEBOOST_cell_22019 ( .a(TIMEBOOST_net_6266), .b(g58655_sb), .o(n_9234) );
in01f02 g52527_u0 ( .a(FE_OFN2243_g52675_p), .o(g52527_sb) );
na02f02 TIMEBOOST_cell_22615 ( .a(TIMEBOOST_net_6564), .b(FE_OFN1565_n_12502), .o(n_12518) );
na02m02 TIMEBOOST_cell_42159 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__Q), .b(n_9677), .o(TIMEBOOST_net_13318) );
na02s01 TIMEBOOST_cell_30989 ( .a(TIMEBOOST_net_9405), .b(g64749_sb), .o(n_3793) );
in01f01 g52528_u0 ( .a(FE_OFN1472_g52675_p), .o(g52528_sb) );
na02m02 TIMEBOOST_cell_43825 ( .a(n_9016), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__Q), .o(TIMEBOOST_net_14151) );
na02s01 TIMEBOOST_cell_40855 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__Q), .b(n_13168), .o(TIMEBOOST_net_12666) );
na02f02 TIMEBOOST_cell_43826 ( .a(TIMEBOOST_net_14151), .b(FE_OFN1407_n_8567), .o(TIMEBOOST_net_12932) );
in01f01 g52529_u0 ( .a(FE_OFN1471_g52675_p), .o(g52529_sb) );
na02s01 TIMEBOOST_cell_31978 ( .a(configuration_pci_err_data_525), .b(wbm_dat_o_24_), .o(TIMEBOOST_net_9900) );
na03s02 TIMEBOOST_cell_5539 ( .a(n_4672), .b(g65084_sb), .c(g65084_db), .o(n_4304) );
na03s02 TIMEBOOST_cell_5540 ( .a(n_4488), .b(g65088_sb), .c(g65088_db), .o(n_4302) );
in01f01 g52530_u0 ( .a(FE_OFN1472_g52675_p), .o(g52530_sb) );
na02s01 TIMEBOOST_cell_30986 ( .a(pci_target_unit_fifos_pcir_data_in_163), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__Q), .o(TIMEBOOST_net_9404) );
na02s02 TIMEBOOST_cell_40854 ( .a(TIMEBOOST_net_12665), .b(FE_OFN1327_n_13547), .o(TIMEBOOST_net_11621) );
na02s01 TIMEBOOST_cell_30985 ( .a(TIMEBOOST_net_9403), .b(g65669_sb), .o(n_2029) );
in01f01 g52531_u0 ( .a(FE_OFN1471_g52675_p), .o(g52531_sb) );
na02s02 TIMEBOOST_cell_31977 ( .a(TIMEBOOST_net_9899), .b(FE_OFN1185_n_3476), .o(TIMEBOOST_net_4880) );
na02s01 TIMEBOOST_cell_42034 ( .a(TIMEBOOST_net_13255), .b(g62480_sb), .o(n_6629) );
na03s02 TIMEBOOST_cell_5542 ( .a(n_4442), .b(g65090_sb), .c(g65090_db), .o(n_4300) );
in01f01 g52532_u0 ( .a(FE_OFN1471_g52675_p), .o(g52532_sb) );
na02s01 TIMEBOOST_cell_31976 ( .a(configuration_pci_err_addr_481), .b(wbm_adr_o_11_), .o(TIMEBOOST_net_9899) );
na02s02 TIMEBOOST_cell_43520 ( .a(TIMEBOOST_net_13998), .b(FE_OFN2064_n_6391), .o(TIMEBOOST_net_12146) );
na03s02 TIMEBOOST_cell_5544 ( .a(n_4444), .b(g65097_sb), .c(g65097_db), .o(n_4295) );
in01f01 g52533_u0 ( .a(FE_OFN1471_g52675_p), .o(g52533_sb) );
na02s02 TIMEBOOST_cell_32017 ( .a(TIMEBOOST_net_9919), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4901) );
na02s01 TIMEBOOST_cell_41786 ( .a(TIMEBOOST_net_13131), .b(g64832_sb), .o(n_4448) );
na02s01 TIMEBOOST_cell_45606 ( .a(TIMEBOOST_net_15041), .b(g65221_sb), .o(n_2666) );
in01f01 g52534_u0 ( .a(FE_OFN1471_g52675_p), .o(g52534_sb) );
na02s02 TIMEBOOST_cell_31975 ( .a(TIMEBOOST_net_9898), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_4879) );
na02s01 TIMEBOOST_cell_38650 ( .a(TIMEBOOST_net_11563), .b(g61812_sb), .o(n_8168) );
na02f02 TIMEBOOST_cell_44230 ( .a(TIMEBOOST_net_14353), .b(FE_OFN1390_n_8567), .o(TIMEBOOST_net_12862) );
ao12f02 g52543_u0 ( .a(pci_target_unit_pci_target_sm_backoff), .b(n_14529), .c(FE_OFN191_n_1193), .o(n_14586) );
no02m02 g52544_u0 ( .a(n_14663), .b(pci_target_unit_wbm_sm_pciw_fifo_control_in), .o(n_14764) );
no02s01 g52545_u0 ( .a(pci_perr_i), .b(out_bckp_perr_en_out), .o(n_14624) );
na02f02 TIMEBOOST_cell_41360 ( .a(TIMEBOOST_net_12918), .b(g57265_sb), .o(n_11487) );
ao12s02 g52547_u0 ( .a(n_8564), .b(n_1185), .c(pci_target_unit_wbm_sm_pciw_fifo_control_in_84), .o(n_14694) );
na02f02 TIMEBOOST_cell_42404 ( .a(TIMEBOOST_net_13440), .b(g57245_sb), .o(n_11512) );
ao12f04 g52549_u0 ( .a(n_8582), .b(n_1101), .c(FE_OFN2198_n_10256), .o(n_10281) );
ao12m03 g52550_u0 ( .a(wishbone_slave_unit_del_sync_req_comp_pending_sample), .b(n_14620), .c(wishbone_slave_unit_del_sync_req_done_reg), .o(n_14623) );
ao22m02 g52551_u0 ( .a(n_671), .b(n_14689), .c(n_14688), .d(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in), .o(n_14691) );
ao22m02 g52552_u0 ( .a(n_661), .b(n_14689), .c(n_14688), .d(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_50), .o(n_14690) );
ao12f02 g52554_u0 ( .a(n_14731), .b(n_14800), .c(wbm_dat_o_0_), .o(n_14802) );
ao12f02 g52556_u0 ( .a(n_14728), .b(n_16306), .c(wbm_dat_o_11_), .o(n_14799) );
ao12f02 g52557_u0 ( .a(n_14727), .b(n_14800), .c(wbm_dat_o_12_), .o(n_14798) );
ao12f02 g52558_u0 ( .a(n_14726), .b(n_16306), .c(wbm_dat_o_13_), .o(n_14797) );
ao12f02 g52559_u0 ( .a(n_14724), .b(n_16306), .c(wbm_dat_o_14_), .o(n_14796) );
ao12m02 g52560_u0 ( .a(n_14670), .b(n_14800), .c(wbm_dat_o_15_), .o(n_14763) );
ao12f02 g52561_u0 ( .a(n_14723), .b(n_14800), .c(wbm_dat_o_16_), .o(n_14794) );
ao12f02 g52562_u0 ( .a(n_14722), .b(n_14800), .c(wbm_dat_o_17_), .o(n_14793) );
ao12f02 g52563_u0 ( .a(n_14669), .b(n_16306), .c(wbm_dat_o_18_), .o(n_14762) );
ao12f02 g52564_u0 ( .a(n_14721), .b(n_16306), .c(wbm_dat_o_19_), .o(n_14792) );
ao12m02 g52565_u0 ( .a(n_14719), .b(n_14800), .c(wbm_dat_o_1_), .o(n_14791) );
ao12f02 g52566_u0 ( .a(n_14717), .b(n_16306), .c(wbm_dat_o_20_), .o(n_14790) );
ao12m02 g52567_u0 ( .a(n_14715), .b(n_14800), .c(wbm_dat_o_21_), .o(n_14789) );
ao12f02 g52569_u0 ( .a(n_14713), .b(n_14800), .c(wbm_dat_o_23_), .o(n_14786) );
ao12f02 g52570_u0 ( .a(n_14711), .b(n_14800), .c(wbm_dat_o_24_), .o(n_14784) );
ao12f02 g52571_u0 ( .a(n_14710), .b(n_16306), .c(wbm_dat_o_25_), .o(n_14783) );
ao12f02 g52572_u0 ( .a(n_14709), .b(n_16306), .c(wbm_dat_o_26_), .o(n_14781) );
ao12m02 g52573_u0 ( .a(n_14708), .b(n_16306), .c(wbm_dat_o_27_), .o(n_14780) );
ao12m02 g52574_u0 ( .a(n_14706), .b(n_16306), .c(wbm_dat_o_28_), .o(n_14778) );
ao12m02 g52575_u0 ( .a(n_14705), .b(n_16306), .c(wbm_dat_o_29_), .o(n_14777) );
ao12f02 g52576_u0 ( .a(n_14703), .b(n_16306), .c(wbm_dat_o_2_), .o(n_14776) );
ao12m02 g52577_u0 ( .a(n_14702), .b(n_16306), .c(wbm_dat_o_30_), .o(n_14775) );
ao12f02 g52578_u0 ( .a(n_14701), .b(n_16306), .c(wbm_dat_o_31_), .o(n_14773) );
ao12f02 g52579_u0 ( .a(n_14700), .b(n_14800), .c(wbm_dat_o_3_), .o(n_14772) );
ao12m02 g52580_u0 ( .a(n_14699), .b(n_14800), .c(wbm_dat_o_4_), .o(n_14770) );
ao12f02 g52581_u0 ( .a(n_14698), .b(n_14800), .c(wbm_dat_o_5_), .o(n_14769) );
ao12f02 g52582_u0 ( .a(n_14697), .b(n_14800), .c(wbm_dat_o_6_), .o(n_14768) );
ao12f02 g52583_u0 ( .a(n_14668), .b(n_16306), .c(wbm_dat_o_7_), .o(n_14761) );
ao12f02 g52584_u0 ( .a(n_14696), .b(n_16306), .c(wbm_dat_o_8_), .o(n_14767) );
ao12f02 g52585_u0 ( .a(n_14695), .b(n_14800), .c(wbm_dat_o_9_), .o(n_14766) );
ao12f02 g52586_u0 ( .a(n_14667), .b(n_16306), .c(wbm_sel_o_0_), .o(n_14760) );
ao12f02 g52587_u0 ( .a(n_14666), .b(n_16306), .c(wbm_sel_o_1_), .o(n_14759) );
ao12f02 g52588_u0 ( .a(n_14665), .b(n_16306), .c(wbm_sel_o_2_), .o(n_14757) );
ao12f02 g52589_u0 ( .a(n_14664), .b(n_16306), .c(wbm_sel_o_3_), .o(n_14756) );
in01s01 g52590_u0 ( .a(n_8757), .o(g52590_sb) );
no02f04 TIMEBOOST_cell_19045 ( .a(TIMEBOOST_net_4779), .b(FE_RN_545_0), .o(TIMEBOOST_net_915) );
na02s02 TIMEBOOST_cell_37830 ( .a(TIMEBOOST_net_11153), .b(g58385_sb), .o(n_9446) );
na02s02 TIMEBOOST_cell_37832 ( .a(TIMEBOOST_net_11154), .b(g58420_sb), .o(n_9427) );
in01s01 g52591_u0 ( .a(n_8757), .o(g52591_sb) );
na02m02 TIMEBOOST_cell_38632 ( .a(TIMEBOOST_net_11554), .b(g59090_sb), .o(n_8716) );
na02s02 TIMEBOOST_cell_37818 ( .a(TIMEBOOST_net_11147), .b(g58177_sb), .o(n_9612) );
na02s02 TIMEBOOST_cell_37800 ( .a(TIMEBOOST_net_11138), .b(g61945_sb), .o(n_7935) );
in01s01 g52592_u0 ( .a(n_8757), .o(g52592_sb) );
na02s01 TIMEBOOST_cell_19028 ( .a(wishbone_slave_unit_pcim_sm_data_in_650), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__Q), .o(TIMEBOOST_net_4771) );
na02s02 g52395_u2 ( .a(n_14674), .b(n_14839), .o(g52395_db) );
na02m02 TIMEBOOST_cell_37792 ( .a(TIMEBOOST_net_11134), .b(g63195_db), .o(n_3460) );
in01s01 g52593_u0 ( .a(n_8757), .o(g52593_sb) );
na02s01 TIMEBOOST_cell_19030 ( .a(wishbone_slave_unit_pcim_sm_data_in_654), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__Q), .o(TIMEBOOST_net_4772) );
na02f02 TIMEBOOST_cell_37128 ( .a(TIMEBOOST_net_10802), .b(n_12580), .o(n_12842) );
na02f02 TIMEBOOST_cell_37092 ( .a(TIMEBOOST_net_10784), .b(FE_OFN1588_n_13736), .o(g53207_p) );
in01m02 g52594_u0 ( .a(n_10256), .o(g52594_sb) );
na02f02 TIMEBOOST_cell_22489 ( .a(TIMEBOOST_net_6501), .b(FE_OFN1581_n_12306), .o(n_12490) );
na02s02 TIMEBOOST_cell_40708 ( .a(TIMEBOOST_net_12592), .b(g62674_sb), .o(n_6191) );
na02s02 TIMEBOOST_cell_43160 ( .a(TIMEBOOST_net_13818), .b(FE_OFN1207_n_6356), .o(TIMEBOOST_net_12130) );
in01f02 g52595_u0 ( .a(FE_OFN2198_n_10256), .o(g52595_sb) );
na02s02 TIMEBOOST_cell_45247 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__Q), .b(n_3619), .o(TIMEBOOST_net_14862) );
na02s02 TIMEBOOST_cell_40798 ( .a(TIMEBOOST_net_12637), .b(g62461_sb), .o(n_6674) );
na02m04 TIMEBOOST_cell_45828 ( .a(TIMEBOOST_net_15152), .b(FE_OFN2134_n_13124), .o(TIMEBOOST_net_14994) );
in01f02 g52596_u0 ( .a(FE_OFN2198_n_10256), .o(g52596_sb) );
na02s02 TIMEBOOST_cell_45021 ( .a(TIMEBOOST_net_1662), .b(g61974_db), .o(TIMEBOOST_net_14749) );
na02s02 TIMEBOOST_cell_40800 ( .a(TIMEBOOST_net_12638), .b(g62455_sb), .o(n_6686) );
na02s02 TIMEBOOST_cell_45248 ( .a(TIMEBOOST_net_14862), .b(FE_OFN1268_n_4095), .o(TIMEBOOST_net_12070) );
in01f01 g52597_u0 ( .a(n_8935), .o(g52597_sb) );
na02f02 TIMEBOOST_cell_41368 ( .a(TIMEBOOST_net_12922), .b(g57211_sb), .o(n_11545) );
na02f01 g52597_u2 ( .a(n_3169), .b(n_8935), .o(g52597_db) );
na02f02 TIMEBOOST_cell_22029 ( .a(TIMEBOOST_net_6271), .b(FE_OFN1596_n_13741), .o(n_14264) );
in01f02 g52598_u0 ( .a(FE_OFN2200_n_10256), .o(g52598_sb) );
na02s01 TIMEBOOST_cell_39554 ( .a(TIMEBOOST_net_12015), .b(g61676_sb), .o(TIMEBOOST_net_10660) );
na02s02 TIMEBOOST_cell_40802 ( .a(TIMEBOOST_net_12639), .b(g62473_sb), .o(n_6644) );
na02s01 TIMEBOOST_cell_30949 ( .a(TIMEBOOST_net_9385), .b(g65087_sb), .o(n_3598) );
in01f02 g52599_u0 ( .a(FE_OFN2200_n_10256), .o(g52599_sb) );
na02f02 TIMEBOOST_cell_44742 ( .a(TIMEBOOST_net_14609), .b(n_11984), .o(n_12514) );
na02s02 TIMEBOOST_cell_40804 ( .a(TIMEBOOST_net_12640), .b(g62403_sb), .o(n_6793) );
na03s02 TIMEBOOST_cell_33791 ( .a(FE_OFN254_n_9825), .b(g58228_sb), .c(g58228_db), .o(n_9561) );
in01f01 g52600_u0 ( .a(n_8935), .o(g52600_sb) );
na02s02 TIMEBOOST_cell_45249 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__Q), .b(n_4194), .o(TIMEBOOST_net_14863) );
na02f01 g52600_u2 ( .a(n_3151), .b(n_8935), .o(g52600_db) );
na03s02 TIMEBOOST_cell_33587 ( .a(TIMEBOOST_net_9556), .b(n_5633), .c(g62090_sb), .o(n_5617) );
in01f02 g52601_u0 ( .a(FE_OFN2200_n_10256), .o(g52601_sb) );
na02f02 TIMEBOOST_cell_44743 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__Q), .b(FE_OFN1579_n_12306), .o(TIMEBOOST_net_14610) );
na02s01 TIMEBOOST_cell_40806 ( .a(TIMEBOOST_net_12641), .b(g62386_sb), .o(n_6828) );
na03s02 TIMEBOOST_cell_5416 ( .a(n_4473), .b(g64884_sb), .c(g64884_db), .o(n_4416) );
in01f02 g52602_u0 ( .a(FE_OFN2200_n_10256), .o(g52602_sb) );
na03s02 TIMEBOOST_cell_33793 ( .a(FE_OFN231_n_9839), .b(g58185_sb), .c(g58185_db), .o(n_9602) );
na02f02 g52602_u2 ( .a(n_4210), .b(FE_OFN2200_n_10256), .o(g52602_db) );
na02s01 TIMEBOOST_cell_30950 ( .a(n_4473), .b(g64848_sb), .o(TIMEBOOST_net_9386) );
in01f02 g52603_u0 ( .a(FE_OFN2200_n_10256), .o(g52603_sb) );
na02s02 TIMEBOOST_cell_41708 ( .a(TIMEBOOST_net_13092), .b(g58779_db), .o(n_9846) );
na02s01 TIMEBOOST_cell_40808 ( .a(TIMEBOOST_net_12642), .b(g62394_sb), .o(n_6809) );
na02s02 TIMEBOOST_cell_43661 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__Q), .b(n_3746), .o(TIMEBOOST_net_14069) );
in01f01 g52604_u0 ( .a(n_10256), .o(g52604_sb) );
na02s02 TIMEBOOST_cell_45250 ( .a(TIMEBOOST_net_14863), .b(FE_OFN1244_n_4092), .o(TIMEBOOST_net_12050) );
na02s02 TIMEBOOST_cell_40710 ( .a(TIMEBOOST_net_12593), .b(g62510_sb), .o(n_6558) );
na02s02 TIMEBOOST_cell_43662 ( .a(TIMEBOOST_net_14069), .b(FE_OFN2063_n_6391), .o(TIMEBOOST_net_12258) );
in01f02 g52605_u0 ( .a(FE_OFN2200_n_10256), .o(g52605_sb) );
na02s02 TIMEBOOST_cell_45251 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__Q), .b(n_3711), .o(TIMEBOOST_net_14864) );
na02s01 TIMEBOOST_cell_40810 ( .a(TIMEBOOST_net_12643), .b(g62372_sb), .o(n_6859) );
na02m02 TIMEBOOST_cell_43777 ( .a(n_9669), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__Q), .o(TIMEBOOST_net_14127) );
in01f01 g52606_u0 ( .a(n_8935), .o(g52606_sb) );
na03s02 TIMEBOOST_cell_33586 ( .a(TIMEBOOST_net_9557), .b(n_5633), .c(g62077_sb), .o(n_5634) );
na02f01 g52606_u2 ( .a(n_3487), .b(n_8935), .o(g52606_db) );
na03s02 TIMEBOOST_cell_33779 ( .a(FE_OFN221_n_9846), .b(g57958_sb), .c(g57958_db), .o(n_9847) );
in01f02 g52607_u0 ( .a(FE_OFN2200_n_10256), .o(g52607_sb) );
na02m04 TIMEBOOST_cell_45829 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_777), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_12__Q), .o(TIMEBOOST_net_15153) );
na02s02 TIMEBOOST_cell_40812 ( .a(TIMEBOOST_net_12644), .b(FE_OFN1310_n_6624), .o(TIMEBOOST_net_11591) );
na02m04 TIMEBOOST_cell_45830 ( .a(TIMEBOOST_net_15153), .b(FE_OFN2134_n_13124), .o(TIMEBOOST_net_14995) );
in01f02 g52608_u0 ( .a(FE_OFN2198_n_10256), .o(g52608_sb) );
na02s02 TIMEBOOST_cell_45252 ( .a(TIMEBOOST_net_14864), .b(FE_OFN1242_n_4092), .o(TIMEBOOST_net_12037) );
na02s02 TIMEBOOST_cell_40814 ( .a(TIMEBOOST_net_12645), .b(FE_OFN1320_n_6436), .o(TIMEBOOST_net_11594) );
na02m04 TIMEBOOST_cell_45831 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_13__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_778), .o(TIMEBOOST_net_15154) );
in01f02 g52609_u0 ( .a(FE_OFN2198_n_10256), .o(g52609_sb) );
na02s02 TIMEBOOST_cell_40840 ( .a(TIMEBOOST_net_12658), .b(FE_OFN1333_n_13547), .o(TIMEBOOST_net_11607) );
na02f02 TIMEBOOST_cell_41382 ( .a(TIMEBOOST_net_12929), .b(g57467_sb), .o(n_11265) );
na02s01 TIMEBOOST_cell_45253 ( .a(n_4914), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__Q), .o(TIMEBOOST_net_14865) );
in01f02 g52610_u0 ( .a(FE_OFN2200_n_10256), .o(g52610_sb) );
na02s01 TIMEBOOST_cell_43161 ( .a(n_3603), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__Q), .o(TIMEBOOST_net_13819) );
na02s02 TIMEBOOST_cell_40816 ( .a(TIMEBOOST_net_12646), .b(g62935_sb), .o(n_6011) );
na02f04 TIMEBOOST_cell_45832 ( .a(TIMEBOOST_net_15154), .b(FE_OFN2134_n_13124), .o(TIMEBOOST_net_14996) );
in01f02 g52611_u0 ( .a(FE_OFN2200_n_10256), .o(g52611_sb) );
na02s04 TIMEBOOST_cell_45833 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_10__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_775), .o(TIMEBOOST_net_15155) );
na02s02 TIMEBOOST_cell_40818 ( .a(TIMEBOOST_net_12647), .b(g63192_sb), .o(n_5772) );
na02s02 TIMEBOOST_cell_39556 ( .a(TIMEBOOST_net_12016), .b(g59797_sb), .o(TIMEBOOST_net_596) );
in01f02 g52612_u0 ( .a(FE_OFN2200_n_10256), .o(g52612_sb) );
na02s02 TIMEBOOST_cell_45254 ( .a(TIMEBOOST_net_14865), .b(FE_OFN1222_n_6391), .o(TIMEBOOST_net_12137) );
na02s02 TIMEBOOST_cell_40820 ( .a(TIMEBOOST_net_12648), .b(g62412_sb), .o(n_6774) );
na02s01 TIMEBOOST_cell_43162 ( .a(TIMEBOOST_net_13819), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_12565) );
oa22m02 g52613_u0 ( .a(FE_OFN2198_n_10256), .b(wbu_addr_in_278), .c(n_10155), .d(n_4208), .o(n_10170) );
in01f01 g52614_u0 ( .a(n_8935), .o(g52614_sb) );
na02f02 TIMEBOOST_cell_44658 ( .a(TIMEBOOST_net_14567), .b(FE_OFN1402_n_8567), .o(TIMEBOOST_net_12789) );
na02f01 g52614_u2 ( .a(n_4890), .b(n_8935), .o(g52614_db) );
na02m02 TIMEBOOST_cell_42241 ( .a(n_9448), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__Q), .o(TIMEBOOST_net_13359) );
oa22f02 g52615_u0 ( .a(FE_OFN2198_n_10256), .b(wbu_addr_in_280), .c(n_10155), .d(n_4196), .o(n_10157) );
in01f02 g52616_u0 ( .a(FE_OFN2198_n_10256), .o(g52616_sb) );
na02m02 TIMEBOOST_cell_40842 ( .a(TIMEBOOST_net_12659), .b(FE_OFN1326_n_13547), .o(TIMEBOOST_net_11614) );
na02f02 TIMEBOOST_cell_22507 ( .a(TIMEBOOST_net_6510), .b(FE_OFN1583_n_12306), .o(n_12741) );
na02s02 TIMEBOOST_cell_43163 ( .a(n_3720), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__Q), .o(TIMEBOOST_net_13820) );
in01f01 g52617_u0 ( .a(n_10256), .o(g52617_sb) );
na02f02 TIMEBOOST_cell_22509 ( .a(TIMEBOOST_net_6511), .b(FE_OFN1579_n_12306), .o(n_12734) );
na02s01 TIMEBOOST_cell_40712 ( .a(TIMEBOOST_net_12594), .b(g63147_sb), .o(n_5846) );
na02s01 TIMEBOOST_cell_42672 ( .a(TIMEBOOST_net_13574), .b(g65419_da), .o(n_4227) );
in01f01 g52618_u0 ( .a(n_10256), .o(g52618_sb) );
na02s02 TIMEBOOST_cell_45255 ( .a(n_4385), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__Q), .o(TIMEBOOST_net_14866) );
na02f02 g52618_u2 ( .a(n_2273), .b(n_10256), .o(g52618_db) );
na02s02 TIMEBOOST_cell_43164 ( .a(TIMEBOOST_net_13820), .b(FE_OFN1224_n_6391), .o(TIMEBOOST_net_12567) );
in01f01 g52619_u0 ( .a(n_10256), .o(g52619_sb) );
na02f02 TIMEBOOST_cell_22513 ( .a(TIMEBOOST_net_6513), .b(FE_OFN1584_n_12306), .o(n_12504) );
na02f02 g52619_u2 ( .a(n_2488), .b(n_10256), .o(g52619_db) );
na02s02 TIMEBOOST_cell_43663 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__Q), .b(n_3662), .o(TIMEBOOST_net_14070) );
in01f02 g52620_u0 ( .a(FE_OFN2198_n_10256), .o(g52620_sb) );
na02s02 TIMEBOOST_cell_40844 ( .a(TIMEBOOST_net_12660), .b(FE_OFN1326_n_13547), .o(TIMEBOOST_net_11612) );
na02s02 TIMEBOOST_cell_45256 ( .a(TIMEBOOST_net_14866), .b(FE_OFN1248_n_4093), .o(TIMEBOOST_net_12601) );
na02s04 TIMEBOOST_cell_45834 ( .a(TIMEBOOST_net_15155), .b(FE_OFN2136_n_13124), .o(TIMEBOOST_net_14997) );
in01f01 g52621_u0 ( .a(n_10256), .o(g52621_sb) );
na02s02 TIMEBOOST_cell_43664 ( .a(TIMEBOOST_net_14070), .b(FE_OFN1230_n_6391), .o(TIMEBOOST_net_12167) );
na02f02 g52621_u2 ( .a(n_2257), .b(n_10256), .o(g52621_db) );
na02f02 TIMEBOOST_cell_22517 ( .a(TIMEBOOST_net_6515), .b(FE_OFN1583_n_12306), .o(n_12625) );
in01f02 g52622_u0 ( .a(FE_OFN2198_n_10256), .o(g52622_sb) );
na02s02 TIMEBOOST_cell_40846 ( .a(TIMEBOOST_net_12661), .b(FE_OFN1333_n_13547), .o(TIMEBOOST_net_11613) );
na02m04 TIMEBOOST_cell_45835 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_11__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_776), .o(TIMEBOOST_net_15156) );
na02s02 TIMEBOOST_cell_43665 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__Q), .b(n_4327), .o(TIMEBOOST_net_14071) );
no02f04 g52623_u0 ( .a(wbu_addr_in_251), .b(FE_OFN2198_n_10256), .o(g52623_p) );
ao12f02 g52623_u1 ( .a(g52623_p), .b(wbu_addr_in_251), .c(FE_OFN2198_n_10256), .o(n_10106) );
in01s01 g52624_u0 ( .a(n_16748), .o(g52624_sb) );
na02s02 g52624_u1 ( .a(pci_target_unit_pcit_if_strd_addr_in_695), .b(g52624_sb), .o(g52624_da) );
na02s01 g52624_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_59), .b(n_16748), .o(g52624_db) );
na02s01 TIMEBOOST_cell_36368 ( .a(TIMEBOOST_net_10422), .b(TIMEBOOST_net_3227), .o(n_1657) );
in01m01 g52625_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52625_sb) );
na02m02 TIMEBOOST_cell_44159 ( .a(n_9626), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__Q), .o(TIMEBOOST_net_14318) );
na02s02 g52625_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_60), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52625_db) );
na02f02 TIMEBOOST_cell_39558 ( .a(n_7543), .b(TIMEBOOST_net_12017), .o(n_8749) );
in01s01 g52626_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52626_sb) );
na02s02 g52626_u1 ( .a(pci_target_unit_pcit_if_strd_addr_in_697), .b(g52626_sb), .o(g52626_da) );
na02f02 TIMEBOOST_cell_44744 ( .a(TIMEBOOST_net_14610), .b(n_16631), .o(n_12658) );
na02f02 TIMEBOOST_cell_38914 ( .a(TIMEBOOST_net_11695), .b(FE_OFN2198_n_10256), .o(TIMEBOOST_net_10701) );
in01s01 g52627_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52627_sb) );
na02f06 TIMEBOOST_cell_36834 ( .a(TIMEBOOST_net_10655), .b(g75160_db), .o(n_16533) );
na02m02 TIMEBOOST_cell_42523 ( .a(TIMEBOOST_net_6361), .b(wbu_addr_in_271), .o(TIMEBOOST_net_13500) );
na02s01 TIMEBOOST_cell_18533 ( .a(TIMEBOOST_net_4523), .b(g63433_sb), .o(n_4932) );
in01m01 g52628_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52628_sb) );
na02s01 TIMEBOOST_cell_9317 ( .a(TIMEBOOST_net_1225), .b(g63548_db), .o(n_4609) );
na02s02 g52628_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_63), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52628_db) );
na02s01 TIMEBOOST_cell_42735 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__Q), .b(n_4525), .o(TIMEBOOST_net_13606) );
in01s01 g52629_u0 ( .a(n_16748), .o(g52629_sb) );
na02s01 TIMEBOOST_cell_38689 ( .a(n_4014), .b(g62808_sb), .o(TIMEBOOST_net_11583) );
na03s02 TIMEBOOST_cell_40325 ( .a(n_4444), .b(FE_OFN636_n_4669), .c(FE_RN_720_0), .o(TIMEBOOST_net_12401) );
na02s01 TIMEBOOST_cell_38652 ( .a(TIMEBOOST_net_11564), .b(n_1600), .o(TIMEBOOST_net_4166) );
in01s02 g52630_u0 ( .a(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52630_sb) );
na02m02 TIMEBOOST_cell_38915 ( .a(n_3465), .b(wbu_addr_in_276), .o(TIMEBOOST_net_11696) );
na02s01 TIMEBOOST_cell_42736 ( .a(TIMEBOOST_net_13606), .b(FE_OFN717_n_8176), .o(TIMEBOOST_net_11099) );
na02s02 TIMEBOOST_cell_38116 ( .a(TIMEBOOST_net_11296), .b(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_4608) );
in01s02 g52631_u0 ( .a(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52631_sb) );
na02s02 g52631_u1 ( .a(pci_target_unit_pcit_if_strd_addr_in_702), .b(g52631_sb), .o(g52631_da) );
na02f02 TIMEBOOST_cell_39135 ( .a(FE_OFN1605_n_13997), .b(TIMEBOOST_net_10179), .o(TIMEBOOST_net_11806) );
na02s01 TIMEBOOST_cell_39310 ( .a(TIMEBOOST_net_11893), .b(g65359_sb), .o(n_4254) );
in01s02 g52632_u0 ( .a(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52632_sb) );
na02s02 g52632_u1 ( .a(pci_target_unit_pcit_if_strd_addr_in_703), .b(g52632_sb), .o(g52632_da) );
na02s02 g52632_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_67), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52632_db) );
na02f02 TIMEBOOST_cell_12615 ( .a(n_13997), .b(TIMEBOOST_net_2874), .o(TIMEBOOST_net_668) );
in01s01 g52633_u0 ( .a(n_16748), .o(g52633_sb) );
na02s01 TIMEBOOST_cell_17868 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__Q), .b(g65314_sb), .o(TIMEBOOST_net_4191) );
na02s01 g52633_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_68), .b(n_16748), .o(g52633_db) );
na02s02 TIMEBOOST_cell_17869 ( .a(TIMEBOOST_net_4191), .b(g65314_db), .o(n_4194) );
in01s01 g52634_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52634_sb) );
na02s01 g52634_u1 ( .a(pci_target_unit_pcit_if_strd_addr_in_705), .b(g52634_sb), .o(g52634_da) );
na03s02 TIMEBOOST_cell_38117 ( .a(g64123_da), .b(g64123_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__Q), .o(TIMEBOOST_net_11297) );
na02s02 TIMEBOOST_cell_38118 ( .a(TIMEBOOST_net_11297), .b(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_4592) );
in01s02 g52635_u0 ( .a(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52635_sb) );
na02s02 g52635_u1 ( .a(pci_target_unit_pcit_if_strd_addr_in_706), .b(g52635_sb), .o(g52635_da) );
na02s02 g52635_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_70), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52635_db) );
na02s02 TIMEBOOST_cell_36288 ( .a(TIMEBOOST_net_10382), .b(n_1365), .o(n_2400) );
in01s01 g52636_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52636_sb) );
na02s01 TIMEBOOST_cell_9954 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_17__Q), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_1544) );
na02s01 g52636_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_71), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52636_db) );
na02s01 TIMEBOOST_cell_9955 ( .a(TIMEBOOST_net_1544), .b(n_13221), .o(TIMEBOOST_net_512) );
in01s02 g52637_u0 ( .a(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52637_sb) );
na02s02 g52637_u1 ( .a(pci_target_unit_pcit_if_strd_addr_in_708), .b(g52637_sb), .o(g52637_da) );
na03s02 TIMEBOOST_cell_38137 ( .a(TIMEBOOST_net_4030), .b(g64231_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__Q), .o(TIMEBOOST_net_11307) );
na02s02 TIMEBOOST_cell_19257 ( .a(TIMEBOOST_net_4885), .b(g60663_sb), .o(n_5656) );
in01s02 g52638_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52638_sb) );
na02s01 TIMEBOOST_cell_18296 ( .a(g61923_sb), .b(g62021_db), .o(TIMEBOOST_net_4405) );
na02s01 g52638_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_73), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52638_db) );
na02s02 TIMEBOOST_cell_38120 ( .a(TIMEBOOST_net_11298), .b(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_4669) );
in01s01 g52639_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52639_sb) );
na02m02 TIMEBOOST_cell_44349 ( .a(n_9559), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__Q), .o(TIMEBOOST_net_14413) );
na02s01 g52639_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_74), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52639_db) );
na02s01 TIMEBOOST_cell_42737 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__Q), .b(n_1648), .o(TIMEBOOST_net_13607) );
na03s02 TIMEBOOST_cell_38119 ( .a(TIMEBOOST_net_4262), .b(g64125_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__Q), .o(TIMEBOOST_net_11298) );
na02s02 TIMEBOOST_cell_18004 ( .a(pci_target_unit_fifos_pciw_cbe_in_152), .b(g64170_sb), .o(TIMEBOOST_net_4259) );
na02s01 TIMEBOOST_cell_39314 ( .a(TIMEBOOST_net_11895), .b(g65840_db), .o(n_2017) );
in01s01 g52641_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52641_sb) );
na02s01 TIMEBOOST_cell_42738 ( .a(TIMEBOOST_net_13607), .b(FE_OFN710_n_8232), .o(TIMEBOOST_net_11089) );
na02s01 g52641_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_76), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52641_db) );
na02f02 TIMEBOOST_cell_42524 ( .a(TIMEBOOST_net_13500), .b(g52606_sb), .o(TIMEBOOST_net_11731) );
in01s01 g52642_u0 ( .a(n_16748), .o(g52642_sb) );
na02s01 TIMEBOOST_cell_17870 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__Q), .b(g65332_sb), .o(TIMEBOOST_net_4192) );
na02s01 g52642_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_77), .b(n_16748), .o(g52642_db) );
na02s01 TIMEBOOST_cell_17871 ( .a(TIMEBOOST_net_4192), .b(g65332_db), .o(n_3553) );
in01s02 g52643_u0 ( .a(n_16748), .o(g52643_sb) );
na02m02 g52643_u1 ( .a(g52643_sb), .b(pci_target_unit_pcit_if_strd_addr_in_714), .o(g52643_da) );
na02s02 g52643_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_78), .b(n_16748), .o(g52643_db) );
na02s02 TIMEBOOST_cell_38122 ( .a(TIMEBOOST_net_11299), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_4567) );
in01m01 g52644_u0 ( .a(n_16748), .o(g52644_sb) );
na02s01 TIMEBOOST_cell_18038 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(g64165_sb), .o(TIMEBOOST_net_4276) );
na02m01 g52644_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_51), .b(n_16748), .o(g52644_db) );
na02s01 TIMEBOOST_cell_37618 ( .a(TIMEBOOST_net_11047), .b(g61788_sb), .o(n_8226) );
in01m01 g52645_u0 ( .a(n_16748), .o(g52645_sb) );
na02s02 TIMEBOOST_cell_39560 ( .a(TIMEBOOST_net_12018), .b(g60407_sb), .o(TIMEBOOST_net_10661) );
na02s02 g52645_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_79), .b(n_16748), .o(g52645_db) );
na02s02 TIMEBOOST_cell_39562 ( .a(TIMEBOOST_net_12019), .b(g60407_sb), .o(TIMEBOOST_net_10662) );
in01m01 g52646_u0 ( .a(n_16748), .o(g52646_sb) );
na02s02 TIMEBOOST_cell_39547 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__Q), .b(g58283_sb), .o(TIMEBOOST_net_12012) );
na02s02 g52646_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_80), .b(n_16748), .o(g52646_db) );
na02s01 TIMEBOOST_cell_39564 ( .a(TIMEBOOST_net_12020), .b(g62610_sb), .o(n_7375) );
in01s01 g52647_u0 ( .a(FE_OFN697_n_16760), .o(g52647_sb) );
na02s02 TIMEBOOST_cell_40438 ( .a(TIMEBOOST_net_12457), .b(g62092_sb), .o(TIMEBOOST_net_11374) );
na02f02 TIMEBOOST_cell_45804 ( .a(TIMEBOOST_net_15140), .b(FE_OFN2179_n_8567), .o(TIMEBOOST_net_14576) );
na02s02 TIMEBOOST_cell_43003 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__Q), .b(g58274_sb), .o(TIMEBOOST_net_13740) );
in01m01 g52648_u0 ( .a(n_16748), .o(g52648_sb) );
na02s01 TIMEBOOST_cell_44897 ( .a(g65738_db), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__Q), .o(TIMEBOOST_net_14687) );
na02m01 g52648_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_53), .b(n_16748), .o(g52648_db) );
na02s02 TIMEBOOST_cell_39566 ( .a(TIMEBOOST_net_12021), .b(g62449_sb), .o(n_6699) );
na02s01 TIMEBOOST_cell_40437 ( .a(parchk_pci_ad_out_in_1188), .b(configuration_wb_err_data_591), .o(TIMEBOOST_net_12457) );
na03s02 TIMEBOOST_cell_517 ( .a(FE_OFN270_n_9836), .b(g57934_sb), .c(g57934_db), .o(n_9875) );
na02s02 TIMEBOOST_cell_42105 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__Q), .b(n_3578), .o(TIMEBOOST_net_13291) );
in01s01 g52650_u0 ( .a(n_16748), .o(g52650_sb) );
na02s02 g52650_u1 ( .a(pci_target_unit_pcit_if_strd_addr_in_691), .b(g52650_sb), .o(g52650_da) );
na02s02 TIMEBOOST_cell_45136 ( .a(TIMEBOOST_net_14806), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_11445) );
na02s01 TIMEBOOST_cell_36496 ( .a(TIMEBOOST_net_10486), .b(g67040_sb), .o(n_2471) );
in01s01 g52651_u0 ( .a(n_16748), .o(g52651_sb) );
na02s01 TIMEBOOST_cell_17876 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__Q), .b(g65338_sb), .o(TIMEBOOST_net_4195) );
na02m01 g52651_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_56), .b(n_16748), .o(g52651_db) );
na02s01 TIMEBOOST_cell_17877 ( .a(TIMEBOOST_net_4195), .b(g65338_db), .o(n_3550) );
in01m01 g52652_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52652_sb) );
na02f02 TIMEBOOST_cell_38916 ( .a(TIMEBOOST_net_11696), .b(FE_OFN2200_n_10256), .o(TIMEBOOST_net_10702) );
na02m01 g52652_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_57), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52652_db) );
na02s01 TIMEBOOST_cell_18301 ( .a(TIMEBOOST_net_4407), .b(FE_OFN2104_g64577_p), .o(n_5136) );
in01m01 g52653_u0 ( .a(n_16748), .o(g52653_sb) );
na02s01 TIMEBOOST_cell_40327 ( .a(n_3741), .b(g64866_db), .o(TIMEBOOST_net_12402) );
na02m01 g52653_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_58), .b(n_16748), .o(g52653_db) );
na02s02 TIMEBOOST_cell_40660 ( .a(TIMEBOOST_net_12568), .b(g62884_sb), .o(n_6109) );
no02f02 g52675_u0 ( .a(n_8872), .b(n_16945), .o(g52675_p) );
na02s02 TIMEBOOST_cell_45257 ( .a(n_4231), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__Q), .o(TIMEBOOST_net_14867) );
na02f02 g52677_u0 ( .a(n_14517), .b(n_14615), .o(n_14629) );
no02f02 g52678_u0 ( .a(n_14725), .b(n_14659), .o(n_14731) );
no02f02 g52679_u0 ( .a(n_14725), .b(n_14658), .o(n_14730) );
no02f02 g52680_u0 ( .a(n_14725), .b(n_14657), .o(n_14728) );
no02f02 g52681_u0 ( .a(n_14725), .b(n_14656), .o(n_14727) );
no02f02 g52682_u0 ( .a(n_14725), .b(n_14655), .o(n_14726) );
no02m02 g52683_u0 ( .a(n_14725), .b(n_14654), .o(n_14724) );
no02f02 g52684_u0 ( .a(n_14725), .b(n_14627), .o(n_14670) );
no02f02 g52685_u0 ( .a(n_14725), .b(n_14653), .o(n_14723) );
no02f02 g52686_u0 ( .a(n_14725), .b(n_14652), .o(n_14722) );
no02f02 g52687_u0 ( .a(n_14725), .b(n_14626), .o(n_14669) );
no02f02 g52688_u0 ( .a(n_14725), .b(n_14651), .o(n_14721) );
no02s02 g52689_u0 ( .a(n_14725), .b(n_14650), .o(n_14719) );
no02s02 g52690_u0 ( .a(n_14725), .b(n_14649), .o(n_14717) );
no02m02 g52691_u0 ( .a(n_14725), .b(n_14648), .o(n_14715) );
no02s02 g52693_u0 ( .a(n_14725), .b(n_14646), .o(n_14713) );
no02f02 g52694_u0 ( .a(n_14725), .b(n_14645), .o(n_14711) );
no02f02 g52695_u0 ( .a(n_14725), .b(n_14644), .o(n_14710) );
no02m02 g52696_u0 ( .a(n_14725), .b(n_14643), .o(n_14709) );
no02s02 g52697_u0 ( .a(n_14725), .b(n_14642), .o(n_14708) );
no02s02 g52698_u0 ( .a(n_14725), .b(n_14641), .o(n_14706) );
no02f02 g52699_u0 ( .a(n_14725), .b(n_14640), .o(n_14705) );
no02f02 g52700_u0 ( .a(n_14725), .b(n_14639), .o(n_14703) );
no02f02 g52701_u0 ( .a(n_14725), .b(n_14638), .o(n_14702) );
no02f02 g52702_u0 ( .a(n_14725), .b(n_14637), .o(n_14701) );
no02f02 g52703_u0 ( .a(n_14725), .b(n_14636), .o(n_14700) );
no02s02 g52704_u0 ( .a(n_14725), .b(n_14635), .o(n_14699) );
no02s02 g52705_u0 ( .a(n_14725), .b(n_14634), .o(n_14698) );
no02f02 g52706_u0 ( .a(n_14725), .b(n_14633), .o(n_14697) );
no02f02 g52707_u0 ( .a(n_14725), .b(n_14625), .o(n_14668) );
no02f02 g52708_u0 ( .a(n_14725), .b(n_14632), .o(n_14696) );
no02f02 g52709_u0 ( .a(n_14725), .b(n_14631), .o(n_14695) );
no02f03 g52710_u0 ( .a(n_16306), .b(pci_target_unit_wbm_sm_pciw_fifo_cbe_in), .o(n_14667) );
no02s04 g52711_u0 ( .a(n_16306), .b(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_81), .o(n_14666) );
no02f03 g52712_u0 ( .a(n_16306), .b(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_82), .o(n_14665) );
no02f03 g52713_u0 ( .a(n_16306), .b(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_83), .o(n_14664) );
na02f02 g52714_u0 ( .a(n_1532), .b(n_14620), .o(g52714_p) );
in01m02 g52714_u1 ( .a(g52714_p), .o(n_14621) );
oa12m01 g52715_u0 ( .a(n_10155), .b(wbs_stb_i), .c(n_779), .o(n_10441) );
na02f02 TIMEBOOST_cell_44350 ( .a(TIMEBOOST_net_14413), .b(FE_OFN1411_n_8567), .o(TIMEBOOST_net_12852) );
na03s02 TIMEBOOST_cell_6321 ( .a(n_4470), .b(g64834_sb), .c(g64834_db), .o(n_4446) );
ao12f02 g52718_u0 ( .a(n_14485), .b(n_13920), .c(n_2285), .o(n_14617) );
oa12m02 g52719_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_control_in_84), .b(n_1541), .c(n_1086), .o(n_14663) );
oa22m01 g52720_u0 ( .a(n_10792), .b(wbs_err_o), .c(wbs_stb_i), .d(n_471), .o(n_8874) );
in01s01 g52778_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in), .o(n_14659) );
in01s01 g52780_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_59), .o(n_14658) );
in01s01 g52782_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_60), .o(n_14657) );
in01s01 g52784_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_61), .o(n_14656) );
in01s01 g52786_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_62), .o(n_14655) );
in01s01 g52788_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_63), .o(n_14654) );
in01s01 g52790_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_64), .o(n_14627) );
in01s01 g52792_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_65), .o(n_14653) );
in01s01 g52794_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_66), .o(n_14652) );
in01s01 g52796_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_67), .o(n_14626) );
in01s01 g52798_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_68), .o(n_14651) );
in01s01 g52800_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_50), .o(n_14650) );
in01s01 g52802_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_69), .o(n_14649) );
in01s01 g52804_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_70), .o(n_14648) );
in01s01 g52808_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_72), .o(n_14646) );
in01s01 g52810_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_73), .o(n_14645) );
in01s01 g52812_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_74), .o(n_14644) );
in01s01 g52814_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_75), .o(n_14643) );
in01s01 g52816_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_76), .o(n_14642) );
in01s01 g52818_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_77), .o(n_14641) );
in01s01 g52820_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_78), .o(n_14640) );
in01s01 g52822_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_51), .o(n_14639) );
in01s01 g52824_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_79), .o(n_14638) );
in01s01 g52826_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_80), .o(n_14637) );
in01s01 g52836_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_52), .o(n_14636) );
in01s01 g52838_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_53), .o(n_14635) );
in01s01 g52840_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_54), .o(n_14634) );
in01s01 g52842_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_55), .o(n_14633) );
in01s01 g52844_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_56), .o(n_14625) );
in01s01 g52846_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_57), .o(n_14632) );
in01s01 g52848_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_58), .o(n_14631) );
in01f10 g52853_u0 ( .a(n_10155), .o(n_10256) );
in01f10 g52862_u0 ( .a(n_8935), .o(n_10155) );
in01f06 g52863_u0 ( .a(n_8872), .o(n_8935) );
no02f06 g52864_u0 ( .a(n_17031), .b(n_17032), .o(n_8872) );
na02f02 g52865_u0 ( .a(n_14074), .b(n_14486), .o(g52865_p) );
in01f02 g52865_u1 ( .a(g52865_p), .o(n_14616) );
in01f01 g52866_u0 ( .a(n_14571), .o(n_14572) );
no02s02 g52867_u0 ( .a(n_14386), .b(parity_checker_pci_perr_en_reg), .o(n_14571) );
na02f02 TIMEBOOST_cell_42160 ( .a(TIMEBOOST_net_13318), .b(FE_OFN1374_n_8567), .o(TIMEBOOST_net_12293) );
no02f02 g52869_u0 ( .a(n_14528), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q), .o(n_14620) );
in01f02 g52870_u0 ( .a(n_14490), .o(n_14531) );
ao12f02 g52871_u0 ( .a(n_14487), .b(FE_OFN1709_n_4868), .c(parchk_pci_ad_out_in_1198), .o(n_14490) );
in01f02 g52872_u0 ( .a(n_14489), .o(n_14530) );
ao12f02 g52873_u0 ( .a(n_14487), .b(FE_OFN1709_n_4868), .c(pci_ad_o_31_), .o(n_14489) );
ao12f02 g52874_u0 ( .a(n_14570), .b(n_14518), .c(n_14898), .o(n_14615) );
ao12f02 g52875_u0 ( .a(n_14385), .b(n_12168), .c(n_2629), .o(n_14529) );
in01s01 g52876_u0 ( .a(FE_OFN1705_n_4868), .o(g52876_sb) );
na02f02 TIMEBOOST_cell_42956 ( .a(TIMEBOOST_net_13716), .b(TIMEBOOST_net_493), .o(n_13464) );
no02m04 TIMEBOOST_cell_19040 ( .a(FE_RN_376_0), .b(n_13784), .o(TIMEBOOST_net_4777) );
na02s01 TIMEBOOST_cell_31055 ( .a(TIMEBOOST_net_9438), .b(g64978_db), .o(n_4367) );
in01s01 g52877_u0 ( .a(FE_OFN1705_n_4868), .o(g52877_sb) );
na02s02 TIMEBOOST_cell_45258 ( .a(TIMEBOOST_net_14867), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_12646) );
no02m04 TIMEBOOST_cell_19042 ( .a(FE_RN_373_0), .b(n_13784), .o(TIMEBOOST_net_4778) );
na02s01 TIMEBOOST_cell_31054 ( .a(n_4645), .b(g64978_sb), .o(TIMEBOOST_net_9438) );
in01s01 g52878_u0 ( .a(FE_OFN1705_n_4868), .o(g52878_sb) );
na02s01 TIMEBOOST_cell_45587 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__Q), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_15032) );
no02m04 TIMEBOOST_cell_19044 ( .a(FE_RN_544_0), .b(n_13784), .o(TIMEBOOST_net_4779) );
na02f02 TIMEBOOST_cell_40988 ( .a(TIMEBOOST_net_12732), .b(g57385_sb), .o(n_11359) );
in01s01 g52879_u0 ( .a(n_14389), .o(g52879_sb) );
in01s01 TIMEBOOST_cell_45921 ( .a(wbm_dat_i_1_), .o(TIMEBOOST_net_15228) );
na02f02 TIMEBOOST_cell_43827 ( .a(n_9059), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__Q), .o(TIMEBOOST_net_14152) );
in01s01 TIMEBOOST_cell_32851 ( .a(TIMEBOOST_net_10352), .o(TIMEBOOST_net_10351) );
in01s01 g52880_u0 ( .a(n_14389), .o(g52880_sb) );
na02s02 TIMEBOOST_cell_43581 ( .a(n_3608), .b(n_3609), .o(TIMEBOOST_net_14029) );
na02s01 TIMEBOOST_cell_41964 ( .a(TIMEBOOST_net_13220), .b(g62683_sb), .o(n_6173) );
na02s01 TIMEBOOST_cell_31053 ( .a(TIMEBOOST_net_9437), .b(g64975_db), .o(n_4368) );
in01s01 g52881_u0 ( .a(n_14389), .o(g52881_sb) );
na02s02 TIMEBOOST_cell_44436 ( .a(TIMEBOOST_net_14456), .b(FE_OFN1306_n_13124), .o(TIMEBOOST_net_13421) );
na02s02 TIMEBOOST_cell_45216 ( .a(TIMEBOOST_net_14846), .b(FE_OFN1259_n_4143), .o(TIMEBOOST_net_12068) );
na02s01 TIMEBOOST_cell_31052 ( .a(n_4488), .b(g64975_sb), .o(TIMEBOOST_net_9437) );
no02f02 g52890_u0 ( .a(n_13843), .b(n_14075), .o(n_14486) );
ao12f04 g52891_u0 ( .a(FE_OFN1709_n_4868), .b(n_13787), .c(n_13286), .o(n_14487) );
na02f02 g52892_u0 ( .a(n_13910), .b(n_1196), .o(n_14385) );
oa12f01 g52893_u0 ( .a(n_14073), .b(n_14484), .c(n_15370), .o(n_14528) );
in01f02 g52894_u0 ( .a(n_14104), .o(n_14384) );
na02f02 g52897_u0 ( .a(n_14357), .b(n_7673), .o(n_14383) );
na02f02 g52898_u0 ( .a(n_14355), .b(n_7672), .o(n_14382) );
na02f02 g52899_u0 ( .a(n_14353), .b(n_7671), .o(n_14381) );
na02f02 g52900_u0 ( .a(n_14351), .b(n_7669), .o(n_14380) );
na02f02 g52901_u0 ( .a(n_7667), .b(n_14085), .o(n_14094) );
na02f02 g52902_u0 ( .a(n_14349), .b(n_7666), .o(n_14379) );
na02f02 g52903_u0 ( .a(n_14083), .b(n_7664), .o(n_14093) );
na02f02 g52904_u0 ( .a(n_14347), .b(n_7663), .o(n_14378) );
na02f02 g52905_u0 ( .a(n_7661), .b(n_14341), .o(n_14377) );
na02f02 g52907_u0 ( .a(n_14343), .b(n_7656), .o(n_14375) );
na02f02 g52908_u0 ( .a(n_14337), .b(n_7655), .o(n_14374) );
na02f02 g52909_u0 ( .a(n_14339), .b(n_7654), .o(n_14373) );
na02f02 g52910_u0 ( .a(n_14335), .b(n_7653), .o(n_14372) );
na02f02 g52911_u0 ( .a(n_7652), .b(n_14081), .o(n_14088) );
na02f02 g52912_u0 ( .a(n_14333), .b(n_7651), .o(n_14371) );
na02f02 g52913_u0 ( .a(n_7650), .b(n_14331), .o(n_14370) );
na02f02 g52914_u0 ( .a(n_14329), .b(n_7649), .o(n_14369) );
na02f02 g52915_u0 ( .a(n_7648), .b(n_14327), .o(n_14368) );
na02f02 g52916_u0 ( .a(n_7647), .b(n_14325), .o(n_14367) );
na02f02 g52917_u0 ( .a(n_14323), .b(n_7528), .o(n_14366) );
na02f02 g52918_u0 ( .a(n_14321), .b(n_7646), .o(n_14365) );
na02s02 TIMEBOOST_cell_45788 ( .a(TIMEBOOST_net_15132), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_12038) );
na02f02 g52920_u0 ( .a(n_14319), .b(n_7636), .o(n_14364) );
na02f02 g52921_u0 ( .a(n_7509), .b(n_14315), .o(n_14363) );
na02m02 g52922_u0 ( .a(n_14317), .b(n_7505), .o(n_14362) );
na02f02 g52923_u0 ( .a(n_14313), .b(n_7522), .o(n_14361) );
na02f02 g52924_u0 ( .a(n_14311), .b(n_7521), .o(n_14360) );
na02f02 g52925_u0 ( .a(n_14309), .b(n_7519), .o(n_14359) );
na02m02 g52926_u0 ( .a(n_14357), .b(n_7629), .o(n_14358) );
na02f02 g52927_u0 ( .a(n_14355), .b(n_7518), .o(n_14356) );
na02f02 g52928_u0 ( .a(n_14353), .b(n_7645), .o(n_14354) );
na02m02 g52929_u0 ( .a(n_14085), .b(n_7517), .o(n_14086) );
na02f02 g52930_u0 ( .a(n_14351), .b(n_7643), .o(n_14352) );
na02f02 g52931_u0 ( .a(n_14349), .b(n_7524), .o(n_14350) );
na02f02 g52932_u0 ( .a(n_14083), .b(n_7516), .o(n_14084) );
na02m02 g52933_u0 ( .a(n_14347), .b(n_7515), .o(n_14348) );
na02m02 g52934_u0 ( .a(n_14345), .b(n_7514), .o(n_14346) );
na02m02 g52935_u0 ( .a(n_14343), .b(n_7640), .o(n_14344) );
na02m02 g52936_u0 ( .a(n_14341), .b(n_7525), .o(n_14342) );
na02m02 g52937_u0 ( .a(n_14339), .b(n_7665), .o(n_14340) );
na02f02 g52938_u0 ( .a(n_14337), .b(n_7639), .o(n_14338) );
na02m02 g52939_u0 ( .a(n_14335), .b(n_7532), .o(n_14336) );
na02m02 g52940_u0 ( .a(n_14081), .b(n_7513), .o(n_14082) );
na02f02 g52941_u0 ( .a(n_14333), .b(n_7512), .o(n_14334) );
na02m02 g52942_u0 ( .a(n_14331), .b(n_7534), .o(n_14332) );
na02f02 g52943_u0 ( .a(n_14329), .b(n_7535), .o(n_14330) );
na02f02 g52944_u0 ( .a(n_7511), .b(n_14327), .o(n_14328) );
na02m02 g52945_u0 ( .a(n_14325), .b(n_7638), .o(n_14326) );
na02f02 g52946_u0 ( .a(n_14323), .b(n_7510), .o(n_14324) );
na02f02 g52947_u0 ( .a(n_14321), .b(n_7637), .o(n_14322) );
na02s01 g52948_u0 ( .a(n_7735), .b(parchk_pci_serr_en_in), .o(n_14080) );
na02f02 g52949_u0 ( .a(n_14319), .b(n_7634), .o(n_14320) );
na02s01 TIMEBOOST_cell_36403 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(g65776_sb), .o(TIMEBOOST_net_10440) );
na02f02 g52951_u0 ( .a(n_14317), .b(n_7632), .o(n_14318) );
na02f02 g52952_u0 ( .a(n_7633), .b(n_14315), .o(n_14316) );
na02f02 g52953_u0 ( .a(n_14313), .b(n_7631), .o(n_14314) );
na02f02 g52954_u0 ( .a(n_14311), .b(n_7630), .o(n_14312) );
na02f02 g52955_u0 ( .a(n_14309), .b(n_7628), .o(n_14310) );
ao12f02 g52956_u0 ( .a(n_8595), .b(n_1979), .c(n_7567), .o(n_10792) );
ao12f02 g52957_u0 ( .a(n_14898), .b(n_14890), .c(n_112), .o(n_14570) );
na03f02 g52966_u0 ( .a(n_16611), .b(n_14283), .c(n_16610), .o(n_14607) );
na02f02 g52990_u0 ( .a(n_14521), .b(n_14539), .o(n_14583) );
na03f02 g52991_u0 ( .a(n_16615), .b(n_14413), .c(n_16614), .o(n_14582) );
na02m02 TIMEBOOST_cell_45789 ( .a(n_4085), .b(n_7618), .o(TIMEBOOST_net_15133) );
na02m20 g52_u0 ( .a(pciu_am1_in_528), .b(pciu_bar1_in_390), .o(g52_p) );
in01f08 g52_u1 ( .a(g52_p), .o(n_15598) );
in01s01 g53004_u0 ( .a(parchk_pci_perr_out_in), .o(n_14079) );
na02f02 g53010_u0 ( .a(n_14484), .b(n_1684), .o(n_14618) );
no02f02 g53011_u0 ( .a(n_13731), .b(FE_OFN1709_n_4868), .o(g53011_p) );
in01f02 g53011_u1 ( .a(g53011_p), .o(n_14085) );
na02s02 TIMEBOOST_cell_42124 ( .a(TIMEBOOST_net_13300), .b(FE_OFN1311_n_6624), .o(TIMEBOOST_net_11593) );
in01f02 g53012_u1 ( .a(g53012_p), .o(n_14341) );
no02f02 g53014_u0 ( .a(n_13776), .b(FE_OFN1710_n_4868), .o(g53014_p) );
in01f02 g53014_u1 ( .a(g53014_p), .o(n_14343) );
no02f02 g53015_u0 ( .a(n_13775), .b(FE_OFN1709_n_4868), .o(g53015_p) );
in01f02 g53015_u1 ( .a(g53015_p), .o(n_14337) );
no02f02 g53016_u0 ( .a(n_13774), .b(FE_OFN1709_n_4868), .o(g53016_p) );
in01f02 g53016_u1 ( .a(g53016_p), .o(n_14339) );
na03s02 TIMEBOOST_cell_5674 ( .a(n_4479), .b(g64807_sb), .c(g64807_db), .o(n_4462) );
in01f02 g53017_u1 ( .a(g53017_p), .o(n_14335) );
no02f02 g53018_u0 ( .a(n_13728), .b(FE_OFN1709_n_4868), .o(g53018_p) );
in01f02 g53018_u1 ( .a(g53018_p), .o(n_14081) );
no02f02 g53019_u0 ( .a(n_14481), .b(n_14302), .o(n_14569) );
no02f02 g53020_u0 ( .a(n_14300), .b(n_14479), .o(n_16594) );
no02f02 g53021_u0 ( .a(n_14298), .b(n_14477), .o(n_14567) );
no02f02 g53022_u0 ( .a(n_13772), .b(FE_OFN1705_n_4868), .o(g53022_p) );
in01f02 g53022_u1 ( .a(g53022_p), .o(n_14333) );
no02f02 g53023_u0 ( .a(n_14295), .b(n_14476), .o(n_14566) );
no02f02 g53024_u0 ( .a(n_14474), .b(n_14293), .o(n_14565) );
no02f02 g53025_u0 ( .a(n_14291), .b(n_14472), .o(n_14564) );
no02f02 g53026_u0 ( .a(n_13756), .b(FE_OFN1705_n_4868), .o(g53026_p) );
in01f02 g53026_u1 ( .a(g53026_p), .o(n_14331) );
no02f02 g53028_u0 ( .a(n_14469), .b(n_14285), .o(n_14563) );
no02f02 g53029_u0 ( .a(n_14284), .b(n_14467), .o(n_16611) );
no02f02 g53031_u0 ( .a(n_13771), .b(FE_OFN1710_n_4868), .o(g53031_p) );
in01f02 g53031_u1 ( .a(g53031_p), .o(n_14329) );
no02f02 g53033_u0 ( .a(n_14462), .b(n_14277), .o(n_14560) );
no02f02 g53034_u0 ( .a(n_14274), .b(n_14461), .o(n_14559) );
no02f02 g53035_u0 ( .a(n_13770), .b(FE_OFN1705_n_4868), .o(g53035_p) );
in01f02 g53035_u1 ( .a(g53035_p), .o(n_14327) );
no02f02 g53036_u0 ( .a(n_14459), .b(n_14458), .o(n_14558) );
no02f02 g53037_u0 ( .a(n_14457), .b(n_14270), .o(n_14557) );
no02f02 g53039_u0 ( .a(n_13755), .b(FE_OFN1705_n_4868), .o(g53039_p) );
in01f02 g53039_u1 ( .a(g53039_p), .o(n_14325) );
no02f02 g53041_u0 ( .a(n_14451), .b(n_14264), .o(n_14554) );
no02f02 g53042_u0 ( .a(n_14448), .b(n_14449), .o(n_16623) );
no02f02 g53044_u0 ( .a(n_14260), .b(n_14447), .o(n_16625) );
no02f02 g53045_u0 ( .a(n_14444), .b(n_14445), .o(n_14551) );
no02f02 g53046_u0 ( .a(n_14256), .b(n_14443), .o(n_14550) );
no02f02 g53047_u0 ( .a(n_14254), .b(n_14441), .o(n_14549) );
no02f02 g53048_u0 ( .a(n_14439), .b(n_14252), .o(n_14548) );
no02f02 g53049_u0 ( .a(n_14437), .b(n_14436), .o(n_14547) );
no02f02 g53051_u0 ( .a(n_14432), .b(n_14514), .o(n_14545) );
no02f02 g53052_u0 ( .a(n_14512), .b(n_14430), .o(n_14544) );
no02f02 g53053_u0 ( .a(n_14510), .b(n_14428), .o(n_14543) );
no02f02 g53056_u0 ( .a(n_14422), .b(n_14508), .o(n_14541) );
no02f02 g53060_u0 ( .a(n_14416), .b(n_14415), .o(n_14521) );
no02f02 g53061_u0 ( .a(n_14414), .b(n_14504), .o(n_16615) );
no02f02 g53063_u0 ( .a(n_14500), .b(n_14410), .o(n_14536) );
no02f02 g53064_u0 ( .a(n_14408), .b(n_14498), .o(n_14535) );
no02f02 g53066_u0 ( .a(n_14403), .b(n_14495), .o(n_14534) );
no02f02 g53067_u0 ( .a(n_14401), .b(n_14493), .o(n_16617) );
no02f02 g53068_u0 ( .a(n_13767), .b(n_13332), .o(n_14386) );
no02f02 g53069_u0 ( .a(n_2446), .b(n_8524), .o(g53069_p) );
in01f02 g53069_u1 ( .a(g53069_p), .o(n_8595) );
na02s01 TIMEBOOST_cell_43273 ( .a(n_3531), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__Q), .o(TIMEBOOST_net_13875) );
no02f03 g53071_u0 ( .a(n_14303), .b(n_14518), .o(g53071_p) );
in01f02 g53071_u1 ( .a(g53071_p), .o(n_14902) );
no02f02 g53072_u0 ( .a(n_14307), .b(n_14518), .o(g53072_p) );
in01f02 g53072_u1 ( .a(g53072_p), .o(n_14517) );
no02f04 g53073_u0 ( .a(n_13764), .b(FE_OFN1708_n_4868), .o(g53073_p) );
in01f02 g53073_u1 ( .a(g53073_p), .o(n_14315) );
no02f04 g53074_u0 ( .a(n_13761), .b(FE_OFN1708_n_4868), .o(g53074_p) );
in01f02 g53074_u1 ( .a(g53074_p), .o(n_14313) );
no02f04 g53075_u0 ( .a(n_13760), .b(FE_OFN1707_n_4868), .o(g53075_p) );
in01f02 g53075_u1 ( .a(g53075_p), .o(n_14311) );
no02f02 g53076_u0 ( .a(n_13759), .b(FE_OFN1706_n_4868), .o(g53076_p) );
in01f02 g53076_u1 ( .a(g53076_p), .o(n_14309) );
na02f02 TIMEBOOST_cell_43771 ( .a(n_9558), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__Q), .o(TIMEBOOST_net_14124) );
in01f02 g53077_u1 ( .a(g53077_p), .o(n_14317) );
na02f02 TIMEBOOST_cell_22617 ( .a(TIMEBOOST_net_6565), .b(FE_OFN1565_n_12502), .o(n_12700) );
in01f02 g53078_u1 ( .a(g53078_p), .o(n_14357) );
no02f02 g53079_u0 ( .a(n_13785), .b(FE_OFN1706_n_4868), .o(g53079_p) );
in01f02 g53079_u1 ( .a(g53079_p), .o(n_14355) );
no02f02 g53080_u0 ( .a(n_13783), .b(FE_OFN1706_n_4868), .o(g53080_p) );
in01f02 g53080_u1 ( .a(g53080_p), .o(n_14353) );
no02f02 g53082_u0 ( .a(n_13780), .b(FE_OFN1706_n_4868), .o(g53082_p) );
in01f02 g53082_u1 ( .a(g53082_p), .o(n_14349) );
no02f02 g53083_u0 ( .a(n_13729), .b(FE_OFN1706_n_4868), .o(g53083_p) );
in01f02 g53083_u1 ( .a(g53083_p), .o(n_14083) );
na02s01 TIMEBOOST_cell_42989 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__Q), .b(n_3205), .o(TIMEBOOST_net_13733) );
in01f02 g53084_u1 ( .a(g53084_p), .o(n_14347) );
na02f02 g53085_u0 ( .a(n_13829), .b(n_7658), .o(n_13831) );
na02f02 g53086_u0 ( .a(n_14076), .b(n_7657), .o(n_14078) );
no02f04 g53087_u0 ( .a(n_13768), .b(FE_OFN1708_n_4868), .o(g53087_p) );
in01f02 g53087_u1 ( .a(g53087_p), .o(n_14321) );
na02m02 g53088_u0 ( .a(n_13753), .b(n_1112), .o(n_14392) );
na02f02 g53089_u0 ( .a(n_13752), .b(n_1108), .o(n_14390) );
na02f02 g53090_u0 ( .a(n_13750), .b(n_1202), .o(n_14387) );
na02f02 g53091_u0 ( .a(n_13907), .b(n_7523), .o(n_13911) );
na02m02 g53092_u0 ( .a(n_13829), .b(n_7642), .o(n_13830) );
na02f02 g53093_u0 ( .a(n_7527), .b(n_14076), .o(n_14077) );
ao12f02 g53094_u0 ( .a(n_1551), .b(n_13749), .c(FE_OCPN1836_n_16798), .o(n_13910) );
na02s01 TIMEBOOST_cell_42990 ( .a(TIMEBOOST_net_13733), .b(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_11444) );
no02s01 g53096_u0 ( .a(n_4796), .b(n_14484), .o(n_14483) );
na02f02 g53097_u0 ( .a(n_13907), .b(n_7635), .o(n_13908) );
no02f02 g53098_u0 ( .a(n_13765), .b(FE_OFN1708_n_4868), .o(g53098_p) );
in01f02 g53098_u1 ( .a(g53098_p), .o(n_14319) );
ao12f02 g53099_u0 ( .a(n_1551), .b(n_2619), .c(n_13819), .o(n_14075) );
ao12f02 g53102_u0 ( .a(n_13592), .b(n_13671), .c(n_13784), .o(n_13785) );
ao12f02 g53103_u0 ( .a(n_13591), .b(n_13670), .c(n_13781), .o(n_13783) );
na03s02 TIMEBOOST_cell_33585 ( .a(TIMEBOOST_net_9558), .b(n_5633), .c(g62134_sb), .o(n_5559) );
na03s02 TIMEBOOST_cell_36287 ( .a(n_1350), .b(n_1433), .c(n_1352), .o(TIMEBOOST_net_10382) );
na03s02 TIMEBOOST_cell_33584 ( .a(TIMEBOOST_net_9559), .b(n_5633), .c(g62132_sb), .o(n_5563) );
ao12f02 g53106_u0 ( .a(n_13587), .b(n_13668), .c(n_13784), .o(n_13780) );
ao12f02 g53107_u0 ( .a(n_13585), .b(n_13562), .c(n_13784), .o(n_13729) );
ao12f02 g53111_u0 ( .a(n_13581), .b(n_13664), .c(FE_OFN1946_n_13784), .o(n_13776) );
ao12f02 g53112_u0 ( .a(n_13579), .b(n_13663), .c(n_13781), .o(n_13775) );
ao12f02 g53113_u0 ( .a(n_13578), .b(n_13662), .c(FE_OFN969_n_13784), .o(n_13774) );
ao12f02 g53115_u0 ( .a(n_13576), .b(n_13560), .c(n_13763), .o(n_13728) );
ao12f02 g53116_u0 ( .a(n_13575), .b(n_13659), .c(FE_OFN1946_n_13784), .o(n_13772) );
ao12f02 g53117_u0 ( .a(n_13574), .b(n_13658), .c(FE_OFN1946_n_13784), .o(n_13771) );
ao12f02 g53118_u0 ( .a(n_13573), .b(n_13657), .c(n_13784), .o(n_13770) );
ao12f01 g53121_u0 ( .a(n_16331), .b(n_13810), .c(n_7310), .o(n_14074) );
na02f02 g53122_u0 ( .a(n_13716), .b(n_13766), .o(n_13767) );
na02f02 g53123_u0 ( .a(n_13716), .b(n_13333), .o(n_13918) );
na02f02 g53124_u0 ( .a(n_13716), .b(n_7396), .o(n_13917) );
no02f02 g53125_u0 ( .a(n_1100), .b(n_13748), .o(n_13828) );
no02s01 g53126_u0 ( .a(n_14305), .b(wbm_cti_o_1_), .o(n_14307) );
ao12f02 g53127_u0 ( .a(n_13569), .b(n_13653), .c(n_13784), .o(n_13765) );
no02s02 g53129_u0 ( .a(n_13844), .b(n_15371), .o(n_14484) );
ao12f02 g53133_u0 ( .a(n_13678), .b(n_13673), .c(n_13784), .o(n_13759) );
ao12f02 g53134_u0 ( .a(n_13680), .b(n_13754), .c(n_13561), .o(n_13829) );
ao12f02 g53135_u0 ( .a(n_13582), .b(n_13754), .c(n_13704), .o(n_14076) );
in01f01 g53136_u0 ( .a(n_13757), .o(n_13758) );
no02f01 g53137_u0 ( .a(n_13715), .b(n_7397), .o(n_13757) );
ao12f02 g53138_u0 ( .a(n_13722), .b(n_13334), .c(n_13721), .o(n_13756) );
ao12f02 g53139_u0 ( .a(FE_OFN1335_n_13720), .b(n_13414), .c(n_13721), .o(n_13755) );
ao12f02 g53140_u0 ( .a(n_1522), .b(n_7043), .c(n_7726), .o(n_8524) );
no02f02 g53141_u0 ( .a(n_13412), .b(n_14305), .o(g53141_p) );
in01f02 g53141_u1 ( .a(g53141_p), .o(n_14306) );
no02f02 g53142_u0 ( .a(n_13411), .b(n_14305), .o(g53142_p) );
in01f02 g53142_u1 ( .a(g53142_p), .o(n_14304) );
na02f02 TIMEBOOST_cell_45805 ( .a(n_9444), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__Q), .o(TIMEBOOST_net_15141) );
oa12s02 g53145_u0 ( .a(n_6941), .b(n_13691), .c(n_13825), .o(n_13827) );
oa12s02 g53146_u0 ( .a(n_6940), .b(n_13689), .c(n_13825), .o(n_13826) );
oa12s02 g53147_u0 ( .a(n_6942), .b(n_13692), .c(n_13825), .o(n_13824) );
oa12m02 g53148_u0 ( .a(n_14305), .b(n_14965), .c(n_3164), .o(n_14303) );
in01m02 g53149_u0 ( .a(n_14890), .o(n_14482) );
ao12m04 g53150_u0 ( .a(n_14305), .b(n_824), .c(wbm_cyc_o_1378), .o(n_14890) );
na02f02 g53152_u0 ( .a(n_14069), .b(n_13906), .o(n_14302) );
na02s02 TIMEBOOST_cell_40857 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__Q), .b(n_13179), .o(TIMEBOOST_net_12667) );
in01f02 g53154_u1 ( .a(g53154_p), .o(n_14301) );
na02f02 TIMEBOOST_cell_41062 ( .a(TIMEBOOST_net_12769), .b(g57228_sb), .o(n_11528) );
in01f02 g53155_u1 ( .a(g53155_p), .o(n_14480) );
na02m02 TIMEBOOST_cell_32444 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__Q), .o(TIMEBOOST_net_10133) );
na02s02 TIMEBOOST_cell_45259 ( .a(n_4278), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__Q), .o(TIMEBOOST_net_14868) );
na02s02 TIMEBOOST_cell_32025 ( .a(TIMEBOOST_net_9923), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4905) );
in01f02 g53158_u1 ( .a(g53158_p), .o(n_16595) );
na02s02 TIMEBOOST_cell_40856 ( .a(TIMEBOOST_net_12666), .b(FE_OFN1327_n_13547), .o(TIMEBOOST_net_11622) );
in01f02 g53159_u1 ( .a(g53159_p), .o(n_14478) );
na02s01 TIMEBOOST_cell_32042 ( .a(configuration_pci_err_addr_499), .b(wbm_adr_o_29_), .o(TIMEBOOST_net_9932) );
na02f02 g53161_u0 ( .a(n_14243), .b(n_14245), .o(n_14477) );
na02s02 TIMEBOOST_cell_40859 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__Q), .b(n_13185), .o(TIMEBOOST_net_12668) );
in01f02 g53163_u1 ( .a(g53163_p), .o(n_14296) );
na02m02 TIMEBOOST_cell_40858 ( .a(TIMEBOOST_net_12667), .b(FE_OFN1331_n_13547), .o(TIMEBOOST_net_11608) );
na02f02 g53165_u0 ( .a(n_14005), .b(n_14007), .o(n_14295) );
na02f02 TIMEBOOST_cell_41056 ( .a(TIMEBOOST_net_12766), .b(g57534_sb), .o(n_11208) );
in01f02 g53167_u1 ( .a(g53167_p), .o(n_14475) );
na02s01 TIMEBOOST_cell_40843 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__Q), .b(n_13173), .o(TIMEBOOST_net_12660) );
na02f02 g53169_u0 ( .a(n_14004), .b(n_14002), .o(n_14293) );
in01f02 g53170_u1 ( .a(g53170_p), .o(n_14292) );
na02m02 TIMEBOOST_cell_32442 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__Q), .o(TIMEBOOST_net_10132) );
in01f02 g53171_u1 ( .a(g53171_p), .o(n_14473) );
in01s01 TIMEBOOST_cell_45946 ( .a(TIMEBOOST_net_15252), .o(TIMEBOOST_net_15253) );
na02f02 g53173_u0 ( .a(n_14061), .b(n_13899), .o(n_14291) );
na02s01 TIMEBOOST_cell_40845 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__Q), .b(n_13186), .o(TIMEBOOST_net_12661) );
in01f02 g53174_u1 ( .a(g53174_p), .o(n_14290) );
na02f02 TIMEBOOST_cell_41058 ( .a(TIMEBOOST_net_12767), .b(g57252_sb), .o(n_11503) );
in01f02 g53175_u1 ( .a(g53175_p), .o(n_14471) );
na02s02 TIMEBOOST_cell_40827 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__Q), .b(n_13170), .o(TIMEBOOST_net_12652) );
na02f02 g53181_u0 ( .a(n_13992), .b(n_13994), .o(n_14285) );
in01f02 g53182_u1 ( .a(g53182_p), .o(n_14286) );
na02m02 TIMEBOOST_cell_32440 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__Q), .o(TIMEBOOST_net_10131) );
in01f02 g53183_u1 ( .a(g53183_p), .o(n_14468) );
na02m02 TIMEBOOST_cell_42525 ( .a(n_16945), .b(n_4078), .o(TIMEBOOST_net_13501) );
na02s01 TIMEBOOST_cell_36290 ( .a(TIMEBOOST_net_10383), .b(g67057_sb), .o(n_1640) );
in01f02 g53187_u1 ( .a(g53187_p), .o(n_16610) );
na02f02 TIMEBOOST_cell_41064 ( .a(TIMEBOOST_net_12770), .b(g57053_sb), .o(n_11683) );
na02f02 g53197_u0 ( .a(n_14225), .b(n_14223), .o(n_14462) );
na02s01 TIMEBOOST_cell_40847 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__Q), .b(n_13183), .o(TIMEBOOST_net_12662) );
in01f02 g53199_u1 ( .a(g53199_p), .o(n_14275) );
na02m02 TIMEBOOST_cell_41838 ( .a(TIMEBOOST_net_13157), .b(g54140_sb), .o(n_13460) );
na02s01 TIMEBOOST_cell_36274 ( .a(TIMEBOOST_net_10375), .b(FE_OFN988_n_574), .o(n_1483) );
na02f02 TIMEBOOST_cell_41060 ( .a(TIMEBOOST_net_12768), .b(g57038_sb), .o(n_11695) );
in01f02 g53203_u1 ( .a(g53203_p), .o(n_14460) );
na02s02 TIMEBOOST_cell_40841 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__Q), .b(n_13163), .o(TIMEBOOST_net_12659) );
na02f02 g53205_u0 ( .a(n_14049), .b(n_14220), .o(n_14458) );
in01f02 g53206_u1 ( .a(g53206_p), .o(n_14272) );
in01s01 TIMEBOOST_cell_45947 ( .a(wbm_dat_i_31_), .o(TIMEBOOST_net_15254) );
in01f02 g53207_u1 ( .a(g53207_p), .o(n_14271) );
na02s02 TIMEBOOST_cell_40831 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__Q), .b(n_13167), .o(TIMEBOOST_net_12654) );
na02f02 g53209_u0 ( .a(n_13973), .b(n_13974), .o(n_14270) );
na02m02 TIMEBOOST_cell_32438 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__Q), .o(TIMEBOOST_net_10130) );
in01f02 g53210_u1 ( .a(g53210_p), .o(n_14456) );
na02f02 TIMEBOOST_cell_41644 ( .a(FE_OFN1436_n_9372), .b(TIMEBOOST_net_13060), .o(TIMEBOOST_net_11673) );
in01f02 g53211_u1 ( .a(g53211_p), .o(n_14269) );
na02s01 TIMEBOOST_cell_30874 ( .a(pci_target_unit_pcit_if_strd_addr_in_711), .b(pci_target_unit_del_sync_addr_in_229), .o(TIMEBOOST_net_9348) );
na02f02 TIMEBOOST_cell_41034 ( .a(TIMEBOOST_net_12755), .b(g57407_sb), .o(n_10366) );
in01f02 g53214_u1 ( .a(g53214_p), .o(n_14454) );
na02m04 TIMEBOOST_cell_32494 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__Q), .o(TIMEBOOST_net_10158) );
na02s02 TIMEBOOST_cell_40830 ( .a(TIMEBOOST_net_12653), .b(FE_OFN1332_n_13547), .o(TIMEBOOST_net_11611) );
na02f02 g53223_u0 ( .a(n_16613), .b(n_16612), .o(g53223_p) );
na02m02 TIMEBOOST_cell_32436 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__Q), .o(TIMEBOOST_net_10129) );
na02s02 TIMEBOOST_cell_36292 ( .a(TIMEBOOST_net_10384), .b(n_1166), .o(n_2231) );
na02m02 TIMEBOOST_cell_32478 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__Q), .o(TIMEBOOST_net_10150) );
in01f02 g53226_u1 ( .a(g53226_p), .o(n_16622) );
na02f02 g53228_u0 ( .a(n_14205), .b(n_14203), .o(n_14447) );
na02s02 TIMEBOOST_cell_40837 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__Q), .b(n_13162), .o(TIMEBOOST_net_12657) );
na02s01 TIMEBOOST_cell_31974 ( .a(configuration_pci_err_data_523), .b(wbm_dat_o_22_), .o(TIMEBOOST_net_9898) );
in01f02 g53230_u1 ( .a(g53230_p), .o(n_16624) );
na02s02 TIMEBOOST_cell_40836 ( .a(TIMEBOOST_net_12656), .b(FE_OFN1330_n_13547), .o(TIMEBOOST_net_11605) );
in01f02 g53231_u1 ( .a(g53231_p), .o(n_14446) );
na02f02 g53232_u0 ( .a(n_14201), .b(n_14202), .o(n_14445) );
na02s02 TIMEBOOST_cell_40850 ( .a(TIMEBOOST_net_12663), .b(FE_OFN1331_n_13547), .o(TIMEBOOST_net_11619) );
na02f02 TIMEBOOST_cell_41092 ( .a(TIMEBOOST_net_12784), .b(g57357_sb), .o(n_10386) );
in01f02 g53234_u1 ( .a(g53234_p), .o(n_14258) );
na02f02 TIMEBOOST_cell_32336 ( .a(n_8527), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(TIMEBOOST_net_10079) );
in01f02 g53235_u1 ( .a(g53235_p), .o(n_14257) );
na02f10 TIMEBOOST_cell_36242 ( .a(TIMEBOOST_net_10359), .b(g67048_db), .o(n_1211) );
in01s01 TIMEBOOST_cell_45948 ( .a(TIMEBOOST_net_15254), .o(TIMEBOOST_net_15255) );
na02s01 TIMEBOOST_cell_32004 ( .a(configuration_pci_err_addr_476), .b(wbm_adr_o_6_), .o(TIMEBOOST_net_9913) );
in01f02 g53238_u1 ( .a(g53238_p), .o(n_14255) );
na02f02 TIMEBOOST_cell_41036 ( .a(TIMEBOOST_net_12756), .b(g57401_sb), .o(n_11342) );
in01f02 g53239_u1 ( .a(g53239_p), .o(n_14442) );
na02s08 TIMEBOOST_cell_36244 ( .a(TIMEBOOST_net_10360), .b(n_1416), .o(TIMEBOOST_net_92) );
na02s02 TIMEBOOST_cell_40716 ( .a(TIMEBOOST_net_12596), .b(g62922_sb), .o(n_6037) );
na02m02 TIMEBOOST_cell_32434 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__Q), .o(TIMEBOOST_net_10128) );
in01f02 g53242_u1 ( .a(g53242_p), .o(n_14440) );
na02f02 TIMEBOOST_cell_41038 ( .a(TIMEBOOST_net_12757), .b(g57110_sb), .o(n_11637) );
in01f02 g53243_u1 ( .a(g53243_p), .o(n_14253) );
na02m02 TIMEBOOST_cell_32472 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__Q), .o(TIMEBOOST_net_10147) );
na02f20 TIMEBOOST_cell_36246 ( .a(TIMEBOOST_net_10361), .b(n_15680), .o(FE_RN_299_0) );
na02s01 TIMEBOOST_cell_40441 ( .a(conf_wb_err_addr_in_969), .b(configuration_wb_err_addr_560), .o(TIMEBOOST_net_12459) );
na02f02 g53249_u0 ( .a(n_14194), .b(n_14195), .o(n_14436) );
na02s02 TIMEBOOST_cell_40440 ( .a(TIMEBOOST_net_12458), .b(g62087_sb), .o(TIMEBOOST_net_11373) );
in01f02 g53250_u1 ( .a(g53250_p), .o(n_14250) );
na02s02 TIMEBOOST_cell_37997 ( .a(pci_target_unit_pcit_if_strd_addr_in_698), .b(g52627_sb), .o(TIMEBOOST_net_11237) );
in01f02 g53251_u1 ( .a(g53251_p), .o(n_14435) );
na02f02 g53253_u0 ( .a(n_14033), .b(n_13878), .o(n_14434) );
na02m02 TIMEBOOST_cell_32432 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__Q), .o(TIMEBOOST_net_10127) );
in01f02 g53254_u1 ( .a(g53254_p), .o(n_14515) );
na02s01 TIMEBOOST_cell_40443 ( .a(conf_wb_err_addr_in_945), .b(configuration_wb_err_addr_536), .o(TIMEBOOST_net_12460) );
in01f02 g53255_u1 ( .a(g53255_p), .o(n_14433) );
na02s02 TIMEBOOST_cell_40442 ( .a(TIMEBOOST_net_12459), .b(g62129_sb), .o(TIMEBOOST_net_11375) );
na02f02 g53257_u0 ( .a(n_13953), .b(n_13954), .o(n_14432) );
na02f02 TIMEBOOST_cell_41066 ( .a(TIMEBOOST_net_12771), .b(g57437_sb), .o(n_11297) );
in01f02 g53258_u1 ( .a(g53258_p), .o(n_14431) );
na02f02 TIMEBOOST_cell_41040 ( .a(TIMEBOOST_net_12758), .b(g57108_sb), .o(n_11638) );
in01f02 g53259_u1 ( .a(g53259_p), .o(n_14513) );
na02f08 TIMEBOOST_cell_36248 ( .a(TIMEBOOST_net_10362), .b(n_16696), .o(n_16286) );
na02s01 TIMEBOOST_cell_44898 ( .a(TIMEBOOST_net_14687), .b(g65738_da), .o(TIMEBOOST_net_10975) );
na02m02 TIMEBOOST_cell_32430 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__Q), .o(TIMEBOOST_net_10126) );
in01f02 g53262_u1 ( .a(g53262_p), .o(n_14511) );
na02f02 TIMEBOOST_cell_41042 ( .a(TIMEBOOST_net_12759), .b(g57414_sb), .o(n_11328) );
in01f02 g53263_u1 ( .a(g53263_p), .o(n_14429) );
na02m02 TIMEBOOST_cell_32428 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__Q), .o(TIMEBOOST_net_10125) );
ao22m02 g53265_u0 ( .a(n_13555), .b(n_13447), .c(FE_OFN1618_n_1787), .d(conf_wb_err_bc_in), .o(n_13753) );
na02f02 g53266_u0 ( .a(n_13875), .b(n_14029), .o(n_14428) );
na02s01 TIMEBOOST_cell_40692 ( .a(TIMEBOOST_net_12584), .b(g62361_sb), .o(n_6876) );
in01f02 g53267_u1 ( .a(g53267_p), .o(n_14427) );
na02s02 TIMEBOOST_cell_40444 ( .a(TIMEBOOST_net_12460), .b(g62135_sb), .o(TIMEBOOST_net_11376) );
in01f02 g53268_u1 ( .a(g53268_p), .o(n_14426) );
na02f02 TIMEBOOST_cell_41044 ( .a(TIMEBOOST_net_12760), .b(g57092_sb), .o(n_11650) );
na02f02 g53274_u0 ( .a(n_13942), .b(n_13943), .o(n_14422) );
na02m02 TIMEBOOST_cell_45790 ( .a(TIMEBOOST_net_15133), .b(g59804_da), .o(n_7620) );
in01f02 g53275_u1 ( .a(g53275_p), .o(n_14421) );
na02m02 TIMEBOOST_cell_32426 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q), .o(TIMEBOOST_net_10124) );
in01f02 g53276_u1 ( .a(g53276_p), .o(n_14420) );
na02f02 TIMEBOOST_cell_32425 ( .a(n_13873), .b(TIMEBOOST_net_10123), .o(TIMEBOOST_net_6271) );
na02m04 TIMEBOOST_cell_32326 ( .a(g57790_sb), .b(TIMEBOOST_net_10324), .o(TIMEBOOST_net_10074) );
ao22f02 g53281_u0 ( .a(n_13554), .b(n_13447), .c(FE_OFN1618_n_1787), .d(conf_wb_err_bc_in_847), .o(n_13752) );
na02f02 g53283_u0 ( .a(n_14177), .b(n_14178), .o(n_14505) );
na02m02 TIMEBOOST_cell_32470 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__Q), .o(TIMEBOOST_net_10146) );
na02s01 TIMEBOOST_cell_36250 ( .a(TIMEBOOST_net_10363), .b(g54160_sb), .o(TIMEBOOST_net_1010) );
na02f02 TIMEBOOST_cell_41068 ( .a(TIMEBOOST_net_12772), .b(g57334_sb), .o(n_10396) );
na03s02 TIMEBOOST_cell_5532 ( .a(n_4470), .b(g65065_sb), .c(g65065_db), .o(n_4315) );
na02s01 TIMEBOOST_cell_44899 ( .a(n_2211), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__Q), .o(TIMEBOOST_net_14688) );
in01f02 g53288_u1 ( .a(g53288_p), .o(n_14413) );
na02m02 TIMEBOOST_cell_39352 ( .a(FE_OFN1150_n_13249), .b(TIMEBOOST_net_11914), .o(TIMEBOOST_net_4288) );
in01f02 g53289_u1 ( .a(g53289_p), .o(n_16614) );
ao22f02 g53290_u0 ( .a(n_13553), .b(n_13447), .c(FE_OFN1618_n_1787), .d(conf_wb_err_bc_in_848), .o(n_13750) );
na02m02 TIMEBOOST_cell_32468 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__16__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__16__Q), .o(TIMEBOOST_net_10145) );
na02f02 g53296_u0 ( .a(n_14020), .b(n_14172), .o(n_14500) );
na02s02 TIMEBOOST_cell_39568 ( .a(TIMEBOOST_net_12022), .b(g62976_sb), .o(n_5930) );
in01f02 g53298_u1 ( .a(g53298_p), .o(n_14499) );
na02f02 g53299_u0 ( .a(n_14170), .b(n_14171), .o(n_14498) );
na02f02 TIMEBOOST_cell_41070 ( .a(TIMEBOOST_net_12773), .b(g57243_sb), .o(n_11515) );
na02s01 TIMEBOOST_cell_44900 ( .a(TIMEBOOST_net_14688), .b(FE_OFN714_n_8140), .o(TIMEBOOST_net_11084) );
in01f02 g53301_u1 ( .a(g53301_p), .o(n_14407) );
na02s02 TIMEBOOST_cell_39570 ( .a(TIMEBOOST_net_12023), .b(g62429_sb), .o(n_6741) );
in01f02 g53302_u1 ( .a(g53302_p), .o(n_14497) );
na02m02 TIMEBOOST_cell_32466 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q), .o(TIMEBOOST_net_10144) );
na02f02 g53308_u0 ( .a(n_14166), .b(n_14167), .o(n_14495) );
in01f02 g53310_u1 ( .a(g53310_p), .o(n_14494) );
na02f02 g53311_u0 ( .a(n_14016), .b(n_13863), .o(n_14401) );
na02m02 TIMEBOOST_cell_32424 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__Q), .o(TIMEBOOST_net_10123) );
in01f02 g53314_u1 ( .a(g53314_p), .o(n_16616) );
na02s02 TIMEBOOST_cell_45607 ( .a(TIMEBOOST_net_9360), .b(FE_OFN789_n_2678), .o(TIMEBOOST_net_15042) );
na02s02 TIMEBOOST_cell_43165 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__Q), .b(n_3750), .o(TIMEBOOST_net_13821) );
na02f02 g53387_u0 ( .a(n_13903), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__Q), .o(n_13906) );
na02f02 g53388_u0 ( .a(FE_OFN1596_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__Q), .o(n_14069) );
na02f02 TIMEBOOST_cell_41046 ( .a(TIMEBOOST_net_12761), .b(g57061_sb), .o(n_10506) );
na02s02 TIMEBOOST_cell_42814 ( .a(TIMEBOOST_net_13645), .b(g65284_db), .o(n_3582) );
na02m02 TIMEBOOST_cell_32422 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__Q), .o(TIMEBOOST_net_10122) );
na02s01 TIMEBOOST_cell_36345 ( .a(TIMEBOOST_net_9299), .b(n_2520), .o(TIMEBOOST_net_10411) );
na02s02 TIMEBOOST_cell_32041 ( .a(TIMEBOOST_net_9931), .b(FE_OFN1183_n_3476), .o(TIMEBOOST_net_4913) );
na02s01 TIMEBOOST_cell_32040 ( .a(configuration_pci_err_data_507), .b(wbm_dat_o_6_), .o(TIMEBOOST_net_9931) );
na02s01 TIMEBOOST_cell_36311 ( .a(parchk_pci_ad_reg_in_1228), .b(g67051_db), .o(TIMEBOOST_net_10394) );
na02f02 g53397_u0 ( .a(FE_OFN1771_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__Q), .o(n_14245) );
na02f02 g53398_u0 ( .a(FE_OFN1774_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__Q), .o(n_14243) );
na02f02 g53399_u0 ( .a(n_13901), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q), .o(n_14957) );
na02f02 g53400_u0 ( .a(FE_OCP_RBN1984_FE_OFN1591_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__Q), .o(n_14956) );
na02s01 TIMEBOOST_cell_36323 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__Q), .b(g65951_sb), .o(TIMEBOOST_net_10400) );
na02f02 TIMEBOOST_cell_40990 ( .a(TIMEBOOST_net_12733), .b(g57410_sb), .o(n_11332) );
na02f02 TIMEBOOST_cell_41072 ( .a(TIMEBOOST_net_12774), .b(g57082_sb), .o(n_11660) );
na02s02 TIMEBOOST_cell_43638 ( .a(TIMEBOOST_net_14057), .b(FE_OFN2064_n_6391), .o(TIMEBOOST_net_12145) );
na02m02 TIMEBOOST_cell_32420 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_0__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_0__Q), .o(TIMEBOOST_net_10121) );
na02f02 g53407_u0 ( .a(FE_OCP_RBN1962_FE_OFN1591_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q), .o(n_14061) );
na02f02 g53408_u0 ( .a(n_13903), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__14__Q), .o(n_13899) );
na02m02 TIMEBOOST_cell_36363 ( .a(wbu_addr_in_271), .b(g58774_sb), .o(TIMEBOOST_net_10420) );
na02f02 TIMEBOOST_cell_40992 ( .a(TIMEBOOST_net_12734), .b(g57190_sb), .o(n_11562) );
na02f02 TIMEBOOST_cell_41048 ( .a(TIMEBOOST_net_12762), .b(g57399_sb), .o(n_10370) );
na02s01 TIMEBOOST_cell_30871 ( .a(TIMEBOOST_net_9346), .b(g57986_db), .o(n_9811) );
na02m06 TIMEBOOST_cell_36299 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_15__Q), .b(FE_OFN2054_n_8831), .o(TIMEBOOST_net_10388) );
na02m02 TIMEBOOST_cell_32418 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_1__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_1__Q), .o(TIMEBOOST_net_10120) );
na02m02 TIMEBOOST_cell_32464 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__Q), .o(TIMEBOOST_net_10143) );
na02s01 TIMEBOOST_cell_36335 ( .a(parchk_pci_ad_reg_in_1229), .b(g67084_db), .o(TIMEBOOST_net_10406) );
na02f02 TIMEBOOST_cell_40994 ( .a(TIMEBOOST_net_12735), .b(g57212_sb), .o(n_10439) );
na02s02 TIMEBOOST_cell_32039 ( .a(TIMEBOOST_net_9930), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_4912) );
na02m02 TIMEBOOST_cell_41108 ( .a(TIMEBOOST_net_12792), .b(g57127_sb), .o(n_11618) );
na02f02 TIMEBOOST_cell_41074 ( .a(TIMEBOOST_net_12775), .b(g57197_sb), .o(n_11556) );
na02f02 g53424_u0 ( .a(FE_OCP_RBN1962_FE_OFN1591_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__Q), .o(n_14056) );
na02s01 TIMEBOOST_cell_36359 ( .a(pci_target_unit_del_sync_bc_in), .b(g66427_db), .o(TIMEBOOST_net_10418) );
na02m02 TIMEBOOST_cell_32416 ( .a(TIMEBOOST_net_996), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_2__Q), .o(TIMEBOOST_net_10119) );
na02f02 g53427_u0 ( .a(FE_OFN1771_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__Q), .o(n_14055) );
na02f02 g53428_u0 ( .a(FE_OFN1774_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__Q), .o(n_14226) );
na02f02 g53429_u0 ( .a(n_13891), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__Q), .o(n_14961) );
na02f02 g53430_u0 ( .a(FE_OCP_RBN1961_FE_OFN1591_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__Q), .o(n_14960) );
na02m02 TIMEBOOST_cell_32462 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__Q), .o(TIMEBOOST_net_10142) );
na02s01 TIMEBOOST_cell_36337 ( .a(parchk_pci_ad_reg_in_1218), .b(g67053_db), .o(TIMEBOOST_net_10407) );
na02f02 g53433_u0 ( .a(FE_OFN1773_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__Q), .o(n_14225) );
na02f02 g53434_u0 ( .a(FE_OFN1769_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__Q), .o(n_14223) );
na02f02 g53435_u0 ( .a(n_13891), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__Q), .o(n_14963) );
na02f02 TIMEBOOST_cell_43742 ( .a(TIMEBOOST_net_14109), .b(FE_OFN1420_n_8567), .o(TIMEBOOST_net_12700) );
na02f02 TIMEBOOST_cell_40996 ( .a(TIMEBOOST_net_12736), .b(g57508_sb), .o(n_11232) );
na02f02 g53439_u0 ( .a(FE_OFN1774_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__Q), .o(n_14220) );
na02f02 g53440_u0 ( .a(FE_OFN1770_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__Q), .o(n_14049) );
na02s02 TIMEBOOST_cell_43639 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__Q), .b(n_3642), .o(TIMEBOOST_net_14058) );
na02m02 TIMEBOOST_cell_32414 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q), .b(n_1225), .o(TIMEBOOST_net_10118) );
na02m02 TIMEBOOST_cell_32532 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__Q), .o(TIMEBOOST_net_10177) );
na02s01 TIMEBOOST_cell_39572 ( .a(TIMEBOOST_net_12024), .b(g62949_sb), .o(n_5983) );
na02f02 g53447_u0 ( .a(n_13903), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__Q), .o(n_13888) );
na02f02 TIMEBOOST_cell_43828 ( .a(TIMEBOOST_net_14152), .b(FE_OFN1380_n_8567), .o(TIMEBOOST_net_12933) );
na02s01 TIMEBOOST_cell_36349 ( .a(pciu_pciif_idsel_reg_in), .b(g67052_db), .o(TIMEBOOST_net_10413) );
na02f02 TIMEBOOST_cell_40998 ( .a(TIMEBOOST_net_12737), .b(g57598_sb), .o(n_10285) );
na02f02 g53451_u0 ( .a(FE_OFN1770_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__Q), .o(n_14212) );
na02f02 g53452_u0 ( .a(FE_OFN1774_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__Q), .o(n_14211) );
na02s02 TIMEBOOST_cell_36343 ( .a(n_2427), .b(n_2237), .o(TIMEBOOST_net_10410) );
na02s02 TIMEBOOST_cell_37996 ( .a(TIMEBOOST_net_11236), .b(n_3814), .o(n_4957) );
na02f02 TIMEBOOST_cell_41118 ( .a(TIMEBOOST_net_12797), .b(g57173_sb), .o(n_11583) );
na02s01 TIMEBOOST_cell_36313 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__Q), .b(g65870_sb), .o(TIMEBOOST_net_10395) );
na02f02 g53457_u0 ( .a(FE_OFN1775_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__Q), .o(n_16613) );
na02f02 g53458_u0 ( .a(FE_OFN1769_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__Q), .o(n_16612) );
na02f02 g53459_u0 ( .a(FE_OFN1774_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__Q), .o(n_14207) );
na02m02 TIMEBOOST_cell_32412 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_2__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_2__Q), .o(TIMEBOOST_net_10117) );
na02m02 TIMEBOOST_cell_32492 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__Q), .o(TIMEBOOST_net_10157) );
na02m02 TIMEBOOST_cell_43743 ( .a(n_9021), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__Q), .o(TIMEBOOST_net_14110) );
na02f02 g53463_u0 ( .a(FE_OFN1774_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__Q), .o(n_14205) );
na02f02 g53464_u0 ( .a(FE_OFN1770_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__Q), .o(n_14203) );
na02s01 TIMEBOOST_cell_36355 ( .a(pci_target_unit_del_sync_addr_in_228), .b(g66412_db), .o(TIMEBOOST_net_10416) );
na02s01 TIMEBOOST_cell_44797 ( .a(g58094_sb), .b(g58094_db), .o(TIMEBOOST_net_14637) );
na02f02 g53467_u0 ( .a(FE_OFN1775_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__28__Q), .o(n_14202) );
na02f02 g53468_u0 ( .a(FE_OFN1769_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__28__Q), .o(n_14201) );
na02m02 TIMEBOOST_cell_32476 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__Q), .o(TIMEBOOST_net_10149) );
na02f02 TIMEBOOST_cell_43744 ( .a(TIMEBOOST_net_14110), .b(FE_OFN1396_n_8567), .o(TIMEBOOST_net_12949) );
na02f02 TIMEBOOST_cell_41094 ( .a(TIMEBOOST_net_12785), .b(g57130_sb), .o(n_10839) );
na03m02 TIMEBOOST_cell_34887 ( .a(TIMEBOOST_net_9993), .b(n_2987), .c(g59382_sb), .o(n_3483) );
na02s02 TIMEBOOST_cell_43666 ( .a(TIMEBOOST_net_14071), .b(FE_OFN1311_n_6624), .o(TIMEBOOST_net_12231) );
na02f02 TIMEBOOST_cell_41000 ( .a(TIMEBOOST_net_12738), .b(g57205_sb), .o(n_10440) );
na02s01 TIMEBOOST_cell_42697 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__Q), .b(FE_OFN652_n_4508), .o(TIMEBOOST_net_13587) );
na02m02 TIMEBOOST_cell_32410 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q), .b(n_971), .o(TIMEBOOST_net_10116) );
na02f02 TIMEBOOST_cell_41002 ( .a(TIMEBOOST_net_12739), .b(g57308_sb), .o(n_11442) );
na02s01 TIMEBOOST_cell_43274 ( .a(TIMEBOOST_net_13875), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_12545) );
na02f02 TIMEBOOST_cell_41076 ( .a(TIMEBOOST_net_12776), .b(g57248_sb), .o(n_11509) );
na02f02 g53480_u0 ( .a(FE_OFN1596_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__Q), .o(n_14035) );
na02f02 g53481_u0 ( .a(FE_OFN1773_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__Q), .o(n_14197) );
na02f02 g53483_u0 ( .a(FE_OFN1775_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__Q), .o(n_14195) );
na02f02 g53484_u0 ( .a(FE_OFN1768_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__Q), .o(n_14194) );
na02s01 TIMEBOOST_cell_36315 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__Q), .b(g65861_sb), .o(TIMEBOOST_net_10396) );
na03f02 TIMEBOOST_cell_31970 ( .a(TIMEBOOST_net_607), .b(g62033_sb), .c(n_2744), .o(TIMEBOOST_net_9896) );
na02f02 g53487_u0 ( .a(n_13903), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q), .o(n_13878) );
na02f02 g53488_u0 ( .a(FE_OFN1596_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__Q), .o(n_14033) );
na02s02 TIMEBOOST_cell_43275 ( .a(n_4245), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__Q), .o(TIMEBOOST_net_13876) );
na02m02 TIMEBOOST_cell_32408 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q), .b(n_829), .o(TIMEBOOST_net_10115) );
na02f02 TIMEBOOST_cell_32551 ( .a(n_12313), .b(TIMEBOOST_net_10186), .o(TIMEBOOST_net_6558) );
na02s01 TIMEBOOST_cell_39574 ( .a(TIMEBOOST_net_12025), .b(g62598_sb), .o(n_6355) );
na02s01 TIMEBOOST_cell_42715 ( .a(g65009_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__Q), .o(TIMEBOOST_net_13596) );
na02f02 TIMEBOOST_cell_41004 ( .a(TIMEBOOST_net_12740), .b(g57578_sb), .o(n_10292) );
na02s01 TIMEBOOST_cell_30813 ( .a(TIMEBOOST_net_9317), .b(TIMEBOOST_net_154), .o(n_8818) );
na02m02 TIMEBOOST_cell_32406 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q), .o(TIMEBOOST_net_10114) );
na02f02 TIMEBOOST_cell_41006 ( .a(TIMEBOOST_net_12741), .b(g57590_sb), .o(n_10289) );
na02s01 TIMEBOOST_cell_30815 ( .a(TIMEBOOST_net_9318), .b(g64810_db), .o(n_3748) );
na02s01 TIMEBOOST_cell_30817 ( .a(TIMEBOOST_net_9319), .b(g64813_db), .o(n_3745) );
na02m02 TIMEBOOST_cell_32404 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q), .b(n_13608), .o(TIMEBOOST_net_10113) );
na02f02 g53501_u0 ( .a(FE_OFN1596_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__Q), .o(n_14029) );
na02f02 g53502_u0 ( .a(n_13903), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__Q), .o(n_13875) );
na02m02 TIMEBOOST_cell_32460 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__22__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q), .o(TIMEBOOST_net_10141) );
na02f02 g53504_u0 ( .a(FE_OFN1593_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__Q), .o(n_14027) );
na02f02 g53505_u0 ( .a(FE_OFN1775_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__Q), .o(n_14186) );
na02f02 g53506_u0 ( .a(FE_OFN1768_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__Q), .o(n_14185) );
na02s01 TIMEBOOST_cell_30819 ( .a(TIMEBOOST_net_9320), .b(g58028_sb), .o(TIMEBOOST_net_1518) );
na02f02 TIMEBOOST_cell_41008 ( .a(TIMEBOOST_net_12742), .b(g57506_sb), .o(n_10815) );
na02m02 TIMEBOOST_cell_32402 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q), .o(TIMEBOOST_net_10112) );
na02s02 TIMEBOOST_cell_45260 ( .a(TIMEBOOST_net_14868), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_13237) );
na02f02 TIMEBOOST_cell_43812 ( .a(TIMEBOOST_net_14144), .b(FE_OFN1382_n_8567), .o(TIMEBOOST_net_12928) );
na02f02 TIMEBOOST_cell_41010 ( .a(TIMEBOOST_net_12743), .b(g57514_sb), .o(n_11228) );
na02f02 g53513_u0 ( .a(n_13901), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__Q), .o(n_13871) );
na02f02 g53514_u0 ( .a(FE_OFN1593_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__Q), .o(n_14025) );
na02f02 g53515_u0 ( .a(FE_OFN1768_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__Q), .o(n_14178) );
na02f02 g53516_u0 ( .a(FE_OFN1775_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__Q), .o(n_14177) );
na02f02 TIMEBOOST_cell_41078 ( .a(TIMEBOOST_net_12777), .b(g57348_sb), .o(n_11402) );
na02f02 g53518_u0 ( .a(FE_OFN1593_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__Q), .o(n_14024) );
na02m02 TIMEBOOST_cell_32458 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q), .o(TIMEBOOST_net_10140) );
no02f08 TIMEBOOST_cell_36317 ( .a(FE_RN_103_0), .b(FE_RN_102_0), .o(TIMEBOOST_net_10397) );
na02m02 TIMEBOOST_cell_43745 ( .a(n_9486), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__Q), .o(TIMEBOOST_net_14111) );
na02m02 TIMEBOOST_cell_32400 ( .a(FE_OCP_RBN2265_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_0__Q), .o(TIMEBOOST_net_10111) );
na02f02 g53523_u0 ( .a(FE_OFN1770_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__Q), .o(n_14174) );
na02f02 TIMEBOOST_cell_41012 ( .a(TIMEBOOST_net_12744), .b(g57335_sb), .o(n_10394) );
na02f02 g53525_u0 ( .a(n_13891), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__Q), .o(n_13868) );
na02f02 g53526_u0 ( .a(FE_OCP_RBN1961_FE_OFN1591_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__Q), .o(n_14022) );
na02f02 TIMEBOOST_cell_32457 ( .a(TIMEBOOST_net_10139), .b(FE_OFN1770_n_14054), .o(TIMEBOOST_net_6253) );
na02f02 TIMEBOOST_cell_43829 ( .a(n_9023), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__Q), .o(TIMEBOOST_net_14153) );
na02f02 g53529_u0 ( .a(FE_OFN1773_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__Q), .o(n_14172) );
na02f02 g53530_u0 ( .a(FE_OFN1769_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__Q), .o(n_14020) );
na02f02 g53531_u0 ( .a(FE_OFN1774_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__Q), .o(n_14171) );
na02f02 g53532_u0 ( .a(FE_OFN1768_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__Q), .o(n_14170) );
na02m02 g53533_u0 ( .a(FE_OFN1593_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__Q), .o(n_14019) );
na02m02 TIMEBOOST_cell_32456 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__Q), .o(TIMEBOOST_net_10139) );
na02f02 g53535_u0 ( .a(n_13903), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__Q), .o(n_13865) );
na02f02 g53536_u0 ( .a(FE_OCP_RBN1961_FE_OFN1591_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__Q), .o(n_14018) );
na02s01 TIMEBOOST_cell_37977 ( .a(g63039_sb), .b(g63039_db), .o(TIMEBOOST_net_11227) );
na02s02 TIMEBOOST_cell_38597 ( .a(TIMEBOOST_net_9938), .b(FE_OFN1181_n_3476), .o(TIMEBOOST_net_11537) );
na02f02 TIMEBOOST_cell_41080 ( .a(TIMEBOOST_net_12778), .b(g57391_sb), .o(n_11352) );
na02f02 TIMEBOOST_cell_43830 ( .a(TIMEBOOST_net_14153), .b(FE_OFN1400_n_8567), .o(TIMEBOOST_net_12963) );
na02f02 g53541_u0 ( .a(FE_OFN1769_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__Q), .o(n_14167) );
na02f02 g53542_u0 ( .a(FE_OFN1775_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__Q), .o(n_14166) );
na02f02 g53543_u0 ( .a(n_13903), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__Q), .o(n_13863) );
na02f02 g53544_u0 ( .a(FE_OCP_RBN1961_FE_OFN1591_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__Q), .o(n_14016) );
na02f02 TIMEBOOST_cell_43746 ( .a(TIMEBOOST_net_14111), .b(FE_OFN1396_n_8567), .o(TIMEBOOST_net_12929) );
na02m02 TIMEBOOST_cell_32398 ( .a(n_13608), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_1__Q), .o(TIMEBOOST_net_10110) );
na02f02 g53547_u0 ( .a(n_13790), .b(n_168), .o(n_14305) );
na02m02 TIMEBOOST_cell_32454 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__14__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__14__Q), .o(TIMEBOOST_net_10138) );
na02s01 TIMEBOOST_cell_42607 ( .a(FE_OFN245_n_9114), .b(g58095_sb), .o(TIMEBOOST_net_13542) );
na02s02 TIMEBOOST_cell_44901 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__Q), .b(n_4520), .o(TIMEBOOST_net_14689) );
na02f02 g53552_u0 ( .a(FE_OFN1588_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__Q), .o(n_14013) );
na02f02 TIMEBOOST_cell_41256 ( .a(TIMEBOOST_net_12866), .b(g57170_sb), .o(n_10453) );
na02s01 TIMEBOOST_cell_30829 ( .a(TIMEBOOST_net_9325), .b(g66397_sb), .o(n_2546) );
na02s02 TIMEBOOST_cell_39576 ( .a(TIMEBOOST_net_12026), .b(g62903_sb), .o(n_6071) );
na02f04 g53556_u0 ( .a(FE_OCP_RBN1997_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__Q), .o(n_14011) );
na02f02 g53557_u0 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__Q), .o(n_13862) );
na02s01 TIMEBOOST_cell_30831 ( .a(TIMEBOOST_net_9326), .b(g66397_sb), .o(n_2540) );
na02f04 TIMEBOOST_cell_39519 ( .a(TIMEBOOST_net_9850), .b(FE_OCPN1911_FE_OFN1152_n_13249), .o(TIMEBOOST_net_11998) );
na02s02 TIMEBOOST_cell_43276 ( .a(TIMEBOOST_net_13876), .b(FE_OFN1225_n_6391), .o(TIMEBOOST_net_12522) );
na02s01 TIMEBOOST_cell_39518 ( .a(TIMEBOOST_net_11997), .b(g58452_db), .o(n_9405) );
na02f02 g53562_u0 ( .a(FE_OCP_RBN1995_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__12__Q), .o(n_14007) );
na02f02 g53563_u0 ( .a(FE_OFN1588_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__12__Q), .o(n_14005) );
no02f04 TIMEBOOST_cell_30835 ( .a(TIMEBOOST_net_9328), .b(FE_RN_505_0), .o(n_2253) );
na02s02 TIMEBOOST_cell_44902 ( .a(TIMEBOOST_net_14689), .b(FE_OFN712_n_8140), .o(TIMEBOOST_net_11086) );
na02f02 g53566_u0 ( .a(FE_OFN1588_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q), .o(n_14004) );
na02f02 g53567_u0 ( .a(n_13993), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q), .o(n_14002) );
na02s01 TIMEBOOST_cell_15832 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_92), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3173) );
na02s02 TIMEBOOST_cell_39578 ( .a(TIMEBOOST_net_12027), .b(g62359_sb), .o(n_6880) );
na02s01 TIMEBOOST_cell_15842 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_75), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3178) );
na02s01 TIMEBOOST_cell_44903 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__Q), .b(n_2162), .o(TIMEBOOST_net_14690) );
na02f02 g53572_u0 ( .a(n_13987), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__15__Q), .o(n_14000) );
na02f02 g53573_u0 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__15__Q), .o(n_13999) );
na02s01 TIMEBOOST_cell_39580 ( .a(TIMEBOOST_net_12028), .b(g62458_sb), .o(n_6680) );
na02s01 TIMEBOOST_cell_15830 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_90), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3172) );
na02s01 TIMEBOOST_cell_44904 ( .a(TIMEBOOST_net_14690), .b(FE_OFN699_n_7845), .o(TIMEBOOST_net_11096) );
na02f02 g53578_u0 ( .a(n_13993), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q), .o(n_13994) );
na02f02 g53579_u0 ( .a(FE_OFN1588_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__16__Q), .o(n_13992) );
na02s01 TIMEBOOST_cell_36339 ( .a(parchk_pci_ad_reg_in_1227), .b(g67088_db), .o(TIMEBOOST_net_10408) );
na02s01 TIMEBOOST_cell_39315 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__Q), .b(g65845_sb), .o(TIMEBOOST_net_11896) );
na02f04 g53582_u0 ( .a(FE_OCP_RBN1997_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__Q), .o(n_13991) );
na02f02 g53583_u0 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__Q), .o(n_13990) );
na02f02 TIMEBOOST_cell_41014 ( .a(TIMEBOOST_net_12745), .b(g57231_sb), .o(n_10433) );
na03s02 TIMEBOOST_cell_36291 ( .a(n_1073), .b(n_1159), .c(n_1164), .o(TIMEBOOST_net_10384) );
na02s01 TIMEBOOST_cell_38124 ( .a(TIMEBOOST_net_11300), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_4603) );
na02s01 TIMEBOOST_cell_36341 ( .a(parchk_pci_ad_reg_in_1214), .b(g67091_db), .o(TIMEBOOST_net_10409) );
na02f02 g53588_u0 ( .a(n_13987), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__Q), .o(n_13982) );
na02s02 TIMEBOOST_cell_30875 ( .a(TIMEBOOST_net_9348), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_3736) );
na02f04 g53590_u0 ( .a(FE_OFN1606_n_13997), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__Q), .o(n_14144) );
na02f02 g53591_u0 ( .a(FE_OFN1600_n_13995), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__Q), .o(n_14142) );
na02f02 g53592_u0 ( .a(FE_OCP_RBN1998_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__1__Q), .o(n_13980) );
na02f02 g53593_u0 ( .a(FE_OFN1587_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q), .o(n_13859) );
na02s01 TIMEBOOST_cell_36361 ( .a(pci_target_unit_del_sync_bc_in_202), .b(g66411_db), .o(TIMEBOOST_net_10419) );
na02s02 TIMEBOOST_cell_39582 ( .a(TIMEBOOST_net_12029), .b(g62946_sb), .o(n_5989) );
na02f02 g53596_u0 ( .a(FE_OFN1606_n_13997), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__Q), .o(n_14140) );
in01s01 TIMEBOOST_cell_45949 ( .a(wbm_dat_i_3_), .o(TIMEBOOST_net_15256) );
na02s01 TIMEBOOST_cell_42628 ( .a(TIMEBOOST_net_13552), .b(g58176_db), .o(n_9613) );
na02s01 TIMEBOOST_cell_37983 ( .a(TIMEBOOST_net_442), .b(g62835_sb), .o(TIMEBOOST_net_11230) );
na02s01 TIMEBOOST_cell_36387 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(g65700_sb), .o(TIMEBOOST_net_10432) );
na02s01 TIMEBOOST_cell_39584 ( .a(TIMEBOOST_net_12030), .b(g62613_sb), .o(n_6331) );
na02s02 TIMEBOOST_cell_41792 ( .a(TIMEBOOST_net_13134), .b(g64213_db), .o(n_3956) );
in01s01 TIMEBOOST_cell_45950 ( .a(TIMEBOOST_net_15256), .o(TIMEBOOST_net_15257) );
na02s01 TIMEBOOST_cell_15863 ( .a(TIMEBOOST_net_3188), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_397), .o(TIMEBOOST_net_58) );
na02s01 TIMEBOOST_cell_39586 ( .a(TIMEBOOST_net_12031), .b(g62424_sb), .o(n_7387) );
na02f02 g53606_u0 ( .a(FE_OFN1588_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__Q), .o(n_13974) );
na02f02 g53607_u0 ( .a(n_13993), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__Q), .o(n_13973) );
na02s01 TIMEBOOST_cell_43277 ( .a(TIMEBOOST_net_4770), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_13877) );
na02f04 g53610_u0 ( .a(FE_OCP_RBN1997_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__Q), .o(n_13972) );
na02f02 g53611_u0 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__Q), .o(n_13857) );
na02m02 TIMEBOOST_cell_32396 ( .a(FE_OCP_RBN2265_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q), .o(TIMEBOOST_net_10109) );
na02s01 TIMEBOOST_cell_36275 ( .a(TIMEBOOST_net_9282), .b(n_574), .o(TIMEBOOST_net_10376) );
na03f02 TIMEBOOST_cell_36199 ( .a(n_12357), .b(TIMEBOOST_net_10296), .c(n_11831), .o(n_12616) );
na02s01 TIMEBOOST_cell_44905 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__Q), .b(n_2164), .o(TIMEBOOST_net_14691) );
na02f01 g53616_u0 ( .a(n_13997), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__Q), .o(n_14128) );
na02m02 TIMEBOOST_cell_43831 ( .a(n_9717), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__Q), .o(TIMEBOOST_net_14154) );
na03f08 TIMEBOOST_cell_36279 ( .a(n_1698), .b(n_1061), .c(n_2648), .o(TIMEBOOST_net_10378) );
na02s02 TIMEBOOST_cell_39588 ( .a(TIMEBOOST_net_12032), .b(g62592_sb), .o(n_6369) );
na02s01 TIMEBOOST_cell_30849 ( .a(TIMEBOOST_net_9335), .b(g65021_db), .o(n_3632) );
na03f10 TIMEBOOST_cell_36283 ( .a(n_1698), .b(n_2648), .c(n_8511), .o(TIMEBOOST_net_10380) );
na02f02 g53623_u0 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__Q), .o(n_13856) );
na02s01 TIMEBOOST_cell_44906 ( .a(TIMEBOOST_net_14691), .b(FE_OFN702_n_7845), .o(TIMEBOOST_net_11057) );
na02s02 TIMEBOOST_cell_41793 ( .a(pci_target_unit_fifos_pciw_addr_data_in_136), .b(g64195_sb), .o(TIMEBOOST_net_13135) );
na02s01 TIMEBOOST_cell_30851 ( .a(TIMEBOOST_net_9336), .b(g65024_db), .o(n_3630) );
na02s02 TIMEBOOST_cell_38618 ( .a(TIMEBOOST_net_11547), .b(g62621_sb), .o(n_6315) );
na02s02 TIMEBOOST_cell_39590 ( .a(TIMEBOOST_net_12033), .b(g62430_sb), .o(n_6738) );
na02m02 TIMEBOOST_cell_42526 ( .a(FE_OFN1438_n_9372), .b(TIMEBOOST_net_13501), .o(TIMEBOOST_net_12336) );
na02s02 TIMEBOOST_cell_41794 ( .a(TIMEBOOST_net_13135), .b(g64195_db), .o(n_3974) );
na02m02 TIMEBOOST_cell_32302 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_2_), .o(TIMEBOOST_net_10062) );
na02s01 TIMEBOOST_cell_15869 ( .a(TIMEBOOST_net_3191), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_404), .o(TIMEBOOST_net_66) );
na02m02 TIMEBOOST_cell_44643 ( .a(n_9077), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__Q), .o(TIMEBOOST_net_14560) );
na02s02 TIMEBOOST_cell_39592 ( .a(TIMEBOOST_net_12034), .b(g62377_sb), .o(n_6849) );
na02f02 g53635_u0 ( .a(FE_OCP_RBN1997_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__Q), .o(n_13960) );
na02s01 TIMEBOOST_cell_15865 ( .a(TIMEBOOST_net_3189), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_399), .o(TIMEBOOST_net_60) );
na02s08 TIMEBOOST_cell_36243 ( .a(n_104), .b(n_247), .o(TIMEBOOST_net_10360) );
na02m02 TIMEBOOST_cell_32300 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_3_), .o(TIMEBOOST_net_10061) );
na02f02 g53639_u0 ( .a(FE_OCP_RBN1996_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__Q), .o(n_13958) );
na02f40 TIMEBOOST_cell_36245 ( .a(wishbone_slave_unit_pci_initiator_sm_cur_state_3_), .b(wishbone_slave_unit_pci_initiator_sm_cur_state_2_), .o(TIMEBOOST_net_10361) );
na02s01 TIMEBOOST_cell_15827 ( .a(TIMEBOOST_net_3170), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_398), .o(TIMEBOOST_net_59) );
na02f02 g53643_u0 ( .a(FE_OFN1587_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__Q), .o(n_13854) );
na02s01 TIMEBOOST_cell_42682 ( .a(TIMEBOOST_net_13579), .b(g64770_db), .o(n_3778) );
na02s02 TIMEBOOST_cell_39594 ( .a(TIMEBOOST_net_12035), .b(g62527_sb), .o(n_6521) );
na02s02 TIMEBOOST_cell_44887 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__Q), .b(FE_OFN644_n_4677), .o(TIMEBOOST_net_14682) );
na02m02 TIMEBOOST_cell_32298 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .o(TIMEBOOST_net_10060) );
na02f01 g53648_u0 ( .a(n_13997), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__Q), .o(n_14111) );
na02s02 TIMEBOOST_cell_45203 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__Q), .b(n_4445), .o(TIMEBOOST_net_14840) );
na02s02 TIMEBOOST_cell_39596 ( .a(TIMEBOOST_net_12036), .b(g62604_sb), .o(n_6344) );
na02m02 TIMEBOOST_cell_44631 ( .a(n_9017), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__Q), .o(TIMEBOOST_net_14554) );
na02m02 TIMEBOOST_cell_32296 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_0_), .o(TIMEBOOST_net_10059) );
na02f02 g53654_u0 ( .a(FE_OFN1586_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__Q), .o(n_13954) );
na02f02 g53655_u0 ( .a(FE_OCP_RBN1999_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__Q), .o(n_13953) );
na02m02 TIMEBOOST_cell_21968 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__Q), .o(TIMEBOOST_net_6241) );
na03f08 TIMEBOOST_cell_36247 ( .a(n_16284), .b(n_16285), .c(conf_w_addr_in_938), .o(TIMEBOOST_net_10362) );
na02s02 TIMEBOOST_cell_39598 ( .a(TIMEBOOST_net_12037), .b(g62542_sb), .o(n_6483) );
na02s01 TIMEBOOST_cell_36249 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_96), .b(wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_10363) );
na02s01 TIMEBOOST_cell_44888 ( .a(TIMEBOOST_net_14682), .b(g65423_sb), .o(TIMEBOOST_net_12415) );
na02f01 g53661_u0 ( .a(n_13997), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__Q), .o(n_13949) );
na02m02 TIMEBOOST_cell_32294 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_), .b(n_1465), .o(TIMEBOOST_net_10058) );
na02s02 TIMEBOOST_cell_43505 ( .a(n_4426), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__Q), .o(TIMEBOOST_net_13991) );
na02s01 TIMEBOOST_cell_39532 ( .a(TIMEBOOST_net_12004), .b(g61708_sb), .o(n_8411) );
na02s01 TIMEBOOST_cell_36253 ( .a(n_9), .b(n_692), .o(TIMEBOOST_net_10365) );
na02f08 TIMEBOOST_cell_36267 ( .a(n_696), .b(n_15331), .o(TIMEBOOST_net_10372) );
na02f02 g53668_u0 ( .a(n_13993), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__Q), .o(n_13943) );
na02f02 g53669_u0 ( .a(FE_OFN1586_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__Q), .o(n_13942) );
na03s02 TIMEBOOST_cell_33992 ( .a(TIMEBOOST_net_4083), .b(g65361_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__Q), .o(TIMEBOOST_net_4795) );
na02s01 TIMEBOOST_cell_36273 ( .a(TIMEBOOST_net_9283), .b(n_574), .o(TIMEBOOST_net_10375) );
na02s02 TIMEBOOST_cell_39600 ( .a(TIMEBOOST_net_12038), .b(g62463_sb), .o(n_6670) );
na02s02 TIMEBOOST_cell_43667 ( .a(n_3669), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__1__Q), .o(TIMEBOOST_net_14072) );
na02f02 g53674_u0 ( .a(FE_OFN1605_n_13997), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__Q), .o(n_13938) );
na02f02 g53675_u0 ( .a(FE_OFN1601_n_13995), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__Q), .o(n_13937) );
no02f08 TIMEBOOST_cell_36257 ( .a(n_16003), .b(n_15924), .o(TIMEBOOST_net_10367) );
na02f02 g53678_u0 ( .a(n_13993), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__Q), .o(n_13936) );
na02f02 TIMEBOOST_cell_36271 ( .a(n_1998), .b(n_2390), .o(TIMEBOOST_net_10374) );
na02f02 TIMEBOOST_cell_41082 ( .a(TIMEBOOST_net_12779), .b(g57129_sb), .o(n_10841) );
na03s02 TIMEBOOST_cell_5531 ( .a(n_4452), .b(g65063_sb), .c(g65063_db), .o(n_4316) );
na02s02 TIMEBOOST_cell_43166 ( .a(TIMEBOOST_net_13821), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_12134) );
na02m02 TIMEBOOST_cell_32290 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_), .b(n_1287), .o(TIMEBOOST_net_10056) );
na02s01 TIMEBOOST_cell_40861 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__Q), .b(n_13541), .o(TIMEBOOST_net_12669) );
na02s01 TIMEBOOST_cell_36251 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_70), .b(wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_10364) );
na02f02 g53687_u0 ( .a(FE_OFN1602_n_13995), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__Q), .o(n_14099) );
na02f02 g53688_u0 ( .a(FE_OCP_RBN1997_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__Q), .o(n_13930) );
na02f02 g53689_u0 ( .a(FE_OFN1587_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__Q), .o(n_13849) );
na02f02 TIMEBOOST_cell_42954 ( .a(TIMEBOOST_net_13715), .b(g54238_sb), .o(n_13436) );
na02f02 TIMEBOOST_cell_32289 ( .a(TIMEBOOST_net_10055), .b(FE_OFN1373_n_8567), .o(TIMEBOOST_net_6058) );
na02s01 TIMEBOOST_cell_42658 ( .a(TIMEBOOST_net_13567), .b(g64328_sb), .o(n_3848) );
na03s02 TIMEBOOST_cell_37935 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__Q), .b(FE_OFN1666_n_9477), .c(FE_OFN270_n_9836), .o(TIMEBOOST_net_11206) );
na02s01 TIMEBOOST_cell_36325 ( .a(parchk_pci_ad_reg_in_1230), .b(g67093_db), .o(TIMEBOOST_net_10401) );
na02s02 TIMEBOOST_cell_39602 ( .a(TIMEBOOST_net_12039), .b(g62390_sb), .o(n_6819) );
na02s02 TIMEBOOST_cell_40860 ( .a(TIMEBOOST_net_12668), .b(FE_OFN1331_n_13547), .o(TIMEBOOST_net_11623) );
na02m02 TIMEBOOST_cell_36261 ( .a(g58789_sb), .b(n_8831), .o(TIMEBOOST_net_10369) );
na02m02 g53698_u0 ( .a(FE_OCPN2218_n_13997), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__Q), .o(n_13926) );
na02f02 TIMEBOOST_cell_37141 ( .a(n_14433), .b(n_14515), .o(TIMEBOOST_net_10809) );
na02f02 g53701_u0 ( .a(FE_OFN1586_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__Q), .o(n_13847) );
na02m02 TIMEBOOST_cell_21974 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__Q), .o(TIMEBOOST_net_6244) );
na02f04 g53706_u0 ( .a(FE_OCP_RBN1997_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__Q), .o(n_13923) );
na02f02 g53707_u0 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__Q), .o(n_13846) );
no02f04 g53708_u0 ( .a(n_13710), .b(n_2629), .o(n_13749) );
no02f01 g53709_u0 ( .a(n_16456), .b(n_13921), .o(g53709_p) );
in01f02 g53709_u1 ( .a(g53709_p), .o(n_13922) );
ao12f02 g53710_u0 ( .a(n_13721), .b(n_13450), .c(n_1789), .o(n_13725) );
ao12f02 g53711_u0 ( .a(n_13721), .b(n_13448), .c(n_1785), .o(n_13722) );
ao12f02 g53712_u0 ( .a(n_13721), .b(n_13444), .c(n_1788), .o(n_13720) );
na03s02 TIMEBOOST_cell_45791 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__6__Q), .b(g64262_da), .c(g64262_db), .o(TIMEBOOST_net_15134) );
ao12f01 g53714_u0 ( .a(n_15347), .b(n_4795), .c(n_13813), .o(n_13844) );
na02f02 g53715_u0 ( .a(n_13681), .b(n_2630), .o(n_13748) );
ao22f02 g53716_u0 ( .a(n_1645), .b(n_7567), .c(n_1523), .d(n_15371), .o(n_7568) );
na02s02 TIMEBOOST_cell_43567 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__Q), .b(n_3625), .o(TIMEBOOST_net_14022) );
in01s02 g53718_u0 ( .a(n_13821), .o(n_13843) );
na02s02 TIMEBOOST_cell_45792 ( .a(TIMEBOOST_net_15134), .b(FE_OFN1094_g64577_p), .o(TIMEBOOST_net_6226) );
ao22f01 g53720_u0 ( .a(n_2629), .b(n_13817), .c(n_13679), .d(n_13820), .o(n_13819) );
in01f02 g53721_u0 ( .a(n_13842), .o(n_13920) );
ao22f02 g53722_u0 ( .a(n_13625), .b(n_13820), .c(n_12167), .d(n_13817), .o(n_13842) );
in01f02 g53723_u0 ( .a(n_13715), .o(n_13716) );
no02f02 g53726_u0 ( .a(n_7093), .b(n_13335), .o(g53726_p) );
ao12f02 g53726_u1 ( .a(g53726_p), .b(n_13335), .c(n_7093), .o(n_13715) );
ao22f01 g53727_u0 ( .a(n_7531), .b(n_13679), .c(n_2764), .d(FE_OCPN1836_n_16798), .o(n_13919) );
no02f02 g53729_u0 ( .a(n_13679), .b(n_2629), .o(g53729_p) );
in01f02 g53729_u1 ( .a(g53729_p), .o(n_13681) );
na02m02 TIMEBOOST_cell_44125 ( .a(n_9018), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__Q), .o(TIMEBOOST_net_14301) );
no02f02 g53731_u0 ( .a(n_13355), .b(n_13784), .o(n_13592) );
no02f02 g53732_u0 ( .a(n_13353), .b(n_13784), .o(n_13591) );
no02f02 g53734_u0 ( .a(n_13350), .b(n_13784), .o(n_13587) );
no02f02 g53735_u0 ( .a(n_13349), .b(n_13784), .o(n_13585) );
na02s02 TIMEBOOST_cell_39604 ( .a(TIMEBOOST_net_12040), .b(g62642_sb), .o(n_6264) );
no02f02 g53738_u0 ( .a(n_13416), .b(FE_OFN1709_n_4868), .o(n_13680) );
no02f02 g53739_u0 ( .a(n_13342), .b(FE_OFN1709_n_4868), .o(n_13582) );
ao12f02 g53740_u0 ( .a(FE_OFN969_n_13784), .b(n_13292), .c(n_7551), .o(n_13581) );
ao12f02 g53741_u0 ( .a(FE_OFN969_n_13784), .b(n_13291), .c(n_7550), .o(n_13579) );
ao12f02 g53742_u0 ( .a(FE_OFN969_n_13784), .b(n_13290), .c(n_7548), .o(n_13578) );
ao12f02 g53744_u0 ( .a(FE_OFN969_n_13784), .b(n_13287), .c(n_7547), .o(n_13576) );
no02f02 g53745_u0 ( .a(n_13339), .b(FE_OFN1946_n_13784), .o(n_13575) );
no02f02 g53746_u0 ( .a(n_13338), .b(FE_OFN1946_n_13784), .o(n_13574) );
no02f02 g53747_u0 ( .a(n_13337), .b(n_13784), .o(n_13573) );
na03s02 TIMEBOOST_cell_5454 ( .a(n_4476), .b(g64789_sb), .c(g64789_db), .o(n_4477) );
in01f01 g53750_u0 ( .a(n_13710), .o(n_13711) );
na02f04 g53751_u0 ( .a(n_15611), .b(n_13679), .o(n_13710) );
na02f01 g53752_u0 ( .a(n_13814), .b(n_13813), .o(g53752_p) );
in01f02 g53752_u1 ( .a(g53752_p), .o(n_13921) );
na02f02 TIMEBOOST_cell_44562 ( .a(TIMEBOOST_net_14519), .b(FE_OFN2182_n_8567), .o(TIMEBOOST_net_13015) );
no02f02 g53754_u0 ( .a(n_13346), .b(n_13784), .o(n_13569) );
na02f02 TIMEBOOST_cell_22519 ( .a(TIMEBOOST_net_6516), .b(FE_OFN1584_n_12306), .o(n_16596) );
na02s01 TIMEBOOST_cell_42991 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__Q), .b(n_3880), .o(TIMEBOOST_net_13734) );
na02s02 TIMEBOOST_cell_39606 ( .a(TIMEBOOST_net_12041), .b(g62689_sb), .o(n_7366) );
na02m02 TIMEBOOST_cell_44321 ( .a(n_9449), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__Q), .o(TIMEBOOST_net_14399) );
no02f02 g53759_u0 ( .a(n_13417), .b(n_13784), .o(n_13678) );
ao12f02 g53760_u0 ( .a(n_13784), .b(n_13295), .c(n_7307), .o(n_13564) );
na02m02 TIMEBOOST_cell_44237 ( .a(n_9816), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__Q), .o(TIMEBOOST_net_14357) );
in01f06 g53762_u0 ( .a(n_13743), .o(n_13903) );
in01f04 g53764_u0 ( .a(n_13743), .o(n_13891) );
in01f02 g53765_u0 ( .a(n_13743), .o(n_13873) );
in01f02 g53769_u0 ( .a(n_13807), .o(n_13987) );
in01f04 g53772_u0 ( .a(n_13807), .o(n_13971) );
in01f02 g53773_u0 ( .a(n_13807), .o(n_13993) );
na02s01 TIMEBOOST_cell_16630 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__Q), .b(g65330_sb), .o(TIMEBOOST_net_3572) );
in01f02 g53787_u0 ( .a(n_13674), .o(n_13741) );
na02f02 g53812_u0 ( .a(n_13467), .b(n_1794), .o(n_13673) );
na02s02 TIMEBOOST_cell_39480 ( .a(TIMEBOOST_net_11978), .b(FE_OFN1174_n_5592), .o(n_5574) );
na02f02 g53814_u0 ( .a(n_13464), .b(n_1786), .o(n_13671) );
na02f02 g53815_u0 ( .a(n_13463), .b(FE_OFN2057_n_2117), .o(n_13670) );
ao12f02 g53817_u0 ( .a(n_3333), .b(n_13273), .c(n_13447), .o(n_13563) );
na02f02 g53818_u0 ( .a(n_13461), .b(FE_OFN2247_n_2113), .o(n_13668) );
na02f02 g53819_u0 ( .a(n_13362), .b(n_2104), .o(n_13562) );
na02s02 TIMEBOOST_cell_38126 ( .a(TIMEBOOST_net_11301), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_4569) );
na02f02 TIMEBOOST_cell_38918 ( .a(TIMEBOOST_net_11697), .b(FE_OFN2200_n_10256), .o(TIMEBOOST_net_10704) );
na02f02 g53823_u0 ( .a(n_13361), .b(n_2108), .o(n_13561) );
na02f02 g53824_u0 ( .a(n_13495), .b(n_2106), .o(n_13704) );
na02f02 g53825_u0 ( .a(n_13455), .b(n_2105), .o(n_13664) );
na02f02 g53826_u0 ( .a(n_13454), .b(n_1793), .o(n_13663) );
na02f02 g53827_u0 ( .a(n_13453), .b(n_2102), .o(n_13662) );
na02f02 TIMEBOOST_cell_38920 ( .a(TIMEBOOST_net_11698), .b(FE_OFN2198_n_10256), .o(TIMEBOOST_net_10085) );
na02f02 g53829_u0 ( .a(n_13360), .b(FE_OFN2249_n_1790), .o(n_13560) );
in01f06 g53839_u0 ( .a(n_13703), .o(n_13997) );
in01f04 g53848_u0 ( .a(n_13701), .o(n_13995) );
in01f02 g53856_u0 ( .a(n_16206), .o(n_13736) );
na02f02 g53858_u0 ( .a(n_13449), .b(n_2110), .o(n_13659) );
na02f02 g53859_u0 ( .a(n_13446), .b(n_2121), .o(n_13658) );
na02f02 g53860_u0 ( .a(n_13445), .b(n_2103), .o(n_13657) );
na02m02 TIMEBOOST_cell_36263 ( .a(n_1381), .b(n_3192), .o(TIMEBOOST_net_10370) );
na02f02 g53863_u0 ( .a(n_13441), .b(n_4692), .o(n_13654) );
na02f02 g53864_u0 ( .a(n_13439), .b(n_2119), .o(n_13653) );
no02f04 TIMEBOOST_cell_19041 ( .a(TIMEBOOST_net_4777), .b(FE_RN_377_0), .o(TIMEBOOST_net_649) );
na02f02 TIMEBOOST_cell_41486 ( .a(TIMEBOOST_net_12981), .b(g57045_sb), .o(n_11689) );
na02s01 TIMEBOOST_cell_38128 ( .a(TIMEBOOST_net_11302), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_4487) );
na02f02 g53868_u0 ( .a(n_13435), .b(FE_OFN1936_n_1781), .o(n_13649) );
oa12m02 g53870_u0 ( .a(n_13434), .b(n_4712), .c(FE_OFN2072_n_15978), .o(n_13648) );
oa12f02 g53871_u0 ( .a(n_13432), .b(n_4200), .c(FE_OFN2072_n_15978), .o(n_13647) );
oa12f02 g53872_u0 ( .a(n_13431), .b(n_4161), .c(FE_OFN1000_n_15978), .o(n_13646) );
oa12m02 g53873_u0 ( .a(n_13430), .b(n_3474), .c(FE_OFN2072_n_15978), .o(n_13645) );
oa12m02 g53874_u0 ( .a(n_13359), .b(n_4206), .c(FE_OFN1000_n_15978), .o(n_13559) );
oa12m02 g53875_u0 ( .a(n_13429), .b(n_4714), .c(FE_OFN2072_n_15978), .o(n_13643) );
oa12m02 g53876_u0 ( .a(n_13428), .b(n_4668), .c(FE_OFN1000_n_15978), .o(n_13642) );
oa12f02 g53877_u0 ( .a(n_13427), .b(n_4201), .c(FE_OFN1000_n_15978), .o(n_13641) );
oa12m02 g53878_u0 ( .a(n_13358), .b(n_4886), .c(FE_OFN1000_n_15978), .o(n_13558) );
oa12m02 g53879_u0 ( .a(n_13490), .b(n_5753), .c(FE_OFN2072_n_15978), .o(n_13695) );
oa12m02 g53880_u0 ( .a(n_13426), .b(n_4862), .c(FE_OFN1000_n_15978), .o(n_13640) );
oa12f02 g53881_u0 ( .a(n_13425), .b(n_4700), .c(FE_OFN2072_n_15978), .o(n_13638) );
oa12m02 g53882_u0 ( .a(n_13424), .b(n_7341), .c(FE_OFN1000_n_15978), .o(n_13636) );
oa12m02 g53883_u0 ( .a(n_13357), .b(n_7362), .c(FE_OFN1000_n_15978), .o(n_13557) );
oa12f02 g53884_u0 ( .a(n_13423), .b(n_5731), .c(FE_OFN1001_n_15978), .o(n_13635) );
oa12m02 g53885_u0 ( .a(n_13422), .b(n_4158), .c(FE_OFN1001_n_15978), .o(n_13634) );
oa12m02 g53886_u0 ( .a(n_13421), .b(n_3477), .c(FE_OFN1001_n_15978), .o(n_13632) );
oa12m02 g53887_u0 ( .a(n_13420), .b(n_3484), .c(FE_OFN1001_n_15978), .o(n_13631) );
oa12m02 g53888_u0 ( .a(n_13419), .b(n_4157), .c(FE_OFN1001_n_15978), .o(n_13629) );
oa12m02 g53889_u0 ( .a(n_13418), .b(n_3479), .c(FE_OFN1000_n_15978), .o(n_13628) );
na02s02 TIMEBOOST_cell_36776 ( .a(TIMEBOOST_net_10626), .b(FE_OFN877_g64577_p), .o(TIMEBOOST_net_4677) );
na02s01 g65679_u1 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(g65679_sb), .o(g65679_da) );
na02s02 TIMEBOOST_cell_36730 ( .a(TIMEBOOST_net_10603), .b(g63608_sb), .o(n_4760) );
na02s01 TIMEBOOST_cell_43278 ( .a(TIMEBOOST_net_13877), .b(g62039_sb), .o(n_7776) );
na02s01 g53891_u2 ( .a(n_13548), .b(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(g53891_db) );
na02s02 TIMEBOOST_cell_38130 ( .a(TIMEBOOST_net_11303), .b(FE_OFN1139_g64577_p), .o(TIMEBOOST_net_4560) );
in01s04 g53892_u0 ( .a(n_692), .o(g53892_sb) );
na02s01 TIMEBOOST_cell_38132 ( .a(TIMEBOOST_net_11304), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_4561) );
na02s01 g53892_u2 ( .a(n_13544), .b(n_692), .o(g53892_db) );
na02s01 TIMEBOOST_cell_18507 ( .a(TIMEBOOST_net_4510), .b(g62810_sb), .o(n_5358) );
na02f02 TIMEBOOST_cell_44238 ( .a(TIMEBOOST_net_14357), .b(FE_OFN1405_n_8567), .o(TIMEBOOST_net_12757) );
na02s01 g53893_u2 ( .a(n_13541), .b(n_692), .o(g53893_db) );
na02s02 TIMEBOOST_cell_18523 ( .a(TIMEBOOST_net_4518), .b(g62834_sb), .o(n_5305) );
ao12s01 g53894_u0 ( .a(n_13494), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__Q), .c(n_1041), .o(n_13692) );
ao12s01 g53895_u0 ( .a(n_13493), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__Q), .c(n_1041), .o(n_13691) );
ao12s01 g53896_u0 ( .a(n_13491), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__Q), .c(n_1041), .o(n_13689) );
in01s03 g53897_u0 ( .a(FE_OFN2072_n_15978), .o(g53897_sb) );
na02s01 TIMEBOOST_cell_43398 ( .a(TIMEBOOST_net_13937), .b(n_6287), .o(TIMEBOOST_net_11578) );
na02f02 TIMEBOOST_cell_41685 ( .a(FE_OFN1759_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q), .o(TIMEBOOST_net_13081) );
na02m02 TIMEBOOST_cell_44563 ( .a(n_9102), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__Q), .o(TIMEBOOST_net_14520) );
in01s01 g53898_u0 ( .a(FE_OFN1330_n_13547), .o(g53898_sb) );
na02s01 TIMEBOOST_cell_36255 ( .a(n_875), .b(n_2235), .o(TIMEBOOST_net_10366) );
na03s02 TIMEBOOST_cell_38061 ( .a(g64291_da), .b(g64291_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__Q), .o(TIMEBOOST_net_11269) );
na03s02 TIMEBOOST_cell_38921 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__Q), .b(FE_OFN1124_g64577_p), .c(n_4009), .o(TIMEBOOST_net_11699) );
in01s01 g53899_u0 ( .a(FE_OFN1330_n_13547), .o(g53899_sb) );
na04f04 TIMEBOOST_cell_36233 ( .a(n_13049), .b(n_12884), .c(n_12785), .d(n_12883), .o(n_13132) );
na02s02 TIMEBOOST_cell_38134 ( .a(TIMEBOOST_net_11305), .b(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_4696) );
na02s01 TIMEBOOST_cell_3890 ( .a(n_14079), .b(parchk_pci_serr_out_in), .o(TIMEBOOST_net_525) );
in01s01 g53900_u0 ( .a(FE_OFN1330_n_13547), .o(g53900_sb) );
na04f04 TIMEBOOST_cell_36235 ( .a(n_13065), .b(n_12932), .c(n_12801), .d(n_12931), .o(n_13142) );
na02s01 TIMEBOOST_cell_3891 ( .a(TIMEBOOST_net_525), .b(n_7739), .o(n_14491) );
na03s02 TIMEBOOST_cell_38107 ( .a(TIMEBOOST_net_4266), .b(g64092_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__Q), .o(TIMEBOOST_net_11292) );
in01m01 g53901_u0 ( .a(FE_OFN1333_n_13547), .o(g53901_sb) );
na02s01 TIMEBOOST_cell_9947 ( .a(TIMEBOOST_net_1540), .b(g65858_sb), .o(n_2577) );
na02f02 TIMEBOOST_cell_12972 ( .a(FE_OFN1746_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__Q), .o(TIMEBOOST_net_3053) );
na02s01 TIMEBOOST_cell_17118 ( .a(pci_target_unit_del_sync_addr_in_216), .b(parchk_pci_ad_reg_in_1217), .o(TIMEBOOST_net_3816) );
in01s01 g53902_u0 ( .a(FE_OFN1331_n_13547), .o(g53902_sb) );
na02s02 TIMEBOOST_cell_36259 ( .a(n_2967), .b(n_940), .o(TIMEBOOST_net_10368) );
na02s01 TIMEBOOST_cell_42602 ( .a(TIMEBOOST_net_13539), .b(g58010_sb), .o(TIMEBOOST_net_11939) );
na02s01 TIMEBOOST_cell_17663 ( .a(TIMEBOOST_net_4088), .b(g65308_db), .o(n_4272) );
in01s01 g53903_u0 ( .a(FE_OFN1326_n_13547), .o(g53903_sb) );
na02s01 TIMEBOOST_cell_9951 ( .a(TIMEBOOST_net_1542), .b(g65858_sb), .o(n_2593) );
na02f02 TIMEBOOST_cell_3897 ( .a(TIMEBOOST_net_528), .b(g54316_sb), .o(n_13010) );
na03s02 TIMEBOOST_cell_43015 ( .a(n_4056), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__Q), .c(FE_OFN1119_g64577_p), .o(TIMEBOOST_net_13746) );
in01s01 g53904_u0 ( .a(FE_OFN1330_n_13547), .o(g53904_sb) );
na02s01 TIMEBOOST_cell_9975 ( .a(TIMEBOOST_net_1554), .b(g65858_sb), .o(n_2588) );
na02s01 TIMEBOOST_cell_44856 ( .a(TIMEBOOST_net_14666), .b(g58384_sb), .o(TIMEBOOST_net_12444) );
na02f02 TIMEBOOST_cell_41110 ( .a(TIMEBOOST_net_12793), .b(g57552_sb), .o(n_10810) );
in01s02 g53905_u0 ( .a(FE_OFN1332_n_13547), .o(g53905_sb) );
na02s01 TIMEBOOST_cell_9945 ( .a(TIMEBOOST_net_1539), .b(g65858_sb), .o(n_2581) );
na02f02 TIMEBOOST_cell_3901 ( .a(TIMEBOOST_net_530), .b(FE_OFN1942_n_3241), .o(n_4879) );
na02s01 TIMEBOOST_cell_43137 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__Q), .b(n_4432), .o(TIMEBOOST_net_13807) );
in01s01 g53906_u0 ( .a(FE_OFN1331_n_13547), .o(g53906_sb) );
na02s01 TIMEBOOST_cell_9977 ( .a(TIMEBOOST_net_1555), .b(g65858_sb), .o(n_2482) );
na02f02 TIMEBOOST_cell_3903 ( .a(TIMEBOOST_net_531), .b(n_3367), .o(n_5232) );
na02s02 TIMEBOOST_cell_38136 ( .a(TIMEBOOST_net_11306), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_4529) );
in01s01 g53907_u0 ( .a(FE_OFN1331_n_13547), .o(g53907_sb) );
na03f02 TIMEBOOST_cell_36201 ( .a(FE_OCP_RBN1973_n_12381), .b(TIMEBOOST_net_10294), .c(n_11831), .o(n_12723) );
na02f02 TIMEBOOST_cell_42406 ( .a(TIMEBOOST_net_13441), .b(g57214_sb), .o(n_10438) );
na02s02 TIMEBOOST_cell_3906 ( .a(g52635_db), .b(n_8757), .o(TIMEBOOST_net_533) );
in01s01 g53908_u0 ( .a(FE_OFN1331_n_13547), .o(g53908_sb) );
na02s01 TIMEBOOST_cell_42659 ( .a(n_3792), .b(g65022_sb), .o(TIMEBOOST_net_13568) );
na02s02 TIMEBOOST_cell_3907 ( .a(TIMEBOOST_net_533), .b(g52635_da), .o(g52401_db) );
na02s02 TIMEBOOST_cell_39343 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__16__Q), .b(g64266_sb), .o(TIMEBOOST_net_11910) );
in01s01 g53909_u0 ( .a(FE_OFN1326_n_13547), .o(g53909_sb) );
na02s01 TIMEBOOST_cell_41840 ( .a(TIMEBOOST_net_13158), .b(FE_OFN563_n_9895), .o(TIMEBOOST_net_9744) );
na02s02 TIMEBOOST_cell_45608 ( .a(TIMEBOOST_net_15042), .b(g65242_sb), .o(n_2640) );
na02s01 TIMEBOOST_cell_38922 ( .a(TIMEBOOST_net_11699), .b(g62789_sb), .o(n_5412) );
in01s01 g53910_u0 ( .a(FE_OFN1332_n_13547), .o(g53910_sb) );
na02s01 TIMEBOOST_cell_15837 ( .a(TIMEBOOST_net_3175), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_411), .o(TIMEBOOST_net_71) );
na03s02 TIMEBOOST_cell_38053 ( .a(g64210_da), .b(g64210_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__Q), .o(TIMEBOOST_net_11265) );
na02f02 TIMEBOOST_cell_36674 ( .a(TIMEBOOST_net_10575), .b(g54318_sb), .o(TIMEBOOST_net_4701) );
in01s01 g53911_u0 ( .a(FE_OFN1327_n_13547), .o(g53911_sb) );
na02s01 TIMEBOOST_cell_42629 ( .a(n_3783), .b(g64898_sb), .o(TIMEBOOST_net_13553) );
na03s02 TIMEBOOST_cell_37999 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__Q), .b(FE_OFN701_n_7845), .c(n_1856), .o(TIMEBOOST_net_11238) );
na02s02 TIMEBOOST_cell_19147 ( .a(TIMEBOOST_net_4830), .b(g60681_sb), .o(TIMEBOOST_net_591) );
in01s01 g53912_u0 ( .a(FE_OFN1333_n_13547), .o(g53912_sb) );
na02s02 TIMEBOOST_cell_45735 ( .a(n_3696), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__Q), .o(TIMEBOOST_net_15106) );
na02s02 TIMEBOOST_cell_38628 ( .a(TIMEBOOST_net_11552), .b(g62488_sb), .o(n_6610) );
na02f02 TIMEBOOST_cell_41026 ( .a(TIMEBOOST_net_12751), .b(g57417_sb), .o(n_11324) );
in01s01 g53913_u0 ( .a(FE_OFN1331_n_13547), .o(g53913_sb) );
na03f02 TIMEBOOST_cell_36205 ( .a(n_12100), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__Q), .c(FE_OFN1757_n_12681), .o(n_12524) );
na03s02 TIMEBOOST_cell_37797 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__Q), .b(FE_OFN2257_n_8060), .c(n_1566), .o(TIMEBOOST_net_11137) );
na02s01 TIMEBOOST_cell_41745 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__Q), .b(g65319_sb), .o(TIMEBOOST_net_13111) );
in01s01 g53914_u0 ( .a(FE_OFN1330_n_13547), .o(g53914_sb) );
na02s01 TIMEBOOST_cell_42939 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__Q), .b(FE_OFN580_n_9531), .o(TIMEBOOST_net_13708) );
na02f02 TIMEBOOST_cell_3919 ( .a(TIMEBOOST_net_539), .b(n_13814), .o(n_7726) );
na02s02 TIMEBOOST_cell_41746 ( .a(TIMEBOOST_net_13111), .b(g65319_db), .o(n_3563) );
in01s01 g53915_u0 ( .a(FE_OFN1331_n_13547), .o(g53915_sb) );
na02s01 TIMEBOOST_cell_42940 ( .a(TIMEBOOST_net_13708), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_11153) );
na02f02 TIMEBOOST_cell_3921 ( .a(TIMEBOOST_net_540), .b(n_8538), .o(n_8659) );
na02s01 TIMEBOOST_cell_18793 ( .a(TIMEBOOST_net_4653), .b(g63175_sb), .o(n_4949) );
in01s02 g53916_u0 ( .a(FE_OFN1326_n_13547), .o(g53916_sb) );
na02f02 TIMEBOOST_cell_3923 ( .a(TIMEBOOST_net_541), .b(n_5232), .o(n_13414) );
na02s01 TIMEBOOST_cell_3924 ( .a(n_2353), .b(n_8498), .o(TIMEBOOST_net_542) );
in01s01 g53917_u0 ( .a(FE_OFN1327_n_13547), .o(g53917_sb) );
na03f02 TIMEBOOST_cell_36213 ( .a(FE_OCP_RBN1976_n_12381), .b(TIMEBOOST_net_10305), .c(FE_OFN1756_n_12681), .o(n_12638) );
na02m02 TIMEBOOST_cell_3925 ( .a(TIMEBOOST_net_542), .b(n_8538), .o(n_8575) );
na02s02 TIMEBOOST_cell_3926 ( .a(n_2367), .b(n_3498), .o(TIMEBOOST_net_543) );
in01s01 g53918_u0 ( .a(FE_OFN1327_n_13547), .o(g53918_sb) );
na02f02 TIMEBOOST_cell_18317 ( .a(TIMEBOOST_net_4415), .b(n_3079), .o(n_4145) );
na02m01 TIMEBOOST_cell_3927 ( .a(TIMEBOOST_net_543), .b(n_8572), .o(n_8573) );
na02f02 TIMEBOOST_cell_44564 ( .a(TIMEBOOST_net_14520), .b(FE_OFN2167_n_8567), .o(TIMEBOOST_net_13496) );
in01s01 g53919_u0 ( .a(FE_OFN1330_n_13547), .o(g53919_sb) );
na02s01 TIMEBOOST_cell_22208 ( .a(g52468_da), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_6361) );
na02s02 TIMEBOOST_cell_19251 ( .a(TIMEBOOST_net_4882), .b(g60659_sb), .o(n_5662) );
na02s02 TIMEBOOST_cell_3930 ( .a(n_4743), .b(n_2742), .o(TIMEBOOST_net_545) );
in01s01 g53920_u0 ( .a(FE_OFN1332_n_13547), .o(g53920_sb) );
na02s01 TIMEBOOST_cell_22272 ( .a(g52462_da), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_6393) );
na02m04 TIMEBOOST_cell_3931 ( .a(TIMEBOOST_net_545), .b(n_7108), .o(n_8468) );
na02s01 TIMEBOOST_cell_3932 ( .a(n_4743), .b(n_2308), .o(TIMEBOOST_net_546) );
in01s01 g53921_u0 ( .a(FE_OFN1331_n_13547), .o(g53921_sb) );
na03f02 TIMEBOOST_cell_36197 ( .a(FE_OCP_RBN1973_n_12381), .b(TIMEBOOST_net_10298), .c(n_11831), .o(n_12665) );
na02m02 TIMEBOOST_cell_3933 ( .a(TIMEBOOST_net_546), .b(n_7108), .o(n_8514) );
na02m02 TIMEBOOST_cell_39161 ( .a(g58796_db), .b(g58783_sb), .o(TIMEBOOST_net_11819) );
in01s01 g53922_u0 ( .a(FE_OFN1331_n_13547), .o(g53922_sb) );
na03f02 TIMEBOOST_cell_36195 ( .a(n_12066), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__Q), .c(n_11831), .o(n_12486) );
na02s02 TIMEBOOST_cell_19253 ( .a(TIMEBOOST_net_4883), .b(g60661_sb), .o(n_5658) );
na02m08 TIMEBOOST_cell_3936 ( .a(n_709), .b(n_1014), .o(TIMEBOOST_net_548) );
in01s02 g53923_u0 ( .a(FE_OFN1327_n_13547), .o(g53923_sb) );
na02s02 TIMEBOOST_cell_45736 ( .a(TIMEBOOST_net_15106), .b(FE_OFN1250_n_4093), .o(TIMEBOOST_net_13266) );
na02f08 TIMEBOOST_cell_3937 ( .a(TIMEBOOST_net_548), .b(n_7705), .o(n_8569) );
na02m02 TIMEBOOST_cell_3938 ( .a(FE_RN_420_0), .b(n_13447), .o(TIMEBOOST_net_549) );
in01s01 g53924_u0 ( .a(FE_OFN1326_n_13547), .o(g53924_sb) );
na02s01 TIMEBOOST_cell_45737 ( .a(n_4523), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__Q), .o(TIMEBOOST_net_15107) );
na02f02 TIMEBOOST_cell_3939 ( .a(TIMEBOOST_net_549), .b(FE_RN_423_0), .o(FE_RN_425_0) );
na02m02 TIMEBOOST_cell_3940 ( .a(n_504), .b(FE_RN_447_0), .o(TIMEBOOST_net_550) );
in01s01 g53925_u0 ( .a(FE_OFN1331_n_13547), .o(g53925_sb) );
na02m02 TIMEBOOST_cell_44209 ( .a(n_9474), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__Q), .o(TIMEBOOST_net_14343) );
na02f02 TIMEBOOST_cell_3941 ( .a(TIMEBOOST_net_550), .b(FE_RN_450_0), .o(FE_RN_452_0) );
na02f04 TIMEBOOST_cell_3942 ( .a(n_15918), .b(n_15908), .o(TIMEBOOST_net_551) );
in01s02 g53926_u0 ( .a(FE_OFN1327_n_13547), .o(g53926_sb) );
na02s01 TIMEBOOST_cell_45738 ( .a(TIMEBOOST_net_15107), .b(FE_OFN706_n_8119), .o(TIMEBOOST_net_11091) );
na02f06 TIMEBOOST_cell_3943 ( .a(FE_RN_895_0), .b(TIMEBOOST_net_551), .o(n_16520) );
na02s01 TIMEBOOST_cell_18659 ( .a(TIMEBOOST_net_4586), .b(g62770_sb), .o(n_5454) );
in01s01 g53927_u0 ( .a(FE_OFN1327_n_13547), .o(g53927_sb) );
na03f02 TIMEBOOST_cell_36185 ( .a(n_12081), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__Q), .c(n_11823), .o(n_12506) );
na02s02 TIMEBOOST_cell_38138 ( .a(TIMEBOOST_net_11307), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_4630) );
na02s02 TIMEBOOST_cell_19263 ( .a(TIMEBOOST_net_4888), .b(g60670_sb), .o(n_5648) );
in01s01 g53928_u0 ( .a(FE_OFN1331_n_13547), .o(g53928_sb) );
na03f02 TIMEBOOST_cell_36183 ( .a(FE_OFN1735_n_16317), .b(TIMEBOOST_net_10285), .c(FE_OFN1739_n_11019), .o(n_12743) );
na02s02 TIMEBOOST_cell_19261 ( .a(TIMEBOOST_net_4887), .b(g60610_sb), .o(n_4844) );
na02s02 TIMEBOOST_cell_19267 ( .a(TIMEBOOST_net_4890), .b(g60619_sb), .o(n_4835) );
in01m01 g53929_u0 ( .a(FE_OFN1333_n_13547), .o(g53929_sb) );
na03f02 TIMEBOOST_cell_36157 ( .a(FE_RN_496_0), .b(FE_OFN1572_n_11027), .c(TIMEBOOST_net_10278), .o(FE_RN_498_0) );
na03s02 TIMEBOOST_cell_38079 ( .a(TIMEBOOST_net_4259), .b(g64170_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__Q), .o(TIMEBOOST_net_11278) );
na02s02 TIMEBOOST_cell_19269 ( .a(TIMEBOOST_net_4891), .b(g60621_sb), .o(n_4833) );
in01s02 g53930_u0 ( .a(FE_OFN1327_n_13547), .o(g53930_sb) );
na03f02 TIMEBOOST_cell_36159 ( .a(FE_OFN2209_n_11027), .b(TIMEBOOST_net_10275), .c(FE_OFN1752_n_12086), .o(n_12758) );
na02s01 TIMEBOOST_cell_39312 ( .a(TIMEBOOST_net_11894), .b(g65894_db), .o(n_1717) );
no02f02 TIMEBOOST_cell_42527 ( .a(TIMEBOOST_net_664), .b(FE_RN_573_0), .o(TIMEBOOST_net_13502) );
in01s01 g53931_u0 ( .a(FE_OFN1331_n_13547), .o(g53931_sb) );
na03f02 TIMEBOOST_cell_36161 ( .a(FE_OFN1753_n_12086), .b(TIMEBOOST_net_10270), .c(FE_OFN1568_n_11027), .o(n_12650) );
na02f02 TIMEBOOST_cell_3953 ( .a(TIMEBOOST_net_556), .b(g54152_da), .o(n_13448) );
na02s02 TIMEBOOST_cell_19279 ( .a(TIMEBOOST_net_4896), .b(g60634_sb), .o(n_5702) );
in01s01 g53932_u0 ( .a(FE_OFN1326_n_13547), .o(g53932_sb) );
na04f02 TIMEBOOST_cell_36163 ( .a(n_11773), .b(n_11040), .c(n_11041), .d(n_11039), .o(n_12530) );
na02s01 TIMEBOOST_cell_37991 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__Q), .b(FE_OFN881_g64577_p), .o(TIMEBOOST_net_11234) );
na02s01 TIMEBOOST_cell_37894 ( .a(TIMEBOOST_net_11185), .b(g58239_sb), .o(n_9552) );
na02f04 TIMEBOOST_cell_22313 ( .a(n_10257), .b(TIMEBOOST_net_6413), .o(n_11869) );
ao22f01 g53934_u0 ( .a(pci_target_unit_wishbone_master_retried), .b(wbm_cyc_o_1378), .c(wbm_ack_i), .d(wbm_stb_o), .o(n_13790) );
na02s02 TIMEBOOST_cell_40874 ( .a(TIMEBOOST_net_12675), .b(g62477_sb), .o(n_6634) );
na02s02 TIMEBOOST_cell_37938 ( .a(TIMEBOOST_net_11207), .b(g58355_sb), .o(n_9467) );
na02s01 TIMEBOOST_cell_43279 ( .a(TIMEBOOST_net_4774), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_13878) );
na02s02 TIMEBOOST_cell_36294 ( .a(TIMEBOOST_net_10385), .b(n_1342), .o(n_2402) );
na02m02 TIMEBOOST_cell_41519 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__Q), .b(n_9639), .o(TIMEBOOST_net_12998) );
na02s02 TIMEBOOST_cell_43506 ( .a(TIMEBOOST_net_13991), .b(FE_OFN1231_n_6391), .o(TIMEBOOST_net_12624) );
in01s01 g53937_u0 ( .a(FE_OFN2072_n_15978), .o(g53937_sb) );
na02m02 TIMEBOOST_cell_12612 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__Q), .o(TIMEBOOST_net_2873) );
na03s02 TIMEBOOST_cell_36761 ( .a(TIMEBOOST_net_4270), .b(g64211_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q), .o(TIMEBOOST_net_10619) );
na02s02 TIMEBOOST_cell_36732 ( .a(TIMEBOOST_net_10604), .b(g63610_sb), .o(n_4758) );
na02s01 TIMEBOOST_cell_3440 ( .a(FE_OFN252_n_9868), .b(g58136_sb), .o(TIMEBOOST_net_300) );
na02s01 g65076_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__Q), .b(FE_OFN662_n_4392), .o(g65076_db) );
na02f02 TIMEBOOST_cell_38654 ( .a(TIMEBOOST_net_11565), .b(n_14618), .o(TIMEBOOST_net_10689) );
in01s01 g53939_u0 ( .a(FE_OFN1001_n_15978), .o(g53939_sb) );
na02f02 TIMEBOOST_cell_43832 ( .a(TIMEBOOST_net_14154), .b(FE_OFN1423_n_8567), .o(TIMEBOOST_net_12951) );
na02m02 TIMEBOOST_cell_43833 ( .a(n_9517), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__Q), .o(TIMEBOOST_net_14155) );
na02f02 TIMEBOOST_cell_43834 ( .a(TIMEBOOST_net_14155), .b(FE_OFN1424_n_8567), .o(TIMEBOOST_net_12823) );
in01s01 g53940_u0 ( .a(FE_OFN1001_n_15978), .o(g53940_sb) );
na02s01 TIMEBOOST_cell_37249 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__Q), .b(n_3792), .o(TIMEBOOST_net_10863) );
na02s02 TIMEBOOST_cell_2903 ( .a(TIMEBOOST_net_31), .b(n_1187), .o(n_2009) );
na02s02 TIMEBOOST_cell_45261 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__Q), .b(n_3564), .o(TIMEBOOST_net_14869) );
na02f04 TIMEBOOST_cell_36296 ( .a(TIMEBOOST_net_10386), .b(FE_RN_600_0), .o(FE_RN_601_0) );
in01s01 TIMEBOOST_cell_45951 ( .a(wbm_dat_i_4_), .o(TIMEBOOST_net_15258) );
na02m02 TIMEBOOST_cell_44505 ( .a(n_9450), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__Q), .o(TIMEBOOST_net_14491) );
na02s02 TIMEBOOST_cell_43057 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__Q), .b(n_3694), .o(TIMEBOOST_net_13767) );
na02s01 TIMEBOOST_cell_41722 ( .a(TIMEBOOST_net_13099), .b(g64829_db), .o(n_3731) );
no02f06 TIMEBOOST_cell_36298 ( .a(TIMEBOOST_net_10387), .b(FE_RN_685_0), .o(TIMEBOOST_net_129) );
na02s02 g53943_u1 ( .a(conf_wb_err_bc_in_847), .b(g53939_sb), .o(g53943_da) );
na02s02 TIMEBOOST_cell_36734 ( .a(TIMEBOOST_net_10605), .b(g63615_sb), .o(n_4753) );
na02s02 g53944_u1 ( .a(conf_wb_err_bc_in_848), .b(g53939_sb), .o(g53944_da) );
na02m02 TIMEBOOST_cell_44351 ( .a(n_9897), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q), .o(TIMEBOOST_net_14414) );
na02s02 TIMEBOOST_cell_37896 ( .a(TIMEBOOST_net_11186), .b(g57992_sb), .o(n_9804) );
na02s02 g53945_u1 ( .a(conf_wb_err_bc_in), .b(g53939_sb), .o(g53945_da) );
na02s02 TIMEBOOST_cell_37926 ( .a(TIMEBOOST_net_11201), .b(FE_OFN1670_n_9477), .o(TIMEBOOST_net_4352) );
in01s01 g53946_u0 ( .a(FE_OFN2072_n_15978), .o(g53946_sb) );
na04f02 TIMEBOOST_cell_36165 ( .a(n_11781), .b(n_11070), .c(n_11069), .d(n_11071), .o(n_12538) );
na02s02 TIMEBOOST_cell_2905 ( .a(TIMEBOOST_net_32), .b(n_1186), .o(n_2007) );
na02s02 TIMEBOOST_cell_45262 ( .a(TIMEBOOST_net_14869), .b(FE_OFN1289_n_4098), .o(TIMEBOOST_net_12062) );
na02s01 g53947_u1 ( .a(wishbone_slave_unit_pci_initiator_if_current_byte_address_36), .b(FE_OFN2071_n_15978), .o(g53947_da) );
na02s02 TIMEBOOST_cell_45263 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__20__Q), .b(n_3690), .o(TIMEBOOST_net_14870) );
na02s02 TIMEBOOST_cell_37898 ( .a(TIMEBOOST_net_11187), .b(g57923_sb), .o(n_9887) );
na02s01 TIMEBOOST_cell_37211 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__Q), .b(g65852_sb), .o(TIMEBOOST_net_10844) );
no02f02 TIMEBOOST_cell_10951 ( .a(FE_RN_542_0), .b(TIMEBOOST_net_2042), .o(TIMEBOOST_net_926) );
na02s01 TIMEBOOST_cell_36370 ( .a(TIMEBOOST_net_10423), .b(TIMEBOOST_net_3229), .o(n_1574) );
na02s01 TIMEBOOST_cell_36372 ( .a(TIMEBOOST_net_10424), .b(TIMEBOOST_net_3228), .o(n_1586) );
na02s01 TIMEBOOST_cell_38002 ( .a(TIMEBOOST_net_11239), .b(g61737_sb), .o(n_8344) );
na02s01 TIMEBOOST_cell_36374 ( .a(TIMEBOOST_net_10425), .b(g65912_db), .o(n_1569) );
na02s02 TIMEBOOST_cell_38004 ( .a(TIMEBOOST_net_11240), .b(g61782_sb), .o(n_8241) );
na02s01 TIMEBOOST_cell_38634 ( .a(TIMEBOOST_net_11555), .b(g59112_sb), .o(n_8701) );
na02f02 TIMEBOOST_cell_45806 ( .a(TIMEBOOST_net_15141), .b(FE_OFN2182_n_8567), .o(TIMEBOOST_net_14575) );
na02m06 TIMEBOOST_cell_36300 ( .a(wbu_addr_in_264), .b(TIMEBOOST_net_10388), .o(TIMEBOOST_net_124) );
na02f04 TIMEBOOST_cell_37130 ( .a(TIMEBOOST_net_10803), .b(n_12560), .o(n_12822) );
na02s01 TIMEBOOST_cell_38006 ( .a(TIMEBOOST_net_11241), .b(g61825_sb), .o(n_8137) );
na02s01 TIMEBOOST_cell_43507 ( .a(n_3577), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__Q), .o(TIMEBOOST_net_13992) );
na03s02 TIMEBOOST_cell_33583 ( .a(TIMEBOOST_net_9560), .b(n_5633), .c(g62101_sb), .o(n_5601) );
na02s02 TIMEBOOST_cell_43508 ( .a(TIMEBOOST_net_13992), .b(FE_OFN1231_n_6391), .o(TIMEBOOST_net_12636) );
na02s02 TIMEBOOST_cell_38008 ( .a(TIMEBOOST_net_11242), .b(g61991_sb), .o(n_7913) );
na03s02 TIMEBOOST_cell_33582 ( .a(TIMEBOOST_net_9561), .b(n_5633), .c(g62094_sb), .o(n_5611) );
na02f02 TIMEBOOST_cell_42408 ( .a(TIMEBOOST_net_13442), .b(g57364_sb), .o(n_11383) );
na02s01 TIMEBOOST_cell_36302 ( .a(TIMEBOOST_net_10389), .b(FE_OFN936_n_2292), .o(TIMEBOOST_net_3311) );
na02s01 TIMEBOOST_cell_43399 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__Q), .b(n_4302), .o(TIMEBOOST_net_13938) );
na02m02 TIMEBOOST_cell_43835 ( .a(n_9829), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__Q), .o(TIMEBOOST_net_14156) );
na02s01 g64856_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__Q), .b(FE_OFN689_n_4438), .o(g64856_db) );
in01f02 g53980_u0 ( .a(n_13679), .o(n_13625) );
na02s02 TIMEBOOST_cell_16821 ( .a(TIMEBOOST_net_3667), .b(g65323_db), .o(n_3560) );
no02f02 TIMEBOOST_cell_37132 ( .a(TIMEBOOST_net_10804), .b(n_14434), .o(FE_RN_847_0) );
na02s01 TIMEBOOST_cell_39450 ( .a(TIMEBOOST_net_11963), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_4606) );
na02f04 TIMEBOOST_cell_37094 ( .a(TIMEBOOST_net_10785), .b(n_12577), .o(n_12839) );
na02s02 TIMEBOOST_cell_2907 ( .a(TIMEBOOST_net_33), .b(n_1186), .o(n_1426) );
na02s02 TIMEBOOST_cell_36890 ( .a(TIMEBOOST_net_10683), .b(g58598_da), .o(n_8855) );
na02s02 TIMEBOOST_cell_38010 ( .a(TIMEBOOST_net_11243), .b(g62017_sb), .o(n_7861) );
no02f02 g53988_u0 ( .a(n_15370), .b(wishbone_slave_unit_wbs_sm_wbr_control_in_190), .o(n_1645) );
na02s01 g53990_u0 ( .a(n_1684), .b(wishbone_slave_unit_wbs_sm_wbr_control_in_190), .o(g53990_p) );
in01s01 g53990_u1 ( .a(g53990_p), .o(n_1979) );
no02s01 g53991_u0 ( .a(n_13329), .b(n_1041), .o(n_13494) );
no02s01 g53992_u0 ( .a(n_13328), .b(n_1041), .o(n_13493) );
no02s01 g53993_u0 ( .a(n_13327), .b(n_1041), .o(n_13491) );
na02s02 TIMEBOOST_cell_43167 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__Q), .b(n_3671), .o(TIMEBOOST_net_13822) );
na02m02 TIMEBOOST_cell_41661 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_27__Q), .o(TIMEBOOST_net_13069) );
na02s01 TIMEBOOST_cell_9061 ( .a(TIMEBOOST_net_1097), .b(g66456_db), .o(n_1532) );
na02f02 TIMEBOOST_cell_22619 ( .a(TIMEBOOST_net_6566), .b(FE_OFN1566_n_12502), .o(n_12660) );
na02s01 TIMEBOOST_cell_43280 ( .a(TIMEBOOST_net_13878), .b(g62053_sb), .o(n_7756) );
na02s02 TIMEBOOST_cell_43168 ( .a(TIMEBOOST_net_13822), .b(FE_OFN1247_n_4093), .o(TIMEBOOST_net_11550) );
in01f08 g53_u0 ( .a(n_15929), .o(n_4743) );
na02f02 TIMEBOOST_cell_22621 ( .a(TIMEBOOST_net_6567), .b(FE_OFN1562_n_12502), .o(n_12655) );
na02s02 TIMEBOOST_cell_38140 ( .a(TIMEBOOST_net_11308), .b(FE_OFN1125_g64577_p), .o(TIMEBOOST_net_4686) );
na02s01 TIMEBOOST_cell_15871 ( .a(TIMEBOOST_net_3192), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_406), .o(TIMEBOOST_net_68) );
na02s02 TIMEBOOST_cell_30891 ( .a(TIMEBOOST_net_9356), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_3742) );
na02s01 TIMEBOOST_cell_30892 ( .a(pci_target_unit_pcit_if_strd_addr_in_705), .b(pci_target_unit_del_sync_addr_in_223), .o(TIMEBOOST_net_9357) );
na02m02 TIMEBOOST_cell_43086 ( .a(TIMEBOOST_net_13781), .b(g54176_da), .o(n_13511) );
na02f02 TIMEBOOST_cell_42510 ( .a(TIMEBOOST_net_13493), .b(g57049_sb), .o(n_11686) );
na02s02 TIMEBOOST_cell_37998 ( .a(TIMEBOOST_net_11237), .b(TIMEBOOST_net_1726), .o(n_14679) );
na02f02 TIMEBOOST_cell_32549 ( .a(FE_OFN1749_n_12004), .b(TIMEBOOST_net_10185), .o(TIMEBOOST_net_6424) );
na02m02 TIMEBOOST_cell_11485 ( .a(n_14390), .b(TIMEBOOST_net_2309), .o(n_14396) );
na02s01 TIMEBOOST_cell_30951 ( .a(TIMEBOOST_net_9386), .b(g64848_db), .o(n_4435) );
na02s01 TIMEBOOST_cell_45126 ( .a(TIMEBOOST_net_14801), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_11398) );
na02s01 TIMEBOOST_cell_15868 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_91), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3191) );
na02s01 TIMEBOOST_cell_37212 ( .a(TIMEBOOST_net_10844), .b(g65852_db), .o(n_1584) );
ao12f02 g54015_u0 ( .a(n_7084), .b(n_13027), .c(n_13354), .o(n_13355) );
ao12f02 g54016_u0 ( .a(n_7083), .b(n_13026), .c(n_7822), .o(n_13353) );
ao12f02 g54018_u0 ( .a(n_7082), .b(n_13022), .c(n_13354), .o(n_13350) );
ao12f02 g54019_u0 ( .a(n_7081), .b(n_13020), .c(n_13354), .o(n_13349) );
ao12f02 g54020_u0 ( .a(n_7080), .b(n_13018), .c(n_13354), .o(n_13348) );
na02s01 g54022_u0 ( .a(n_2027), .b(wbm_cyc_o), .o(n_13789) );
ao12f02 g54023_u0 ( .a(n_7320), .b(n_12985), .c(n_7822), .o(n_13346) );
in01s02 g54024_u0 ( .a(n_13813), .o(n_13732) );
no02m02 g54025_u0 ( .a(wishbone_slave_unit_wbs_sm_wbr_control_in_190), .b(wishbone_slave_unit_wbs_sm_wbr_control_in), .o(n_13813) );
ao12f02 g54029_u0 ( .a(n_7707), .b(n_13098), .c(n_13354), .o(n_13417) );
in01s02 g54030_u0 ( .a(n_12595), .o(g54030_sb) );
no02f02 TIMEBOOST_cell_42528 ( .a(TIMEBOOST_net_13502), .b(TIMEBOOST_net_2890), .o(TIMEBOOST_net_6240) );
no02f02 TIMEBOOST_cell_11466 ( .a(FE_OFN1706_n_4868), .b(FE_RN_361_0), .o(TIMEBOOST_net_2300) );
na02s01 TIMEBOOST_cell_43281 ( .a(TIMEBOOST_net_4772), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_13879) );
ao22f02 g54031_u0 ( .a(n_7338), .b(n_13415), .c(n_13102), .d(n_13341), .o(n_13416) );
ao22f02 g54032_u0 ( .a(n_7504), .b(n_13415), .c(n_13012), .d(n_13341), .o(n_13342) );
ao22f02 g54033_u0 ( .a(n_12986), .b(n_13341), .c(n_8488), .d(n_13415), .o(n_13340) );
ao12f02 g54034_u0 ( .a(n_7046), .b(n_12998), .c(n_13354), .o(n_13339) );
ao12f02 g54035_u0 ( .a(n_7045), .b(n_12994), .c(n_13354), .o(n_13338) );
ao12f02 g54036_u0 ( .a(n_7075), .b(n_12992), .c(n_13354), .o(n_13337) );
in01s01 g54038_u0 ( .a(parchk_pci_par_en_in), .o(g54038_sb) );
na03s02 TIMEBOOST_cell_38385 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__Q), .b(FE_OFN1134_g64577_p), .c(n_4026), .o(TIMEBOOST_net_11431) );
na02s01 g54038_u2 ( .a(pci_par_i), .b(parchk_pci_par_en_in), .o(g54038_db) );
na02s01 TIMEBOOST_cell_18023 ( .a(TIMEBOOST_net_4268), .b(g63538_db), .o(n_4617) );
in01s01 g54039_u0 ( .a(n_12595), .o(g54039_sb) );
na02s02 TIMEBOOST_cell_37928 ( .a(TIMEBOOST_net_11202), .b(g57979_sb), .o(n_9820) );
na02s01 TIMEBOOST_cell_38636 ( .a(TIMEBOOST_net_11556), .b(g59110_sb), .o(n_8708) );
na02f02 g54039_u3 ( .a(g54039_da), .b(g54039_db), .o(n_13334) );
in01m02 g54040_u0 ( .a(n_7822), .o(g54040_sb) );
na02f02 TIMEBOOST_cell_44352 ( .a(TIMEBOOST_net_14414), .b(FE_OFN1385_n_8567), .o(TIMEBOOST_net_12853) );
na02s02 TIMEBOOST_cell_43466 ( .a(TIMEBOOST_net_13971), .b(FE_OFN1235_n_6391), .o(TIMEBOOST_net_12159) );
na02s02 TIMEBOOST_cell_45264 ( .a(TIMEBOOST_net_14870), .b(FE_OFN1207_n_6356), .o(TIMEBOOST_net_12109) );
in01s01 g54044_u0 ( .a(wbm_cyc_o_1378), .o(wbm_cyc_o) );
na02f02 TIMEBOOST_cell_38842 ( .a(TIMEBOOST_net_11659), .b(g58475_sb), .o(n_9366) );
na02f02 g54118_u0 ( .a(n_13010), .b(n_12595), .o(n_13292) );
na02s01 TIMEBOOST_cell_36498 ( .a(TIMEBOOST_net_10487), .b(g66415_sb), .o(n_2510) );
in01s01 TIMEBOOST_cell_32826 ( .a(TIMEBOOST_net_10327), .o(wbs_dat_i_5_) );
na02s01 TIMEBOOST_cell_42739 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__Q), .b(n_1581), .o(TIMEBOOST_net_13608) );
na02s02 TIMEBOOST_cell_43668 ( .a(TIMEBOOST_net_14072), .b(FE_OFN1231_n_6391), .o(TIMEBOOST_net_12631) );
na02f03 g54123_u0 ( .a(n_13000), .b(n_13341), .o(n_13286) );
in01s01 g54125_u0 ( .a(n_13332), .o(n_13333) );
na02s01 TIMEBOOST_cell_40406 ( .a(g63605_da), .b(TIMEBOOST_net_12441), .o(n_7165) );
ao12f02 g54127_u0 ( .a(n_13306), .b(n_13486), .c(wbm_sel_o_0_), .o(n_13488) );
ao12f02 g54128_u0 ( .a(n_13305), .b(n_13486), .c(wbm_sel_o_1_), .o(n_13487) );
ao12f02 g54129_u0 ( .a(n_13303), .b(n_13486), .c(wbm_sel_o_2_), .o(n_13485) );
ao12f02 g54130_u0 ( .a(n_13302), .b(n_13486), .c(wbm_sel_o_3_), .o(n_13484) );
in01f02 g54131_u0 ( .a(FE_OFN2125_n_16497), .o(g54131_sb) );
na02f04 g54131_u1 ( .a(n_13145), .b(g54131_sb), .o(g54131_da) );
na02f02 TIMEBOOST_cell_43836 ( .a(TIMEBOOST_net_14156), .b(FE_OFN1400_n_8567), .o(TIMEBOOST_net_12824) );
na02s02 TIMEBOOST_cell_41808 ( .a(TIMEBOOST_net_13142), .b(g64870_sb), .o(n_4424) );
in01m01 g54132_u0 ( .a(FE_OFN1150_n_13249), .o(g54132_sb) );
na02f02 TIMEBOOST_cell_39103 ( .a(TIMEBOOST_net_10211), .b(FE_OFN1513_n_14987), .o(TIMEBOOST_net_11790) );
na02s02 TIMEBOOST_cell_36800 ( .a(TIMEBOOST_net_10638), .b(FE_OFN877_g64577_p), .o(TIMEBOOST_net_4492) );
na02s01 TIMEBOOST_cell_39452 ( .a(TIMEBOOST_net_11964), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_4541) );
in01f02 g54133_u0 ( .a(FE_OFN1150_n_13249), .o(g54133_sb) );
na03s02 TIMEBOOST_cell_38371 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__Q), .b(FE_OFN1130_g64577_p), .c(n_3953), .o(TIMEBOOST_net_11424) );
na02s02 TIMEBOOST_cell_45609 ( .a(TIMEBOOST_net_9367), .b(FE_OFN789_n_2678), .o(TIMEBOOST_net_15043) );
na02s01 TIMEBOOST_cell_38066 ( .a(TIMEBOOST_net_11271), .b(FE_OFN877_g64577_p), .o(TIMEBOOST_net_4568) );
in01f01 g54134_u0 ( .a(FE_OFN1151_n_13249), .o(g54134_sb) );
na02f02 TIMEBOOST_cell_44565 ( .a(n_9129), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__Q), .o(TIMEBOOST_net_14521) );
in01s01 TIMEBOOST_cell_45952 ( .a(TIMEBOOST_net_15258), .o(TIMEBOOST_net_15259) );
in01m01 g54135_u0 ( .a(FE_OFN1149_n_13249), .o(g54135_sb) );
na02s02 TIMEBOOST_cell_10544 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_23__Q), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_1839) );
no02f10 TIMEBOOST_cell_44760 ( .a(TIMEBOOST_net_14618), .b(n_16290), .o(TIMEBOOST_net_10373) );
na02s01 TIMEBOOST_cell_36376 ( .a(TIMEBOOST_net_10426), .b(g65853_sb), .o(n_1567) );
in01f02 g54137_u0 ( .a(FE_OFN1148_n_13249), .o(g54137_sb) );
na02f02 g54137_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_384), .b(g54137_sb), .o(g54137_da) );
na02f02 g54137_u2 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__Q), .b(FE_OFN1148_n_13249), .o(g54137_db) );
na02f02 g54137_u3 ( .a(g54137_da), .b(g54137_db), .o(n_13273) );
in01f01 g54138_u0 ( .a(FE_OFN1149_n_13249), .o(g54138_sb) );
na02m02 TIMEBOOST_cell_10546 ( .a(FE_OFN1000_n_15978), .b(wishbone_slave_unit_del_sync_addr_out_reg_27__Q), .o(TIMEBOOST_net_1840) );
na02f02 TIMEBOOST_cell_39488 ( .a(TIMEBOOST_net_11982), .b(n_3237), .o(TIMEBOOST_net_510) );
na02f02 TIMEBOOST_cell_37974 ( .a(TIMEBOOST_net_11225), .b(FE_OFN1071_n_15729), .o(n_3084) );
na02f02 g54139_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_404), .b(FE_OCPN1910_FE_OFN1152_n_13249), .o(g54139_da) );
na03s02 TIMEBOOST_cell_38419 ( .a(n_3862), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q), .c(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_11448) );
no02f06 TIMEBOOST_cell_37170 ( .a(TIMEBOOST_net_10823), .b(FE_RN_678_0), .o(TIMEBOOST_net_128) );
in01m02 g54140_u0 ( .a(FE_OFN1150_n_13249), .o(g54140_sb) );
na02s01 TIMEBOOST_cell_39608 ( .a(TIMEBOOST_net_12042), .b(g62685_sb), .o(n_6168) );
na02s02 TIMEBOOST_cell_40397 ( .a(pci_target_unit_pcit_if_strd_addr_in_704), .b(g52633_sb), .o(TIMEBOOST_net_12437) );
na02s02 TIMEBOOST_cell_38064 ( .a(TIMEBOOST_net_11270), .b(FE_OFN1140_g64577_p), .o(TIMEBOOST_net_4610) );
in01m02 g54141_u0 ( .a(FE_OFN1151_n_13249), .o(g54141_sb) );
na02s01 TIMEBOOST_cell_43282 ( .a(TIMEBOOST_net_13879), .b(g62045_sb), .o(n_7767) );
na02s01 TIMEBOOST_cell_18438 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__Q), .b(g58369_sb), .o(TIMEBOOST_net_4476) );
na02s02 TIMEBOOST_cell_38656 ( .a(TIMEBOOST_net_11566), .b(g62655_sb), .o(n_6234) );
in01m01 g54143_u0 ( .a(FE_OCPN1911_FE_OFN1152_n_13249), .o(g54143_sb) );
na02f02 TIMEBOOST_cell_42410 ( .a(TIMEBOOST_net_13443), .b(g57541_sb), .o(n_10813) );
na02s02 TIMEBOOST_cell_43583 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__Q), .b(n_4306), .o(TIMEBOOST_net_14030) );
na02s02 TIMEBOOST_cell_43669 ( .a(TIMEBOOST_net_10004), .b(FE_OFN1333_n_13547), .o(TIMEBOOST_net_14073) );
in01f01 g54144_u0 ( .a(FE_OFN1147_n_13249), .o(g54144_sb) );
na03s02 TIMEBOOST_cell_38155 ( .a(TIMEBOOST_net_3553), .b(g64363_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__Q), .o(TIMEBOOST_net_11316) );
na02s01 TIMEBOOST_cell_40389 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__Q), .b(g65278_sb), .o(TIMEBOOST_net_12433) );
na02s01 TIMEBOOST_cell_36304 ( .a(TIMEBOOST_net_10390), .b(g67051_sb), .o(n_1495) );
in01m01 g54145_u0 ( .a(FE_OFN1149_n_13249), .o(g54145_sb) );
na02s02 TIMEBOOST_cell_10550 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_5__Q), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_1842) );
na03s02 TIMEBOOST_cell_40393 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__8__Q), .b(FE_OFN2256_n_8060), .c(n_1866), .o(TIMEBOOST_net_12435) );
na02f02 TIMEBOOST_cell_37134 ( .a(TIMEBOOST_net_10805), .b(n_12575), .o(n_12837) );
in01m01 g54146_u0 ( .a(FE_OFN1150_n_13249), .o(g54146_sb) );
na03s02 TIMEBOOST_cell_38373 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__Q), .b(FE_OFN1127_g64577_p), .c(g62744_sb), .o(TIMEBOOST_net_11425) );
na03s02 TIMEBOOST_cell_40395 ( .a(n_1855), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__Q), .c(FE_OFN716_n_8176), .o(TIMEBOOST_net_12436) );
na02f02 TIMEBOOST_cell_39096 ( .a(TIMEBOOST_net_11786), .b(FE_OFN1588_n_13736), .o(n_14260) );
in01m01 g54147_u0 ( .a(FE_OFN1149_n_13249), .o(g54147_sb) );
na02s01 TIMEBOOST_cell_10552 ( .a(wishbone_slave_unit_del_sync_bc_out_reg_1__Q), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_1843) );
na02f02 g54147_u2 ( .a(FE_OFN1150_n_13249), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__Q), .o(g54147_db) );
na02f02 TIMEBOOST_cell_37136 ( .a(n_16251), .b(TIMEBOOST_net_10806), .o(n_16254) );
in01f02 g54148_u0 ( .a(FE_OCPN1911_FE_OFN1152_n_13249), .o(g54148_sb) );
na02s02 TIMEBOOST_cell_45610 ( .a(TIMEBOOST_net_15043), .b(g65241_sb), .o(n_2641) );
na02f02 TIMEBOOST_cell_42412 ( .a(TIMEBOOST_net_13444), .b(g57284_sb), .o(n_11470) );
na02s02 TIMEBOOST_cell_45611 ( .a(TIMEBOOST_net_9365), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_15044) );
in01f01 g54149_u0 ( .a(FE_OFN1151_n_13249), .o(g54149_sb) );
na02s01 TIMEBOOST_cell_39305 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__Q), .b(g65836_sb), .o(TIMEBOOST_net_11891) );
na02s01 TIMEBOOST_cell_39492 ( .a(TIMEBOOST_net_11984), .b(g62756_sb), .o(n_6125) );
na02s02 TIMEBOOST_cell_43509 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__22__Q), .b(n_3525), .o(TIMEBOOST_net_13993) );
in01f02 g54150_u0 ( .a(FE_OFN1150_n_13249), .o(g54150_sb) );
na02f02 g54150_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_414), .b(g54150_sb), .o(g54150_da) );
na02f02 TIMEBOOST_cell_38653 ( .a(TIMEBOOST_net_626), .b(FE_OFN1189_n_5742), .o(TIMEBOOST_net_11565) );
na02s02 TIMEBOOST_cell_39454 ( .a(TIMEBOOST_net_11965), .b(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_4564) );
in01f02 g54151_u0 ( .a(FE_OCPN1911_FE_OFN1152_n_13249), .o(g54151_sb) );
na02s02 TIMEBOOST_cell_37993 ( .a(TIMEBOOST_net_9675), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_11235) );
na02f02 TIMEBOOST_cell_42414 ( .a(TIMEBOOST_net_13445), .b(g57379_sb), .o(n_11369) );
na02s02 TIMEBOOST_cell_45612 ( .a(TIMEBOOST_net_15044), .b(g65217_sb), .o(n_2670) );
in01f02 g54152_u0 ( .a(FE_OCPN1911_FE_OFN1152_n_13249), .o(g54152_sb) );
na02f02 g54152_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_387), .b(g54152_sb), .o(g54152_da) );
na02f02 TIMEBOOST_cell_38571 ( .a(FE_OFN1813_n_2919), .b(g54039_sb), .o(TIMEBOOST_net_11524) );
na02f02 TIMEBOOST_cell_42416 ( .a(TIMEBOOST_net_13446), .b(g57449_sb), .o(n_10348) );
in01f01 g54153_u0 ( .a(FE_OFN1148_n_13249), .o(g54153_sb) );
na02s02 TIMEBOOST_cell_10556 ( .a(pci_cbe_o_0_), .b(n_14389), .o(TIMEBOOST_net_1845) );
na02s01 TIMEBOOST_cell_18292 ( .a(g61880_sb), .b(g61979_db), .o(TIMEBOOST_net_4403) );
na02f02 TIMEBOOST_cell_12553 ( .a(n_16966), .b(TIMEBOOST_net_2843), .o(TIMEBOOST_net_650) );
in01f02 g54154_u0 ( .a(FE_OFN1148_n_13249), .o(g54154_sb) );
in01s01 TIMEBOOST_cell_45924 ( .a(TIMEBOOST_net_15230), .o(TIMEBOOST_net_15231) );
na02s02 TIMEBOOST_cell_38579 ( .a(TIMEBOOST_net_9907), .b(FE_OFN1180_n_3476), .o(TIMEBOOST_net_11528) );
na02s01 TIMEBOOST_cell_36306 ( .a(TIMEBOOST_net_10391), .b(g67040_sb), .o(n_1501) );
in01f02 g54155_u0 ( .a(FE_OFN1151_n_13249), .o(g54155_sb) );
na02f02 g54155_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_390), .b(g54155_sb), .o(g54155_da) );
na03s02 TIMEBOOST_cell_38111 ( .a(TIMEBOOST_net_4240), .b(g64218_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__Q), .o(TIMEBOOST_net_11294) );
na02m02 TIMEBOOST_cell_43837 ( .a(n_9111), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__Q), .o(TIMEBOOST_net_14157) );
in01f01 g54157_u0 ( .a(FE_OFN1151_n_13249), .o(g54157_sb) );
na02f02 g54157_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_392), .b(g54157_sb), .o(g54157_da) );
na02s02 TIMEBOOST_cell_38575 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .b(n_4658), .o(TIMEBOOST_net_11526) );
na02s01 TIMEBOOST_cell_38142 ( .a(TIMEBOOST_net_11309), .b(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_4519) );
in01m01 g54158_u0 ( .a(FE_OFN1147_n_13249), .o(g54158_sb) );
na02s02 TIMEBOOST_cell_45613 ( .a(TIMEBOOST_net_9358), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_15045) );
na02m02 TIMEBOOST_cell_18260 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_30__Q), .b(n_12595), .o(TIMEBOOST_net_4387) );
na02s02 TIMEBOOST_cell_45595 ( .a(TIMEBOOST_net_9363), .b(FE_OFN784_n_2678), .o(TIMEBOOST_net_15036) );
in01s01 g54159_u0 ( .a(n_13548), .o(n_13329) );
in01s03 g54160_u0 ( .a(wishbone_slave_unit_pci_initiator_if_data_source), .o(g54160_sb) );
na02s01 TIMEBOOST_cell_44907 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__Q), .b(n_2185), .o(TIMEBOOST_net_14692) );
na02s01 TIMEBOOST_cell_41747 ( .a(n_3777), .b(g64844_sb), .o(TIMEBOOST_net_13112) );
in01s01 g54161_u0 ( .a(FE_OFN1147_n_13249), .o(g54161_sb) );
na02s02 TIMEBOOST_cell_10562 ( .a(pci_cbe_o_1_), .b(n_14389), .o(TIMEBOOST_net_1848) );
na02s02 TIMEBOOST_cell_43610 ( .a(TIMEBOOST_net_14043), .b(FE_OFN1314_n_6624), .o(TIMEBOOST_net_12223) );
na02f02 TIMEBOOST_cell_44506 ( .a(TIMEBOOST_net_14491), .b(FE_OFN2168_n_8567), .o(TIMEBOOST_net_13452) );
in01s01 g54162_u0 ( .a(n_13544), .o(n_13328) );
na02s02 TIMEBOOST_cell_45137 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__Q), .b(n_3988), .o(TIMEBOOST_net_14807) );
na02s02 TIMEBOOST_cell_43058 ( .a(TIMEBOOST_net_13767), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_12079) );
na03s02 TIMEBOOST_cell_6699 ( .a(FE_OFN262_n_9851), .b(g58047_sb), .c(g58047_db), .o(n_9742) );
in01m01 g54164_u0 ( .a(FE_OFN1147_n_13249), .o(g54164_sb) );
na03s02 TIMEBOOST_cell_34255 ( .a(TIMEBOOST_net_9820), .b(FE_OFN1165_n_5615), .c(g62084_sb), .o(n_5625) );
na02s02 TIMEBOOST_cell_43611 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__Q), .b(n_3704), .o(TIMEBOOST_net_14044) );
na02s02 TIMEBOOST_cell_43059 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__Q), .b(n_4375), .o(TIMEBOOST_net_13768) );
in01s01 g54165_u0 ( .a(n_13541), .o(n_13327) );
na02s01 TIMEBOOST_cell_40283 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__Q), .b(n_8407), .o(TIMEBOOST_net_12380) );
na02s02 TIMEBOOST_cell_45614 ( .a(TIMEBOOST_net_15045), .b(g65214_sb), .o(n_2673) );
na02s02 TIMEBOOST_cell_39610 ( .a(TIMEBOOST_net_12043), .b(g62417_sb), .o(n_6763) );
in01s01 g54167_u0 ( .a(FE_OFN2119_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54167_sb) );
na02s01 TIMEBOOST_cell_42083 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__Q), .b(n_3515), .o(TIMEBOOST_net_13280) );
na03m04 TIMEBOOST_cell_32956 ( .a(n_539), .b(g58791_db), .c(g58791_sb), .o(n_9830) );
na02m02 TIMEBOOST_cell_18991 ( .a(TIMEBOOST_net_4752), .b(g54143_sb), .o(n_13361) );
in01s02 g54168_u0 ( .a(FE_OFN1083_n_13221), .o(g54168_sb) );
na02f02 TIMEBOOST_cell_42418 ( .a(TIMEBOOST_net_13447), .b(g57377_sb), .o(n_10378) );
na02f02 TIMEBOOST_cell_44250 ( .a(TIMEBOOST_net_14363), .b(FE_OFN1407_n_8567), .o(TIMEBOOST_net_12918) );
in01s02 g54169_u0 ( .a(FE_OFN1083_n_13221), .o(g54169_sb) );
na03s02 TIMEBOOST_cell_38135 ( .a(TIMEBOOST_net_4031), .b(g64235_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q), .o(TIMEBOOST_net_11306) );
na02m02 TIMEBOOST_cell_44325 ( .a(n_9460), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__Q), .o(TIMEBOOST_net_14401) );
na02s01 TIMEBOOST_cell_43670 ( .a(TIMEBOOST_net_14073), .b(g53912_sb), .o(n_13529) );
in01s02 g54170_u0 ( .a(FE_OFN1083_n_13221), .o(g54170_sb) );
na02s01 TIMEBOOST_cell_44908 ( .a(TIMEBOOST_net_14692), .b(FE_OFN699_n_7845), .o(TIMEBOOST_net_11058) );
na02s02 TIMEBOOST_cell_45615 ( .a(TIMEBOOST_net_9370), .b(FE_OFN787_n_2678), .o(TIMEBOOST_net_15046) );
na02f02 TIMEBOOST_cell_22523 ( .a(TIMEBOOST_net_6518), .b(FE_OFN1756_n_12681), .o(n_12496) );
in01s01 g54171_u0 ( .a(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54171_sb) );
na02f02 TIMEBOOST_cell_44160 ( .a(TIMEBOOST_net_14318), .b(FE_OFN1417_n_8567), .o(TIMEBOOST_net_12799) );
na02s01 TIMEBOOST_cell_41789 ( .a(n_4672), .b(g64991_db), .o(TIMEBOOST_net_13133) );
na02s01 TIMEBOOST_cell_43169 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__Q), .b(n_3546), .o(TIMEBOOST_net_13823) );
in01s01 g54172_u0 ( .a(FE_OFN1082_n_13221), .o(g54172_sb) );
na02m04 TIMEBOOST_cell_39019 ( .a(wbs_wbb3_2_wbb2_dat_o_i_126), .b(wbs_dat_o_27_), .o(TIMEBOOST_net_11748) );
na02s02 TIMEBOOST_cell_37834 ( .a(TIMEBOOST_net_11155), .b(g58450_sb), .o(n_9406) );
na02s01 TIMEBOOST_cell_39313 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__Q), .b(g65840_sb), .o(TIMEBOOST_net_11895) );
in01s01 g54173_u0 ( .a(FE_OFN1082_n_13221), .o(g54173_sb) );
na02m04 TIMEBOOST_cell_39041 ( .a(wbs_wbb3_2_wbb2_dat_o_i_112), .b(wbs_dat_o_13_), .o(TIMEBOOST_net_11759) );
na02s01 TIMEBOOST_cell_44860 ( .a(TIMEBOOST_net_14668), .b(g58434_sb), .o(TIMEBOOST_net_11934) );
na02m02 TIMEBOOST_cell_44353 ( .a(n_9604), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__Q), .o(TIMEBOOST_net_14415) );
in01s01 g54174_u0 ( .a(n_13221), .o(g54174_sb) );
na02s02 g54174_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_385), .b(g54174_sb), .o(g54174_da) );
na02s01 TIMEBOOST_cell_18302 ( .a(g61923_sb), .b(g61923_db), .o(TIMEBOOST_net_4408) );
no02f04 TIMEBOOST_cell_44776 ( .a(TIMEBOOST_net_14626), .b(FE_RN_628_0), .o(TIMEBOOST_net_151) );
in01s01 g54175_u0 ( .a(n_13221), .o(g54175_sb) );
na02s01 TIMEBOOST_cell_37692 ( .a(TIMEBOOST_net_11084), .b(g61706_sb), .o(n_8415) );
na02s01 g54175_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_12__Q), .b(n_13221), .o(g54175_db) );
na03s02 TIMEBOOST_cell_37693 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__Q), .b(FE_OFN710_n_8232), .c(n_1895), .o(TIMEBOOST_net_11085) );
in01s02 g54176_u0 ( .a(FE_OFN1085_n_13221), .o(g54176_sb) );
na02s06 g54176_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_396), .b(g54176_sb), .o(g54176_da) );
na02f02 TIMEBOOST_cell_42420 ( .a(TIMEBOOST_net_13448), .b(g57242_sb), .o(n_11516) );
na02s02 TIMEBOOST_cell_43558 ( .a(TIMEBOOST_net_14017), .b(FE_OFN1313_n_6624), .o(TIMEBOOST_net_12226) );
in01s02 g54177_u0 ( .a(FE_OFN1082_n_13221), .o(g54177_sb) );
na03f02 TIMEBOOST_cell_1988 ( .a(n_4199), .b(g52444_sb), .c(g52444_db), .o(n_14848) );
na02m02 TIMEBOOST_cell_32518 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__Q), .o(TIMEBOOST_net_10170) );
na02f02 TIMEBOOST_cell_43838 ( .a(TIMEBOOST_net_14157), .b(FE_OFN1381_n_8567), .o(TIMEBOOST_net_12845) );
in01s02 g54178_u0 ( .a(FE_OFN1082_n_13221), .o(g54178_sb) );
na02s01 TIMEBOOST_cell_44798 ( .a(TIMEBOOST_net_14637), .b(FE_OFN243_n_9116), .o(n_9082) );
na02s02 g54178_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_15__Q), .b(FE_OFN1084_n_13221), .o(g54178_db) );
na02s02 TIMEBOOST_cell_37948 ( .a(TIMEBOOST_net_11212), .b(g58244_sb), .o(n_9548) );
in01s02 g54179_u0 ( .a(FE_OFN1084_n_13221), .o(g54179_sb) );
na02s01 TIMEBOOST_cell_44799 ( .a(FE_OFN245_n_9114), .b(g58165_sb), .o(TIMEBOOST_net_14638) );
na02s01 TIMEBOOST_cell_43087 ( .a(n_4322), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__Q), .o(TIMEBOOST_net_13782) );
na02f02 TIMEBOOST_cell_22626 ( .a(FE_OFN2202_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__20__Q), .o(TIMEBOOST_net_6570) );
in01s01 g54180_u0 ( .a(n_13221), .o(g54180_sb) );
na02s01 g54180_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_400), .b(g54180_sb), .o(g54180_da) );
na02s02 TIMEBOOST_cell_36802 ( .a(TIMEBOOST_net_10639), .b(FE_OFN877_g64577_p), .o(TIMEBOOST_net_4571) );
na04f04 TIMEBOOST_cell_35282 ( .a(n_9216), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__Q), .c(FE_OFN1416_n_8567), .d(g57434_sb), .o(n_10821) );
in01s02 g54181_u0 ( .a(FE_OFN1084_n_13221), .o(g54181_sb) );
na02m02 g54181_u1 ( .a(g54181_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_401), .o(g54181_da) );
na02s01 TIMEBOOST_cell_45616 ( .a(TIMEBOOST_net_15046), .b(g65215_sb), .o(n_2672) );
in01s01 g54182_u0 ( .a(n_13221), .o(g54182_sb) );
na02s01 TIMEBOOST_cell_39612 ( .a(TIMEBOOST_net_12044), .b(g62608_sb), .o(n_6337) );
na02s01 g54182_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_19__Q), .b(n_13221), .o(g54182_db) );
na02s01 g64939_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__Q), .b(FE_OFN659_n_4392), .o(g64939_db) );
in01s01 g54183_u0 ( .a(FE_OFN1084_n_13221), .o(g54183_sb) );
na02m02 TIMEBOOST_cell_44311 ( .a(n_9470), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__Q), .o(TIMEBOOST_net_14394) );
na02m02 TIMEBOOST_cell_43839 ( .a(n_9734), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__Q), .o(TIMEBOOST_net_14158) );
in01s01 g54184_u0 ( .a(n_13221), .o(g54184_sb) );
na02f02 TIMEBOOST_cell_38789 ( .a(n_9691), .b(g57395_sb), .o(TIMEBOOST_net_11633) );
na02s01 g54184_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_21__Q), .b(n_13221), .o(g54184_db) );
na02s02 TIMEBOOST_cell_42368 ( .a(TIMEBOOST_net_13422), .b(g54363_sb), .o(n_13079) );
in01s01 g54185_u0 ( .a(n_13221), .o(g54185_sb) );
na02s02 g54185_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_386), .b(g54185_sb), .o(g54185_da) );
na02s01 TIMEBOOST_cell_18304 ( .a(g61880_sb), .b(g61971_db), .o(TIMEBOOST_net_4409) );
na02f02 TIMEBOOST_cell_43840 ( .a(TIMEBOOST_net_14158), .b(FE_OFN1387_n_8567), .o(TIMEBOOST_net_12891) );
in01s02 g54186_u0 ( .a(FE_OFN1084_n_13221), .o(g54186_sb) );
na02s01 TIMEBOOST_cell_44800 ( .a(TIMEBOOST_net_14638), .b(g58165_db), .o(n_9064) );
na02f02 TIMEBOOST_cell_41120 ( .a(TIMEBOOST_net_12798), .b(g57384_sb), .o(n_11361) );
na02s01 TIMEBOOST_cell_30967 ( .a(TIMEBOOST_net_9394), .b(g64929_db), .o(n_3679) );
in01s02 g54187_u0 ( .a(FE_OFN1085_n_13221), .o(g54187_sb) );
na03s02 TIMEBOOST_cell_37963 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__Q), .b(FE_OFN710_n_8232), .c(n_1889), .o(TIMEBOOST_net_11220) );
na02s01 TIMEBOOST_cell_43088 ( .a(TIMEBOOST_net_13782), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_12529) );
na02s01 TIMEBOOST_cell_43400 ( .a(TIMEBOOST_net_13938), .b(n_6319), .o(TIMEBOOST_net_11574) );
in01s01 g54188_u0 ( .a(n_13221), .o(g54188_sb) );
na02s02 TIMEBOOST_cell_39614 ( .a(TIMEBOOST_net_12045), .b(g62548_sb), .o(n_6470) );
na02s01 g54188_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_24__Q), .b(n_13221), .o(g54188_db) );
na02m02 TIMEBOOST_cell_43841 ( .a(n_9005), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__Q), .o(TIMEBOOST_net_14159) );
in01s01 g54189_u0 ( .a(n_13221), .o(g54189_sb) );
na02s01 TIMEBOOST_cell_38620 ( .a(TIMEBOOST_net_11548), .b(g63158_sb), .o(n_5822) );
na02s01 g54189_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_25__Q), .b(n_13221), .o(g54189_db) );
na02s03 TIMEBOOST_cell_45757 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__Q), .b(n_13184), .o(TIMEBOOST_net_15117) );
in01s02 g54190_u0 ( .a(FE_OFN1085_n_13221), .o(g54190_sb) );
na02s02 TIMEBOOST_cell_19129 ( .a(TIMEBOOST_net_4821), .b(g59096_sb), .o(TIMEBOOST_net_586) );
na02f02 TIMEBOOST_cell_42422 ( .a(TIMEBOOST_net_13449), .b(g57207_sb), .o(n_11549) );
na02f02 TIMEBOOST_cell_41520 ( .a(TIMEBOOST_net_12998), .b(FE_OFN2191_n_8567), .o(TIMEBOOST_net_11640) );
in01s02 g54191_u0 ( .a(FE_OFN1085_n_13221), .o(g54191_sb) );
na02m02 TIMEBOOST_cell_19127 ( .a(TIMEBOOST_net_4820), .b(g58843_sb), .o(TIMEBOOST_net_609) );
na02s02 TIMEBOOST_cell_45617 ( .a(TIMEBOOST_net_9343), .b(FE_OFN784_n_2678), .o(TIMEBOOST_net_15047) );
na02f02 TIMEBOOST_cell_41668 ( .a(TIMEBOOST_net_13072), .b(n_13621), .o(TIMEBOOST_net_11765) );
in01s02 g54192_u0 ( .a(FE_OFN1082_n_13221), .o(g54192_sb) );
na02s02 TIMEBOOST_cell_19125 ( .a(TIMEBOOST_net_4819), .b(g62067_sb), .o(TIMEBOOST_net_595) );
na02s02 TIMEBOOST_cell_41748 ( .a(TIMEBOOST_net_13112), .b(g64844_db), .o(n_3725) );
na02s02 TIMEBOOST_cell_45618 ( .a(TIMEBOOST_net_15047), .b(g65249_sb), .o(n_2633) );
in01s02 g54193_u0 ( .a(FE_OFN1084_n_13221), .o(g54193_sb) );
na02f02 TIMEBOOST_cell_37973 ( .a(configuration_wb_err_data_571), .b(n_2388), .o(TIMEBOOST_net_11225) );
na02s02 TIMEBOOST_cell_43089 ( .a(n_3791), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__Q), .o(TIMEBOOST_net_13783) );
na02f02 TIMEBOOST_cell_32573 ( .a(FE_OCPN1825_n_12030), .b(TIMEBOOST_net_10197), .o(TIMEBOOST_net_6564) );
in01s01 g54194_u0 ( .a(n_13221), .o(g54194_sb) );
na02f02 TIMEBOOST_cell_38924 ( .a(TIMEBOOST_net_11700), .b(g52596_sb), .o(TIMEBOOST_net_10703) );
na02s01 TIMEBOOST_cell_36378 ( .a(TIMEBOOST_net_10427), .b(g65865_db), .o(n_1708) );
na02s01 TIMEBOOST_cell_36380 ( .a(TIMEBOOST_net_10428), .b(g65853_db), .o(n_1583) );
in01s02 g54195_u0 ( .a(FE_OFN1082_n_13221), .o(g54195_sb) );
na02s01 TIMEBOOST_cell_44801 ( .a(FE_OFN245_n_9114), .b(g58224_sb), .o(TIMEBOOST_net_14639) );
na02m02 TIMEBOOST_cell_32516 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__Q), .o(TIMEBOOST_net_10169) );
na02m02 TIMEBOOST_cell_32572 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__Q), .o(TIMEBOOST_net_10197) );
in01m01 g54196_u0 ( .a(n_13221), .o(g54196_sb) );
na02s02 TIMEBOOST_cell_39616 ( .a(TIMEBOOST_net_12046), .b(g63168_sb), .o(n_5802) );
na02m01 g54196_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_4__Q), .b(n_13221), .o(g54196_db) );
na02s02 TIMEBOOST_cell_41723 ( .a(FE_OFN205_n_9140), .b(g57899_sb), .o(TIMEBOOST_net_13100) );
in01m02 g54197_u0 ( .a(FE_OFN1082_n_13221), .o(g54197_sb) );
na02s01 TIMEBOOST_cell_44802 ( .a(TIMEBOOST_net_14639), .b(g58224_db), .o(n_9049) );
na02s02 TIMEBOOST_cell_41749 ( .a(n_3747), .b(g65061_sb), .o(TIMEBOOST_net_13113) );
na02f02 TIMEBOOST_cell_41122 ( .a(TIMEBOOST_net_12799), .b(g57299_sb), .o(n_11452) );
in01m01 g54198_u0 ( .a(n_13221), .o(g54198_sb) );
no02f02 TIMEBOOST_cell_43671 ( .a(TIMEBOOST_net_2039), .b(FE_RN_371_0), .o(TIMEBOOST_net_14074) );
na02m01 g54198_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_6__Q), .b(n_13221), .o(g54198_db) );
na02s02 TIMEBOOST_cell_40446 ( .a(TIMEBOOST_net_12461), .b(g62088_sb), .o(TIMEBOOST_net_11378) );
in01s01 g54199_u0 ( .a(n_13221), .o(g54199_sb) );
na02f02 TIMEBOOST_cell_39099 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__Q), .o(TIMEBOOST_net_11788) );
na02s01 g54199_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_7__Q), .b(n_13221), .o(g54199_db) );
na02s02 TIMEBOOST_cell_41750 ( .a(TIMEBOOST_net_13113), .b(g65061_db), .o(n_3612) );
in01s01 g54200_u0 ( .a(FE_OFN1082_n_13221), .o(g54200_sb) );
na02f02 TIMEBOOST_cell_3889 ( .a(TIMEBOOST_net_524), .b(n_3229), .o(n_4786) );
na02s01 g54200_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_8__Q), .b(FE_OFN1082_n_13221), .o(g54200_db) );
na02s02 TIMEBOOST_cell_37825 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__Q), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_11151) );
in01s01 g54201_u0 ( .a(n_13221), .o(g54201_sb) );
na02s01 TIMEBOOST_cell_42740 ( .a(TIMEBOOST_net_13608), .b(FE_OFN710_n_8232), .o(TIMEBOOST_net_11065) );
na02s01 g54201_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_9__Q), .b(n_13221), .o(g54201_db) );
na02s01 TIMEBOOST_cell_18815 ( .a(TIMEBOOST_net_4664), .b(g63116_sb), .o(n_5023) );
in01s02 g54202_u0 ( .a(FE_OFN1084_n_13221), .o(g54202_sb) );
na02s02 g54202_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_393), .b(g54202_sb), .o(g54202_da) );
na02s02 TIMEBOOST_cell_43090 ( .a(TIMEBOOST_net_13783), .b(FE_OFN1222_n_6391), .o(TIMEBOOST_net_12573) );
na02s02 TIMEBOOST_cell_30933 ( .a(TIMEBOOST_net_9377), .b(g64794_sb), .o(n_3760) );
in01s01 g54203_u0 ( .a(n_13221), .o(g54203_sb) );
na02s02 TIMEBOOST_cell_38144 ( .a(TIMEBOOST_net_11310), .b(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_4534) );
na02s01 TIMEBOOST_cell_44909 ( .a(TIMEBOOST_net_9511), .b(FE_OFN1043_n_2037), .o(TIMEBOOST_net_14693) );
na02m02 TIMEBOOST_cell_41627 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_26__Q), .b(FE_OFN231_n_9839), .o(TIMEBOOST_net_13052) );
na02s02 TIMEBOOST_cell_43170 ( .a(TIMEBOOST_net_13823), .b(FE_OFN1285_n_4097), .o(TIMEBOOST_net_12136) );
na02s01 TIMEBOOST_cell_37277 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__Q), .b(FE_OFN517_n_9697), .o(TIMEBOOST_net_10877) );
in01s01 g54205_u0 ( .a(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54205_sb) );
na02f02 TIMEBOOST_cell_44686 ( .a(TIMEBOOST_net_14581), .b(g57540_sb), .o(n_11202) );
na02s04 TIMEBOOST_cell_45807 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_8__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_773), .o(TIMEBOOST_net_15142) );
na02s03 TIMEBOOST_cell_45770 ( .a(TIMEBOOST_net_15123), .b(FE_OFN1327_n_13547), .o(TIMEBOOST_net_14958) );
na02m02 TIMEBOOST_cell_44687 ( .a(n_9217), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__Q), .o(TIMEBOOST_net_14582) );
na02s02 TIMEBOOST_cell_43004 ( .a(TIMEBOOST_net_13740), .b(g58274_db), .o(n_9035) );
in01s01 g54207_u0 ( .a(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54207_sb) );
in01s01 TIMEBOOST_cell_45883 ( .a(n_8576), .o(TIMEBOOST_net_15190) );
na04s02 TIMEBOOST_cell_6754 ( .a(configuration_wb_err_data_580), .b(FE_OFN1169_n_5592), .c(parchk_pci_ad_out_in_1177), .d(g62080_sb), .o(n_5630) );
na02s01 TIMEBOOST_cell_37276 ( .a(TIMEBOOST_net_10876), .b(g64778_sb), .o(TIMEBOOST_net_223) );
na02s01 TIMEBOOST_cell_31043 ( .a(TIMEBOOST_net_9432), .b(g64932_db), .o(n_4387) );
na02s02 TIMEBOOST_cell_40376 ( .a(TIMEBOOST_net_12426), .b(g58353_db), .o(n_9468) );
in01s01 g54209_u0 ( .a(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54209_sb) );
na02s02 TIMEBOOST_cell_39618 ( .a(TIMEBOOST_net_12047), .b(g62452_sb), .o(n_6693) );
na02s01 TIMEBOOST_cell_41724 ( .a(TIMEBOOST_net_13100), .b(g57899_db), .o(n_9138) );
na03f02 TIMEBOOST_cell_22266 ( .a(n_16840), .b(n_10002), .c(n_10007), .o(TIMEBOOST_net_6390) );
na02s02 TIMEBOOST_cell_40378 ( .a(TIMEBOOST_net_12427), .b(FE_OFN233_n_9876), .o(TIMEBOOST_net_10045) );
na02f02 TIMEBOOST_cell_42522 ( .a(TIMEBOOST_net_13499), .b(g52600_sb), .o(TIMEBOOST_net_11764) );
na02f02 TIMEBOOST_cell_22267 ( .a(TIMEBOOST_net_6390), .b(n_16841), .o(n_12140) );
na02s02 TIMEBOOST_cell_39620 ( .a(TIMEBOOST_net_12048), .b(g62568_sb), .o(n_6420) );
na02m02 TIMEBOOST_cell_43521 ( .a(n_14743), .b(n_14839), .o(TIMEBOOST_net_13999) );
na03f02 TIMEBOOST_cell_22268 ( .a(n_16834), .b(n_10048), .c(n_16835), .o(TIMEBOOST_net_6391) );
na02s01 TIMEBOOST_cell_43140 ( .a(TIMEBOOST_net_13808), .b(FE_OFN1241_n_4092), .o(TIMEBOOST_net_12126) );
na02s01 TIMEBOOST_cell_42616 ( .a(TIMEBOOST_net_13546), .b(g58003_db), .o(n_9105) );
na02s01 TIMEBOOST_cell_37279 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__31__Q), .b(FE_OFN671_n_4505), .o(TIMEBOOST_net_10878) );
na02f02 TIMEBOOST_cell_42424 ( .a(TIMEBOOST_net_13450), .b(g57268_sb), .o(n_11484) );
na02s02 TIMEBOOST_cell_39622 ( .a(TIMEBOOST_net_12049), .b(g63157_sb), .o(n_5824) );
na02s01 TIMEBOOST_cell_37278 ( .a(TIMEBOOST_net_10877), .b(g58147_sb), .o(TIMEBOOST_net_370) );
na02s02 TIMEBOOST_cell_43171 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__Q), .b(n_3512), .o(TIMEBOOST_net_13824) );
na02f02 TIMEBOOST_cell_43842 ( .a(TIMEBOOST_net_14159), .b(FE_OFN1412_n_8567), .o(TIMEBOOST_net_12936) );
na02s02 TIMEBOOST_cell_43401 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__Q), .b(n_3595), .o(TIMEBOOST_net_13939) );
na02s01 TIMEBOOST_cell_45619 ( .a(n_4493), .b(g65002_sb), .o(TIMEBOOST_net_15048) );
na02s01 TIMEBOOST_cell_37281 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__Q), .b(FE_OFN670_n_4505), .o(TIMEBOOST_net_10879) );
in01s01 g54216_u0 ( .a(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54216_sb) );
na02s02 TIMEBOOST_cell_37280 ( .a(TIMEBOOST_net_10878), .b(g64787_sb), .o(TIMEBOOST_net_224) );
na02f02 TIMEBOOST_cell_42256 ( .a(TIMEBOOST_net_13366), .b(FE_OFN1425_n_8567), .o(TIMEBOOST_net_12325) );
na02s01 TIMEBOOST_cell_41751 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__Q), .b(g65883_sb), .o(TIMEBOOST_net_13114) );
na02f02 TIMEBOOST_cell_42426 ( .a(TIMEBOOST_net_13451), .b(g57573_sb), .o(n_11178) );
na02s02 TIMEBOOST_cell_43105 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__Q), .b(n_3772), .o(TIMEBOOST_net_13791) );
na02s03 TIMEBOOST_cell_45771 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__Q), .b(n_13177), .o(TIMEBOOST_net_15124) );
na02s01 TIMEBOOST_cell_43016 ( .a(TIMEBOOST_net_13746), .b(g62743_sb), .o(n_5493) );
na02f02 TIMEBOOST_cell_42257 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__Q), .b(n_9761), .o(TIMEBOOST_net_13367) );
na02s01 TIMEBOOST_cell_37283 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__Q), .b(FE_OFN516_n_9697), .o(TIMEBOOST_net_10880) );
in01s01 g54219_u0 ( .a(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54219_sb) );
na02s01 TIMEBOOST_cell_37282 ( .a(TIMEBOOST_net_10879), .b(g64773_sb), .o(TIMEBOOST_net_204) );
na02f02 TIMEBOOST_cell_42258 ( .a(TIMEBOOST_net_13367), .b(FE_OFN1384_n_8567), .o(TIMEBOOST_net_12295) );
na02s01 TIMEBOOST_cell_37285 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__Q), .b(FE_OFN670_n_4505), .o(TIMEBOOST_net_10881) );
na02f02 TIMEBOOST_cell_44296 ( .a(TIMEBOOST_net_14386), .b(FE_OFN1399_n_8567), .o(TIMEBOOST_net_12849) );
no02f02 TIMEBOOST_cell_43672 ( .a(TIMEBOOST_net_14074), .b(TIMEBOOST_net_944), .o(TIMEBOOST_net_3027) );
na02s01 TIMEBOOST_cell_31262 ( .a(pci_target_unit_fifos_pcir_data_in_187), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__Q), .o(TIMEBOOST_net_9542) );
na02s01 TIMEBOOST_cell_37284 ( .a(TIMEBOOST_net_10880), .b(g58153_sb), .o(TIMEBOOST_net_375) );
na02s01 TIMEBOOST_cell_42016 ( .a(TIMEBOOST_net_13246), .b(g62590_sb), .o(n_6372) );
na02s01 TIMEBOOST_cell_37287 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__Q), .b(n_3744), .o(TIMEBOOST_net_10882) );
na02s01 TIMEBOOST_cell_37286 ( .a(TIMEBOOST_net_10881), .b(g64775_sb), .o(TIMEBOOST_net_222) );
na02s02 TIMEBOOST_cell_45265 ( .a(n_4225), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__Q), .o(TIMEBOOST_net_14871) );
na03s02 TIMEBOOST_cell_33276 ( .a(FE_OFN227_n_9841), .b(g58183_sb), .c(g58183_db), .o(n_9604) );
na02s01 TIMEBOOST_cell_15872 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_97), .b(FE_OFN2119_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3193) );
na02f02 TIMEBOOST_cell_44220 ( .a(TIMEBOOST_net_14348), .b(FE_OFN1404_n_8567), .o(TIMEBOOST_net_13414) );
na02s02 TIMEBOOST_cell_31042 ( .a(n_4493), .b(g64932_sb), .o(TIMEBOOST_net_9432) );
na02s01 TIMEBOOST_cell_15873 ( .a(TIMEBOOST_net_3193), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_410), .o(TIMEBOOST_net_70) );
na02f02 TIMEBOOST_cell_37096 ( .a(TIMEBOOST_net_10786), .b(n_12584), .o(n_12846) );
na02s02 TIMEBOOST_cell_45138 ( .a(TIMEBOOST_net_14807), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_11410) );
na02s01 TIMEBOOST_cell_41752 ( .a(TIMEBOOST_net_13114), .b(g65883_db), .o(n_1575) );
na02m02 TIMEBOOST_cell_32490 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__Q), .o(TIMEBOOST_net_10156) );
na02f02 TIMEBOOST_cell_41681 ( .a(FE_OCP_RBN1996_n_13971), .b(TIMEBOOST_net_10227), .o(TIMEBOOST_net_13079) );
na02f02 g54940_u0 ( .a(n_12328), .b(n_12327), .o(n_12761) );
na02f02 TIMEBOOST_cell_41096 ( .a(TIMEBOOST_net_12786), .b(g57164_sb), .o(n_10838) );
na02s01 TIMEBOOST_cell_15864 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_86), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3189) );
na02f02 TIMEBOOST_cell_42276 ( .a(TIMEBOOST_net_13376), .b(g57063_sb), .o(n_10503) );
na02s02 TIMEBOOST_cell_38146 ( .a(TIMEBOOST_net_11311), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_4664) );
na02s01 TIMEBOOST_cell_43122 ( .a(TIMEBOOST_net_13799), .b(FE_OFN1196_n_4090), .o(TIMEBOOST_net_12092) );
na02s02 TIMEBOOST_cell_40448 ( .a(TIMEBOOST_net_12462), .b(g62082_sb), .o(TIMEBOOST_net_11377) );
na02s03 TIMEBOOST_cell_45772 ( .a(TIMEBOOST_net_15124), .b(FE_OFN1327_n_13547), .o(TIMEBOOST_net_14959) );
na02s02 TIMEBOOST_cell_41974 ( .a(TIMEBOOST_net_13225), .b(g62343_sb), .o(n_6913) );
na02s01 g54229_u2 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_76), .b(wishbone_slave_unit_pci_initiator_if_data_source), .o(g54229_db) );
na02s01 TIMEBOOST_cell_41899 ( .a(g62821_sb), .b(g62821_db), .o(TIMEBOOST_net_13188) );
na02f02 TIMEBOOST_cell_44688 ( .a(TIMEBOOST_net_14582), .b(FE_OFN1377_n_8567), .o(TIMEBOOST_net_13029) );
na02s01 TIMEBOOST_cell_41717 ( .a(FE_OFN205_n_9140), .b(g58262_sb), .o(TIMEBOOST_net_13097) );
na02s01 TIMEBOOST_cell_15843 ( .a(TIMEBOOST_net_3178), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_388), .o(TIMEBOOST_net_79) );
na03s02 TIMEBOOST_cell_33625 ( .a(TIMEBOOST_net_3671), .b(g65327_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__Q), .o(TIMEBOOST_net_4801) );
na02s01 TIMEBOOST_cell_41718 ( .a(TIMEBOOST_net_13097), .b(g58262_db), .o(n_9039) );
na02s01 TIMEBOOST_cell_37289 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__Q), .b(n_3739), .o(TIMEBOOST_net_10883) );
na02s02 TIMEBOOST_cell_42084 ( .a(TIMEBOOST_net_13280), .b(n_6287), .o(TIMEBOOST_net_11570) );
na02s02 TIMEBOOST_cell_41719 ( .a(n_3764), .b(g64783_sb), .o(TIMEBOOST_net_13098) );
na02s01 TIMEBOOST_cell_37288 ( .a(TIMEBOOST_net_10882), .b(FE_OFN662_n_4392), .o(TIMEBOOST_net_9385) );
na02s01 TIMEBOOST_cell_41917 ( .a(FE_OFN201_n_9230), .b(g57891_sb), .o(TIMEBOOST_net_13197) );
na02m02 TIMEBOOST_cell_44299 ( .a(n_9622), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__Q), .o(TIMEBOOST_net_14388) );
in01m02 g54234_u0 ( .a(FE_OFN1148_n_13249), .o(g54234_sb) );
na02s01 TIMEBOOST_cell_38658 ( .a(TIMEBOOST_net_11567), .b(g62435_sb), .o(n_6726) );
na02s02 TIMEBOOST_cell_43612 ( .a(TIMEBOOST_net_14044), .b(FE_OFN1313_n_6624), .o(TIMEBOOST_net_12246) );
na02s01 TIMEBOOST_cell_41725 ( .a(n_3744), .b(g64847_sb), .o(TIMEBOOST_net_13101) );
in01m01 g54235_u0 ( .a(FE_OFN1150_n_13249), .o(g54235_sb) );
na02f02 TIMEBOOST_cell_38926 ( .a(TIMEBOOST_net_11701), .b(n_9177), .o(n_9180) );
na02s02 TIMEBOOST_cell_44419 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_794), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_29__Q), .o(TIMEBOOST_net_14448) );
na02s02 TIMEBOOST_cell_38012 ( .a(TIMEBOOST_net_11244), .b(g61941_sb), .o(n_7941) );
in01m01 g54236_u0 ( .a(FE_OFN1151_n_13249), .o(g54236_sb) );
na02f02 TIMEBOOST_cell_39098 ( .a(TIMEBOOST_net_11787), .b(FE_OFN1588_n_13736), .o(n_14274) );
na02m02 TIMEBOOST_cell_44161 ( .a(n_9462), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q), .o(TIMEBOOST_net_14319) );
no02f02 TIMEBOOST_cell_37138 ( .a(TIMEBOOST_net_10807), .b(n_16233), .o(n_16234) );
in01f02 g54237_u0 ( .a(FE_OCPN1911_FE_OFN1152_n_13249), .o(g54237_sb) );
na02s02 TIMEBOOST_cell_45266 ( .a(TIMEBOOST_net_14871), .b(FE_OFN1223_n_6391), .o(TIMEBOOST_net_13242) );
na02f02 TIMEBOOST_cell_38569 ( .a(TIMEBOOST_net_4855), .b(n_3290), .o(TIMEBOOST_net_11523) );
na02s01 TIMEBOOST_cell_42945 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__Q), .b(FE_OFN584_n_9692), .o(TIMEBOOST_net_13711) );
in01f02 g54238_u0 ( .a(FE_OFN1149_n_13249), .o(g54238_sb) );
na02s01 TIMEBOOST_cell_18623 ( .a(TIMEBOOST_net_4568), .b(g63067_sb), .o(n_5116) );
na02f02 TIMEBOOST_cell_43782 ( .a(TIMEBOOST_net_14129), .b(FE_OFN1404_n_8567), .o(n_10411) );
na02f02 TIMEBOOST_cell_37098 ( .a(TIMEBOOST_net_10787), .b(n_12442), .o(n_12775) );
in01f01 g54239_u0 ( .a(FE_OFN1150_n_13249), .o(g54239_sb) );
na02s01 TIMEBOOST_cell_18054 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__Q), .b(g65367_sb), .o(TIMEBOOST_net_4284) );
na02s02 TIMEBOOST_cell_38014 ( .a(TIMEBOOST_net_11245), .b(g62024_sb), .o(n_7849) );
in01f01 g54244_u0 ( .a(FE_OFN1306_n_13124), .o(g54244_sb) );
na02m02 TIMEBOOST_cell_12614 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__Q), .o(TIMEBOOST_net_2874) );
na03f02 TIMEBOOST_cell_36153 ( .a(FE_OFN1583_n_12306), .b(TIMEBOOST_net_10256), .c(FE_OFN1762_n_10780), .o(n_12598) );
na03f04 TIMEBOOST_cell_37109 ( .a(n_10627), .b(n_10922), .c(n_10630), .o(TIMEBOOST_net_10793) );
na02f02 g54265_u0 ( .a(n_13410), .b(wbm_cti_o_0_), .o(n_13412) );
na02f02 g54266_u0 ( .a(n_13410), .b(wbm_cti_o_2_), .o(n_13411) );
no02f02 g54267_u0 ( .a(n_13486), .b(n_8757), .o(n_13624) );
na02f02 g54269_u0 ( .a(n_13317), .b(n_13068), .o(n_13409) );
na02f02 g54271_u0 ( .a(n_13315), .b(n_12963), .o(n_13407) );
na02f02 g54273_u0 ( .a(n_13314), .b(n_13063), .o(n_13406) );
na02f02 g54274_u0 ( .a(n_13313), .b(n_13066), .o(n_13405) );
na02f02 g54283_u0 ( .a(n_16413), .b(n_13056), .o(n_13404) );
na02f02 g54289_u0 ( .a(n_13311), .b(n_12958), .o(n_13403) );
na02f02 g54290_u0 ( .a(n_13310), .b(n_13052), .o(n_13402) );
oa12f02 g54294_u0 ( .a(n_13620), .b(n_13621), .c(pci_target_unit_fifos_pciw_outTransactionCount_1_), .o(n_13623) );
oa12f02 g54295_u0 ( .a(n_13620), .b(n_13621), .c(pci_target_unit_fifos_outGreyCount_0_), .o(n_13622) );
na02f02 g54297_u0 ( .a(n_13309), .b(n_13048), .o(n_13401) );
na02f02 g54298_u0 ( .a(n_13308), .b(n_13047), .o(n_13400) );
na02f02 g54303_u0 ( .a(n_16401), .b(n_13042), .o(n_13399) );
in01f02 g54304_u0 ( .a(FE_OFN2128_n_16497), .o(g54304_sb) );
na02s01 TIMEBOOST_cell_39177 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__Q), .b(FE_OFN577_n_9902), .o(TIMEBOOST_net_11827) );
na02s02 TIMEBOOST_cell_38595 ( .a(TIMEBOOST_net_9941), .b(FE_OFN1179_n_3476), .o(TIMEBOOST_net_11536) );
na02f02 g64457_u0 ( .a(n_3290), .b(pciu_bar0_in_376), .o(n_3287) );
in01f01 g54305_u0 ( .a(FE_OFN2128_n_16497), .o(g54305_sb) );
na02f02 g54305_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_782), .b(g54305_sb), .o(g54305_da) );
na02f02 g54305_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_17__Q), .b(FE_OFN2126_n_16497), .o(g54305_db) );
na02f02 g54305_u3 ( .a(g54305_da), .b(g54305_db), .o(n_13027) );
in01f01 g54306_u0 ( .a(FE_OFN2128_n_16497), .o(g54306_sb) );
na02f02 g54306_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_783), .b(g54306_sb), .o(g54306_da) );
na02f02 g54306_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_18__Q), .b(FE_OFN2128_n_16497), .o(g54306_db) );
na02f02 g54306_u3 ( .a(g54306_da), .b(g54306_db), .o(n_13026) );
ao12f02 g54308_u0 ( .a(n_13073), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_1__Q), .c(FE_OCPN1909_n_16497), .o(n_13127) );
in01f01 g54309_u0 ( .a(FE_OFN2128_n_16497), .o(g54309_sb) );
na02f02 g54309_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_785), .b(g54309_sb), .o(g54309_da) );
na02f02 g54309_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_20__Q), .b(FE_OFN2128_n_16497), .o(g54309_db) );
na02f02 g54309_u3 ( .a(g54309_da), .b(g54309_db), .o(n_13022) );
in01f01 g54310_u0 ( .a(FE_OFN2128_n_16497), .o(g54310_sb) );
na02f02 g54310_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_786), .b(g54310_sb), .o(g54310_da) );
na02f02 g54310_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_21__Q), .b(FE_OFN2128_n_16497), .o(g54310_db) );
na02f02 g54310_u3 ( .a(g54310_da), .b(g54310_db), .o(n_13020) );
in01m01 g54311_u0 ( .a(FE_OFN2126_n_16497), .o(g54311_sb) );
na02m02 g54311_u1 ( .a(g54311_sb), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_787), .o(g54311_da) );
na02f01 g54311_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_22__Q), .b(FE_OFN2126_n_16497), .o(g54311_db) );
na02f02 g54311_u3 ( .a(g54311_da), .b(g54311_db), .o(n_13018) );
in01m01 g54312_u0 ( .a(FE_OFN2127_n_16497), .o(g54312_sb) );
na02s02 g54312_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_788), .b(g54312_sb), .o(g54312_da) );
na02f01 g54312_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_23__Q), .b(FE_OFN2127_n_16497), .o(g54312_db) );
na02m02 TIMEBOOST_cell_38844 ( .a(TIMEBOOST_net_11660), .b(g58470_sb), .o(n_9377) );
in01f01 g54314_u0 ( .a(FE_OFN2126_n_16497), .o(g54314_sb) );
na02f02 g54314_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_790), .b(g54314_sb), .o(g54314_da) );
na02f01 g54314_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_25__Q), .b(FE_OFN2126_n_16497), .o(g54314_db) );
na02f02 g54314_u3 ( .a(g54314_da), .b(g54314_db), .o(n_13102) );
in01f01 g54315_u0 ( .a(FE_OFN2126_n_16497), .o(g54315_sb) );
na02f02 g54315_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_791), .b(g54315_sb), .o(g54315_da) );
na02f01 g54315_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_26__Q), .b(FE_OFN2125_n_16497), .o(g54315_db) );
na02f02 g54315_u3 ( .a(g54315_da), .b(g54315_db), .o(n_13012) );
in01f02 g54316_u0 ( .a(FE_OCPN1909_n_16497), .o(g54316_sb) );
na02s01 TIMEBOOST_cell_37214 ( .a(TIMEBOOST_net_10845), .b(FE_OFN2095_n_2520), .o(TIMEBOOST_net_9325) );
na02s02 TIMEBOOST_cell_17662 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__Q), .b(g65308_sb), .o(TIMEBOOST_net_4088) );
na02s02 TIMEBOOST_cell_38148 ( .a(TIMEBOOST_net_11312), .b(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_4552) );
in01f01 g54317_u0 ( .a(FE_OFN2127_n_16497), .o(g54317_sb) );
na02f02 g54317_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_793), .b(g54317_sb), .o(g54317_da) );
na02f02 g54317_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_28__Q), .b(FE_OFN2127_n_16497), .o(g54317_db) );
na02m02 TIMEBOOST_cell_38846 ( .a(TIMEBOOST_net_11661), .b(g58465_sb), .o(n_9385) );
in01f01 g54318_u0 ( .a(FE_OFN2127_n_16497), .o(g54318_sb) );
na02s02 TIMEBOOST_cell_44420 ( .a(TIMEBOOST_net_14448), .b(FE_OFN1306_n_13124), .o(TIMEBOOST_net_13424) );
na02f02 g54318_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_29__Q), .b(FE_OCPN1909_n_16497), .o(g54318_db) );
na02s01 TIMEBOOST_cell_22308 ( .a(g52477_da), .b(FE_OFN8_n_11877), .o(TIMEBOOST_net_6411) );
in01f02 g54319_u0 ( .a(FE_OCPN1909_n_16497), .o(g54319_sb) );
na02f02 g54319_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_767), .b(g54319_sb), .o(g54319_da) );
na02s02 TIMEBOOST_cell_39624 ( .a(TIMEBOOST_net_12050), .b(g62927_sb), .o(n_6027) );
na02f02 TIMEBOOST_cell_44326 ( .a(TIMEBOOST_net_14401), .b(FE_OFN1417_n_8567), .o(TIMEBOOST_net_12901) );
in01f02 g54320_u0 ( .a(FE_OCPN1909_n_16497), .o(g54320_sb) );
na02f02 g54320_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_795), .b(g54320_sb), .o(g54320_da) );
na02s01 TIMEBOOST_cell_39626 ( .a(TIMEBOOST_net_12051), .b(g62944_sb), .o(n_5993) );
na02s01 TIMEBOOST_cell_44910 ( .a(TIMEBOOST_net_14693), .b(g65826_sb), .o(TIMEBOOST_net_326) );
in01f01 g54321_u0 ( .a(FE_OCPN1909_n_16497), .o(g54321_sb) );
na02s01 TIMEBOOST_cell_44861 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__Q), .b(FE_OFN1657_n_9502), .o(TIMEBOOST_net_14669) );
na02m02 g54321_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_31__Q), .b(FE_OCPN1909_n_16497), .o(g54321_db) );
na02s02 TIMEBOOST_cell_19301 ( .a(TIMEBOOST_net_4907), .b(g60660_sb), .o(n_5660) );
in01f02 g54322_u0 ( .a(FE_OCPN1909_n_16497), .o(g54322_sb) );
na02f02 g54322_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_768), .b(g54322_sb), .o(g54322_da) );
na02f02 g54322_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_3__Q), .b(FE_OCPN1909_n_16497), .o(g54322_db) );
na02f02 g54322_u3 ( .a(g54322_da), .b(g54322_db), .o(n_12998) );
in01f01 g54323_u0 ( .a(FE_OFN2127_n_16497), .o(g54323_sb) );
na02f02 g54323_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_769), .b(g54323_sb), .o(g54323_da) );
na03s02 TIMEBOOST_cell_39437 ( .a(TIMEBOOST_net_3965), .b(g64337_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__Q), .o(TIMEBOOST_net_11957) );
na03m02 TIMEBOOST_cell_1453 ( .a(n_3425), .b(g52448_sb), .c(g52448_db), .o(n_14844) );
in01f02 g54324_u0 ( .a(FE_OCPN1909_n_16497), .o(g54324_sb) );
na02f02 g54324_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_770), .b(g54324_sb), .o(g54324_da) );
na02f02 g54324_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_5__Q), .b(FE_OCPN1909_n_16497), .o(g54324_db) );
na02f02 g54324_u3 ( .a(g54324_da), .b(g54324_db), .o(n_12994) );
in01f02 g54325_u0 ( .a(FE_OFN2125_n_16497), .o(g54325_sb) );
na02f02 g54325_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_771), .b(g54325_sb), .o(g54325_da) );
na02f02 g54325_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_6__Q), .b(FE_OFN2125_n_16497), .o(g54325_db) );
na02f02 g54325_u3 ( .a(g54325_da), .b(g54325_db), .o(n_12992) );
in01f02 g54326_u0 ( .a(FE_OFN2127_n_16497), .o(g54326_sb) );
na03s02 TIMEBOOST_cell_38415 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_), .b(FE_OFN1117_g64577_p), .c(n_2057), .o(TIMEBOOST_net_11446) );
na02s02 TIMEBOOST_cell_17664 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__31__Q), .b(g65412_sb), .o(TIMEBOOST_net_4089) );
na02s02 TIMEBOOST_cell_22309 ( .a(n_10170), .b(TIMEBOOST_net_6411), .o(n_11856) );
in01f02 g54328_u0 ( .a(FE_OFN2126_n_16497), .o(g54328_sb) );
na02f02 TIMEBOOST_cell_37097 ( .a(FE_RN_191_0), .b(n_10105), .o(TIMEBOOST_net_10787) );
na02s01 TIMEBOOST_cell_43054 ( .a(TIMEBOOST_net_13765), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_11541) );
na02s02 TIMEBOOST_cell_39349 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__12__Q), .b(g64308_sb), .o(TIMEBOOST_net_11913) );
no02f02 g54329_u0 ( .a(pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q), .b(n_13621), .o(g54329_p) );
ao12f01 g54329_u1 ( .a(g54329_p), .b(pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q), .c(n_13621), .o(n_13483) );
in01f01 g54330_u0 ( .a(FE_OCPN1909_n_16497), .o(g54330_sb) );
na02s01 TIMEBOOST_cell_45620 ( .a(TIMEBOOST_net_15048), .b(g65002_db), .o(n_4353) );
na02m02 g54330_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_0__Q), .b(FE_OCPN1909_n_16497), .o(g54330_db) );
na02s02 TIMEBOOST_cell_19303 ( .a(TIMEBOOST_net_4908), .b(g60607_sb), .o(n_4847) );
in01f01 g54331_u0 ( .a(FE_OFN2126_n_16497), .o(g54331_sb) );
na02f02 g54331_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_775), .b(g54331_sb), .o(g54331_da) );
na02f02 g54331_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_10__Q), .b(FE_OFN2126_n_16497), .o(g54331_db) );
na02f02 g54331_u3 ( .a(g54331_da), .b(g54331_db), .o(n_12985) );
in01f02 g54332_u0 ( .a(FE_OFN2128_n_16497), .o(g54332_sb) );
na03s02 TIMEBOOST_cell_38379 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__Q), .b(FE_OFN1132_g64577_p), .c(n_7217), .o(TIMEBOOST_net_11428) );
na02s01 TIMEBOOST_cell_18306 ( .a(g61880_sb), .b(g61975_db), .o(TIMEBOOST_net_4410) );
na02f02 TIMEBOOST_cell_38928 ( .a(TIMEBOOST_net_11702), .b(n_9177), .o(n_9179) );
in01f02 g54333_u0 ( .a(FE_OFN2128_n_16497), .o(g54333_sb) );
na02f02 TIMEBOOST_cell_18454 ( .a(n_3233), .b(n_4880), .o(TIMEBOOST_net_4484) );
na02s02 TIMEBOOST_cell_38720 ( .a(TIMEBOOST_net_11598), .b(g62484_sb), .o(n_6620) );
na02m02 TIMEBOOST_cell_18061 ( .a(TIMEBOOST_net_4287), .b(g54132_sb), .o(n_13467) );
in01f02 g54334_u0 ( .a(FE_OFN2128_n_16497), .o(g54334_sb) );
na02s02 TIMEBOOST_cell_45202 ( .a(TIMEBOOST_net_14839), .b(FE_OFN1260_n_4143), .o(TIMEBOOST_net_12103) );
na02s02 TIMEBOOST_cell_43613 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__Q), .b(n_3584), .o(TIMEBOOST_net_14045) );
na02s01 TIMEBOOST_cell_38542 ( .a(TIMEBOOST_net_11509), .b(g62061_sb), .o(n_7749) );
in01f02 g54335_u0 ( .a(FE_OFN2126_n_16497), .o(g54335_sb) );
na02s02 TIMEBOOST_cell_42741 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q), .b(g65394_sb), .o(TIMEBOOST_net_13609) );
na02s02 TIMEBOOST_cell_43614 ( .a(TIMEBOOST_net_14045), .b(FE_OFN1313_n_6624), .o(TIMEBOOST_net_12225) );
na02s01 TIMEBOOST_cell_38544 ( .a(TIMEBOOST_net_11510), .b(g62064_sb), .o(n_7745) );
in01f01 g54336_u0 ( .a(FE_OFN2128_n_16497), .o(g54336_sb) );
na02f02 g54336_u1 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_780), .b(g54336_sb), .o(g54336_da) );
na02f02 g54336_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_15__Q), .b(FE_OFN2128_n_16497), .o(g54336_db) );
na02f02 g54336_u3 ( .a(g54336_da), .b(g54336_db), .o(n_13098) );
in01f01 g54337_u0 ( .a(n_13621), .o(g54337_sb) );
na02s01 TIMEBOOST_cell_45621 ( .a(FE_OFN213_n_9124), .b(g58143_sb), .o(TIMEBOOST_net_15049) );
na02f02 TIMEBOOST_cell_22525 ( .a(FE_OFN1577_n_12028), .b(TIMEBOOST_net_6519), .o(n_12749) );
na02s02 TIMEBOOST_cell_43172 ( .a(TIMEBOOST_net_13824), .b(FE_OFN1260_n_4143), .o(TIMEBOOST_net_12060) );
in01m01 g54338_u0 ( .a(FE_OFN1305_n_13124), .o(g54338_sb) );
na02s01 TIMEBOOST_cell_18308 ( .a(g61885_sb), .b(g61980_db), .o(TIMEBOOST_net_4411) );
na02s01 TIMEBOOST_cell_36308 ( .a(TIMEBOOST_net_10392), .b(g67040_sb), .o(n_1649) );
na02f02 TIMEBOOST_cell_37119 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_10176), .o(TIMEBOOST_net_10798) );
in01s02 g54339_u0 ( .a(FE_OFN2136_n_13124), .o(g54339_sb) );
no02f04 TIMEBOOST_cell_12916 ( .a(FE_RN_806_0), .b(FE_RN_805_0), .o(TIMEBOOST_net_3025) );
na02f01 TIMEBOOST_cell_4077 ( .a(n_16444), .b(TIMEBOOST_net_618), .o(n_9154) );
na04f02 TIMEBOOST_cell_36167 ( .a(n_11078), .b(n_11075), .c(n_11076), .d(n_11077), .o(n_12540) );
in01m02 g54340_u0 ( .a(FE_OFN2134_n_13124), .o(g54340_sb) );
na02s01 TIMEBOOST_cell_17416 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__Q), .b(g64337_sb), .o(TIMEBOOST_net_3965) );
na03f02 TIMEBOOST_cell_36142 ( .a(FE_RN_194_0), .b(n_10731), .c(n_12583), .o(n_12845) );
na02s02 TIMEBOOST_cell_45267 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__Q), .b(n_4314), .o(TIMEBOOST_net_14872) );
in01s02 g54341_u0 ( .a(FE_OFN2134_n_13124), .o(g54341_sb) );
na02s02 TIMEBOOST_cell_39402 ( .a(TIMEBOOST_net_11939), .b(FE_OFN260_n_9860), .o(n_9783) );
na02m01 TIMEBOOST_cell_4081 ( .a(TIMEBOOST_net_620), .b(n_15517), .o(n_8853) );
na02s01 TIMEBOOST_cell_32012 ( .a(configuration_pci_err_data_514), .b(wbm_dat_o_13_), .o(TIMEBOOST_net_9917) );
in01m02 g54342_u0 ( .a(FE_OFN2134_n_13124), .o(g54342_sb) );
na02s01 TIMEBOOST_cell_18003 ( .a(TIMEBOOST_net_4258), .b(g64111_db), .o(n_4741) );
na02m01 TIMEBOOST_cell_4083 ( .a(n_9173), .b(TIMEBOOST_net_621), .o(n_8877) );
na02s01 TIMEBOOST_cell_42617 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__Q), .b(FE_OFN541_n_9690), .o(TIMEBOOST_net_13547) );
in01m02 g54343_u0 ( .a(FE_OFN2136_n_13124), .o(g54343_sb) );
na02f06 TIMEBOOST_cell_38481 ( .a(FE_OCPN1909_n_16497), .b(TIMEBOOST_net_4380), .o(TIMEBOOST_net_11479) );
na02m02 TIMEBOOST_cell_38848 ( .a(TIMEBOOST_net_11662), .b(g58841_sb), .o(n_8673) );
na02s01 TIMEBOOST_cell_45576 ( .a(TIMEBOOST_net_15026), .b(g64937_db), .o(n_4383) );
in01s02 g54344_u0 ( .a(FE_OFN2134_n_13124), .o(g54344_sb) );
na02s02 TIMEBOOST_cell_45740 ( .a(TIMEBOOST_net_15108), .b(FE_OFN709_n_8232), .o(TIMEBOOST_net_11092) );
na02m01 TIMEBOOST_cell_4087 ( .a(TIMEBOOST_net_623), .b(n_15515), .o(n_8852) );
na02s01 TIMEBOOST_cell_43113 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__23__Q), .b(n_3639), .o(TIMEBOOST_net_13795) );
in01m02 g54345_u0 ( .a(FE_OFN2134_n_13124), .o(g54345_sb) );
na02s01 TIMEBOOST_cell_18310 ( .a(g61923_sb), .b(g61985_db), .o(TIMEBOOST_net_4412) );
na02f06 TIMEBOOST_cell_4089 ( .a(TIMEBOOST_net_624), .b(n_16161), .o(n_16167) );
na02f03 TIMEBOOST_cell_4090 ( .a(n_1538), .b(n_7568), .o(TIMEBOOST_net_625) );
in01s02 g54346_u0 ( .a(FE_OFN2134_n_13124), .o(g54346_sb) );
na02s02 TIMEBOOST_cell_42968 ( .a(TIMEBOOST_net_13722), .b(g54198_db), .o(n_13420) );
na02f01 TIMEBOOST_cell_4113 ( .a(TIMEBOOST_net_636), .b(n_12858), .o(n_14693) );
na02s01 TIMEBOOST_cell_40511 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__Q), .b(wishbone_slave_unit_pcim_sm_data_in_636), .o(TIMEBOOST_net_12494) );
in01s02 g54347_u0 ( .a(FE_OFN2134_n_13124), .o(g54347_sb) );
na02s01 TIMEBOOST_cell_38445 ( .a(FE_OFN201_n_9230), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q), .o(TIMEBOOST_net_11461) );
na02f04 TIMEBOOST_cell_4091 ( .a(TIMEBOOST_net_625), .b(n_16459), .o(n_17031) );
na02f01 TIMEBOOST_cell_4092 ( .a(n_7399), .b(FE_OCPN1875_n_14526), .o(TIMEBOOST_net_626) );
in01s02 g54348_u0 ( .a(FE_OFN2135_n_13124), .o(g54348_sb) );
na02s02 TIMEBOOST_cell_18090 ( .a(n_1953), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__Q), .o(TIMEBOOST_net_4302) );
na02s01 TIMEBOOST_cell_36375 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__Q), .b(g65918_db), .o(TIMEBOOST_net_10426) );
in01s01 TIMEBOOST_cell_32825 ( .a(TIMEBOOST_net_10326), .o(TIMEBOOST_net_10325) );
in01m01 g54349_u0 ( .a(FE_OFN1306_n_13124), .o(g54349_sb) );
na03s02 TIMEBOOST_cell_36755 ( .a(g64131_da), .b(g64131_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__Q), .o(TIMEBOOST_net_10616) );
na02m02 TIMEBOOST_cell_12884 ( .a(FE_OFN9_n_11877), .b(FE_RN_122_0), .o(TIMEBOOST_net_3009) );
na02f02 TIMEBOOST_cell_37105 ( .a(FE_RN_101_0), .b(n_11717), .o(TIMEBOOST_net_10791) );
in01s02 g54350_u0 ( .a(FE_OFN2134_n_13124), .o(g54350_sb) );
na02s02 TIMEBOOST_cell_41924 ( .a(TIMEBOOST_net_13200), .b(g58413_db), .o(n_9204) );
na02f08 TIMEBOOST_cell_4095 ( .a(TIMEBOOST_net_627), .b(n_8801), .o(n_9177) );
na02f02 TIMEBOOST_cell_44302 ( .a(TIMEBOOST_net_14389), .b(FE_OFN1391_n_8567), .o(TIMEBOOST_net_12730) );
in01s02 g54351_u0 ( .a(FE_OFN2134_n_13124), .o(g54351_sb) );
in01s01 TIMEBOOST_cell_45877 ( .a(n_8576), .o(TIMEBOOST_net_15184) );
no02f02 TIMEBOOST_cell_36892 ( .a(TIMEBOOST_net_10684), .b(FE_RN_565_0), .o(TIMEBOOST_net_664) );
na02s02 TIMEBOOST_cell_38582 ( .a(TIMEBOOST_net_11529), .b(g60666_sb), .o(n_5652) );
in01s02 g54352_u0 ( .a(FE_OFN2135_n_13124), .o(g54352_sb) );
na03s02 TIMEBOOST_cell_38367 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__Q), .b(FE_OFN1129_g64577_p), .c(n_3831), .o(TIMEBOOST_net_11422) );
na02s02 TIMEBOOST_cell_20113 ( .a(TIMEBOOST_net_5313), .b(n_13625), .o(TIMEBOOST_net_610) );
na03f02 TIMEBOOST_cell_4100 ( .a(n_2830), .b(n_3232), .c(n_2857), .o(TIMEBOOST_net_630) );
in01m01 g54353_u0 ( .a(FE_OFN1305_n_13124), .o(g54353_sb) );
na02m02 TIMEBOOST_cell_12618 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__13__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__13__Q), .o(TIMEBOOST_net_2876) );
na02s01 TIMEBOOST_cell_38660 ( .a(TIMEBOOST_net_11568), .b(g62370_sb), .o(n_6863) );
na02s01 TIMEBOOST_cell_37694 ( .a(TIMEBOOST_net_11085), .b(g61876_sb), .o(n_8079) );
in01m01 g54354_u0 ( .a(FE_OFN1305_n_13124), .o(g54354_sb) );
na02m02 TIMEBOOST_cell_12620 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__16__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__16__Q), .o(TIMEBOOST_net_2877) );
na02s01 TIMEBOOST_cell_45139 ( .a(n_852), .b(pci_target_unit_fifos_inGreyCount_reg_1__Q), .o(TIMEBOOST_net_14808) );
na03s02 TIMEBOOST_cell_33271 ( .a(FE_OFN227_n_9841), .b(g58244_sb), .c(g58245_db), .o(n_9547) );
in01s02 g54355_u0 ( .a(FE_OFN2136_n_13124), .o(g54355_sb) );
na02s01 TIMEBOOST_cell_36391 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(g65802_sb), .o(TIMEBOOST_net_10434) );
na02f02 TIMEBOOST_cell_4101 ( .a(TIMEBOOST_net_630), .b(n_3424), .o(n_5643) );
in01s01 TIMEBOOST_cell_45953 ( .a(wbm_dat_i_5_), .o(TIMEBOOST_net_15260) );
in01s02 g54356_u0 ( .a(FE_OFN2136_n_13124), .o(g54356_sb) );
na02s02 TIMEBOOST_cell_42969 ( .a(TIMEBOOST_net_4370), .b(g54196_sb), .o(TIMEBOOST_net_13723) );
na02s02 TIMEBOOST_cell_39628 ( .a(TIMEBOOST_net_12052), .b(g62522_sb), .o(n_6532) );
na02s01 TIMEBOOST_cell_9199 ( .a(TIMEBOOST_net_1166), .b(g65774_db), .o(n_2193) );
in01m01 g54357_u0 ( .a(FE_OFN1306_n_13124), .o(g54357_sb) );
na02m02 TIMEBOOST_cell_41631 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_4__Q), .b(FE_OFN243_n_9116), .o(TIMEBOOST_net_13054) );
no02f02 TIMEBOOST_cell_39179 ( .a(FE_RN_609_0), .b(FE_RN_621_0), .o(TIMEBOOST_net_11828) );
na02s02 TIMEBOOST_cell_43515 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__Q), .b(n_4316), .o(TIMEBOOST_net_13996) );
in01m01 g54358_u0 ( .a(FE_OFN1305_n_13124), .o(g54358_sb) );
na02s02 TIMEBOOST_cell_37930 ( .a(TIMEBOOST_net_11203), .b(g58441_sb), .o(n_9410) );
na02m02 TIMEBOOST_cell_44211 ( .a(n_9848), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__Q), .o(TIMEBOOST_net_14344) );
na02f06 TIMEBOOST_cell_4038 ( .a(n_7398), .b(n_16914), .o(TIMEBOOST_net_599) );
in01m01 g54359_u0 ( .a(FE_OFN1306_n_13124), .o(g54359_sb) );
na02f06 TIMEBOOST_cell_4039 ( .a(TIMEBOOST_net_599), .b(n_15442), .o(n_16438) );
na04f02 TIMEBOOST_cell_36169 ( .a(n_10788), .b(n_11124), .c(n_11123), .d(n_11122), .o(n_12551) );
na02s02 TIMEBOOST_cell_16802 ( .a(n_3770), .b(g65025_sb), .o(TIMEBOOST_net_3658) );
in01f01 g54360_u0 ( .a(FE_OFN1306_n_13124), .o(g54360_sb) );
na03f02 TIMEBOOST_cell_36909 ( .a(n_3044), .b(n_2824), .c(n_2614), .o(TIMEBOOST_net_10693) );
na03f02 TIMEBOOST_cell_36181 ( .a(FE_OFN1733_n_16317), .b(TIMEBOOST_net_10291), .c(FE_OFN1738_n_11019), .o(n_12634) );
na02s02 TIMEBOOST_cell_4042 ( .a(n_4743), .b(n_2742), .o(TIMEBOOST_net_601) );
in01m01 g54361_u0 ( .a(FE_OFN1306_n_13124), .o(g54361_sb) );
na02m04 TIMEBOOST_cell_4043 ( .a(TIMEBOOST_net_601), .b(n_7110), .o(n_8465) );
na02s01 TIMEBOOST_cell_36310 ( .a(TIMEBOOST_net_10393), .b(g67040_sb), .o(n_1641) );
na02s01 TIMEBOOST_cell_4044 ( .a(n_4743), .b(n_2308), .o(TIMEBOOST_net_602) );
in01m01 g54362_u0 ( .a(FE_OFN1305_n_13124), .o(g54362_sb) );
na02m02 TIMEBOOST_cell_4045 ( .a(TIMEBOOST_net_602), .b(n_7110), .o(n_8512) );
na02s01 TIMEBOOST_cell_36312 ( .a(TIMEBOOST_net_10394), .b(g67051_sb), .o(n_1503) );
na02s02 TIMEBOOST_cell_4046 ( .a(n_13745), .b(n_15405), .o(TIMEBOOST_net_603) );
in01m01 g54363_u0 ( .a(FE_OFN1306_n_13124), .o(g54363_sb) );
na02f04 g53828_u0 ( .a(n_13452), .b(n_2120), .o(n_13661) );
na02s01 TIMEBOOST_cell_36314 ( .a(TIMEBOOST_net_10395), .b(g65870_db), .o(n_2300) );
na02s01 TIMEBOOST_cell_42834 ( .a(TIMEBOOST_net_13655), .b(g65351_db), .o(n_4257) );
in01m01 g54364_u0 ( .a(FE_OFN1305_n_13124), .o(g54364_sb) );
na02m02 TIMEBOOST_cell_4049 ( .a(n_13625), .b(TIMEBOOST_net_604), .o(n_13821) );
na02s01 TIMEBOOST_cell_44803 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(g65779_sb), .o(TIMEBOOST_net_14640) );
na02s01 TIMEBOOST_cell_4050 ( .a(n_7530), .b(n_7044), .o(TIMEBOOST_net_605) );
in01m01 g54365_u0 ( .a(FE_OFN1306_n_13124), .o(g54365_sb) );
na02f02 TIMEBOOST_cell_4051 ( .a(TIMEBOOST_net_605), .b(n_13625), .o(n_13810) );
na02s01 TIMEBOOST_cell_36316 ( .a(TIMEBOOST_net_10396), .b(g65861_db), .o(n_2183) );
no02f04 TIMEBOOST_cell_4052 ( .a(FE_RN_284_0), .b(FE_RN_285_0), .o(TIMEBOOST_net_606) );
in01m01 g54366_u0 ( .a(FE_OFN1305_n_13124), .o(g54366_sb) );
no02f04 TIMEBOOST_cell_4053 ( .a(TIMEBOOST_net_606), .b(g59129_p), .o(n_7094) );
na02s02 TIMEBOOST_cell_45729 ( .a(n_3762), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__Q), .o(TIMEBOOST_net_15103) );
na02s02 TIMEBOOST_cell_39630 ( .a(TIMEBOOST_net_12053), .b(g62573_sb), .o(n_6407) );
in01f01 g54367_u0 ( .a(FE_OFN1305_n_13124), .o(g54367_sb) );
na02s01 TIMEBOOST_cell_18723 ( .a(TIMEBOOST_net_4618), .b(g62854_sb), .o(n_5260) );
no02f02 TIMEBOOST_cell_12908 ( .a(FE_RN_817_0), .b(FE_RN_818_0), .o(TIMEBOOST_net_3021) );
na02s02 TIMEBOOST_cell_37900 ( .a(TIMEBOOST_net_11188), .b(g58272_sb), .o(n_9529) );
in01s02 g54368_u0 ( .a(FE_OFN2135_n_13124), .o(g54368_sb) );
na02s01 TIMEBOOST_cell_38016 ( .a(TIMEBOOST_net_11246), .b(g62023_sb), .o(n_7851) );
na02s01 TIMEBOOST_cell_36500 ( .a(TIMEBOOST_net_10488), .b(g66415_sb), .o(n_2505) );
na02f02 TIMEBOOST_cell_41296 ( .a(TIMEBOOST_net_12886), .b(g57121_sb), .o(n_10476) );
in01m02 g54369_u0 ( .a(FE_OFN2135_n_13124), .o(g54369_sb) );
na03s02 TIMEBOOST_cell_38427 ( .a(n_3907), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__16__Q), .c(FE_OFN2106_g64577_p), .o(TIMEBOOST_net_11452) );
na02f04 TIMEBOOST_cell_22363 ( .a(TIMEBOOST_net_6438), .b(n_12441), .o(n_12774) );
na02f06 TIMEBOOST_cell_4108 ( .a(FE_RN_500_0), .b(n_7712), .o(TIMEBOOST_net_634) );
no02f02 g54408_u0 ( .a(n_13041), .b(n_12759), .o(n_13317) );
no02f02 g54410_u0 ( .a(n_17028), .b(n_17029), .o(n_13315) );
no02f02 g54411_u0 ( .a(n_16600), .b(n_16601), .o(n_13314) );
no02f02 g54412_u0 ( .a(n_16602), .b(n_16603), .o(n_13313) );
no02f02 g54414_u0 ( .a(n_15440), .b(n_15441), .o(n_13311) );
no02f02 g54415_u0 ( .a(n_16589), .b(n_16588), .o(n_13310) );
no02f02 g54416_u0 ( .a(n_15438), .b(n_15439), .o(n_13309) );
no02f02 g54417_u0 ( .a(n_16591), .b(n_16592), .o(n_13308) );
na02f04 g54419_u0 ( .a(n_998), .b(n_13621), .o(n_13620) );
na02f02 g54420_u0 ( .a(FE_OFN2163_n_16301), .b(wbm_dat_o_0_), .o(n_13398) );
na02f02 g54422_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_11_), .o(n_13395) );
na02f02 g54423_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_12_), .o(n_13394) );
na02f02 g54424_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_13_), .o(n_13393) );
na02f02 g54425_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_14_), .o(n_13392) );
na02f02 g54426_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_15_), .o(n_13391) );
na02f02 g54427_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_16_), .o(n_13390) );
na02f02 g54428_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_17_), .o(n_13389) );
na02f02 g54429_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_18_), .o(n_13388) );
na02f02 g54430_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_19_), .o(n_13387) );
na02f02 g54431_u0 ( .a(FE_OFN2163_n_16301), .b(wbm_dat_o_1_), .o(n_13386) );
na02f02 g54432_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_20_), .o(n_13384) );
na02f02 g54433_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_21_), .o(n_13383) );
na02f02 g54435_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_23_), .o(n_13381) );
na02f02 g54436_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_24_), .o(n_13380) );
na02f02 g54437_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_25_), .o(n_13379) );
na02f02 g54438_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_26_), .o(n_13378) );
na02f02 g54439_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_27_), .o(n_13377) );
na02f02 g54440_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_28_), .o(n_13376) );
na02f02 g54441_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_29_), .o(n_13375) );
na02f02 g54442_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_2_), .o(n_13374) );
na02f02 g54443_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_30_), .o(n_13373) );
na02f02 g54444_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_31_), .o(n_13372) );
na02f02 g54445_u0 ( .a(FE_OFN2163_n_16301), .b(wbm_dat_o_3_), .o(n_13371) );
na02f02 g54446_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_4_), .o(n_13370) );
na02f02 g54447_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_5_), .o(n_13369) );
na02f02 g54448_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_6_), .o(n_13368) );
na02f02 g54449_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_7_), .o(n_13367) );
na02f02 g54450_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_8_), .o(n_13366) );
na02f02 g54451_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_9_), .o(n_13365) );
no02f02 g54452_u0 ( .a(n_12952), .b(FE_OCPN1909_n_16497), .o(n_13073) );
na02f01 g54453_u0 ( .a(n_16495), .b(pci_target_unit_pcit_if_pcir_fifo_control_in_637), .o(g54453_p) );
in01f02 g54453_u1 ( .a(g54453_p), .o(n_13145) );
in01f03 g54454_u0 ( .a(n_13410), .o(n_14518) );
no02f02 g54456_u0 ( .a(n_16299), .b(n_13122), .o(g54456_p) );
in01f02 g54456_u1 ( .a(g54456_p), .o(n_14898) );
no02f08 g54457_u0 ( .a(FE_OFN1705_n_4868), .b(n_13721), .o(n_13754) );
na02f02 g54458_u0 ( .a(n_16299), .b(n_12956), .o(g54458_p) );
in01f04 g54458_u1 ( .a(g54458_p), .o(n_13486) );
no02f02 g54459_u0 ( .a(n_13304), .b(pci_target_unit_del_sync_be_out_reg_0__Q), .o(n_13306) );
na02f02 g54460_u0 ( .a(n_14967), .b(n_13122), .o(n_14895) );
no02f02 g54461_u0 ( .a(n_13304), .b(pci_target_unit_del_sync_be_out_reg_1__Q), .o(n_13305) );
no02f02 g54462_u0 ( .a(n_13304), .b(pci_target_unit_del_sync_be_out_reg_2__Q), .o(n_13303) );
no02f02 g54463_u0 ( .a(n_13304), .b(pci_target_unit_del_sync_be_out_reg_3__Q), .o(n_13302) );
no02m02 g54464_u0 ( .a(FE_OFN969_n_13784), .b(n_12595), .o(n_13415) );
na02s02 g54465_u0 ( .a(n_12776), .b(n_12595), .o(g54465_p) );
in01s02 g54465_u1 ( .a(g54465_p), .o(n_13341) );
no02f02 g54466_u0 ( .a(FE_OFN2165_n_16301), .b(n_8757), .o(n_13481) );
na02f02 TIMEBOOST_cell_42428 ( .a(TIMEBOOST_net_13452), .b(g57522_sb), .o(n_11219) );
in01s01 g54468_u0 ( .a(n_12855), .o(n_12954) );
no02s01 g54470_u0 ( .a(n_13721), .b(n_14905), .o(n_12855) );
in01f01 g54471_u0 ( .a(n_13617), .o(g54471_sb) );
in01s01 TIMEBOOST_cell_32824 ( .a(TIMEBOOST_net_10325), .o(n_1064) );
na02f02 TIMEBOOST_cell_22527 ( .a(FE_OFN1577_n_12028), .b(TIMEBOOST_net_6520), .o(n_12631) );
in01f01 g54472_u0 ( .a(n_13617), .o(g54472_sb) );
in01s02 TIMEBOOST_cell_32823 ( .a(TIMEBOOST_net_10323), .o(TIMEBOOST_net_10324) );
na02s02 TIMEBOOST_cell_45268 ( .a(TIMEBOOST_net_14872), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_12117) );
na02f02 TIMEBOOST_cell_44566 ( .a(TIMEBOOST_net_14521), .b(FE_OFN2167_n_8567), .o(TIMEBOOST_net_13469) );
in01f01 g54474_u0 ( .a(n_16967), .o(n_13479) );
in01f01 g54480_u0 ( .a(n_16205), .o(n_13475) );
in01f01 g54484_u0 ( .a(n_13617), .o(g54484_sb) );
na02m02 TIMEBOOST_cell_32562 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__Q), .o(TIMEBOOST_net_10192) );
na02s02 TIMEBOOST_cell_31065 ( .a(TIMEBOOST_net_9443), .b(g64996_db), .o(n_4355) );
na02s01 TIMEBOOST_cell_43674 ( .a(TIMEBOOST_net_14075), .b(g58634_db), .o(n_8846) );
in01f01 g54485_u0 ( .a(n_13617), .o(g54485_sb) );
na03s01 TIMEBOOST_cell_34800 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__Q), .b(g63199_sb), .c(g63199_db), .o(n_5766) );
na02s02 TIMEBOOST_cell_45269 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__Q), .b(n_4311), .o(TIMEBOOST_net_14873) );
na02s02 TIMEBOOST_cell_43173 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__Q), .b(n_3674), .o(TIMEBOOST_net_13825) );
in01f02 g54486_u0 ( .a(n_13617), .o(g54486_sb) );
na02f02 TIMEBOOST_cell_21829 ( .a(TIMEBOOST_net_6171), .b(n_8582), .o(n_8583) );
na02s02 TIMEBOOST_cell_45270 ( .a(TIMEBOOST_net_14873), .b(FE_OFN1285_n_4097), .o(TIMEBOOST_net_12071) );
in01f01 g54487_u0 ( .a(n_13617), .o(g54487_sb) );
na02f02 TIMEBOOST_cell_41124 ( .a(TIMEBOOST_net_12800), .b(g57223_sb), .o(n_10436) );
na02m02 TIMEBOOST_cell_43747 ( .a(n_9703), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__Q), .o(TIMEBOOST_net_14112) );
na02s02 TIMEBOOST_cell_45271 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__Q), .b(n_4368), .o(TIMEBOOST_net_14874) );
in01f01 g54488_u0 ( .a(n_13617), .o(g54488_sb) );
na02m02 TIMEBOOST_cell_32448 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__Q), .o(TIMEBOOST_net_10135) );
na02s01 TIMEBOOST_cell_30816 ( .a(n_3744), .b(g64813_sb), .o(TIMEBOOST_net_9319) );
na02s02 TIMEBOOST_cell_45022 ( .a(TIMEBOOST_net_14749), .b(FE_OFN2021_n_4778), .o(TIMEBOOST_net_13741) );
in01f01 g54489_u0 ( .a(n_13617), .o(g54489_sb) );
in01s02 TIMEBOOST_cell_32822 ( .a(parchk_pci_cbe_en_in), .o(TIMEBOOST_net_10323) );
na02f02 TIMEBOOST_cell_22537 ( .a(TIMEBOOST_net_6525), .b(FE_OFN1577_n_12028), .o(n_12659) );
na02s01 TIMEBOOST_cell_30822 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__Q), .o(TIMEBOOST_net_9322) );
in01f01 g54490_u0 ( .a(n_13617), .o(g54490_sb) );
na02m02 TIMEBOOST_cell_32530 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__Q), .o(TIMEBOOST_net_10176) );
na02f02 TIMEBOOST_cell_44354 ( .a(TIMEBOOST_net_14415), .b(FE_OFN1424_n_8567), .o(TIMEBOOST_net_12923) );
na02s02 TIMEBOOST_cell_45272 ( .a(TIMEBOOST_net_14874), .b(FE_OFN1293_n_4098), .o(TIMEBOOST_net_12125) );
in01f01 g54491_u0 ( .a(n_13617), .o(g54491_sb) );
na02s02 TIMEBOOST_cell_41771 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__Q), .b(g58279_sb), .o(TIMEBOOST_net_13124) );
na02s01 TIMEBOOST_cell_45023 ( .a(TIMEBOOST_net_4205), .b(g61964_db), .o(TIMEBOOST_net_14750) );
na02s02 TIMEBOOST_cell_44415 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_770), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_5__Q), .o(TIMEBOOST_net_14446) );
in01f01 g54492_u0 ( .a(n_13617), .o(g54492_sb) );
na02s02 TIMEBOOST_cell_41772 ( .a(TIMEBOOST_net_13124), .b(g58279_db), .o(n_9523) );
na02s01 TIMEBOOST_cell_43283 ( .a(TIMEBOOST_net_4769), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_13880) );
na02f02 TIMEBOOST_cell_22541 ( .a(TIMEBOOST_net_6527), .b(FE_OFN1577_n_12028), .o(n_12603) );
in01f01 g54493_u0 ( .a(n_13617), .o(g54493_sb) );
na02f02 TIMEBOOST_cell_41126 ( .a(TIMEBOOST_net_12801), .b(g57250_sb), .o(n_11507) );
na02f02 TIMEBOOST_cell_43772 ( .a(TIMEBOOST_net_14124), .b(FE_OFN1414_n_8567), .o(TIMEBOOST_net_12930) );
na02s01 TIMEBOOST_cell_43284 ( .a(TIMEBOOST_net_13880), .b(g62034_sb), .o(n_7782) );
in01f01 g54494_u0 ( .a(n_13617), .o(g54494_sb) );
na02f02 TIMEBOOST_cell_41206 ( .a(TIMEBOOST_net_12841), .b(g57453_sb), .o(n_11281) );
na02s01 TIMEBOOST_cell_45024 ( .a(TIMEBOOST_net_14750), .b(FE_OFN2021_n_4778), .o(TIMEBOOST_net_13657) );
na02f02 TIMEBOOST_cell_22543 ( .a(TIMEBOOST_net_6528), .b(FE_OFN1736_n_16317), .o(n_12487) );
in01f01 g54495_u0 ( .a(n_13617), .o(g54495_sb) );
na02m02 TIMEBOOST_cell_32590 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q), .o(TIMEBOOST_net_10206) );
na02s02 TIMEBOOST_cell_43174 ( .a(TIMEBOOST_net_13825), .b(FE_OFN1242_n_4092), .o(TIMEBOOST_net_12075) );
na02s02 TIMEBOOST_cell_45273 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__Q), .b(n_4446), .o(TIMEBOOST_net_14875) );
oa12f01 g54496_u0 ( .a(n_13474), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q), .c(n_13617), .o(n_13682) );
in01s02 g54504_u0 ( .a(n_13784), .o(n_13721) );
in01s02 g54510_u0 ( .a(n_12776), .o(n_13763) );
in01s01 g54511_u0 ( .a(n_12776), .o(n_13781) );
in01m06 g54512_u0 ( .a(FE_OFN969_n_13784), .o(n_12776) );
in01s01 g54519_u0 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_766), .o(n_12952) );
na02f02 g54549_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q), .b(n_13617), .o(n_13474) );
no02f02 g54567_u0 ( .a(n_12819), .b(n_12764), .o(n_12964) );
na02f02 g54568_u0 ( .a(n_12756), .b(n_12946), .o(g54568_p) );
in01f02 g54568_u1 ( .a(g54568_p), .o(n_13068) );
na02f02 g54569_u0 ( .a(n_12943), .b(n_12528), .o(g54569_p) );
in01f02 g54569_u1 ( .a(g54569_p), .o(n_13067) );
no02f02 g54570_u0 ( .a(n_12806), .b(n_12818), .o(n_12963) );
no02f02 g54571_u0 ( .a(n_12817), .b(n_12741), .o(n_12962) );
na02f02 g54572_u0 ( .a(n_12936), .b(n_12736), .o(g54572_p) );
in01f02 g54572_u1 ( .a(g54572_p), .o(n_13063) );
na02f02 g54573_u0 ( .a(n_12933), .b(n_12731), .o(g54573_p) );
in01f02 g54573_u1 ( .a(g54573_p), .o(n_13066) );
na02f02 g54574_u0 ( .a(n_12930), .b(n_12725), .o(g54574_p) );
in01f02 g54574_u1 ( .a(g54574_p), .o(n_13065) );
in01f02 g54575_u0 ( .a(n_13064), .o(n_13120) );
na02f02 g54576_u0 ( .a(n_12927), .b(n_12519), .o(n_13064) );
na02f02 g54579_u0 ( .a(n_12921), .b(n_12709), .o(g54579_p) );
in01f02 g54579_u1 ( .a(g54579_p), .o(n_13059) );
na02f02 g54580_u0 ( .a(n_12919), .b(n_12705), .o(g54580_p) );
in01f02 g54580_u1 ( .a(g54580_p), .o(n_13061) );
na02f02 g54581_u0 ( .a(n_12916), .b(n_12699), .o(g54581_p) );
in01f02 g54581_u1 ( .a(g54581_p), .o(n_13060) );
in01f02 g54582_u0 ( .a(n_12961), .o(n_13058) );
na02f02 g54583_u0 ( .a(n_12693), .b(n_12815), .o(n_12961) );
in01f02 g54584_u0 ( .a(n_13057), .o(n_13118) );
na02f02 g54585_u0 ( .a(n_12688), .b(n_12911), .o(n_13057) );
na02f02 g54586_u0 ( .a(n_12908), .b(n_12682), .o(g54586_p) );
in01f02 g54586_u1 ( .a(g54586_p), .o(n_13056) );
na02f02 g54587_u0 ( .a(n_12905), .b(n_12503), .o(g54587_p) );
in01f02 g54587_u1 ( .a(g54587_p), .o(n_13055) );
no02f02 g54588_u0 ( .a(n_12813), .b(n_12676), .o(n_12960) );
no02f02 g54589_u0 ( .a(n_12901), .b(n_12672), .o(n_13054) );
no02f02 g54590_u0 ( .a(n_12898), .b(n_12667), .o(n_13053) );
na02f02 g54591_u0 ( .a(n_12812), .b(n_12662), .o(g54591_p) );
in01f02 g54591_u1 ( .a(g54591_p), .o(n_12959) );
no02f02 g54592_u0 ( .a(n_12811), .b(n_12788), .o(n_12958) );
na02f02 g54593_u0 ( .a(n_12891), .b(n_12495), .o(g54593_p) );
in01f02 g54593_u1 ( .a(g54593_p), .o(n_13052) );
na02f02 g54594_u0 ( .a(n_12888), .b(n_12647), .o(g54594_p) );
in01f02 g54594_u1 ( .a(g54594_p), .o(n_13051) );
na02f02 g54595_u0 ( .a(n_12885), .b(n_12642), .o(g54595_p) );
in01f02 g54595_u1 ( .a(g54595_p), .o(n_13050) );
na02f02 g54596_u0 ( .a(n_12882), .b(n_12636), .o(g54596_p) );
in01f02 g54596_u1 ( .a(g54596_p), .o(n_13049) );
na02f02 g54597_u0 ( .a(n_13116), .b(pci_target_unit_wbm_sm_pciw_fifo_control_in), .o(g54597_p) );
in01f04 g54597_u1 ( .a(g54597_p), .o(n_13621) );
no02f02 g54598_u0 ( .a(n_12810), .b(n_12784), .o(n_12957) );
no02f02 g54599_u0 ( .a(n_12783), .b(n_12877), .o(n_13048) );
no02f02 g54600_u0 ( .a(n_12874), .b(n_12623), .o(n_13047) );
na02f02 g54601_u0 ( .a(n_12871), .b(n_12619), .o(g54601_p) );
in01f02 g54601_u1 ( .a(g54601_p), .o(n_13046) );
no02f02 g54602_u0 ( .a(n_12868), .b(n_12614), .o(n_13045) );
na02f02 g54603_u0 ( .a(n_12865), .b(n_12484), .o(g54603_p) );
in01f02 g54603_u1 ( .a(g54603_p), .o(n_13044) );
in01f02 g54604_u0 ( .a(n_13043), .o(n_13117) );
na02f02 g54605_u0 ( .a(n_12602), .b(n_12862), .o(n_13043) );
na02f02 g54606_u0 ( .a(n_12859), .b(n_12480), .o(g54606_p) );
in01f02 g54606_u1 ( .a(g54606_p), .o(n_13042) );
in01f08 g54610_u0 ( .a(n_13363), .o(n_14725) );
in01f06 g54616_u0 ( .a(n_13363), .o(n_14800) );
na02s01 TIMEBOOST_cell_45622 ( .a(TIMEBOOST_net_15049), .b(g58143_db), .o(n_9069) );
na02f02 TIMEBOOST_cell_41586 ( .a(TIMEBOOST_net_13031), .b(FE_OFN1440_n_9372), .o(TIMEBOOST_net_11651) );
in01f02 g54665_u0 ( .a(n_13122), .o(n_13304) );
in01f02 g54666_u0 ( .a(n_12956), .o(n_13122) );
na02f02 TIMEBOOST_cell_42268 ( .a(TIMEBOOST_net_13372), .b(FE_OFN1382_n_8567), .o(TIMEBOOST_net_12306) );
oa12f02 g54669_u0 ( .a(n_8727), .b(n_8730), .c(n_10825), .o(n_12170) );
na02f02 g54670_u0 ( .a(n_12947), .b(n_12948), .o(n_13041) );
na02f02 g54672_u0 ( .a(n_12941), .b(n_12942), .o(n_17028) );
na02f02 g54673_u0 ( .a(n_12938), .b(n_12937), .o(n_16600) );
na02f02 g54674_u0 ( .a(n_12934), .b(n_12935), .o(n_16602) );
no02f02 g54677_u0 ( .a(n_12814), .b(n_12904), .o(n_13034) );
na02f02 g54678_u0 ( .a(n_12894), .b(n_12895), .o(n_15440) );
na02f02 g54679_u0 ( .a(n_12892), .b(n_12893), .o(n_16588) );
na02f02 g54680_u0 ( .a(n_12878), .b(n_12879), .o(n_15438) );
na02f02 g54681_u0 ( .a(n_12875), .b(n_12876), .o(n_16591) );
no02f02 g54716_u0 ( .a(n_12166), .b(n_11014), .o(n_12591) );
no02f02 g54717_u0 ( .a(n_12165), .b(n_11741), .o(n_12590) );
no02f03 g54718_u0 ( .a(n_12164), .b(n_11740), .o(n_12589) );
no02f02 g54719_u0 ( .a(n_12163), .b(n_10987), .o(n_12588) );
no02f02 g54720_u0 ( .a(n_12162), .b(n_10764), .o(n_12587) );
no02f02 g54721_u0 ( .a(n_12161), .b(n_10978), .o(n_12586) );
no02f02 g54722_u0 ( .a(n_12160), .b(n_10976), .o(n_12585) );
no02f02 g54723_u0 ( .a(n_12159), .b(n_10975), .o(n_12584) );
no02f02 g54724_u0 ( .a(n_12158), .b(n_10971), .o(n_12583) );
no02f02 g54726_u0 ( .a(n_12156), .b(n_10963), .o(n_12581) );
no02f02 g54727_u0 ( .a(n_10962), .b(n_12155), .o(n_12580) );
no02f02 g54728_u0 ( .a(n_12154), .b(n_10952), .o(n_12579) );
no02f02 g54729_u0 ( .a(n_11847), .b(n_11738), .o(n_12442) );
no02f02 g54730_u0 ( .a(n_12153), .b(n_10943), .o(n_12578) );
no02f02 g54731_u0 ( .a(n_17042), .b(n_17041), .o(n_12577) );
no02f04 g54733_u0 ( .a(n_11846), .b(n_10932), .o(n_12441) );
no02f02 g54734_u0 ( .a(n_12439), .b(n_11736), .o(n_12772) );
no02f02 g54735_u0 ( .a(n_12148), .b(n_10923), .o(n_12575) );
no02f02 g54736_u0 ( .a(n_12147), .b(n_10638), .o(n_12574) );
no02f02 g54737_u0 ( .a(n_12146), .b(n_10631), .o(n_12573) );
no02f02 g54738_u0 ( .a(n_12145), .b(n_10919), .o(n_12572) );
no02f03 g54739_u0 ( .a(n_11845), .b(n_10917), .o(n_12440) );
no02f02 g54740_u0 ( .a(n_12144), .b(n_10913), .o(n_12571) );
no02f02 g54741_u0 ( .a(n_11734), .b(n_12143), .o(n_12570) );
no02f02 g54742_u0 ( .a(n_12141), .b(n_10906), .o(n_12569) );
no02f02 g54743_u0 ( .a(n_12140), .b(n_11731), .o(n_12568) );
no02f02 g54744_u0 ( .a(n_12139), .b(n_11727), .o(n_12567) );
no02f02 g54745_u0 ( .a(n_12137), .b(n_11880), .o(n_12566) );
no02f02 g54746_u0 ( .a(n_12135), .b(n_11724), .o(n_12565) );
no02f03 g54747_u0 ( .a(n_12134), .b(n_10882), .o(n_12564) );
no02f02 g54748_u0 ( .a(n_12133), .b(n_10876), .o(n_12563) );
no02f02 g54749_u0 ( .a(n_12132), .b(n_10867), .o(n_12562) );
no02f02 g54750_u0 ( .a(n_11718), .b(n_12130), .o(n_12561) );
no02f03 g54751_u0 ( .a(n_12129), .b(n_10860), .o(n_12560) );
no02f02 g54752_u0 ( .a(n_12128), .b(n_10856), .o(n_12559) );
no02f02 g54754_u0 ( .a(n_12767), .b(n_12768), .o(n_12950) );
no02f02 g54755_u0 ( .a(n_12765), .b(n_12766), .o(n_12949) );
no02f02 g54757_u0 ( .a(n_12762), .b(n_12763), .o(n_12948) );
no02f02 g54758_u0 ( .a(n_12761), .b(n_12760), .o(n_12947) );
no02f02 g54759_u0 ( .a(n_12757), .b(n_12758), .o(n_12946) );
no02f02 g54762_u0 ( .a(n_12750), .b(n_12751), .o(n_12943) );
no02f02 g54763_u0 ( .a(n_12748), .b(n_12749), .o(n_12942) );
no02f02 g54764_u0 ( .a(n_12747), .b(n_12746), .o(n_12941) );
no02f02 g54766_u0 ( .a(n_12744), .b(n_12745), .o(n_12940) );
no02f02 g54767_u0 ( .a(n_12742), .b(n_12743), .o(n_12939) );
no02f02 g54769_u0 ( .a(n_17036), .b(n_17035), .o(n_12938) );
no02f02 g54770_u0 ( .a(n_12738), .b(n_12527), .o(n_12937) );
no02f02 g54771_u0 ( .a(n_12526), .b(n_12737), .o(n_12936) );
no02f02 g54772_u0 ( .a(n_12734), .b(n_12735), .o(n_12935) );
no02f02 g54773_u0 ( .a(n_12733), .b(n_12525), .o(n_12934) );
no02f02 g54774_u0 ( .a(n_12524), .b(n_12732), .o(n_12933) );
no02f02 g54775_u0 ( .a(n_12729), .b(n_12523), .o(n_12932) );
no02f02 g54776_u0 ( .a(n_12728), .b(n_12727), .o(n_12931) );
no02f02 g54777_u0 ( .a(n_12522), .b(n_12726), .o(n_12930) );
no02f02 g54778_u0 ( .a(n_12723), .b(n_12724), .o(n_12929) );
no02f02 g54779_u0 ( .a(n_12521), .b(n_12722), .o(n_12928) );
no02f02 g54780_u0 ( .a(n_12520), .b(n_12720), .o(n_12927) );
no02f02 g54783_u0 ( .a(n_12715), .b(n_12518), .o(n_12924) );
no02f02 g54784_u0 ( .a(n_12517), .b(n_12713), .o(n_12923) );
no02f02 g54785_u0 ( .a(n_12712), .b(n_12711), .o(n_12922) );
no02f02 g54786_u0 ( .a(n_12516), .b(n_12710), .o(n_12921) );
no02f02 g54789_u0 ( .a(n_12515), .b(n_12706), .o(n_12919) );
no02f02 g54790_u0 ( .a(n_12703), .b(n_12704), .o(n_12918) );
no02f02 g54791_u0 ( .a(n_12702), .b(n_12701), .o(n_12917) );
no02f02 g54792_u0 ( .a(n_12514), .b(n_12700), .o(n_12916) );
no02f02 g54793_u0 ( .a(n_12513), .b(n_12697), .o(n_12915) );
no02f02 g54794_u0 ( .a(n_12696), .b(n_12512), .o(n_12914) );
no02f02 g54795_u0 ( .a(n_12510), .b(n_12511), .o(n_12815) );
no02f02 g54796_u0 ( .a(n_12509), .b(n_12692), .o(n_12913) );
no02f02 g54798_u0 ( .a(n_12689), .b(n_12508), .o(n_12911) );
no02f02 g54801_u0 ( .a(n_12684), .b(n_12683), .o(n_12908) );
no02f02 g54802_u0 ( .a(n_12506), .b(n_12680), .o(n_12907) );
no02f02 g54803_u0 ( .a(n_12505), .b(n_12679), .o(n_12906) );
no02f02 g54804_u0 ( .a(n_12678), .b(n_12504), .o(n_12905) );
na02m02 TIMEBOOST_cell_41942 ( .a(TIMEBOOST_net_13209), .b(TIMEBOOST_net_9880), .o(n_13499) );
no02f02 g54808_u0 ( .a(n_12500), .b(n_12675), .o(n_12903) );
no02f02 g54809_u0 ( .a(n_12673), .b(n_12674), .o(n_12902) );
na04f04 g54810_u0 ( .a(n_12116), .b(n_12243), .c(n_12244), .d(n_12372), .o(n_12901) );
no02f02 g54811_u0 ( .a(n_12671), .b(n_12670), .o(n_12900) );
no02f02 g54812_u0 ( .a(n_12669), .b(n_12668), .o(n_12899) );
na04f04 g54813_u0 ( .a(n_12238), .b(n_12237), .c(n_12369), .d(n_12115), .o(n_12898) );
no02f02 g54814_u0 ( .a(n_12665), .b(n_12666), .o(n_12897) );
no02f02 g54815_u0 ( .a(n_12664), .b(n_12663), .o(n_12896) );
no02f02 g54816_u0 ( .a(n_12499), .b(n_12498), .o(n_12812) );
no02f02 g54817_u0 ( .a(n_12661), .b(n_12660), .o(n_12895) );
no02f02 g54818_u0 ( .a(n_12658), .b(n_12659), .o(n_12894) );
na04f04 g54819_u0 ( .a(n_11937), .b(n_11814), .c(n_11938), .d(n_12075), .o(n_12811) );
no02f02 g54820_u0 ( .a(n_12656), .b(n_12655), .o(n_12893) );
no02f02 g54821_u0 ( .a(n_12653), .b(n_12654), .o(n_12892) );
no02f02 g54822_u0 ( .a(n_12652), .b(n_12496), .o(n_12891) );
no02f02 g54823_u0 ( .a(n_12494), .b(n_12651), .o(n_12890) );
no02f02 g54824_u0 ( .a(n_12649), .b(n_12650), .o(n_12889) );
no02f02 g54825_u0 ( .a(n_12493), .b(n_12648), .o(n_12888) );
no02f02 g54826_u0 ( .a(n_12646), .b(n_12492), .o(n_12887) );
no02f02 g54827_u0 ( .a(n_12645), .b(n_12644), .o(n_12886) );
no02f02 g54828_u0 ( .a(n_12491), .b(n_12643), .o(n_12885) );
no02f02 g54829_u0 ( .a(n_12640), .b(n_12641), .o(n_12884) );
no02f02 g54830_u0 ( .a(n_12638), .b(n_12639), .o(n_12883) );
no02f02 g54831_u0 ( .a(n_12637), .b(n_12490), .o(n_12882) );
no02f02 g54832_u0 ( .a(n_15759), .b(FE_OFN186_n_15768), .o(n_11450) );
in01f02 TIMEBOOST_cell_32821 ( .a(TIMEBOOST_net_10322), .o(TIMEBOOST_net_10321) );
in01f06 g54834_u0 ( .a(n_13116), .o(n_13617) );
in01m06 g54838_u0 ( .a(n_16981), .o(n_13116) );
no02f02 g54840_u0 ( .a(n_12489), .b(n_12635), .o(n_12881) );
no02f02 g54841_u0 ( .a(n_12633), .b(n_12634), .o(n_12880) );
no02f02 g54843_u0 ( .a(n_12630), .b(n_12631), .o(n_12879) );
no02f02 g54844_u0 ( .a(n_12628), .b(n_12629), .o(n_12878) );
no02f02 g54846_u0 ( .a(n_12625), .b(n_12626), .o(n_12876) );
no02f02 g54847_u0 ( .a(n_12624), .b(n_12488), .o(n_12875) );
no02f02 g54849_u0 ( .a(n_12622), .b(n_12487), .o(n_12873) );
no02f02 g54850_u0 ( .a(n_12486), .b(n_12621), .o(n_12872) );
no02f02 g54851_u0 ( .a(n_12485), .b(n_12620), .o(n_12871) );
no02f02 g54852_u0 ( .a(n_12618), .b(n_12617), .o(n_12870) );
no02f02 g54853_u0 ( .a(n_12616), .b(n_12615), .o(n_12869) );
no02f02 g54855_u0 ( .a(n_12612), .b(n_12613), .o(n_12867) );
no02f02 g54856_u0 ( .a(n_12610), .b(n_12611), .o(n_12866) );
no02f02 g54857_u0 ( .a(n_16597), .b(n_16596), .o(n_12865) );
no02f02 g54858_u0 ( .a(n_12606), .b(n_12607), .o(n_12864) );
no02f02 g54859_u0 ( .a(n_12604), .b(n_12605), .o(n_12863) );
no02f02 g54860_u0 ( .a(n_12483), .b(n_12603), .o(n_12862) );
no02f02 g54863_u0 ( .a(n_12481), .b(n_12596), .o(n_12859) );
in01f02 g54864_u0 ( .a(n_12167), .o(n_12168) );
in01f02 g54865_u0 ( .a(n_15611), .o(n_12167) );
na04f04 g54868_u0 ( .a(n_11796), .b(n_11153), .c(n_11147), .d(n_11155), .o(n_12557) );
na02s01 TIMEBOOST_cell_43175 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__Q), .b(n_4249), .o(TIMEBOOST_net_13826) );
na04f04 g54870_u0 ( .a(n_11142), .b(n_11143), .c(n_11146), .d(n_11145), .o(n_12555) );
na04f04 g54872_u0 ( .a(n_11135), .b(n_11134), .c(n_11131), .d(n_11132), .o(n_12553) );
na02m02 TIMEBOOST_cell_44355 ( .a(n_9092), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__Q), .o(TIMEBOOST_net_14416) );
na04f04 g54877_u0 ( .a(n_16583), .b(n_11115), .c(n_11113), .d(n_16584), .o(n_12549) );
na04f04 g54878_u0 ( .a(n_11111), .b(n_11110), .c(n_11108), .d(n_11109), .o(n_12548) );
na04f04 g54883_u0 ( .a(n_11086), .b(n_11786), .c(n_11087), .d(n_10784), .o(n_12770) );
na02s02 TIMEBOOST_cell_43176 ( .a(TIMEBOOST_net_13826), .b(FE_OFN1295_n_4098), .o(TIMEBOOST_net_12064) );
na04f04 g54885_u0 ( .a(n_11085), .b(n_11784), .c(n_11084), .d(n_11083), .o(n_12542) );
na04f04 g54886_u0 ( .a(n_16586), .b(n_16585), .c(n_11079), .d(n_11081), .o(n_12541) );
na02s02 TIMEBOOST_cell_43177 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__Q), .b(n_4451), .o(TIMEBOOST_net_13827) );
na04f04 g54888_u0 ( .a(n_11782), .b(n_11783), .c(n_11072), .d(n_11073), .o(n_12539) );
na02s02 TIMEBOOST_cell_43178 ( .a(TIMEBOOST_net_13827), .b(FE_OFN1204_n_4090), .o(TIMEBOOST_net_12518) );
na04f04 g54891_u0 ( .a(n_11063), .b(n_11780), .c(n_11064), .d(n_11778), .o(n_12536) );
na04f04 g54893_u0 ( .a(n_11776), .b(n_11059), .c(n_11057), .d(n_11058), .o(n_12534) );
na04f04 g54895_u0 ( .a(n_11050), .b(n_11049), .c(n_11051), .d(n_11048), .o(n_12532) );
na04f04 g54896_u0 ( .a(n_11775), .b(n_11044), .c(n_11047), .d(n_11046), .o(n_12531) );
na04f04 g54897_u0 ( .a(n_10781), .b(n_11043), .c(n_11774), .d(n_11042), .o(n_12769) );
na04f04 g54899_u0 ( .a(n_11038), .b(n_11034), .c(n_11037), .d(n_11036), .o(n_12529) );
in01f01 g54903_u0 ( .a(n_16131), .o(n_12858) );
in01f02 g54907_u0 ( .a(n_15301), .o(n_10825) );
na02m02 TIMEBOOST_cell_41645 ( .a(wbu_sel_in_313), .b(wishbone_slave_unit_fifos_wbr_be_in_265), .o(TIMEBOOST_net_13061) );
na02s02 TIMEBOOST_cell_37498 ( .a(TIMEBOOST_net_10987), .b(FE_OFN1807_n_4501), .o(TIMEBOOST_net_9640) );
na02m02 TIMEBOOST_cell_44567 ( .a(n_9034), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__Q), .o(TIMEBOOST_net_14522) );
na02s01 TIMEBOOST_cell_30888 ( .a(pci_target_unit_pcit_if_strd_addr_in_707), .b(pci_target_unit_del_sync_addr_in_225), .o(TIMEBOOST_net_9355) );
ao12f02 g54936_u0 ( .a(n_12479), .b(FE_OFN1553_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__Q), .o(n_12809) );
na02f02 g54937_u0 ( .a(n_12331), .b(n_12051), .o(n_12764) );
na02s01 TIMEBOOST_cell_42920 ( .a(TIMEBOOST_net_13698), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_11149) );
na02s01 TIMEBOOST_cell_37802 ( .a(TIMEBOOST_net_11139), .b(g61881_sb), .o(n_8068) );
na02s01 TIMEBOOST_cell_30956 ( .a(n_3744), .b(g64883_sb), .o(TIMEBOOST_net_9389) );
na02s01 TIMEBOOST_cell_37159 ( .a(n_15330), .b(n_2092), .o(TIMEBOOST_net_10818) );
na02f02 g54942_u0 ( .a(n_12326), .b(n_12325), .o(n_12759) );
na02f02 TIMEBOOST_cell_44568 ( .a(TIMEBOOST_net_14522), .b(FE_OFN2169_n_8567), .o(TIMEBOOST_net_13470) );
na02f02 g54944_u0 ( .a(n_12323), .b(n_12047), .o(n_12757) );
ao12f02 g54945_u0 ( .a(n_12417), .b(FE_OFN1757_n_12681), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__Q), .o(n_12756) );
na02m02 TIMEBOOST_cell_43344 ( .a(TIMEBOOST_net_13910), .b(g59118_sb), .o(n_8692) );
na02s04 TIMEBOOST_cell_37158 ( .a(TIMEBOOST_net_10817), .b(n_531), .o(n_1410) );
na02s01 TIMEBOOST_cell_36641 ( .a(parchk_pci_ad_reg_in_1219), .b(g65813_sb), .o(TIMEBOOST_net_10559) );
na02f02 TIMEBOOST_cell_44130 ( .a(TIMEBOOST_net_14303), .b(FE_OFN1411_n_8567), .o(TIMEBOOST_net_12747) );
na02f02 g54952_u0 ( .a(n_12318), .b(n_12045), .o(n_12750) );
ao12f02 g54953_u0 ( .a(n_12044), .b(FE_OFN1749_n_12004), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__Q), .o(n_12528) );
na02s01 TIMEBOOST_cell_42921 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__Q), .b(FE_OFN526_n_9899), .o(TIMEBOOST_net_13699) );
no02f08 TIMEBOOST_cell_37161 ( .a(n_15998), .b(FE_RN_709_0), .o(TIMEBOOST_net_10819) );
na02m02 TIMEBOOST_cell_43843 ( .a(n_9534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__Q), .o(TIMEBOOST_net_14160) );
na02s01 TIMEBOOST_cell_37160 ( .a(TIMEBOOST_net_10818), .b(TIMEBOOST_net_1006), .o(n_2093) );
na02f02 g54958_u0 ( .a(n_12471), .b(n_11840), .o(n_17029) );
na02f02 g54959_u0 ( .a(n_12469), .b(n_12413), .o(n_12806) );
na02s01 TIMEBOOST_cell_44804 ( .a(TIMEBOOST_net_14640), .b(g65779_db), .o(TIMEBOOST_net_274) );
na02f02 g54961_u0 ( .a(n_12309), .b(n_12035), .o(n_12744) );
na02s01 TIMEBOOST_cell_42922 ( .a(TIMEBOOST_net_13699), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_11173) );
na02s01 TIMEBOOST_cell_31784 ( .a(configuration_wb_err_addr_561), .b(conf_wb_err_addr_in_970), .o(TIMEBOOST_net_9803) );
ao12f04 g54964_u0 ( .a(n_12478), .b(FE_OFN1553_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__Q), .o(n_12805) );
na02s02 TIMEBOOST_cell_45728 ( .a(TIMEBOOST_net_15102), .b(FE_OFN1250_n_4093), .o(TIMEBOOST_net_13260) );
na02s02 TIMEBOOST_cell_43488 ( .a(TIMEBOOST_net_13982), .b(FE_OFN1236_n_6391), .o(TIMEBOOST_net_12613) );
na02s01 TIMEBOOST_cell_42923 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__Q), .b(FE_OFN560_n_9895), .o(TIMEBOOST_net_13700) );
na02f02 TIMEBOOST_cell_43844 ( .a(TIMEBOOST_net_14160), .b(FE_OFN1396_n_8567), .o(TIMEBOOST_net_12838) );
na03s02 TIMEBOOST_cell_31856 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__Q), .b(FE_OFN1129_g64577_p), .c(g63138_sb), .o(TIMEBOOST_net_9839) );
na02s01 TIMEBOOST_cell_30922 ( .a(pci_target_unit_pcit_if_strd_addr_in_702), .b(pci_target_unit_del_sync_addr_in_220), .o(TIMEBOOST_net_9372) );
na02s01 TIMEBOOST_cell_41925 ( .a(FE_OFN201_n_9230), .b(g57897_sb), .o(TIMEBOOST_net_13201) );
na02s01 TIMEBOOST_cell_37291 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__Q), .b(n_3792), .o(TIMEBOOST_net_10884) );
ao12f02 g54973_u0 ( .a(n_12300), .b(FE_OFN1734_n_16317), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__Q), .o(n_12736) );
na02m02 TIMEBOOST_cell_43845 ( .a(n_9505), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__Q), .o(TIMEBOOST_net_14161) );
na02s01 TIMEBOOST_cell_31737 ( .a(TIMEBOOST_net_9779), .b(FE_OFN258_n_9862), .o(n_9785) );
na02s01 TIMEBOOST_cell_45274 ( .a(TIMEBOOST_net_14875), .b(FE_OFN1260_n_4143), .o(TIMEBOOST_net_12102) );
na02s01 TIMEBOOST_cell_37457 ( .a(pci_target_unit_del_sync_addr_in_228), .b(parchk_pci_ad_reg_in_1229), .o(TIMEBOOST_net_10967) );
na02f02 g54978_u0 ( .a(n_12466), .b(n_12408), .o(n_16603) );
na02s02 TIMEBOOST_cell_37950 ( .a(TIMEBOOST_net_11213), .b(g58238_sb), .o(n_9553) );
na02s02 TIMEBOOST_cell_45275 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__Q), .b(n_3702), .o(TIMEBOOST_net_14876) );
ao12f02 g54981_u0 ( .a(n_12294), .b(FE_OFN1734_n_16317), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__Q), .o(n_12731) );
na02s02 TIMEBOOST_cell_45276 ( .a(TIMEBOOST_net_14876), .b(FE_OFN1285_n_4097), .o(TIMEBOOST_net_12132) );
na02s02 TIMEBOOST_cell_41812 ( .a(TIMEBOOST_net_13144), .b(FE_OFN1104_g64577_p), .o(TIMEBOOST_net_4305) );
na02s02 TIMEBOOST_cell_37500 ( .a(TIMEBOOST_net_10988), .b(g58356_db), .o(n_9466) );
na02f02 g54985_u0 ( .a(n_12292), .b(n_12011), .o(n_12727) );
ao12f02 g54986_u0 ( .a(n_12476), .b(FE_OFN1552_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__Q), .o(n_12801) );
na03s02 TIMEBOOST_cell_31854 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__Q), .b(FE_OFN1129_g64577_p), .c(g63096_sb), .o(TIMEBOOST_net_9838) );
na02f02 g54989_u0 ( .a(n_12008), .b(n_12009), .o(n_12522) );
na02f02 g54990_u0 ( .a(n_12097), .b(n_12402), .o(n_12724) );
na02s01 TIMEBOOST_cell_31782 ( .a(conf_wb_err_addr_in_948), .b(configuration_wb_err_addr_539), .o(TIMEBOOST_net_9802) );
na02f02 g54992_u0 ( .a(n_12289), .b(n_12007), .o(n_12722) );
na02s01 TIMEBOOST_cell_44805 ( .a(FE_OFN250_n_9789), .b(g57931_sb), .o(TIMEBOOST_net_14641) );
na02s01 TIMEBOOST_cell_45741 ( .a(n_1981), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__Q), .o(TIMEBOOST_net_15109) );
ao12f02 g54996_u0 ( .a(n_12003), .b(FE_OFN1562_n_12502), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__Q), .o(n_12519) );
na02s02 TIMEBOOST_cell_42125 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__Q), .b(n_3679), .o(TIMEBOOST_net_13301) );
na02s02 TIMEBOOST_cell_41900 ( .a(TIMEBOOST_net_13188), .b(n_4741), .o(n_7130) );
na02f02 g55001_u0 ( .a(n_12000), .b(n_12282), .o(n_12716) );
na02s02 TIMEBOOST_cell_45277 ( .a(n_424), .b(n_4912), .o(TIMEBOOST_net_14877) );
na02s01 TIMEBOOST_cell_31853 ( .a(TIMEBOOST_net_9837), .b(n_4660), .o(n_5713) );
ao12f02 g55005_u0 ( .a(n_12280), .b(FE_OFN1759_n_10780), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q), .o(n_12714) );
na02s01 TIMEBOOST_cell_37437 ( .a(TIMEBOOST_net_1492), .b(n_3423), .o(TIMEBOOST_net_10957) );
na03m02 TIMEBOOST_cell_36122 ( .a(n_14013), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__Q), .c(FE_OCP_RBN1995_n_13971), .o(n_14300) );
na02s01 TIMEBOOST_cell_30890 ( .a(pci_target_unit_pcit_if_strd_addr_in_696), .b(pci_target_unit_del_sync_addr_in_214), .o(TIMEBOOST_net_9356) );
na02s02 TIMEBOOST_cell_37952 ( .a(TIMEBOOST_net_11214), .b(g58229_sb), .o(n_9560) );
na02s01 TIMEBOOST_cell_42683 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(g64151_sb), .o(TIMEBOOST_net_13580) );
na02s01 TIMEBOOST_cell_37804 ( .a(TIMEBOOST_net_11140), .b(g61875_sb), .o(n_8082) );
na02s01 g65240_u1 ( .a(n_8511), .b(g65240_sb), .o(g65240_da) );
na02s02 TIMEBOOST_cell_31961 ( .a(TIMEBOOST_net_9891), .b(FE_OFN1698_n_5751), .o(TIMEBOOST_net_4829) );
na02s02 TIMEBOOST_cell_45278 ( .a(TIMEBOOST_net_14877), .b(FE_OFN1200_n_4090), .o(TIMEBOOST_net_12020) );
ao12f02 g55018_u0 ( .a(n_12271), .b(FE_OFN1735_n_16317), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__Q), .o(n_12705) );
na02s02 TIMEBOOST_cell_43584 ( .a(TIMEBOOST_net_14030), .b(FE_OFN1311_n_6624), .o(TIMEBOOST_net_12234) );
na02s02 TIMEBOOST_cell_41905 ( .a(TIMEBOOST_net_9831), .b(g54194_sb), .o(TIMEBOOST_net_13191) );
na02s02 TIMEBOOST_cell_45279 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__Q), .b(n_3718), .o(TIMEBOOST_net_14878) );
na02s01 TIMEBOOST_cell_37290 ( .a(TIMEBOOST_net_10883), .b(FE_OFN661_n_4392), .o(TIMEBOOST_net_9395) );
ao12f02 g55023_u0 ( .a(n_12459), .b(FE_OCP_RBN2013_FE_OCPN1895_FE_OFN1559_n_12042), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__Q), .o(n_12797) );
na02s02 TIMEBOOST_cell_45280 ( .a(TIMEBOOST_net_14878), .b(FE_OFN1260_n_4143), .o(TIMEBOOST_net_12052) );
na02f02 TIMEBOOST_cell_41656 ( .a(TIMEBOOST_net_13066), .b(g55851_sb), .o(TIMEBOOST_net_11701) );
ao12f02 g55026_u0 ( .a(n_12430), .b(FE_OFN1552_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__Q), .o(n_12699) );
na02s02 TIMEBOOST_cell_45281 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__Q), .b(n_4318), .o(TIMEBOOST_net_14879) );
na02s02 TIMEBOOST_cell_31960 ( .a(n_740), .b(wbm_adr_o_3_), .o(TIMEBOOST_net_9891) );
na02s02 TIMEBOOST_cell_45282 ( .a(TIMEBOOST_net_14879), .b(FE_OFN1258_n_4143), .o(TIMEBOOST_net_12085) );
na02f02 TIMEBOOST_cell_21981 ( .a(TIMEBOOST_net_6247), .b(n_13901), .o(TIMEBOOST_net_3018) );
ao12f02 g55031_u0 ( .a(n_12266), .b(FE_OFN1761_n_10780), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__Q), .o(n_12695) );
na02s02 TIMEBOOST_cell_41906 ( .a(TIMEBOOST_net_13191), .b(FE_OFN1085_n_13221), .o(n_13357) );
na02s01 TIMEBOOST_cell_37293 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__Q), .b(n_3761), .o(TIMEBOOST_net_10885) );
ao12f02 g55034_u0 ( .a(n_12264), .b(FE_OFN1558_n_12042), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q), .o(n_12693) );
na02s01 g65236_u1 ( .a(n_2648), .b(g65236_sb), .o(g65236_da) );
na02s01 TIMEBOOST_cell_41813 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q), .b(g65335_sb), .o(TIMEBOOST_net_13145) );
na02s01 TIMEBOOST_cell_37292 ( .a(TIMEBOOST_net_10884), .b(FE_OFN661_n_4392), .o(TIMEBOOST_net_9393) );
na02s01 TIMEBOOST_cell_45283 ( .a(n_4354), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__Q), .o(TIMEBOOST_net_14880) );
ao12f02 g55042_u0 ( .a(n_12258), .b(FE_OFN1760_n_10780), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__Q), .o(n_12688) );
na02m02 TIMEBOOST_cell_37794 ( .a(TIMEBOOST_net_11135), .b(g58605_sb), .o(TIMEBOOST_net_337) );
na02s01 TIMEBOOST_cell_41907 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__Q), .b(g58418_sb), .o(TIMEBOOST_net_13192) );
na02s01 TIMEBOOST_cell_37217 ( .a(parchk_pci_ad_reg_in_1219), .b(pci_target_unit_del_sync_addr_in_218), .o(TIMEBOOST_net_10847) );
na02s02 TIMEBOOST_cell_45284 ( .a(TIMEBOOST_net_14880), .b(FE_OFN1250_n_4093), .o(TIMEBOOST_net_12600) );
na02s01 TIMEBOOST_cell_37294 ( .a(TIMEBOOST_net_10885), .b(FE_OFN662_n_4392), .o(TIMEBOOST_net_9392) );
ao12f02 g55050_u0 ( .a(n_12382), .b(FE_OFN1757_n_12681), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__Q), .o(n_12682) );
na02m02 TIMEBOOST_cell_44287 ( .a(n_9207), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__Q), .o(TIMEBOOST_net_14382) );
na02s01 g65216_u1 ( .a(n_3030), .b(g65216_sb), .o(g65216_da) );
na02m02 TIMEBOOST_cell_31959 ( .a(TIMEBOOST_net_9890), .b(FE_OFN1697_n_5751), .o(TIMEBOOST_net_4828) );
na02s02 TIMEBOOST_cell_45285 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__Q), .b(n_4381), .o(TIMEBOOST_net_14881) );
ao12f02 g55055_u0 ( .a(n_12475), .b(FE_OFN1553_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__Q), .o(n_12792) );
na02s01 g64827_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__Q), .b(FE_OFN1810_n_4454), .o(g64827_db) );
na02s02 TIMEBOOST_cell_37216 ( .a(TIMEBOOST_net_10846), .b(n_1826), .o(n_1827) );
ao12f02 g55058_u0 ( .a(n_11964), .b(FE_OFN1562_n_12502), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__31__Q), .o(n_12503) );
in01f02 g55059_u0 ( .a(n_12501), .o(n_12677) );
na02m02 TIMEBOOST_cell_44569 ( .a(n_9427), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q), .o(TIMEBOOST_net_14523) );
na02f02 g55061_u0 ( .a(n_12376), .b(n_12375), .o(n_12676) );
na02f02 TIMEBOOST_cell_41596 ( .a(FE_OFN1436_n_9372), .b(TIMEBOOST_net_13036), .o(TIMEBOOST_net_11670) );
na02f02 g55063_u0 ( .a(n_12245), .b(n_11953), .o(n_12675) );
na02f02 g55064_u0 ( .a(n_16338), .b(n_12374), .o(n_12674) );
na02s01 TIMEBOOST_cell_37502 ( .a(TIMEBOOST_net_10989), .b(FE_OFN239_n_9832), .o(n_9594) );
ao12f02 g55066_u0 ( .a(n_12455), .b(FE_OFN1563_n_12502), .c(n_7373), .o(n_12791) );
na02f02 g55067_u0 ( .a(n_12242), .b(n_11952), .o(n_12672) );
na02s01 TIMEBOOST_cell_37297 ( .a(n_3780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q), .o(TIMEBOOST_net_10887) );
na02f02 g55069_u0 ( .a(n_12371), .b(n_12078), .o(n_12670) );
na02s01 TIMEBOOST_cell_42861 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__Q), .b(FE_OFN517_n_9697), .o(TIMEBOOST_net_13669) );
na02s01 TIMEBOOST_cell_31780 ( .a(configuration_wb_err_data_600), .b(parchk_pci_ad_out_in_1197), .o(TIMEBOOST_net_9801) );
na02f02 g55073_u0 ( .a(n_12236), .b(n_11949), .o(n_12667) );
na02f02 g55074_u0 ( .a(n_12235), .b(n_11948), .o(n_12666) );
na02m02 TIMEBOOST_cell_44205 ( .a(n_8990), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__Q), .o(TIMEBOOST_net_14341) );
na02s02 TIMEBOOST_cell_31958 ( .a(n_1675), .b(wbm_adr_o_4_), .o(TIMEBOOST_net_9890) );
na04f02 TIMEBOOST_cell_35970 ( .a(wbu_addr_in_254), .b(g52618_sb), .c(g52618_db), .d(TIMEBOOST_net_6329), .o(n_11852) );
ao12f02 g55078_u0 ( .a(n_12452), .b(FE_OFN1564_n_12502), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__Q), .o(n_12789) );
na02s01 TIMEBOOST_cell_37219 ( .a(parchk_pci_ad_reg_in_1227), .b(pci_target_unit_del_sync_addr_in_226), .o(TIMEBOOST_net_10848) );
na02s01 TIMEBOOST_cell_41842 ( .a(TIMEBOOST_net_13159), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_9724) );
ao12f02 g55081_u0 ( .a(n_12429), .b(FE_OFN1552_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__Q), .o(n_12662) );
na02s02 TIMEBOOST_cell_45286 ( .a(TIMEBOOST_net_14881), .b(FE_OFN1283_n_4097), .o(TIMEBOOST_net_12577) );
na02s01 TIMEBOOST_cell_37218 ( .a(TIMEBOOST_net_10847), .b(FE_OFN2096_n_2520), .o(TIMEBOOST_net_3417) );
na02s01 TIMEBOOST_cell_37596 ( .a(TIMEBOOST_net_11036), .b(g61799_sb), .o(n_8198) );
na02m02 TIMEBOOST_cell_41393 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q), .b(n_9562), .o(TIMEBOOST_net_12935) );
na02f02 g55087_u0 ( .a(n_12464), .b(n_12363), .o(n_12788) );
na02s02 TIMEBOOST_cell_45287 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__Q), .b(n_4226), .o(TIMEBOOST_net_14882) );
na02s01 TIMEBOOST_cell_31844 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_392), .b(FE_OFN2070_n_15978), .o(TIMEBOOST_net_9833) );
na02s02 TIMEBOOST_cell_37504 ( .a(TIMEBOOST_net_10990), .b(g58306_sb), .o(n_9505) );
na02s02 TIMEBOOST_cell_45288 ( .a(TIMEBOOST_net_14882), .b(FE_OFN1270_n_4095), .o(TIMEBOOST_net_12606) );
na02f02 g55092_u0 ( .a(n_11933), .b(n_11932), .o(n_16589) );
na02s02 TIMEBOOST_cell_45289 ( .a(n_4464), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q), .o(TIMEBOOST_net_14883) );
na03f02 TIMEBOOST_cell_35291 ( .a(TIMEBOOST_net_10060), .b(FE_OFN1369_n_8567), .c(g58621_sb), .o(n_9181) );
ao12f02 g55095_u0 ( .a(n_12073), .b(FE_OCP_RBN2272_n_10268), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__Q), .o(n_12495) );
na02s02 TIMEBOOST_cell_45290 ( .a(TIMEBOOST_net_14883), .b(FE_OFN1284_n_4097), .o(TIMEBOOST_net_12598) );
na02f04 TIMEBOOST_cell_37296 ( .a(TIMEBOOST_net_10886), .b(n_15927), .o(n_15928) );
na02m02 TIMEBOOST_cell_31957 ( .a(TIMEBOOST_net_9889), .b(FE_OFN1697_n_5751), .o(TIMEBOOST_net_4827) );
na02f02 g55099_u0 ( .a(n_12222), .b(n_11929), .o(n_12649) );
ao12f02 g55100_u0 ( .a(n_12474), .b(FE_OFN1552_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__Q), .o(n_12787) );
na02s02 TIMEBOOST_cell_37598 ( .a(TIMEBOOST_net_11037), .b(g61786_sb), .o(n_8231) );
na02s01 TIMEBOOST_cell_45291 ( .a(n_4443), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__28__Q), .o(TIMEBOOST_net_14884) );
na02s01 TIMEBOOST_cell_45292 ( .a(TIMEBOOST_net_14884), .b(FE_OFN1275_n_4096), .o(TIMEBOOST_net_12578) );
na02s01 TIMEBOOST_cell_31778 ( .a(configuration_wb_err_addr_534), .b(conf_wb_err_addr_in_943), .o(TIMEBOOST_net_9800) );
na02f02 g55107_u0 ( .a(n_12070), .b(n_12356), .o(n_12644) );
ao12f02 g55108_u0 ( .a(n_12451), .b(FE_OFN1556_n_12042), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__Q), .o(n_12786) );
na03f02 TIMEBOOST_cell_35289 ( .a(TIMEBOOST_net_10062), .b(FE_OFN1369_n_8567), .c(g58618_sb), .o(n_9184) );
ao12f02 g55110_u0 ( .a(n_12425), .b(FE_OFN1552_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__Q), .o(n_12642) );
na02s01 TIMEBOOST_cell_45293 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__Q), .b(n_4190), .o(TIMEBOOST_net_14885) );
na02m02 TIMEBOOST_cell_31956 ( .a(n_2259), .b(wbm_adr_o_8_), .o(TIMEBOOST_net_9889) );
na02s02 TIMEBOOST_cell_45294 ( .a(TIMEBOOST_net_14885), .b(FE_OFN1270_n_4095), .o(TIMEBOOST_net_12603) );
na03s02 TIMEBOOST_cell_34468 ( .a(wbm_adr_o_17_), .b(FE_OFN1699_n_5751), .c(g59230_sb), .o(TIMEBOOST_net_589) );
na03f02 TIMEBOOST_cell_36110 ( .a(FE_RN_92_0), .b(n_10977), .c(n_12586), .o(n_12848) );
ao12f02 g55116_u0 ( .a(n_12450), .b(FE_OFN1564_n_12502), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__Q), .o(n_12785) );
na02s02 TIMEBOOST_cell_31842 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_389), .b(FE_OFN2070_n_15978), .o(TIMEBOOST_net_9832) );
na02s01 TIMEBOOST_cell_9748 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__Q), .b(g65868_sb), .o(TIMEBOOST_net_1441) );
na02f02 TIMEBOOST_cell_44235 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__Q), .b(n_8995), .o(TIMEBOOST_net_14356) );
na02f02 TIMEBOOST_cell_42430 ( .a(TIMEBOOST_net_13453), .b(g57521_sb), .o(n_10316) );
na02s01 TIMEBOOST_cell_45623 ( .a(FE_OFN239_n_9832), .b(g58059_sb), .o(TIMEBOOST_net_15050) );
na03s02 TIMEBOOST_cell_33360 ( .a(n_4482), .b(n_6), .c(g64852_sb), .o(TIMEBOOST_net_277) );
na02f02 TIMEBOOST_cell_44356 ( .a(TIMEBOOST_net_14416), .b(FE_OFN1382_n_8567), .o(TIMEBOOST_net_12851) );
na02f02 TIMEBOOST_cell_44262 ( .a(TIMEBOOST_net_14369), .b(FE_OFN1381_n_8567), .o(TIMEBOOST_net_12934) );
na03s01 TIMEBOOST_cell_34018 ( .a(TIMEBOOST_net_972), .b(g62111_sb), .c(g62111_db), .o(n_5587) );
na03s02 TIMEBOOST_cell_33359 ( .a(n_4672), .b(g65005_sb), .c(g65005_db), .o(n_4351) );
na04f04 g55132_u0 ( .a(n_10956), .b(n_9296), .c(n_10120), .d(n_9297), .o(n_12154) );
na02s02 TIMEBOOST_cell_41984 ( .a(TIMEBOOST_net_13230), .b(g62883_sb), .o(n_6111) );
na03s01 TIMEBOOST_cell_34019 ( .a(TIMEBOOST_net_976), .b(g62114_sb), .c(g62114_db), .o(n_5582) );
na02f02 TIMEBOOST_cell_42432 ( .a(TIMEBOOST_net_13454), .b(g57258_sb), .o(n_10421) );
na02s01 TIMEBOOST_cell_45624 ( .a(TIMEBOOST_net_15050), .b(g58059_db), .o(n_9731) );
na02m02 TIMEBOOST_cell_45781 ( .a(n_3385), .b(n_7618), .o(TIMEBOOST_net_15129) );
na02f02 TIMEBOOST_cell_42502 ( .a(TIMEBOOST_net_13489), .b(g57109_sb), .o(n_10478) );
na02s01 TIMEBOOST_cell_45625 ( .a(FE_OFN233_n_9876), .b(g58186_sb), .o(TIMEBOOST_net_15051) );
na03s02 TIMEBOOST_cell_33357 ( .a(n_4476), .b(g64882_sb), .c(g64882_db), .o(n_4418) );
na02m02 TIMEBOOST_cell_45782 ( .a(TIMEBOOST_net_15129), .b(g59807_da), .o(n_7616) );
na03s02 TIMEBOOST_cell_33355 ( .a(n_4442), .b(g64910_sb), .c(g64910_db), .o(n_4402) );
na03s02 TIMEBOOST_cell_33353 ( .a(n_4442), .b(g64934_sb), .c(g64934_db), .o(n_4385) );
na02f02 TIMEBOOST_cell_44703 ( .a(TIMEBOOST_net_10099), .b(FE_OFN1472_g52675_p), .o(TIMEBOOST_net_14590) );
na02f02 TIMEBOOST_cell_44204 ( .a(TIMEBOOST_net_14340), .b(FE_OFN1402_n_8567), .o(TIMEBOOST_net_12736) );
na02f02 TIMEBOOST_cell_41562 ( .a(TIMEBOOST_net_13019), .b(g57387_sb), .o(n_11357) );
na03s02 TIMEBOOST_cell_33350 ( .a(n_4465), .b(g64980_sb), .c(g64980_db), .o(n_4365) );
na02f02 TIMEBOOST_cell_44704 ( .a(TIMEBOOST_net_14590), .b(g52527_sb), .o(n_13694) );
na02f02 TIMEBOOST_cell_41632 ( .a(TIMEBOOST_net_13054), .b(FE_OFN1438_n_9372), .o(TIMEBOOST_net_11676) );
na02s01 TIMEBOOST_cell_9746 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__Q), .b(g65816_sb), .o(TIMEBOOST_net_1440) );
na02m02 TIMEBOOST_cell_31955 ( .a(TIMEBOOST_net_9888), .b(FE_OFN1697_n_5751), .o(TIMEBOOST_net_4826) );
na02s01 TIMEBOOST_cell_9744 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q), .b(g65814_sb), .o(TIMEBOOST_net_1439) );
na02s02 TIMEBOOST_cell_37600 ( .a(TIMEBOOST_net_11038), .b(g61787_sb), .o(n_8229) );
ao12f02 g55161_u0 ( .a(n_12212), .b(FE_OFN1759_n_10780), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__Q), .o(n_12632) );
na02f02 g55162_u0 ( .a(n_12473), .b(n_12351), .o(n_12784) );
na02s02 TIMEBOOST_cell_41844 ( .a(TIMEBOOST_net_13160), .b(FE_OFN262_n_9851), .o(n_9421) );
na02s02 TIMEBOOST_cell_43179 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__30__Q), .b(n_3790), .o(TIMEBOOST_net_13828) );
na02s01 TIMEBOOST_cell_37506 ( .a(TIMEBOOST_net_10991), .b(TIMEBOOST_net_3509), .o(n_8255) );
na02s02 TIMEBOOST_cell_45295 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__Q), .b(n_3728), .o(TIMEBOOST_net_14886) );
na02f02 g55167_u0 ( .a(n_12208), .b(n_12207), .o(n_15439) );
na02f02 g55168_u0 ( .a(n_12463), .b(n_12348), .o(n_12783) );
na02f02 TIMEBOOST_cell_43846 ( .a(TIMEBOOST_net_14161), .b(FE_OFN1422_n_8567), .o(TIMEBOOST_net_12937) );
na02m02 TIMEBOOST_cell_43847 ( .a(n_9495), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__Q), .o(TIMEBOOST_net_14162) );
na02s02 TIMEBOOST_cell_45296 ( .a(TIMEBOOST_net_14886), .b(FE_OFN1261_n_4143), .o(TIMEBOOST_net_12607) );
na03s02 TIMEBOOST_cell_37585 ( .a(n_1590), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__Q), .c(FE_OFN714_n_8140), .o(TIMEBOOST_net_11031) );
na02f02 g55173_u0 ( .a(n_12462), .b(n_12346), .o(n_16592) );
na02f02 g55174_u0 ( .a(n_12202), .b(n_12201), .o(n_12623) );
na03s02 TIMEBOOST_cell_34469 ( .a(pci_target_unit_wishbone_master_bc_register_reg_3__Q), .b(g52593_sb), .c(TIMEBOOST_net_882), .o(n_14683) );
na02s02 TIMEBOOST_cell_45297 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__Q), .b(n_4250), .o(TIMEBOOST_net_14887) );
na03f02 TIMEBOOST_cell_35290 ( .a(TIMEBOOST_net_10061), .b(FE_OFN1369_n_8567), .c(g58619_sb), .o(n_9183) );
na02f02 TIMEBOOST_cell_43848 ( .a(TIMEBOOST_net_14162), .b(FE_OFN1391_n_8567), .o(TIMEBOOST_net_12895) );
ao12f02 g55179_u0 ( .a(n_12449), .b(FE_OCP_RBN2013_FE_OCPN1895_FE_OFN1559_n_12042), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__Q), .o(n_12781) );
na02s02 TIMEBOOST_cell_45298 ( .a(TIMEBOOST_net_14887), .b(FE_OFN1295_n_4098), .o(TIMEBOOST_net_12519) );
na02s01 TIMEBOOST_cell_37584 ( .a(TIMEBOOST_net_11030), .b(g61769_sb), .o(n_8271) );
ao12f02 g55182_u0 ( .a(n_12423), .b(FE_OFN1552_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__Q), .o(n_12619) );
na02s02 TIMEBOOST_cell_31954 ( .a(n_2271), .b(wbm_adr_o_5_), .o(TIMEBOOST_net_9888) );
na02f02 g55184_u0 ( .a(n_12198), .b(n_11897), .o(n_12617) );
na02s01 TIMEBOOST_cell_31776 ( .a(configuration_wb_err_cs_bit_565), .b(conf_wb_err_bc_in_847), .o(TIMEBOOST_net_9799) );
na02f02 g55186_u0 ( .a(n_11896), .b(n_12197), .o(n_12615) );
ao12f02 g55187_u0 ( .a(n_12448), .b(FE_OFN1565_n_12502), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__Q), .o(n_12780) );
na02f02 g55188_u0 ( .a(n_12194), .b(n_11895), .o(n_12614) );
na04f02 TIMEBOOST_cell_14749 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__Q), .b(FE_OFN1394_n_8567), .c(n_8562), .d(g58586_sb), .o(n_8959) );
na02s02 TIMEBOOST_cell_45299 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__Q), .b(n_3664), .o(TIMEBOOST_net_14888) );
na02s01 TIMEBOOST_cell_42924 ( .a(TIMEBOOST_net_13700), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_11176) );
na02s01 TIMEBOOST_cell_37508 ( .a(TIMEBOOST_net_10992), .b(g64265_db), .o(n_3908) );
ao12f02 g55193_u0 ( .a(n_12447), .b(FE_OCP_RBN2013_FE_OCPN1895_FE_OFN1559_n_12042), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__14__Q), .o(n_12779) );
na02s01 TIMEBOOST_cell_37299 ( .a(n_3747), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__Q), .o(TIMEBOOST_net_10888) );
na02s02 TIMEBOOST_cell_45300 ( .a(TIMEBOOST_net_14888), .b(FE_OFN1249_n_4093), .o(TIMEBOOST_net_12592) );
ao12f02 g55196_u0 ( .a(n_11891), .b(FE_OFN1565_n_12502), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__14__Q), .o(n_12484) );
na04f02 TIMEBOOST_cell_14751 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__Q), .b(FE_OFN1394_n_8567), .c(n_8554), .d(g58594_sb), .o(n_8902) );
na02s01 TIMEBOOST_cell_30924 ( .a(pci_target_unit_pcit_if_strd_addr_in_710), .b(pci_target_unit_del_sync_addr_in_228), .o(TIMEBOOST_net_9373) );
na02s03 TIMEBOOST_cell_45773 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__Q), .b(n_13178), .o(TIMEBOOST_net_15125) );
na02s02 TIMEBOOST_cell_37440 ( .a(TIMEBOOST_net_10958), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(n_14738) );
na02s01 TIMEBOOST_cell_30936 ( .a(n_3752), .b(g64986_sb), .o(TIMEBOOST_net_9379) );
na02s01 TIMEBOOST_cell_45045 ( .a(n_1945), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__Q), .o(TIMEBOOST_net_14761) );
ao12f02 g55204_u0 ( .a(n_12186), .b(FE_OFN1760_n_10780), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__Q), .o(n_12602) );
na02s01 TIMEBOOST_cell_37298 ( .a(TIMEBOOST_net_10887), .b(FE_OFN636_n_4669), .o(TIMEBOOST_net_3626) );
na03f02 TIMEBOOST_cell_35293 ( .a(TIMEBOOST_net_10058), .b(FE_OFN1369_n_8567), .c(g58620_sb), .o(n_9182) );
na02s02 TIMEBOOST_cell_41846 ( .a(TIMEBOOST_net_13161), .b(FE_OFN272_n_9828), .o(n_9541) );
na02s01 TIMEBOOST_cell_37586 ( .a(TIMEBOOST_net_11031), .b(g61803_sb), .o(n_8189) );
na02m02 TIMEBOOST_cell_31953 ( .a(TIMEBOOST_net_9887), .b(FE_OFN1699_n_5751), .o(TIMEBOOST_net_4824) );
na02s02 TIMEBOOST_cell_45301 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__Q), .b(n_3670), .o(TIMEBOOST_net_14889) );
ao12f02 g55212_u0 ( .a(n_11885), .b(FE_OFN1749_n_12004), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__Q), .o(n_12480) );
no02f04 g55217_u0 ( .a(n_15001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__56), .o(n_12479) );
na03s02 TIMEBOOST_cell_37589 ( .a(n_1859), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__Q), .c(FE_OFN709_n_8232), .o(TIMEBOOST_net_11033) );
na02s02 TIMEBOOST_cell_38018 ( .a(TIMEBOOST_net_11247), .b(g61815_sb), .o(n_8161) );
na02m02 TIMEBOOST_cell_30739 ( .a(wbu_addr_in_258), .b(TIMEBOOST_net_9280), .o(TIMEBOOST_net_126) );
no02f04 g55221_u0 ( .a(n_15001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__59), .o(n_12478) );
na02m02 TIMEBOOST_cell_43849 ( .a(n_9519), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__Q), .o(TIMEBOOST_net_14163) );
na02f02 g55223_u0 ( .a(FE_OFN1513_n_14987), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__Q), .o(n_12433) );
no02f01 g55224_u0 ( .a(FE_OCP_RBN1922_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__62), .o(n_12476) );
na02f02 TIMEBOOST_cell_43778 ( .a(TIMEBOOST_net_14127), .b(FE_OFN1386_n_8567), .o(TIMEBOOST_net_12942) );
na02f02 g55226_u0 ( .a(FE_OCP_RBN1980_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__Q), .o(n_12124) );
na02m02 TIMEBOOST_cell_44357 ( .a(n_8996), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__Q), .o(TIMEBOOST_net_14417) );
na02f02 g55228_u0 ( .a(FE_OCPN1827_n_14995), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__Q), .o(n_12122) );
no02f02 g55229_u0 ( .a(FE_OCP_RBN1922_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__67), .o(n_12430) );
na02s01 TIMEBOOST_cell_42673 ( .a(n_4444), .b(g65037_sb), .o(TIMEBOOST_net_13575) );
na02s02 TIMEBOOST_cell_37588 ( .a(TIMEBOOST_net_11032), .b(g62015_sb), .o(n_7865) );
na02f02 TIMEBOOST_cell_22072 ( .a(n_13873), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__Q), .o(TIMEBOOST_net_6293) );
no02f04 g55233_u0 ( .a(n_15001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__70), .o(n_12475) );
na02f02 g55234_u0 ( .a(FE_OCP_RBN1979_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__Q), .o(n_12117) );
na02f02 g55235_u0 ( .a(FE_OCPN1827_n_14995), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q), .o(n_12116) );
na02f02 g55236_u0 ( .a(FE_OCPN1827_n_14995), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__Q), .o(n_12115) );
no02f02 g55237_u0 ( .a(FE_OCP_RBN1922_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__43), .o(n_12429) );
na02f02 g55238_u0 ( .a(FE_OFN1513_n_14987), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__5__Q), .o(n_12427) );
na02s02 TIMEBOOST_cell_30747 ( .a(TIMEBOOST_net_9284), .b(wishbone_slave_unit_pcim_if_wbw_cbe_in_416), .o(TIMEBOOST_net_1029) );
no02f02 g55240_u0 ( .a(FE_OCP_RBN1922_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__46), .o(n_12474) );
no02f02 g55241_u0 ( .a(FE_OCP_RBN1922_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__47), .o(n_12425) );
na03s02 TIMEBOOST_cell_37591 ( .a(n_1610), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__Q), .c(FE_OFN716_n_8176), .o(TIMEBOOST_net_11034) );
na02s02 g55243_u0 ( .a(FE_OCPN1827_n_14995), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q), .o(n_12473) );
na02s01 TIMEBOOST_cell_30863 ( .a(TIMEBOOST_net_9342), .b(FE_OFN227_n_9841), .o(n_9670) );
na02f02 g55245_u0 ( .a(FE_OFN1513_n_14987), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__Q), .o(n_12113) );
no02f02 g55246_u0 ( .a(FE_OCP_RBN1922_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__51), .o(n_12423) );
na02f02 g55247_u0 ( .a(FE_OCP_RBN1924_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__Q), .o(n_12112) );
na02f02 TIMEBOOST_cell_41370 ( .a(TIMEBOOST_net_12923), .b(g57324_sb), .o(n_11425) );
na02s02 TIMEBOOST_cell_30935 ( .a(TIMEBOOST_net_9378), .b(g64878_sb), .o(n_3709) );
na02s01 TIMEBOOST_cell_37590 ( .a(TIMEBOOST_net_11033), .b(g61913_sb), .o(n_7995) );
na02s01 TIMEBOOST_cell_31774 ( .a(parchk_pci_ad_out_in_1186), .b(configuration_wb_err_data_589), .o(TIMEBOOST_net_9798) );
na02s02 TIMEBOOST_cell_43676 ( .a(TIMEBOOST_net_14076), .b(g58635_db), .o(n_8847) );
na02m02 TIMEBOOST_cell_31952 ( .a(wbm_adr_o_7_), .b(n_2224), .o(TIMEBOOST_net_9887) );
na03f02 TIMEBOOST_cell_36177 ( .a(n_11816), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__Q), .c(FE_OCPN1866_n_12377), .o(n_12668) );
na03f02 TIMEBOOST_cell_36155 ( .a(FE_OFN1583_n_12306), .b(TIMEBOOST_net_10249), .c(FE_OFN1762_n_10780), .o(n_12763) );
na02f02 TIMEBOOST_cell_45857 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__15__Q), .b(FE_OCP_RBN1979_n_10273), .o(TIMEBOOST_net_15167) );
no02f02 g55257_u0 ( .a(n_12381), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__330), .o(n_12417) );
na03s02 TIMEBOOST_cell_37677 ( .a(n_1909), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__Q), .c(FE_OFN714_n_8140), .o(TIMEBOOST_net_11077) );
na02s01 TIMEBOOST_cell_43036 ( .a(TIMEBOOST_net_13756), .b(g57906_db), .o(n_9221) );
na02s02 TIMEBOOST_cell_43180 ( .a(TIMEBOOST_net_13828), .b(FE_OFN1282_n_4097), .o(TIMEBOOST_net_12061) );
na02s01 TIMEBOOST_cell_37620 ( .a(TIMEBOOST_net_11048), .b(g61791_sb), .o(n_8218) );
na02s02 TIMEBOOST_cell_31830 ( .a(g53940_sb), .b(FE_OFN2072_n_15978), .o(TIMEBOOST_net_9826) );
na02f02 g55263_u0 ( .a(FE_OCP_RBN1976_n_12381), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__Q), .o(n_12471) );
na02f02 g55264_u0 ( .a(FE_OFN2209_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__Q), .o(n_12469) );
na02f02 g55265_u0 ( .a(n_12362), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__Q), .o(n_12413) );
na02s02 TIMEBOOST_cell_36830 ( .a(TIMEBOOST_net_10653), .b(g62607_db), .o(n_6338) );
na02m02 TIMEBOOST_cell_31949 ( .a(TIMEBOOST_net_9885), .b(FE_OFN1697_n_5751), .o(TIMEBOOST_net_4822) );
na02s01 TIMEBOOST_cell_37510 ( .a(TIMEBOOST_net_10993), .b(g64347_db), .o(n_3830) );
na02s02 TIMEBOOST_cell_36685 ( .a(FE_OFN272_n_9828), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__Q), .o(TIMEBOOST_net_10581) );
na02s02 TIMEBOOST_cell_30921 ( .a(TIMEBOOST_net_9371), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_3765) );
na02f02 g55271_u0 ( .a(FE_OFN2209_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__Q), .o(n_12468) );
na02f01 g55272_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__Q), .o(n_12101) );
na02f02 TIMEBOOST_cell_41208 ( .a(TIMEBOOST_net_12842), .b(g57389_sb), .o(n_10376) );
na02f02 g55274_u0 ( .a(FE_OFN1572_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__Q), .o(n_12466) );
na02f02 g55275_u0 ( .a(n_12362), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__Q), .o(n_12408) );
na02f01 g55276_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__Q), .o(n_12100) );
na02f02 g55277_u0 ( .a(FE_OFN2210_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__23__Q), .o(n_12406) );
na02f02 TIMEBOOST_cell_41298 ( .a(TIMEBOOST_net_12887), .b(g57151_sb), .o(n_11599) );
na02s01 TIMEBOOST_cell_31772 ( .a(configuration_wb_err_cs_bit31_24), .b(conf_wb_err_bc_in), .o(TIMEBOOST_net_9797) );
na02f02 g55280_u0 ( .a(FE_OFN1753_n_12086), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__Q), .o(n_12097) );
na02s01 TIMEBOOST_cell_37512 ( .a(TIMEBOOST_net_10994), .b(g64232_db), .o(n_3940) );
na02f02 g55282_u0 ( .a(FE_OFN1568_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__Q), .o(n_12402) );
na02s02 TIMEBOOST_cell_43481 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__Q), .b(n_1850), .o(TIMEBOOST_net_13979) );
na02s01 TIMEBOOST_cell_31770 ( .a(configuration_wb_err_addr_540), .b(conf_wb_err_addr_in_949), .o(TIMEBOOST_net_9796) );
na02s01 TIMEBOOST_cell_42660 ( .a(TIMEBOOST_net_13568), .b(g65022_db), .o(n_3631) );
na02s01 TIMEBOOST_cell_45742 ( .a(TIMEBOOST_net_15109), .b(FE_OFN716_n_8176), .o(TIMEBOOST_net_11054) );
na02f02 TIMEBOOST_cell_41210 ( .a(TIMEBOOST_net_12843), .b(g57597_sb), .o(n_10795) );
na02s01 TIMEBOOST_cell_41901 ( .a(g61698_sb), .b(g61698_db), .o(TIMEBOOST_net_13189) );
na02s02 TIMEBOOST_cell_43181 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__Q), .b(n_3659), .o(TIMEBOOST_net_13829) );
na02m02 TIMEBOOST_cell_31948 ( .a(wbm_adr_o_9_), .b(n_2739), .o(TIMEBOOST_net_9885) );
na02f02 TIMEBOOST_cell_42529 ( .a(TIMEBOOST_net_6242), .b(n_135), .o(TIMEBOOST_net_13503) );
na02f02 g55292_u0 ( .a(FE_OFN1553_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__Q), .o(n_12393) );
na02s01 TIMEBOOST_cell_44889 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(g65766_sb), .o(TIMEBOOST_net_14683) );
na03s02 TIMEBOOST_cell_37955 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__Q), .b(FE_OFN589_n_9692), .c(FE_OFN270_n_9836), .o(TIMEBOOST_net_11216) );
na02f01 g55295_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__Q), .o(n_12090) );
na02s02 TIMEBOOST_cell_41908 ( .a(TIMEBOOST_net_13192), .b(g58418_db), .o(n_8998) );
na02f02 g55297_u0 ( .a(FE_OFN2210_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q), .o(n_12389) );
na02f02 TIMEBOOST_cell_41300 ( .a(TIMEBOOST_net_12888), .b(g57147_sb), .o(n_11603) );
na02m01 g55299_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__Q), .o(n_12088) );
na02s01 TIMEBOOST_cell_37954 ( .a(TIMEBOOST_net_11215), .b(g58139_sb), .o(n_9657) );
na02s01 TIMEBOOST_cell_41787 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__Q), .b(g58267_sb), .o(TIMEBOOST_net_13132) );
na02s02 TIMEBOOST_cell_45727 ( .a(n_3758), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__Q), .o(TIMEBOOST_net_15102) );
na02m01 g55303_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__Q), .o(n_12084) );
na02s02 TIMEBOOST_cell_41909 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__Q), .b(g58370_sb), .o(TIMEBOOST_net_13193) );
na02s01 TIMEBOOST_cell_42914 ( .a(TIMEBOOST_net_13695), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_11183) );
na02f02 g55308_u0 ( .a(FE_OFN2209_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__Q), .o(n_12465) );
na02f02 g55309_u0 ( .a(n_12362), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__Q), .o(n_12383) );
no02f02 g55310_u0 ( .a(n_12381), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__342), .o(n_12382) );
na02f01 g55311_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__Q), .o(n_12081) );
na02s02 TIMEBOOST_cell_41910 ( .a(TIMEBOOST_net_13193), .b(g58370_db), .o(n_9011) );
na02s02 TIMEBOOST_cell_44806 ( .a(TIMEBOOST_net_14641), .b(g57943_db), .o(n_9870) );
na02f02 g55314_u0 ( .a(FE_OFN1551_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__Q), .o(n_12379) );
na02f02 g55315_u0 ( .a(FE_OCP_RBN1975_n_12381), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__Q), .o(n_12378) );
na02f02 g55316_u0 ( .a(FE_OFN1572_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__Q), .o(n_12376) );
na02f02 g55317_u0 ( .a(n_12362), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__Q), .o(n_12375) );
na02f02 g55318_u0 ( .a(FE_OCP_RBN2272_n_10268), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__Q), .o(n_12374) );
na02s01 TIMEBOOST_cell_37514 ( .a(TIMEBOOST_net_10995), .b(g64237_db), .o(n_3935) );
na02f02 g55321_u0 ( .a(FE_OFN1551_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__Q), .o(n_12372) );
na02f02 g55322_u0 ( .a(FE_OFN1572_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__Q), .o(n_12371) );
na02f02 g55323_u0 ( .a(FE_OFN1751_n_12086), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__Q), .o(n_12078) );
na02s01 TIMEBOOST_cell_31768 ( .a(configuration_wb_err_data_596), .b(parchk_pci_ad_out_in_1193), .o(TIMEBOOST_net_9795) );
na02f02 g55325_u0 ( .a(FE_OFN1551_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__Q), .o(n_12369) );
na02s02 TIMEBOOST_cell_41911 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__Q), .b(g58344_sb), .o(TIMEBOOST_net_13194) );
na02f02 g55327_u0 ( .a(FE_OFN1568_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__Q), .o(n_12366) );
na02s01 TIMEBOOST_cell_37956 ( .a(TIMEBOOST_net_11216), .b(g58187_sb), .o(n_9598) );
na02f02 TIMEBOOST_cell_41212 ( .a(TIMEBOOST_net_12844), .b(g57583_sb), .o(n_10291) );
na02f02 g55330_u0 ( .a(FE_OFN1572_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__Q), .o(n_12464) );
na02f02 g55331_u0 ( .a(n_12362), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__Q), .o(n_12363) );
na02f01 g55332_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__Q), .o(n_12075) );
na02s02 TIMEBOOST_cell_37516 ( .a(TIMEBOOST_net_10996), .b(g64339_db), .o(n_3839) );
na03f02 TIMEBOOST_cell_36109 ( .a(FE_RN_182_0), .b(n_10870), .c(n_12563), .o(n_12825) );
no02f02 g55335_u0 ( .a(FE_OCPN1907_n_11767), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_2__6), .o(n_12073) );
na02m01 g55336_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__Q), .o(n_12072) );
na02s01 TIMEBOOST_cell_22060 ( .a(FE_OFN1025_n_11877), .b(g52484_da), .o(TIMEBOOST_net_6287) );
na02f04 TIMEBOOST_cell_31943 ( .a(TIMEBOOST_net_9882), .b(n_17030), .o(n_15188) );
na02s01 TIMEBOOST_cell_31766 ( .a(configuration_wb_err_cs_bit_566), .b(conf_wb_err_bc_in_848), .o(TIMEBOOST_net_9794) );
na02f02 g55340_u0 ( .a(FE_OFN1753_n_12086), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__8__Q), .o(n_12070) );
na02f02 g55341_u0 ( .a(FE_OFN1568_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__Q), .o(n_12356) );
na02s01 TIMEBOOST_cell_41902 ( .a(TIMEBOOST_net_13189), .b(n_4617), .o(n_5716) );
na02s01 TIMEBOOST_cell_39293 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(g65736_sb), .o(TIMEBOOST_net_11885) );
na02m02 TIMEBOOST_cell_44633 ( .a(n_9701), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__Q), .o(TIMEBOOST_net_14555) );
na02f02 TIMEBOOST_cell_41214 ( .a(TIMEBOOST_net_12845), .b(g57107_sb), .o(n_10479) );
na02f01 g55346_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__Q), .o(n_12068) );
na02s01 TIMEBOOST_cell_44807 ( .a(pci_target_unit_fifos_pcir_data_in_165), .b(g65746_sb), .o(TIMEBOOST_net_14642) );
na02f02 g55348_u0 ( .a(FE_OFN1568_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__Q), .o(n_12352) );
na02f02 g55349_u0 ( .a(FE_OFN1552_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__0__Q), .o(n_12351) );
na02s01 TIMEBOOST_cell_37518 ( .a(TIMEBOOST_net_10997), .b(g64242_sb), .o(TIMEBOOST_net_442) );
na02f02 TIMEBOOST_cell_41362 ( .a(TIMEBOOST_net_12919), .b(g57326_sb), .o(n_11424) );
na02f02 g55352_u0 ( .a(FE_OFN2209_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__Q), .o(n_12463) );
na02f02 g55353_u0 ( .a(n_12362), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__Q), .o(n_12348) );
na02f02 TIMEBOOST_cell_41216 ( .a(TIMEBOOST_net_12846), .b(g57500_sb), .o(n_11238) );
na02f02 g55355_u0 ( .a(FE_OFN2209_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__Q), .o(n_12462) );
na02f02 g55356_u0 ( .a(n_12362), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__Q), .o(n_12346) );
na02f02 TIMEBOOST_cell_41364 ( .a(TIMEBOOST_net_12920), .b(g57330_sb), .o(n_10397) );
na02f01 g55358_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__Q), .o(n_12066) );
na02s01 TIMEBOOST_cell_22062 ( .a(g52466_da), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_6288) );
na03f02 TIMEBOOST_cell_36111 ( .a(FE_RN_468_0), .b(n_11002), .c(n_12590), .o(n_12852) );
na02f02 TIMEBOOST_cell_43850 ( .a(TIMEBOOST_net_14163), .b(FE_OFN1419_n_8567), .o(TIMEBOOST_net_12825) );
na02s01 TIMEBOOST_cell_41777 ( .a(FE_OFN247_n_9112), .b(g58035_sb), .o(TIMEBOOST_net_13127) );
na02s01 TIMEBOOST_cell_31764 ( .a(configuration_wb_err_data_595), .b(parchk_pci_ad_out_in_1192), .o(TIMEBOOST_net_9793) );
na02f02 g55364_u0 ( .a(FE_OFN1553_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__Q), .o(n_12341) );
na03m02 TIMEBOOST_cell_34531 ( .a(TIMEBOOST_net_9878), .b(g54200_db), .c(TIMEBOOST_net_4766), .o(n_13505) );
na02s01 TIMEBOOST_cell_18082 ( .a(n_1598), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__Q), .o(TIMEBOOST_net_4298) );
na02s01 TIMEBOOST_cell_37520 ( .a(TIMEBOOST_net_10998), .b(g64187_sb), .o(TIMEBOOST_net_443) );
na02f02 g55368_u0 ( .a(FE_OFN1553_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__Q), .o(n_12338) );
na02f02 g55369_u0 ( .a(FE_OFN1572_n_11027), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__Q), .o(n_12337) );
na02s02 TIMEBOOST_cell_30923 ( .a(TIMEBOOST_net_9372), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_3764) );
na02f02 TIMEBOOST_cell_43851 ( .a(n_9100), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__Q), .o(TIMEBOOST_net_14164) );
na02s02 g55372_u0 ( .a(FE_OFN1554_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__15__Q), .o(n_12061) );
na02s01 TIMEBOOST_cell_42925 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__Q), .b(FE_OFN576_n_9902), .o(TIMEBOOST_net_13701) );
na03f02 TIMEBOOST_cell_36079 ( .a(n_11968), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__Q), .c(FE_OFN1748_n_12004), .o(n_12505) );
na02s01 TIMEBOOST_cell_44808 ( .a(TIMEBOOST_net_14642), .b(g65746_db), .o(TIMEBOOST_net_270) );
na02f01 g55376_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__Q), .o(n_12058) );
no03f02 TIMEBOOST_cell_44763 ( .a(FE_RN_343_0), .b(FE_RN_338_0), .c(FE_RN_348_0), .o(TIMEBOOST_net_14620) );
na02f02 g55378_u0 ( .a(FE_OFN1741_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__Q), .o(n_12334) );
na02f02 TIMEBOOST_cell_41936 ( .a(TIMEBOOST_net_13206), .b(g54151_sb), .o(n_13449) );
na02s02 TIMEBOOST_cell_30887 ( .a(TIMEBOOST_net_9354), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_3734) );
na02f02 g55381_u0 ( .a(n_12010), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__Q), .o(n_12056) );
na02f02 g55382_u0 ( .a(FE_OCPN1825_n_12030), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__Q), .o(n_12055) );
na02f02 g55383_u0 ( .a(FE_OFN1565_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__Q), .o(n_12054) );
na02f02 g55384_u0 ( .a(FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__Q), .o(n_12053) );
na02f02 g55385_u0 ( .a(FE_OFN1559_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__17__Q), .o(n_12052) );
na02f02 g55386_u0 ( .a(FE_OFN1762_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__Q), .o(n_12051) );
na02f02 g55387_u0 ( .a(FE_OFN1584_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__Q), .o(n_12331) );
na02f02 TIMEBOOST_cell_44358 ( .a(TIMEBOOST_net_14417), .b(FE_OFN1389_n_8567), .o(TIMEBOOST_net_12893) );
na02s01 TIMEBOOST_cell_42943 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__Q), .b(FE_OFN881_g64577_p), .o(TIMEBOOST_net_13710) );
na02s01 TIMEBOOST_cell_41726 ( .a(TIMEBOOST_net_13101), .b(g64847_db), .o(n_3724) );
na02f02 g55391_u0 ( .a(FE_OFN1566_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__18__Q), .o(n_12049) );
na02s01 TIMEBOOST_cell_30955 ( .a(TIMEBOOST_net_9388), .b(g64880_sb), .o(n_3707) );
na02f02 g55393_u0 ( .a(FE_OFN2202_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__Q), .o(n_12327) );
na02f02 g55394_u0 ( .a(n_12228), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__Q), .o(n_12326) );
na02f02 g55395_u0 ( .a(FE_OFN1749_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__Q), .o(n_12325) );
na02f02 g55396_u0 ( .a(FE_OFN1735_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__Q), .o(n_12047) );
na02f02 g55397_u0 ( .a(FE_OFN1741_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__Q), .o(n_12323) );
na02s01 TIMEBOOST_cell_37301 ( .a(n_3761), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__Q), .o(TIMEBOOST_net_10889) );
na02s02 TIMEBOOST_cell_45007 ( .a(pci_target_unit_fifos_pciw_addr_data_in_125), .b(g64097_sb), .o(TIMEBOOST_net_14742) );
na03s02 TIMEBOOST_cell_36683 ( .a(TIMEBOOST_net_1235), .b(g64122_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__Q), .o(TIMEBOOST_net_10580) );
na02s01 TIMEBOOST_cell_30749 ( .a(TIMEBOOST_net_9285), .b(g65270_sb), .o(TIMEBOOST_net_19) );
na03f02 TIMEBOOST_cell_35292 ( .a(TIMEBOOST_net_10059), .b(FE_OFN1369_n_8567), .c(g58616_sb), .o(n_9187) );
na02s01 TIMEBOOST_cell_42926 ( .a(TIMEBOOST_net_13701), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_11171) );
na02f02 g55404_u0 ( .a(FE_OFN1757_n_12681), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__Q), .o(n_11841) );
na02f02 g55405_u0 ( .a(FE_OFN1741_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__Q), .o(n_12318) );
na02f02 g55406_u0 ( .a(FE_OFN1735_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__Q), .o(n_12045) );
no02f02 g55407_u0 ( .a(FE_OCPN1834_n_11884), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__487), .o(n_12044) );
na02s01 TIMEBOOST_cell_42927 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__Q), .b(FE_OFN1648_n_9428), .o(TIMEBOOST_net_13702) );
na02s01 TIMEBOOST_cell_42609 ( .a(g58081_sb), .b(g58081_db), .o(TIMEBOOST_net_13543) );
na02s01 TIMEBOOST_cell_41727 ( .a(FE_OFN205_n_9140), .b(g58414_sb), .o(TIMEBOOST_net_13102) );
na02f02 g55411_u0 ( .a(FE_OFN1566_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__1__Q), .o(n_12041) );
na02f02 TIMEBOOST_cell_41308 ( .a(TIMEBOOST_net_12892), .b(g57114_sb), .o(n_11632) );
na02s01 TIMEBOOST_cell_30953 ( .a(TIMEBOOST_net_9387), .b(g64879_sb), .o(n_3708) );
na02f02 g55414_u0 ( .a(FE_OFN1757_n_12681), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__Q), .o(n_11840) );
na02f02 g55415_u0 ( .a(FE_OFN1735_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__Q), .o(n_12038) );
na02f02 g55416_u0 ( .a(FE_OFN1741_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__Q), .o(n_12310) );
na02f02 g55417_u0 ( .a(n_12001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__Q), .o(n_12037) );
na02f02 g55418_u0 ( .a(FE_OFN1749_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__Q), .o(n_12036) );
na02f02 g55419_u0 ( .a(n_11977), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__Q), .o(n_12035) );
na02f02 g55420_u0 ( .a(FE_OFN1748_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__Q), .o(n_12309) );
na02s01 TIMEBOOST_cell_42928 ( .a(TIMEBOOST_net_13702), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_11155) );
na02m02 TIMEBOOST_cell_30751 ( .a(TIMEBOOST_net_9286), .b(g66457_db), .o(n_1134) );
na02f02 g55423_u0 ( .a(FE_OFN1757_n_12681), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__Q), .o(n_11839) );
na02f02 g55424_u0 ( .a(FE_OFN1566_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__20__Q), .o(n_12032) );
na02f04 g55425_u0 ( .a(FE_OCPN1825_n_12030), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__20__Q), .o(n_12031) );
na02s02 TIMEBOOST_cell_30957 ( .a(TIMEBOOST_net_9389), .b(g64883_db), .o(n_3705) );
na02s01 TIMEBOOST_cell_41778 ( .a(TIMEBOOST_net_13127), .b(g58035_db), .o(n_9096) );
na02s01 TIMEBOOST_cell_42929 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__Q), .b(FE_OFN601_n_9687), .o(TIMEBOOST_net_13703) );
na02s02 TIMEBOOST_cell_30753 ( .a(TIMEBOOST_net_9287), .b(wishbone_slave_unit_pcim_if_wbw_cbe_in), .o(TIMEBOOST_net_1068) );
na03s02 TIMEBOOST_cell_36681 ( .a(TIMEBOOST_net_3706), .b(g64271_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q), .o(TIMEBOOST_net_10579) );
na02f02 g55431_u0 ( .a(FE_OFN1566_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__Q), .o(n_11838) );
na02m02 g55432_u0 ( .a(FE_OFN1760_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__Q), .o(n_12024) );
na02s01 TIMEBOOST_cell_30959 ( .a(TIMEBOOST_net_9390), .b(g64887_sb), .o(n_3703) );
na02f02 g55435_u0 ( .a(FE_OFN2202_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__Q), .o(n_12022) );
na02s01 TIMEBOOST_cell_42661 ( .a(n_3764), .b(g64897_sb), .o(TIMEBOOST_net_13569) );
na02s01 TIMEBOOST_cell_41926 ( .a(TIMEBOOST_net_13201), .b(g57897_db), .o(n_9227) );
na02s02 TIMEBOOST_cell_45702 ( .a(TIMEBOOST_net_15089), .b(FE_OFN1258_n_4143), .o(TIMEBOOST_net_12569) );
no02f04 g55439_u0 ( .a(n_12293), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__177), .o(n_12300) );
na02s01 TIMEBOOST_cell_30961 ( .a(TIMEBOOST_net_9391), .b(g64894_sb), .o(n_3699) );
na02f02 g55441_u0 ( .a(FE_OFN2202_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__Q), .o(n_12020) );
na02s01 TIMEBOOST_cell_37300 ( .a(TIMEBOOST_net_10888), .b(FE_OFN640_n_4669), .o(TIMEBOOST_net_3651) );
na02s01 TIMEBOOST_cell_42630 ( .a(TIMEBOOST_net_13553), .b(g64898_db), .o(n_3695) );
na02s01 TIMEBOOST_cell_41728 ( .a(TIMEBOOST_net_13102), .b(g58414_db), .o(n_9000) );
na02s02 TIMEBOOST_cell_30755 ( .a(TIMEBOOST_net_9288), .b(wishbone_slave_unit_pcim_if_wbw_cbe_in_417), .o(TIMEBOOST_net_1030) );
na02s01 TIMEBOOST_cell_42930 ( .a(TIMEBOOST_net_13703), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_11148) );
na02s01 TIMEBOOST_cell_44809 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(g65762_sb), .o(TIMEBOOST_net_14643) );
na02f02 TIMEBOOST_cell_41422 ( .a(TIMEBOOST_net_12949), .b(g57474_sb), .o(n_10340) );
no02f02 g55449_u0 ( .a(n_12293), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__178), .o(n_12294) );
na02s02 TIMEBOOST_cell_43182 ( .a(TIMEBOOST_net_13829), .b(FE_OFN1244_n_4092), .o(TIMEBOOST_net_12110) );
na02f02 TIMEBOOST_cell_43852 ( .a(TIMEBOOST_net_14164), .b(FE_OFN1380_n_8567), .o(TIMEBOOST_net_12896) );
na02s01 TIMEBOOST_cell_42903 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__Q), .b(FE_OFN516_n_9697), .o(TIMEBOOST_net_13690) );
na02f02 g55453_u0 ( .a(n_12010), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__23__Q), .o(n_12011) );
na02f02 g55454_u0 ( .a(FE_OFN1747_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__Q), .o(n_12292) );
na02s01 TIMEBOOST_cell_42877 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__Q), .b(FE_OFN596_n_9694), .o(TIMEBOOST_net_13677) );
na02s01 TIMEBOOST_cell_22144 ( .a(FE_OFN9_n_11877), .b(g52481_da), .o(TIMEBOOST_net_6329) );
na02f02 g55457_u0 ( .a(FE_OFN1759_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__Q), .o(n_12009) );
na02f02 g55458_u0 ( .a(FE_OFN1584_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__Q), .o(n_12008) );
no02f02 g55459_u0 ( .a(FE_OCP_RBN2291_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__374), .o(n_12290) );
na02s01 TIMEBOOST_cell_41927 ( .a(FE_OFN203_n_9228), .b(g57895_sb), .o(TIMEBOOST_net_13202) );
na02f02 g55461_u0 ( .a(FE_OFN1738_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__Q), .o(n_12289) );
na02f02 g55462_u0 ( .a(FE_OFN1733_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__Q), .o(n_12007) );
na02s01 TIMEBOOST_cell_42662 ( .a(TIMEBOOST_net_13569), .b(g64897_db), .o(n_3696) );
na02s01 TIMEBOOST_cell_41779 ( .a(FE_OFN247_n_9112), .b(g58004_sb), .o(TIMEBOOST_net_13128) );
na02f04 TIMEBOOST_cell_37022 ( .a(TIMEBOOST_net_10749), .b(g52521_sb), .o(n_13698) );
na02s02 TIMEBOOST_cell_43560 ( .a(TIMEBOOST_net_14018), .b(FE_OFN1314_n_6624), .o(TIMEBOOST_net_12221) );
no02f02 g55468_u0 ( .a(FE_OCP_RBN2286_FE_RN_494_0), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__258), .o(n_12003) );
na02f02 g55469_u0 ( .a(n_12001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__25__Q), .o(n_12002) );
na02f02 g55470_u0 ( .a(FE_OFN1747_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__Q), .o(n_12283) );
na02s01 TIMEBOOST_cell_42631 ( .a(FE_OFN245_n_9114), .b(g58255_sb), .o(TIMEBOOST_net_13554) );
na02f02 g55472_u0 ( .a(FE_OFN1742_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__Q), .o(n_12282) );
na02f02 g55473_u0 ( .a(FE_OFN1736_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__Q), .o(n_12000) );
no02f02 g55474_u0 ( .a(FE_OCP_RBN2292_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__376), .o(n_12461) );
na02s01 TIMEBOOST_cell_42878 ( .a(TIMEBOOST_net_13677), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_11217) );
no02f04 g55477_u0 ( .a(n_16587), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__532), .o(n_12280) );
na03m02 TIMEBOOST_cell_34425 ( .a(n_2699), .b(g59368_sb), .c(g59368_db), .o(n_7541) );
na02f02 g55479_u0 ( .a(FE_OFN1736_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__26__Q), .o(n_11996) );
na02m02 TIMEBOOST_cell_44359 ( .a(n_9660), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q), .o(TIMEBOOST_net_14418) );
na02f02 g55481_u0 ( .a(n_12010), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__Q), .o(n_11995) );
na02s02 TIMEBOOST_cell_30889 ( .a(TIMEBOOST_net_9355), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_3735) );
no02f02 g55483_u0 ( .a(n_12453), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__260), .o(n_12460) );
na02f02 TIMEBOOST_cell_41310 ( .a(TIMEBOOST_net_12893), .b(g57575_sb), .o(n_10294) );
na02s02 TIMEBOOST_cell_45302 ( .a(TIMEBOOST_net_14889), .b(FE_OFN1249_n_4093), .o(TIMEBOOST_net_12552) );
no02f02 g55486_u0 ( .a(FE_OCP_RBN2292_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__377), .o(n_12277) );
na02f02 g55487_u0 ( .a(n_11881), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__Q), .o(n_12276) );
na02f02 g55488_u0 ( .a(FE_OFN1562_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__Q), .o(n_11992) );
na02f02 g55489_u0 ( .a(FE_OFN2202_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__Q), .o(n_12275) );
na02f02 g55490_u0 ( .a(FE_OFN1577_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__Q), .o(n_12274) );
na02f02 g55491_u0 ( .a(FE_OFN1762_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__Q), .o(n_11991) );
na02f02 g55492_u0 ( .a(FE_OFN1583_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__Q), .o(n_11990) );
na02s02 g55493_u0 ( .a(n_12228), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__Q), .o(n_12273) );
na03f02 TIMEBOOST_cell_36057 ( .a(FE_OFN1601_n_13995), .b(TIMEBOOST_net_10175), .c(FE_OFN1605_n_13997), .o(n_16210) );
no02f02 g55495_u0 ( .a(n_12293), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__183), .o(n_12271) );
na02f02 TIMEBOOST_cell_41384 ( .a(TIMEBOOST_net_12930), .b(g57376_sb), .o(n_11372) );
na02f02 g55497_u0 ( .a(n_12001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__28__Q), .o(n_11988) );
na02s01 TIMEBOOST_cell_38074 ( .a(TIMEBOOST_net_11275), .b(FE_OFN1135_g64577_p), .o(TIMEBOOST_net_4520) );
na02s03 TIMEBOOST_cell_30761 ( .a(TIMEBOOST_net_9291), .b(n_1689), .o(TIMEBOOST_net_183) );
na02s01 TIMEBOOST_cell_31717 ( .a(TIMEBOOST_net_9769), .b(FE_OFN262_n_9851), .o(n_9716) );
na02s01 TIMEBOOST_cell_45025 ( .a(TIMEBOOST_net_4206), .b(g61969_db), .o(TIMEBOOST_net_14751) );
no02f02 g55502_u0 ( .a(FE_OCP_RBN2292_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__379), .o(n_12459) );
na02f02 TIMEBOOST_cell_41386 ( .a(TIMEBOOST_net_12931), .b(g57034_sb), .o(n_11698) );
na02f02 g55504_u0 ( .a(FE_OFN1761_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__Q), .o(n_11984) );
na02f04 TIMEBOOST_cell_37024 ( .a(TIMEBOOST_net_10750), .b(g52522_sb), .o(n_13735) );
na02f02 TIMEBOOST_cell_44360 ( .a(TIMEBOOST_net_14418), .b(FE_OFN1420_n_8567), .o(TIMEBOOST_net_12696) );
na02f02 TIMEBOOST_cell_41388 ( .a(TIMEBOOST_net_12932), .b(g57494_sb), .o(n_10331) );
na02f02 g55508_u0 ( .a(FE_OFN1739_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__Q), .o(n_12267) );
na02f02 TIMEBOOST_cell_41448 ( .a(TIMEBOOST_net_12962), .b(g57339_sb), .o(n_11413) );
na02s01 TIMEBOOST_cell_42663 ( .a(FE_OFN217_n_9889), .b(g58103_sb), .o(TIMEBOOST_net_13570) );
na02s01 TIMEBOOST_cell_32000 ( .a(configuration_pci_err_addr_501), .b(wbm_adr_o_31_), .o(TIMEBOOST_net_9911) );
no02f04 g55512_u0 ( .a(FE_OCP_RBN2293_FE_OFN1581_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__536), .o(n_12266) );
na02s01 TIMEBOOST_cell_37522 ( .a(TIMEBOOST_net_10999), .b(g64985_sb), .o(TIMEBOOST_net_9979) );
na02f02 g55514_u0 ( .a(FE_OFN1562_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__Q), .o(n_11822) );
no02f04 g55515_u0 ( .a(FE_OCP_RBN2292_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__380), .o(n_12264) );
na02s01 g65240_u3 ( .a(g65240_da), .b(g65240_db), .o(n_2643) );
na02f02 g55517_u0 ( .a(n_11977), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__Q), .o(n_11978) );
na03f02 TIMEBOOST_cell_14616 ( .a(TIMEBOOST_net_2412), .b(n_4205), .c(TIMEBOOST_net_586), .o(n_14817) );
no02f02 g55521_u0 ( .a(n_12453), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__236), .o(n_12457) );
na02f02 TIMEBOOST_cell_41424 ( .a(TIMEBOOST_net_12950), .b(g57203_sb), .o(n_10444) );
na02f02 g55523_u0 ( .a(FE_OFN1559_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__Q), .o(n_12259) );
no02f02 g55524_u0 ( .a(n_11762), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__509), .o(n_12258) );
na02f02 g55525_u0 ( .a(FE_OFN1762_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__Q), .o(n_11975) );
na02f02 g55526_u0 ( .a(FE_OFN1583_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__Q), .o(n_12257) );
na03f02 TIMEBOOST_cell_35294 ( .a(TIMEBOOST_net_10056), .b(FE_OFN1369_n_8567), .c(g58576_sb), .o(n_9192) );
na02s01 g65236_u3 ( .a(g65236_da), .b(g65236_db), .o(n_2649) );
na02s01 TIMEBOOST_cell_31818 ( .a(parchk_pci_ad_out_in_1181), .b(configuration_wb_err_data_584), .o(TIMEBOOST_net_9820) );
na02f02 g55530_u0 ( .a(FE_OFN1566_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__30__Q), .o(n_11973) );
na02f02 g55531_u0 ( .a(n_12010), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__Q), .o(n_11972) );
na02f02 TIMEBOOST_cell_41168 ( .a(TIMEBOOST_net_12822), .b(g57498_sb), .o(n_11240) );
na02s01 TIMEBOOST_cell_31695 ( .a(TIMEBOOST_net_9758), .b(g57952_sb), .o(n_9837) );
na02s01 TIMEBOOST_cell_42684 ( .a(TIMEBOOST_net_13580), .b(g64151_db), .o(n_4014) );
na02s01 TIMEBOOST_cell_41815 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__Q), .b(g58276_sb), .o(TIMEBOOST_net_13146) );
na02s01 g65235_u3 ( .a(g65235_da), .b(g65235_db), .o(n_2652) );
na02s02 g55537_u0 ( .a(FE_OFN1734_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__Q), .o(n_11970) );
na02f02 TIMEBOOST_cell_41170 ( .a(TIMEBOOST_net_12823), .b(g57423_sb), .o(n_11314) );
na02f02 g55539_u0 ( .a(n_12010), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__Q), .o(n_11968) );
na02s01 g65216_u3 ( .a(g65216_da), .b(g65216_db), .o(n_3031) );
na02s01 TIMEBOOST_cell_42664 ( .a(TIMEBOOST_net_13570), .b(g58103_db), .o(n_9693) );
na02f02 g55542_u0 ( .a(FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__31__Q), .o(n_12250) );
na02s02 TIMEBOOST_cell_37524 ( .a(TIMEBOOST_net_11000), .b(FE_OFN713_n_8140), .o(TIMEBOOST_net_4169) );
no02f02 g55544_u0 ( .a(FE_OCP_RBN2286_FE_RN_494_0), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__265), .o(n_11964) );
na02m02 g55545_u0 ( .a(FE_OFN1760_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__Q), .o(n_11962) );
na02f02 g55546_u0 ( .a(FE_OFN1579_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__Q), .o(n_11961) );
na02f02 g55547_u0 ( .a(FE_OFN2204_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__Q), .o(n_12248) );
na02f02 g55548_u0 ( .a(FE_OFN1559_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__Q), .o(n_12246) );
na02f02 g55549_u0 ( .a(FE_OCPN1825_n_12030), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__Q), .o(n_11960) );
na02f02 g55550_u0 ( .a(FE_OFN1563_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__Q), .o(n_11819) );
na03s02 TIMEBOOST_cell_31694 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__Q), .b(FE_OFN556_n_9864), .c(FE_OFN270_n_9836), .o(TIMEBOOST_net_9758) );
na02s02 TIMEBOOST_cell_45596 ( .a(TIMEBOOST_net_15036), .b(g65224_sb), .o(n_2663) );
na02f02 g55553_u0 ( .a(n_11823), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__Q), .o(n_11818) );
na02f02 g55554_u0 ( .a(FE_OFN1748_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__Q), .o(n_11957) );
na02f02 g55555_u0 ( .a(n_12001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__Q), .o(n_11956) );
na02s02 TIMEBOOST_cell_45703 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__Q), .b(n_4352), .o(TIMEBOOST_net_15090) );
na02s02 g55557_u0 ( .a(FE_OFN1734_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__Q), .o(n_11954) );
na02f02 g55558_u0 ( .a(n_11977), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__Q), .o(n_11953) );
na02f02 g55559_u0 ( .a(FE_OFN1749_n_12004), .b(n_395), .o(n_12245) );
na03s02 TIMEBOOST_cell_6318 ( .a(n_3761), .b(g64827_sb), .c(g64827_db), .o(n_3732) );
no02f02 g55561_u0 ( .a(n_12453), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__271), .o(n_12455) );
na02f02 g55562_u0 ( .a(FE_OFN1574_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__Q), .o(n_12244) );
na02f02 g55563_u0 ( .a(FE_OFN1559_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__Q), .o(n_12243) );
na02f02 g55564_u0 ( .a(FE_OFN1761_n_10780), .b(n_323), .o(n_11952) );
na02f02 g55565_u0 ( .a(FE_OFN1579_n_12306), .b(n_263), .o(n_12242) );
na02f02 TIMEBOOST_cell_42530 ( .a(TIMEBOOST_net_13503), .b(n_14971), .o(TIMEBOOST_net_11703) );
na02s02 g55567_u0 ( .a(FE_OFN1734_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__Q), .o(n_11951) );
na02s01 TIMEBOOST_cell_42665 ( .a(FE_OFN219_n_9853), .b(g58236_sb), .o(TIMEBOOST_net_13571) );
na02s01 TIMEBOOST_cell_42931 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__Q), .b(FE_OFN601_n_9687), .o(TIMEBOOST_net_13704) );
na02f02 g55570_u0 ( .a(FE_OFN1756_n_12681), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__Q), .o(n_11816) );
no02f02 g55571_u0 ( .a(n_12453), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__237), .o(n_12454) );
na02f02 g55572_u0 ( .a(FE_OFN1574_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__Q), .o(n_12238) );
na02f02 g55573_u0 ( .a(FE_OFN1559_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__Q), .o(n_12237) );
na02f02 g55574_u0 ( .a(FE_OFN1760_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__Q), .o(n_11949) );
na02f02 g55575_u0 ( .a(FE_OFN1579_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__Q), .o(n_12236) );
na02f02 g55576_u0 ( .a(n_12001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__Q), .o(n_11948) );
na02f02 g55577_u0 ( .a(FE_OFN1746_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__Q), .o(n_12235) );
na02s01 TIMEBOOST_cell_43285 ( .a(TIMEBOOST_net_4768), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_13881) );
na02s03 TIMEBOOST_cell_45759 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__Q), .b(n_13105), .o(TIMEBOOST_net_15118) );
na02s01 TIMEBOOST_cell_43286 ( .a(TIMEBOOST_net_13881), .b(g62038_sb), .o(n_7777) );
no02f02 g55581_u0 ( .a(n_12453), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__238), .o(n_12452) );
na02f02 TIMEBOOST_cell_41390 ( .a(TIMEBOOST_net_12933), .b(g57325_sb), .o(n_10399) );
na02s01 TIMEBOOST_cell_31816 ( .a(configuration_wb_err_data_578), .b(parchk_pci_ad_out_in_1175), .o(TIMEBOOST_net_9819) );
na02s02 TIMEBOOST_cell_41848 ( .a(TIMEBOOST_net_13162), .b(FE_OFN268_n_9880), .o(n_9712) );
na02s01 TIMEBOOST_cell_30775 ( .a(TIMEBOOST_net_9298), .b(n_2651), .o(TIMEBOOST_net_3274) );
na02s01 TIMEBOOST_cell_43183 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__Q), .b(n_3553), .o(TIMEBOOST_net_13830) );
na02s02 TIMEBOOST_cell_37526 ( .a(TIMEBOOST_net_11001), .b(FE_OFN704_n_8069), .o(TIMEBOOST_net_4149) );
na02s01 TIMEBOOST_cell_43287 ( .a(TIMEBOOST_net_4767), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_13882) );
na02s01 TIMEBOOST_cell_31814 ( .a(configuration_wb_err_data_577), .b(parchk_pci_ad_out_in_1174), .o(TIMEBOOST_net_9818) );
na02f02 g55590_u0 ( .a(FE_OFN1760_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__Q), .o(n_16631) );
na02f02 TIMEBOOST_cell_41392 ( .a(TIMEBOOST_net_12934), .b(g57375_sb), .o(n_10380) );
na02s03 TIMEBOOST_cell_45760 ( .a(TIMEBOOST_net_15118), .b(FE_OFN1326_n_13547), .o(TIMEBOOST_net_14951) );
na02s01 TIMEBOOST_cell_42666 ( .a(TIMEBOOST_net_13571), .b(g58236_db), .o(n_9555) );
na02f02 g55594_u0 ( .a(FE_OFN1739_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__Q), .o(n_11938) );
na02m02 g55595_u0 ( .a(FE_OFN1734_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__Q), .o(n_11937) );
na02f02 g55596_u0 ( .a(FE_OFN1757_n_12681), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__Q), .o(n_11814) );
na02f02 g55597_u0 ( .a(FE_OFN1574_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__Q), .o(n_12227) );
na02f02 TIMEBOOST_cell_41304 ( .a(TIMEBOOST_net_12890), .b(g57593_sb), .o(n_11161) );
na02s02 TIMEBOOST_cell_37528 ( .a(TIMEBOOST_net_11002), .b(FE_OFN2257_n_8060), .o(TIMEBOOST_net_4096) );
na02s02 TIMEBOOST_cell_43184 ( .a(TIMEBOOST_net_13830), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_12080) );
na02f02 g55601_u0 ( .a(FE_OFN1761_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__Q), .o(n_11934) );
na02f02 TIMEBOOST_cell_41394 ( .a(TIMEBOOST_net_12935), .b(g57370_sb), .o(TIMEBOOST_net_11642) );
na02f02 g55603_u0 ( .a(FE_OFN1740_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__Q), .o(n_11933) );
na02f02 g55604_u0 ( .a(FE_OFN1734_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__Q), .o(n_11932) );
na02f02 TIMEBOOST_cell_41198 ( .a(TIMEBOOST_net_12837), .b(g57553_sb), .o(n_10807) );
na02f01 g55606_u0 ( .a(n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__Q), .o(n_12224) );
na02s01 TIMEBOOST_cell_37303 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__22__Q), .b(n_3749), .o(TIMEBOOST_net_10890) );
na02f02 TIMEBOOST_cell_41396 ( .a(TIMEBOOST_net_12936), .b(g57538_sb), .o(n_10311) );
in01s01 TIMEBOOST_cell_45939 ( .a(wbm_dat_i_28_), .o(TIMEBOOST_net_15246) );
na02s02 g55610_u0 ( .a(FE_OFN1733_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__Q), .o(n_11930) );
na02f02 g55611_u0 ( .a(n_12010), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__Q), .o(n_11929) );
na02f02 g55612_u0 ( .a(FE_OFN1746_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__Q), .o(n_12222) );
na02s01 TIMEBOOST_cell_31812 ( .a(configuration_wb_err_data_592), .b(parchk_pci_ad_out_in_1189), .o(TIMEBOOST_net_9817) );
na02s02 TIMEBOOST_cell_43185 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__Q), .b(n_4386), .o(TIMEBOOST_net_13831) );
na02f02 TIMEBOOST_cell_41312 ( .a(TIMEBOOST_net_12894), .b(g57488_sb), .o(n_11249) );
na02f02 g55616_u0 ( .a(FE_OFN1581_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__Q), .o(n_11927) );
no02f02 g55617_u0 ( .a(FE_OCP_RBN2291_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__358), .o(n_12220) );
na02s02 TIMEBOOST_cell_45783 ( .a(n_1883), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__Q), .o(TIMEBOOST_net_15130) );
na02m02 g55619_u0 ( .a(FE_OFN1736_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q), .o(n_11925) );
na02f02 g55620_u0 ( .a(n_11977), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q), .o(n_11924) );
na02f02 TIMEBOOST_cell_41172 ( .a(TIMEBOOST_net_12824), .b(g57100_sb), .o(n_11647) );
na02s02 TIMEBOOST_cell_41850 ( .a(TIMEBOOST_net_13163), .b(FE_OFN260_n_9860), .o(n_9721) );
no02f04 g55623_u0 ( .a(FE_OCP_RBN2291_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__359), .o(n_12451) );
na02s02 TIMEBOOST_cell_41888 ( .a(TIMEBOOST_net_13182), .b(TIMEBOOST_net_4265), .o(TIMEBOOST_net_4512) );
na02s02 TIMEBOOST_cell_31727 ( .a(TIMEBOOST_net_9774), .b(FE_OFN262_n_9851), .o(n_9580) );
na02f02 g55626_u0 ( .a(FE_OFN1581_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__Q), .o(n_11923) );
na02f02 TIMEBOOST_cell_41314 ( .a(TIMEBOOST_net_12895), .b(g57455_sb), .o(n_11279) );
na02f02 g55628_u0 ( .a(n_11977), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__Q), .o(n_11921) );
na02f02 TIMEBOOST_cell_41174 ( .a(TIMEBOOST_net_12825), .b(g57420_sb), .o(n_11318) );
na03s02 TIMEBOOST_cell_34470 ( .a(pci_target_unit_wishbone_master_bc_register_reg_1__Q), .b(g52591_sb), .c(TIMEBOOST_net_880), .o(n_14686) );
na02f02 g55631_u0 ( .a(FE_OFN1733_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__Q), .o(n_11920) );
na02m02 TIMEBOOST_cell_43741 ( .a(n_9827), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__Q), .o(TIMEBOOST_net_14109) );
no02f04 g55633_u0 ( .a(n_12453), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__243), .o(n_12450) );
na02s01 TIMEBOOST_cell_30781 ( .a(TIMEBOOST_net_9301), .b(FE_OFN989_n_574), .o(TIMEBOOST_net_3279) );
na03f02 TIMEBOOST_cell_35997 ( .a(TIMEBOOST_net_10113), .b(n_13617), .c(g54485_sb), .o(n_13614) );
no02f02 g55636_u0 ( .a(FE_OCP_RBN2291_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__360), .o(n_12215) );
na02s01 TIMEBOOST_cell_9749 ( .a(TIMEBOOST_net_1441), .b(g65868_db), .o(n_2054) );
na02s01 TIMEBOOST_cell_9747 ( .a(TIMEBOOST_net_1440), .b(g65816_db), .o(n_1900) );
na02s01 TIMEBOOST_cell_42655 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__Q), .b(pci_target_unit_fifos_pcir_data_in_188), .o(TIMEBOOST_net_13566) );
na02f02 g55641_u0 ( .a(n_12010), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__Q), .o(n_11916) );
na02s01 TIMEBOOST_cell_43288 ( .a(TIMEBOOST_net_13882), .b(g62042_sb), .o(n_7771) );
no02f04 g55643_u0 ( .a(FE_OCP_RBN2293_FE_OFN1581_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13_), .o(n_12212) );
na02f02 g55644_u0 ( .a(FE_OCPN1825_n_12030), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__Q), .o(n_11915) );
na02f02 g55645_u0 ( .a(FE_OFN1564_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__Q), .o(n_11914) );
na02s02 g55646_u0 ( .a(FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__Q), .o(n_11913) );
na02f02 g55647_u0 ( .a(FE_OFN1556_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__Q), .o(n_11912) );
na02s01 TIMEBOOST_cell_9745 ( .a(TIMEBOOST_net_1439), .b(g65814_db), .o(n_2032) );
na02m02 TIMEBOOST_cell_43678 ( .a(TIMEBOOST_net_14077), .b(g58631_db), .o(n_8850) );
na02s02 TIMEBOOST_cell_37530 ( .a(TIMEBOOST_net_11003), .b(FE_OFN712_n_8140), .o(TIMEBOOST_net_4161) );
na02f02 g55651_u0 ( .a(FE_OFN1566_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__Q), .o(n_11910) );
na02f02 g55652_u0 ( .a(FE_OFN1762_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__Q), .o(n_16629) );
na02f02 TIMEBOOST_cell_41398 ( .a(TIMEBOOST_net_12937), .b(g57443_sb), .o(n_11290) );
na02f02 g55654_u0 ( .a(n_12228), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__Q), .o(n_12208) );
na02f02 g55655_u0 ( .a(FE_OFN1749_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__Q), .o(n_12207) );
na02f02 g55656_u0 ( .a(FE_OFN1741_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__Q), .o(n_12206) );
na02f02 g55657_u0 ( .a(FE_OFN1735_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__Q), .o(n_11908) );
na02f02 g55658_u0 ( .a(FE_OFN1757_n_12681), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__Q), .o(n_11806) );
na02s01 TIMEBOOST_cell_30963 ( .a(TIMEBOOST_net_9392), .b(g64918_sb), .o(n_3685) );
na02f02 g55660_u0 ( .a(FE_OFN2202_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q), .o(n_11907) );
na02m02 TIMEBOOST_cell_41597 ( .a(wbu_sel_in), .b(wishbone_slave_unit_fifos_wbr_be_in), .o(TIMEBOOST_net_13037) );
na02m02 TIMEBOOST_cell_30785 ( .a(n_2229), .b(TIMEBOOST_net_9303), .o(TIMEBOOST_net_144) );
na02s01 TIMEBOOST_cell_31810 ( .a(configuration_wb_err_cs_bit_568), .b(parchk_pci_cbe_out_in_1202), .o(TIMEBOOST_net_9816) );
na02s01 TIMEBOOST_cell_43186 ( .a(TIMEBOOST_net_13831), .b(FE_OFN1268_n_4095), .o(TIMEBOOST_net_11545) );
na02f02 g55665_u0 ( .a(FE_OFN1741_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__Q), .o(n_12203) );
na02f02 g55666_u0 ( .a(FE_OFN1735_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__Q), .o(n_11903) );
na02f02 g55667_u0 ( .a(FE_OFN1757_n_12681), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__Q), .o(n_11805) );
na02f02 g55668_u0 ( .a(n_12228), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__Q), .o(n_12202) );
na02f02 g55669_u0 ( .a(FE_OFN1749_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__Q), .o(n_12201) );
na03s02 TIMEBOOST_cell_34471 ( .a(pci_target_unit_wishbone_master_bc_register_reg_2__Q), .b(g52592_sb), .c(TIMEBOOST_net_881), .o(n_14685) );
na02s01 TIMEBOOST_cell_41851 ( .a(g62858_sb), .b(g62858_db), .o(TIMEBOOST_net_13164) );
na02f02 g55672_u0 ( .a(n_11977), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__Q), .o(n_11900) );
na02f02 TIMEBOOST_cell_41176 ( .a(TIMEBOOST_net_12826), .b(g57513_sb), .o(n_11229) );
na02s02 TIMEBOOST_cell_37302 ( .a(TIMEBOOST_net_10889), .b(FE_OFN640_n_4669), .o(TIMEBOOST_net_3652) );
no02f02 g55675_u0 ( .a(FE_OCP_RBN2291_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__363), .o(n_12449) );
na02f02 TIMEBOOST_cell_41316 ( .a(TIMEBOOST_net_12896), .b(g57156_sb), .o(n_10462) );
na02f02 g55677_u0 ( .a(FE_OFN1584_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q), .o(n_11898) );
na02s02 TIMEBOOST_cell_37532 ( .a(TIMEBOOST_net_11004), .b(FE_OFN2257_n_8060), .o(TIMEBOOST_net_4131) );
na02s02 TIMEBOOST_cell_43187 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__Q), .b(n_3624), .o(TIMEBOOST_net_13832) );
na02m02 g55680_u0 ( .a(FE_OFN1736_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__Q), .o(n_11897) );
na02f02 g55681_u0 ( .a(FE_OFN1741_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__Q), .o(n_12198) );
na02s01 TIMEBOOST_cell_42904 ( .a(TIMEBOOST_net_13690), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_11194) );
na02f02 g55683_u0 ( .a(n_12010), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__Q), .o(n_11896) );
na02f02 g55684_u0 ( .a(FE_OFN1747_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__Q), .o(n_12197) );
no02f02 g55685_u0 ( .a(n_12453), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__247), .o(n_12448) );
na02f02 g55686_u0 ( .a(FE_OFN1559_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__13__Q), .o(n_12196) );
na02f02 g55687_u0 ( .a(FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__Q), .o(n_12195) );
na02f02 g55688_u0 ( .a(FE_OFN1761_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__Q), .o(n_11895) );
na02f02 g55689_u0 ( .a(FE_OFN1584_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__Q), .o(n_12194) );
na03f02 TIMEBOOST_cell_34472 ( .a(FE_RN_566_0), .b(FE_RN_568_0), .c(FE_RN_567_0), .o(FE_RN_569_0) );
na02s01 TIMEBOOST_cell_43289 ( .a(TIMEBOOST_net_4773), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_13883) );
na02f02 TIMEBOOST_cell_41178 ( .a(TIMEBOOST_net_12827), .b(g57116_sb), .o(n_11630) );
na02f02 g55693_u0 ( .a(n_11977), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__Q), .o(n_11893) );
na02s01 TIMEBOOST_cell_30965 ( .a(TIMEBOOST_net_9393), .b(g64923_sb), .o(n_3682) );
no02f02 g55695_u0 ( .a(FE_OCP_RBN2292_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__365), .o(n_12447) );
na02m02 TIMEBOOST_cell_43853 ( .a(n_9457), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__Q), .o(TIMEBOOST_net_14165) );
na02s02 TIMEBOOST_cell_45008 ( .a(TIMEBOOST_net_14742), .b(g64097_db), .o(n_4058) );
no02f02 g55698_u0 ( .a(FE_OCP_RBN2286_FE_RN_494_0), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__248), .o(n_11891) );
na04f02 TIMEBOOST_cell_14750 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__Q), .b(FE_OFN1394_n_8567), .c(n_8556), .d(g58592_sb), .o(n_8906) );
na02s02 g55700_u0 ( .a(FE_OFN1734_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__Q), .o(n_11890) );
na02s01 TIMEBOOST_cell_42667 ( .a(g64096_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__22__Q), .o(TIMEBOOST_net_13572) );
na02s01 TIMEBOOST_cell_42905 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__Q), .b(FE_OFN533_n_9823), .o(TIMEBOOST_net_13691) );
na02f02 TIMEBOOST_cell_41426 ( .a(TIMEBOOST_net_12951), .b(g57217_sb), .o(n_11540) );
no02f02 g55704_u0 ( .a(n_12453), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__249), .o(n_12446) );
na02s01 TIMEBOOST_cell_45009 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__Q), .b(g64311_sb), .o(TIMEBOOST_net_14743) );
na02s01 TIMEBOOST_cell_31808 ( .a(configuration_wb_err_data_597), .b(parchk_pci_ad_out_in_1194), .o(TIMEBOOST_net_9815) );
no02f02 g55707_u0 ( .a(n_11762), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__522), .o(n_12186) );
na02s01 TIMEBOOST_cell_41852 ( .a(TIMEBOOST_net_13164), .b(n_3993), .o(n_5251) );
na02f02 TIMEBOOST_cell_43854 ( .a(TIMEBOOST_net_14165), .b(FE_OFN1409_n_8567), .o(TIMEBOOST_net_12826) );
na02s01 TIMEBOOST_cell_37305 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__Q), .b(n_3783), .o(TIMEBOOST_net_10891) );
na02m02 TIMEBOOST_cell_44507 ( .a(n_9110), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__Q), .o(TIMEBOOST_net_14492) );
na03f02 TIMEBOOST_cell_35999 ( .a(TIMEBOOST_net_10111), .b(n_13617), .c(g54487_sb), .o(n_13611) );
na02s01 TIMEBOOST_cell_42685 ( .a(pci_target_unit_fifos_pciw_addr_data_in_141), .b(g64184_sb), .o(TIMEBOOST_net_13581) );
na02m02 g55714_u0 ( .a(FE_OFN1741_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__Q), .o(n_11887) );
na02s01 TIMEBOOST_cell_37304 ( .a(TIMEBOOST_net_10890), .b(FE_OFN615_n_4501), .o(TIMEBOOST_net_9473) );
na02f02 TIMEBOOST_cell_41428 ( .a(TIMEBOOST_net_12952), .b(g57451_sb), .o(n_11283) );
no02f02 g55717_u0 ( .a(FE_OCPN1834_n_11884), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__484), .o(n_11885) );
ao22f02 g55720_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__Q), .c(FE_OFN1466_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__Q), .o(n_11157) );
ao22f02 g55721_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__Q), .c(FE_OFN1444_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__Q), .o(n_17016) );
ao22f02 g55722_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__Q), .o(n_11155) );
ao22f02 g55723_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__Q), .o(n_11153) );
ao22f02 g55725_u0 ( .a(FE_OFN1461_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__Q), .o(n_11793) );
ao22f02 g55726_u0 ( .a(FE_OFN1478_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__Q), .c(FE_OFN1449_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__Q), .o(n_11152) );
ao22f02 g55727_u0 ( .a(FE_OFN1431_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__Q), .c(FE_OFN1444_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__Q), .o(n_11149) );
ao22f02 g55728_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__Q), .o(n_11148) );
ao22f02 g55729_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__Q), .o(n_11147) );
ao22f02 g55730_u0 ( .a(FE_OFN1477_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__Q), .c(FE_OFN1449_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__Q), .o(n_11146) );
ao22f02 g55731_u0 ( .a(FE_OFN1461_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__Q), .o(n_11145) );
ao22f02 g55732_u0 ( .a(FE_OFN1478_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__Q), .c(FE_OFN2193_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__Q), .o(n_11144) );
ao22f02 g55733_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__Q), .o(n_11143) );
ao22f02 g55734_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__Q), .o(n_11142) );
ao22f02 g55735_u0 ( .a(FE_OFN1478_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__Q), .c(FE_OFN2193_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__Q), .o(n_11140) );
ao22f02 g55738_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__Q), .o(n_11136) );
ao22f02 g55739_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__Q), .o(n_11135) );
ao22f02 g55740_u0 ( .a(FE_OCP_RBN2010_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__Q), .o(n_11134) );
ao22f02 g55741_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__Q), .o(n_11132) );
ao22f02 g55742_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__Q), .o(n_11131) );
ao22f02 g55744_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__Q), .c(FE_OFN1444_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__Q), .o(n_11792) );
ao22f02 g55745_u0 ( .a(FE_OFN1477_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__Q), .c(FE_OFN1449_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__Q), .o(n_11130) );
ao22f02 g55746_u0 ( .a(FE_OFN1461_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__Q), .o(n_11791) );
ao22f02 g55747_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__Q), .c(FE_OFN1466_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__Q), .o(n_16582) );
ao22f02 g55748_u0 ( .a(FE_OFN1462_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__Q), .c(FE_OFN1457_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__Q), .o(n_11129) );
ao22f02 g55749_u0 ( .a(FE_OFN1478_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__Q), .c(FE_OFN2193_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__Q), .o(n_16581) );
ao22f02 g55750_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__Q), .o(n_11126) );
ao22f02 g55751_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__Q), .c(FE_OFN1466_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__Q), .o(n_10788) );
ao22f02 g55752_u0 ( .a(FE_OFN1462_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__Q), .c(FE_OFN1457_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__Q), .o(n_11124) );
ao22f02 g55753_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__Q), .o(n_11123) );
ao22f02 g55754_u0 ( .a(FE_OFN1478_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__Q), .c(FE_OFN2193_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__Q), .o(n_11122) );
ao22f02 g55755_u0 ( .a(FE_OFN1462_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__Q), .c(FE_OFN1457_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__Q), .o(n_11121) );
ao22f02 g55756_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__Q), .c(FE_OFN1466_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__Q), .o(n_11120) );
ao22f02 g55757_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__Q), .o(n_11119) );
ao22f02 g55759_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__Q), .o(n_16584) );
ao22f02 g55760_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__Q), .o(n_11115) );
ao22f02 g55761_u0 ( .a(FE_OFN1477_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__Q), .c(FE_OFN1450_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__Q), .o(n_16583) );
ao22f02 g55763_u0 ( .a(FE_OFN1477_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__Q), .c(FE_OFN1450_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__Q), .o(n_11111) );
ao22f02 g55764_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__Q), .o(n_11110) );
ao22f02 g55765_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__Q), .c(n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__Q), .o(n_11109) );
ao22f02 g55766_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__Q), .o(n_11108) );
ao22f02 g55767_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__Q), .o(n_11790) );
ao22f02 g55771_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__Q), .c(FE_OFN2193_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__Q), .o(n_11102) );
ao22f02 g55772_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__Q), .o(n_11101) );
ao22f02 g55773_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__Q), .c(FE_OFN1466_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__Q), .o(n_11100) );
ao22f02 g55774_u0 ( .a(FE_OFN1462_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__Q), .c(FE_OFN1457_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__Q), .o(n_11099) );
ao22f02 g55775_u0 ( .a(FE_OFN1431_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__Q), .c(FE_OFN1444_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__Q), .o(n_11788) );
ao22f02 g55776_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q), .c(FE_OFN1449_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__22__Q), .o(n_11097) );
ao22f02 g55777_u0 ( .a(FE_OFN1461_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__Q), .o(n_11096) );
ao22f02 g55778_u0 ( .a(FE_OFN1716_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__Q), .o(n_11095) );
ao22f02 g55779_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__Q), .o(n_11094) );
ao22f02 g55781_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__Q), .o(n_11092) );
ao22f02 g55783_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__Q), .o(n_10785) );
ao22f02 g55784_u0 ( .a(FE_OFN2208_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__Q), .c(FE_OFN1455_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__Q), .o(n_11090) );
ao22f02 g55785_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__Q), .o(n_11089) );
ao22s02 g55786_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__Q), .o(n_11088) );
ao22f02 g55787_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__Q), .c(FE_OFN1466_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__Q), .o(n_10784) );
ao22f02 g55788_u0 ( .a(FE_OFN1461_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__Q), .o(n_11786) );
ao22f02 g55789_u0 ( .a(FE_OFN1478_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__Q), .c(FE_OFN2193_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__Q), .o(n_11087) );
ao22f02 g55790_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__Q), .o(n_11086) );
ao22f02 g55791_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__Q), .o(n_11784) );
ao22f02 g55792_u0 ( .a(FE_OFN2208_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__Q), .c(FE_OFN1455_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__Q), .o(n_11085) );
ao22f02 g55793_u0 ( .a(FE_OFN1477_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__Q), .c(FE_OFN1450_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__Q), .o(n_11084) );
ao22f02 g55794_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__Q), .o(n_11083) );
ao22f02 g55795_u0 ( .a(FE_OCP_RBN2010_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__Q), .o(n_16586) );
ao22f02 g55796_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__Q), .o(n_11081) );
ao22f02 g55797_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__Q), .o(n_16585) );
ao22f02 g55798_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__Q), .o(n_11079) );
ao22f02 g55799_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__Q), .o(n_11078) );
ao22f02 g55801_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__Q), .o(n_11076) );
ao22f02 g55802_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__Q), .o(n_11075) );
ao22f02 g55803_u0 ( .a(FE_OFN2208_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__Q), .c(FE_OFN1455_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__Q), .o(n_11783) );
ao22f02 g55804_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__Q), .o(n_11782) );
ao22f02 g55806_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__Q), .o(n_11072) );
ao22f02 g55807_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__Q), .o(n_11781) );
ao22f02 g55808_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__Q), .o(n_11071) );
ao22f02 g55809_u0 ( .a(FE_OFN2208_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__Q), .c(FE_OFN1455_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__Q), .o(n_11070) );
ao22f02 g55810_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__Q), .o(n_11069) );
ao22f02 g55811_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__Q), .o(n_10782) );
ao22f02 g55812_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__Q), .o(n_11067) );
ao22f02 g55813_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__Q), .o(n_11066) );
ao22f02 g55814_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__Q), .o(n_11065) );
ao22f02 g55815_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__Q), .o(n_11780) );
ao22f02 g55816_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__Q), .o(n_11778) );
ao22f02 g55817_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__Q), .o(n_11064) );
ao22f02 g55818_u0 ( .a(FE_OCP_RBN2010_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__Q), .o(n_11063) );
ao22f02 g55820_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__Q), .o(n_11062) );
ao22f02 g55821_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__Q), .o(n_11061) );
ao22f02 g55822_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__Q), .o(n_11060) );
ao22f02 g55823_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__Q), .o(n_11776) );
ao22f02 g55826_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__Q), .o(n_11057) );
ao22f02 g55827_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__Q), .o(n_11056) );
ao22f02 g55828_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__Q), .o(n_11055) );
ao22f02 g55829_u0 ( .a(FE_OFN2208_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__Q), .c(FE_OFN1455_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__Q), .o(n_11054) );
ao22f02 g55830_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__Q), .o(n_11053) );
ao22f02 g55832_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__Q), .o(n_11050) );
ao22f02 g55833_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__Q), .o(n_11049) );
ao22f02 g55835_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__Q), .o(n_11775) );
ao22f02 g55836_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__Q), .o(n_11047) );
ao22f02 g55837_u0 ( .a(FE_OCP_RBN2010_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__Q), .o(n_11046) );
ao22f02 g55838_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__Q), .c(FE_OFN2195_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__Q), .o(n_11044) );
ao22f02 g55839_u0 ( .a(FE_OCP_RBN2010_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__Q), .o(n_10781) );
ao22f02 g55840_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__Q), .o(n_11043) );
ao22f02 g55841_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__Q), .o(n_11042) );
ao22f02 g55842_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__Q), .o(n_11774) );
ao22f02 g55843_u0 ( .a(FE_OFN1431_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__Q), .c(FE_OFN1444_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__Q), .o(n_11773) );
ao22f02 g55844_u0 ( .a(FE_OFN1716_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__Q), .o(n_11041) );
ao22f02 g55845_u0 ( .a(FE_OFN1461_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__Q), .o(n_11040) );
ao22m02 g55846_u0 ( .a(FE_OFN1477_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__8__Q), .c(FE_OFN1449_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q), .o(n_11039) );
ao22f02 g55847_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__Q), .c(FE_OFN2196_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__Q), .o(n_11038) );
ao22m02 g55848_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__Q), .o(n_11037) );
ao22f02 g55849_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__Q), .o(n_11036) );
ao22f02 g55850_u0 ( .a(FE_OFN1462_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__Q), .c(FE_OFN1457_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__Q), .o(n_11034) );
in01f02 g55851_u0 ( .a(n_9177), .o(g55851_sb) );
na02s02 TIMEBOOST_cell_43599 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__Q), .b(n_3647), .o(TIMEBOOST_net_14038) );
na02s01 TIMEBOOST_cell_37307 ( .a(n_3744), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__Q), .o(TIMEBOOST_net_10892) );
na02s01 TIMEBOOST_cell_37306 ( .a(TIMEBOOST_net_10891), .b(FE_OFN1659_n_4490), .o(TIMEBOOST_net_9461) );
in01f02 g55852_u0 ( .a(n_9177), .o(g55852_sb) );
na02f02 TIMEBOOST_cell_32571 ( .a(FE_OCPN1825_n_12030), .b(TIMEBOOST_net_10196), .o(TIMEBOOST_net_6562) );
na02s01 TIMEBOOST_cell_37309 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__Q), .b(n_3783), .o(TIMEBOOST_net_10893) );
na02s01 TIMEBOOST_cell_37308 ( .a(TIMEBOOST_net_10892), .b(FE_OFN640_n_4669), .o(TIMEBOOST_net_3625) );
in01f02 g55853_u0 ( .a(n_9177), .o(g55853_sb) );
na03s02 TIMEBOOST_cell_34279 ( .a(TIMEBOOST_net_9804), .b(FE_OFN1173_n_5592), .c(g62086_sb), .o(n_5622) );
na02m02 TIMEBOOST_cell_44361 ( .a(n_9735), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__Q), .o(TIMEBOOST_net_14419) );
no02s02 g56438_u0 ( .a(n_4697), .b(FE_OFN778_n_4152), .o(n_5744) );
no02m02 g56439_u0 ( .a(n_4800), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8579) );
in01f02 g56450_u0 ( .a(n_9338), .o(n_10780) );
na02f02 g56451_u0 ( .a(FE_OCP_RBN2226_g75174_p), .b(n_16313), .o(n_9338) );
na02f02 g56461_u0 ( .a(n_16334), .b(n_16445), .o(n_10273) );
in01f04 g56466_u0 ( .a(n_12381), .o(n_12357) );
in01f08 g56468_u0 ( .a(n_12099), .o(n_12381) );
in01f04 g56469_u0 ( .a(n_10270), .o(n_12099) );
na02f02 g56470_u0 ( .a(n_10258), .b(n_16334), .o(n_10270) );
in01f04 g56471_u0 ( .a(FE_OCPN1890_n_16553), .o(n_11831) );
in01f04 g56472_u0 ( .a(FE_OCPN1890_n_16553), .o(n_11823) );
in01f02 g56473_u0 ( .a(n_16553), .o(n_12681) );
na02f02 g56485_u0 ( .a(n_16552), .b(n_16445), .o(n_10268) );
in01f04 g56491_u0 ( .a(FE_OCPN1907_n_11767), .o(n_12362) );
in01f02 g56509_u0 ( .a(n_10261), .o(n_12004) );
na02f02 g56510_u0 ( .a(FE_OCP_RBN2226_g75174_p), .b(FE_OCP_RBN2282_g74996_p), .o(n_10261) );
in01f02 g56516_u0 ( .a(FE_OFN1584_n_12306), .o(n_16587) );
in01f02 g56517_u0 ( .a(FE_OFN1579_n_12306), .o(n_11762) );
na02f02 g56522_u0 ( .a(n_10258), .b(n_16313), .o(n_10259) );
in01f02 g56529_u0 ( .a(n_9336), .o(n_12502) );
na02f02 g56530_u0 ( .a(n_16313), .b(n_16364), .o(n_9336) );
in01f02 g56554_u0 ( .a(n_10254), .o(n_12104) );
na02f02 g56555_u0 ( .a(FE_OCP_RBN2281_g74996_p), .b(n_16445), .o(n_10254) );
in01f04 g56556_u0 ( .a(FE_OFN1739_n_11019), .o(n_12293) );
in01f02 g56564_u0 ( .a(n_10252), .o(n_11019) );
na02f02 g56565_u0 ( .a(n_16552), .b(n_16364), .o(n_10252) );
in01f04 g56566_u0 ( .a(n_11884), .o(n_12010) );
in01f02 g56567_u0 ( .a(n_11884), .o(n_11977) );
in01f04 g56568_u0 ( .a(FE_OCPN1834_n_11884), .o(n_12228) );
in01f02 g56572_u0 ( .a(n_11884), .o(n_12001) );
na02f04 g56575_u0 ( .a(n_10258), .b(FE_OCP_RBN2283_g74996_p), .o(n_11884) );
in01f08 g56577_u0 ( .a(FE_OCP_RBN2286_FE_RN_494_0), .o(n_12313) );
in01f08 g56580_u0 ( .a(n_11881), .o(n_12453) );
in01f06 g56582_u0 ( .a(FE_OCP_RBN2286_FE_RN_494_0), .o(n_11881) );
in01f02 g56598_u0 ( .a(n_10244), .o(n_12028) );
na02f02 g56599_u0 ( .a(n_10258), .b(n_16552), .o(n_10244) );
ao22f02 g56600_u0 ( .a(FE_OCPN1879_FE_OFN470_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__Q), .c(FE_OFN1528_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__Q), .o(n_16987) );
ao22f02 g56601_u0 ( .a(FE_OFN1511_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__Q), .o(n_9335) );
ao22f02 g56602_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q), .o(n_9334) );
ao22f02 g56603_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__Q), .c(FE_OCPN1872_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__Q), .o(n_16986) );
in01f02 g56604_u0 ( .a(n_10777), .o(n_11014) );
ao22f02 g56605_u0 ( .a(FE_OFN1493_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__Q), .o(n_10777) );
ao22f02 g56606_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q), .c(FE_OFN2206_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__Q), .o(n_10774) );
ao22f02 g56607_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__Q), .o(n_10771) );
ao22f02 g56608_u0 ( .a(FE_OFN2216_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__Q), .o(n_11013) );
ao22f02 g56609_u0 ( .a(FE_OFN2147_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__Q), .c(FE_OFN1523_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__Q), .o(n_11008) );
ao22f02 g56611_u0 ( .a(FE_OFN2146_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__Q), .c(FE_OFN1547_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__Q), .o(n_9331) );
ao22f02 g56612_u0 ( .a(FE_OCP_RBN1969_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__Q), .c(n_10232), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__Q), .o(n_10235) );
in01f02 g56613_u0 ( .a(n_11005), .o(n_11741) );
ao22f02 g56614_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__10__Q), .c(FE_OCPN1873_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q), .o(n_11005) );
ao22f02 g56615_u0 ( .a(n_10680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__Q), .o(n_10768) );
ao22f02 g56616_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q), .c(FE_OFN1498_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__10__Q), .o(n_10230) );
ao22f02 g56617_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__Q), .o(n_11002) );
ao22f02 g56619_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__Q), .o(n_9330) );
ao22f02 g56621_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__Q), .c(FE_OCP_RBN1932_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__Q), .o(n_9329) );
in01f02 g56622_u0 ( .a(n_10994), .o(n_11740) );
ao22f02 g56623_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__Q), .c(FE_OCPN1888_FE_OFN473_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__Q), .o(n_10994) );
ao22f02 g56624_u0 ( .a(FE_OCPN1886_FE_OFN1508_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__Q), .o(n_10221) );
ao22f02 g56625_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__Q), .c(FE_OFN1502_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__Q), .o(n_10216) );
ao22f02 g56626_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__Q), .o(n_10991) );
ao22f01 g56627_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__Q), .c(n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__Q), .o(n_16843) );
ao22f01 g56629_u0 ( .a(n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__Q), .o(n_16842) );
ao22f01 g56630_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__Q), .c(n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__Q), .o(n_9325) );
in01f02 g56631_u0 ( .a(n_10765), .o(n_10987) );
ao22f02 g56632_u0 ( .a(FE_OFN1538_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__Q), .c(FE_OCPN1915_FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__Q), .o(n_10765) );
ao22f02 g56633_u0 ( .a(FE_OFN1491_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__Q), .c(n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__Q), .o(n_10205) );
ao22f02 g56634_u0 ( .a(FE_OFN1728_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__Q), .c(FE_OCP_RBN1933_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__Q), .o(n_10202) );
ao22f01 g56635_u0 ( .a(n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__Q), .o(n_10986) );
ao22f02 g56636_u0 ( .a(FE_OFN2149_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__Q), .c(FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__Q), .o(n_10985) );
ao22f02 g56637_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__Q), .c(FE_OCP_RBN2005_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__Q), .o(n_9322) );
ao22f02 g56638_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__Q), .o(n_9321) );
ao22f02 g56639_u0 ( .a(FE_OCP_RBN1969_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__Q), .c(FE_OCPN2015_n_10195), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__Q), .o(n_10198) );
in01f02 g56640_u0 ( .a(n_10193), .o(n_10764) );
ao22f02 g56641_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__Q), .c(FE_OFN1498_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__Q), .o(n_10193) );
ao22f02 g56642_u0 ( .a(n_10680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__Q), .o(n_10763) );
ao22f02 g56644_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__Q), .o(n_10981) );
ao22f02 g56647_u0 ( .a(FE_OFN2147_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__Q), .c(FE_OFN1523_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__Q), .o(n_10183) );
in01f02 g56648_u0 ( .a(n_10755), .o(n_10978) );
ao22f02 g56650_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__Q), .c(FE_OCP_RBN2006_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__Q), .o(n_9315) );
ao22f02 g56652_u0 ( .a(n_10680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__Q), .o(n_10754) );
ao22f02 g56653_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__Q), .o(n_10977) );
ao22f02 g56654_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__Q), .c(FE_OCP_RBN2005_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__Q), .o(n_9312) );
ao22f02 g56655_u0 ( .a(FE_OCP_RBN1968_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__Q), .c(n_10185), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__Q), .o(n_10176) );
in01f02 g56658_u0 ( .a(n_10753), .o(n_10976) );
ao22f02 g56659_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__15__Q), .c(n_10693), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__15__Q), .o(n_10753) );
ao22f02 g56660_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__Q), .o(n_10750) );
ao22f02 g56661_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__Q), .c(FE_OCPN1873_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__Q), .o(n_10747) );
ao22f02 g56662_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__Q), .o(n_10744) );
ao22f02 g56663_u0 ( .a(FE_OFN1511_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__Q), .o(n_9309) );
ao22f02 g56664_u0 ( .a(n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__Q), .o(n_16849) );
ao22f02 g56665_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__Q), .c(FE_OFN2143_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__Q), .o(n_16848) );
ao22f02 g56666_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__Q), .o(n_10163) );
in01f02 g56667_u0 ( .a(n_10741), .o(n_10975) );
ao22f02 g56669_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__Q), .c(FE_OFN2206_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__Q), .o(n_10738) );
ao22f02 g56670_u0 ( .a(FE_OFN2216_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q), .o(n_10974) );
ao22f02 g56671_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__Q), .c(FE_OCP_RBN2006_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__Q), .o(n_10160) );
ao22f02 g56672_u0 ( .a(FE_OFN1508_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__Q), .o(n_9307) );
ao22f02 g56673_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__Q), .c(FE_OFN2139_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__Q), .o(n_10154) );
ao22f02 g56674_u0 ( .a(n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q), .c(FE_OFN1500_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q), .o(n_9306) );
ao22f02 g56675_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__Q), .o(n_10151) );
in01f02 g56676_u0 ( .a(n_10734), .o(n_10971) );
ao22f02 g56677_u0 ( .a(FE_OFN2149_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__Q), .c(FE_OCPN1915_FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__Q), .o(n_10734) );
ao22f02 g56678_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__Q), .o(n_10970) );
ao22f02 g56679_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__Q), .o(n_10731) );
ao22f02 g56680_u0 ( .a(FE_OCPN1892_FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__Q), .c(FE_OCP_RBN1932_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__Q), .o(n_10147) );
ao22f02 g56681_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__Q), .o(n_9305) );
ao22f02 g56683_u0 ( .a(FE_OCP_RBN1969_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__Q), .c(n_10141), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__Q), .o(n_10144) );
in01f02 g56685_u0 ( .a(n_10967), .o(n_11739) );
ao22f02 g56686_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__Q), .c(FE_OCPN1888_FE_OFN473_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__Q), .o(n_10967) );
ao22f02 g56690_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__Q), .c(FE_OCP_RBN1934_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__Q), .o(n_17051) );
ao22f02 g56691_u0 ( .a(FE_OFN1490_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__Q), .c(FE_OFN1545_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__Q), .o(n_9301) );
ao22f02 g56692_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__Q), .o(n_17050) );
ao22f02 g56693_u0 ( .a(FE_OFN1538_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__Q), .c(FE_OCPN1915_FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__Q), .o(n_10134) );
in01f02 g56694_u0 ( .a(n_10715), .o(n_10963) );
ao22f02 g56695_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__Q), .o(n_10715) );
ao22f02 g56696_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__Q), .c(FE_OFN1502_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__Q), .o(n_10131) );
ao22f02 g56697_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__Q), .o(n_10711) );
ao22f02 g56698_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__Q), .o(n_10708) );
ao22f02 g56699_u0 ( .a(FE_OCPN1879_FE_OFN470_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__Q), .c(FE_OFN1528_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__Q), .o(n_10127) );
ao22f02 g56700_u0 ( .a(n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__Q), .o(n_9299) );
ao22f02 g56701_u0 ( .a(FE_OFN1511_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__Q), .o(n_9298) );
ao22f02 g56702_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__Q), .c(FE_OCPN1872_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__Q), .o(n_10124) );
in01f02 g56703_u0 ( .a(n_10705), .o(n_10962) );
ao22f02 g56704_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__Q), .o(n_10705) );
ao22f02 g56706_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__Q), .c(FE_OFN2206_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__Q), .o(n_10699) );
ao22f02 g56707_u0 ( .a(FE_OFN2216_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q), .o(n_10961) );
ao22f02 g56708_u0 ( .a(FE_OFN2147_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__Q), .c(FE_OFN1523_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__Q), .o(n_10956) );
ao22f02 g56710_u0 ( .a(FE_OCP_RBN1968_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__Q), .c(n_10232), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__Q), .o(n_10120) );
ao22f02 g56711_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q), .c(FE_OCP_RBN2005_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__Q), .o(n_9296) );
in01f02 g56712_u0 ( .a(n_10696), .o(n_10952) );
ao22f02 g56713_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__Q), .c(n_10693), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__Q), .o(n_10696) );
ao22f02 g56715_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__Q), .c(FE_OCPN1873_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__Q), .o(n_10691) );
ao22f02 g56716_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__Q), .o(n_10688) );
ao22f02 g56717_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__Q), .o(n_10116) );
ao22f02 g56718_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__Q), .o(n_10112) );
ao22f02 g56719_u0 ( .a(n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__Q), .c(FE_OFN1501_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__Q), .o(n_9295) );
ao22f02 g56720_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q), .c(FE_OFN1723_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__Q), .o(n_9294) );
in01f02 g56721_u0 ( .a(n_10947), .o(n_11738) );
ao22f02 g56723_u0 ( .a(FE_OFN1728_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__Q), .c(FE_OCP_RBN1933_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__Q), .o(n_10109) );
ao22f02 g56724_u0 ( .a(FE_OFN1539_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__Q), .c(FE_OFN1521_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__Q), .o(n_10685) );
ao22f02 g56725_u0 ( .a(FE_OFN1490_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__Q), .o(n_10105) );
ao22f02 g56726_u0 ( .a(FE_OFN2148_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__Q), .c(FE_OFN1523_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__Q), .o(n_10944) );
ao22m02 g56727_u0 ( .a(FE_OCP_RBN1969_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__Q), .c(n_10185), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__Q), .o(n_10102) );
ao22f02 g56728_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__Q), .c(FE_OCP_RBN2005_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__Q), .o(n_9293) );
ao22f02 g56729_u0 ( .a(FE_OFN2146_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__Q), .c(FE_OFN1547_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__Q), .o(n_9290) );
in01f02 g56730_u0 ( .a(n_10682), .o(n_10943) );
ao22f02 g56731_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__22__Q), .c(FE_OCPN1888_FE_OFN473_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__22__Q), .o(n_10682) );
ao22f02 g56732_u0 ( .a(n_10680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__Q), .o(n_10681) );
ao22f02 g56733_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__Q), .c(n_15568), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__Q), .o(n_10679) );
ao22f02 g56734_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__Q), .o(n_10676) );
ao22f02 g56735_u0 ( .a(FE_OFN2149_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__Q), .c(FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__Q), .o(n_10942) );
ao22f02 g56737_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__Q), .c(n_10141), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__Q), .o(n_10099) );
ao22f02 g56738_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__Q), .c(FE_OCP_RBN1932_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__Q), .o(n_9286) );
in01f02 g56739_u0 ( .a(n_10939), .o(n_17042) );
ao22f02 g56740_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__Q), .o(n_10939) );
ao22f02 g56741_u0 ( .a(FE_OCPN1886_FE_OFN1508_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__Q), .o(n_10096) );
ao22f02 g56742_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__Q), .c(n_15568), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__Q), .o(n_10675) );
ao22f02 g56743_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__Q), .o(n_10672) );
ao22f02 g56744_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__Q), .c(FE_OCP_RBN1932_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__Q), .o(n_9285) );
ao22f02 g56745_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__Q), .o(n_9284) );
ao22f02 g56746_u0 ( .a(FE_OFN2149_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__Q), .c(FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__Q), .o(n_10093) );
ao22f02 g56747_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__Q), .c(FE_OCPN2015_n_10195), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__Q), .o(n_10090) );
in01f02 g56748_u0 ( .a(n_10087), .o(n_10669) );
ao22f02 g56749_u0 ( .a(FE_OCPN1886_FE_OFN1508_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__Q), .o(n_10087) );
ao22f01 g56753_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__Q), .o(n_10084) );
ao22f01 g56754_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__Q), .o(n_10081) );
ao22f02 g56755_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__Q), .o(n_9283) );
ao22f02 g56756_u0 ( .a(n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__Q), .c(FE_OFN1500_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__Q), .o(n_9280) );
in01f02 g56757_u0 ( .a(n_10662), .o(n_10932) );
ao22f02 g56758_u0 ( .a(FE_OFN1538_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__Q), .c(FE_OCPN1915_FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__Q), .o(n_10662) );
ao22f02 g56759_u0 ( .a(FE_OFN1728_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__Q), .c(FE_OCP_RBN1933_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__Q), .o(n_10661) );
ao22f02 g56761_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__Q), .c(n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__Q), .o(n_10660) );
ao22f02 g56762_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__Q), .o(n_9277) );
ao22f02 g56764_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__Q), .c(FE_OCP_RBN1932_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__Q), .o(n_9276) );
in01f02 g56766_u0 ( .a(n_10927), .o(n_11736) );
ao22f02 g56767_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__Q), .o(n_10927) );
ao22f02 g56768_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__Q), .c(FE_OFN1502_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__Q), .o(n_10075) );
ao22f02 g56769_u0 ( .a(n_10680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__Q), .o(n_10659) );
ao22f02 g56770_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__Q), .c(FE_OCPN1888_FE_OFN473_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__Q), .o(n_10656) );
ao22f02 g56772_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__Q), .o(n_9274) );
ao22f02 g56773_u0 ( .a(FE_OCP_RBN1969_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__Q), .c(n_10141), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__Q), .o(n_17043) );
ao22f02 g56774_u0 ( .a(FE_OFN2149_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__Q), .c(FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__Q), .o(n_10069) );
in01f02 g56775_u0 ( .a(n_10653), .o(n_10923) );
ao22f02 g56776_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__Q), .c(FE_OCPN1888_FE_OFN473_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__Q), .o(n_10653) );
ao22f02 g56777_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__Q), .o(n_10650) );
ao22f02 g56778_u0 ( .a(n_10680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__Q), .o(n_10647) );
ao22f02 g56779_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q), .c(n_15568), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q), .o(n_10644) );
ao22f02 g56780_u0 ( .a(FE_OFN2146_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__Q), .c(FE_OFN1547_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__Q), .o(n_9272) );
ao22f02 g56781_u0 ( .a(FE_OFN2147_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__Q), .c(FE_OFN1523_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__Q), .o(n_10641) );
ao22f02 g56782_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__Q), .c(FE_OCP_RBN2005_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__Q), .o(n_9271) );
ao22f02 g56783_u0 ( .a(FE_OCP_RBN1968_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__Q), .c(n_10232), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__Q), .o(n_10066) );
in01f02 g56784_u0 ( .a(n_10063), .o(n_10638) );
ao22f02 g56785_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__Q), .o(n_10063) );
ao22f02 g56786_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__Q), .o(n_10637) );
ao22f02 g56787_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q), .c(FE_OFN1498_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q), .o(n_10060) );
ao22f02 g56788_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__Q), .c(FE_OCPN1863_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__Q), .o(n_10634) );
ao22f02 g56789_u0 ( .a(FE_OCP_RBN1969_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__Q), .c(n_10185), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__Q), .o(n_10057) );
ao22f02 g56790_u0 ( .a(FE_OFN2146_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q), .c(FE_OFN1547_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__29__Q), .o(n_9270) );
in01f02 g56792_u0 ( .a(n_10051), .o(n_10631) );
ao22f02 g56793_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__Q), .o(n_10051) );
ao22f02 g56794_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__Q), .c(FE_OCP_RBN2005_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__Q), .o(n_9269) );
ao22f02 g56795_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__Q), .c(FE_OCPN1863_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__Q), .o(n_10922) );
ao22f02 g56796_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__Q), .o(n_10630) );
ao22f02 g56797_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__29__Q), .c(n_15568), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q), .o(n_10627) );
ao22f02 g56798_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__Q), .c(FE_OFN1723_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__Q), .o(n_16835) );
ao22f02 g56799_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q), .o(n_10048) );
in01f02 g56801_u0 ( .a(n_10624), .o(n_10919) );
ao22f02 g56802_u0 ( .a(FE_OFN1539_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__Q), .c(FE_OFN1521_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__Q), .o(n_10624) );
ao22f02 g56804_u0 ( .a(FE_OFN1728_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__Q), .c(FE_OCP_RBN1933_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__Q), .o(n_10041) );
ao22f02 g56805_u0 ( .a(FE_OFN1490_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__Q), .c(n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__Q), .o(n_10038) );
ao22f02 g56806_u0 ( .a(FE_OFN1535_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__Q), .o(n_10918) );
ao22f02 g56807_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__Q), .o(n_10035) );
ao22f02 g56808_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__Q), .c(FE_OFN2140_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__Q), .o(n_10032) );
ao22f02 g56809_u0 ( .a(n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__Q), .o(n_9262) );
in01f02 g56810_u0 ( .a(n_10622), .o(n_10917) );
ao22f02 g56811_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__Q), .o(n_10622) );
ao22f02 g56812_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__Q), .o(n_9261) );
ao22f02 g56813_u0 ( .a(FE_OFN1539_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__Q), .c(FE_OFN1521_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__Q), .o(n_10617) );
ao22f02 g56814_u0 ( .a(FE_OFN1490_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__Q), .o(n_10029) );
ao22f02 g56815_u0 ( .a(FE_OFN1535_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__Q), .o(n_10916) );
ao22f02 g56816_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__Q), .c(FE_OCP_RBN2006_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__Q), .o(n_9260) );
ao22f02 g56818_u0 ( .a(FE_OFN2147_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__Q), .c(FE_OFN1523_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__Q), .o(n_10614) );
in01f02 g56820_u0 ( .a(n_10611), .o(n_10913) );
ao22f02 g56821_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__Q), .o(n_10611) );
ao22f02 g56822_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__Q), .o(n_11735) );
ao22f02 g56823_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q), .c(FE_OCPN1863_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__Q), .o(n_10912) );
ao22f02 g56824_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__31__Q), .c(FE_OFN1498_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__31__Q), .o(n_10608) );
ao22f02 g56825_u0 ( .a(FE_OFN1511_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__Q), .o(n_10020) );
ao22f02 g56826_u0 ( .a(FE_OCPN1879_FE_OFN470_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__Q), .c(FE_OFN1528_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__Q), .o(n_10605) );
ao22f02 g56827_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__Q), .o(n_10017) );
ao22f02 g56828_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__Q), .c(FE_OCPN1872_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__Q), .o(n_10602) );
in01f02 g56829_u0 ( .a(n_10909), .o(n_11734) );
ao22f02 g56830_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__Q), .c(FE_OFN2207_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__Q), .o(n_10909) );
ao22f02 g56831_u0 ( .a(FE_OFN1493_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__Q), .o(n_10908) );
ao22f02 g56833_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__Q), .o(n_10907) );
ao22f02 g56835_u0 ( .a(FE_OFN2146_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__Q), .c(FE_OFN1547_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__Q), .o(n_10014) );
ao22f02 g56837_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__Q), .c(FE_OCP_RBN2006_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__Q), .o(n_10010) );
in01f02 g56838_u0 ( .a(n_10592), .o(n_10906) );
ao22f02 g56839_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__Q), .c(FE_OFN1498_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__Q), .o(n_10592) );
ao22f02 g56840_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q), .c(FE_OCPN1873_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q), .o(n_11732) );
ao22f02 g56841_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__Q), .o(n_10905) );
ao22f02 g56842_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__Q), .o(n_10904) );
ao22f02 g56843_u0 ( .a(FE_OFN2131_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__Q), .c(FE_OFN1528_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__Q), .o(n_16841) );
ao22f02 g56844_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__Q), .c(FE_OFN2142_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__Q), .o(n_16840) );
ao22f02 g56845_u0 ( .a(FE_OFN1511_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__34__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q), .o(n_10007) );
in01f02 g56846_u0 ( .a(n_10903), .o(n_11731) );
ao22f02 g56849_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__Q), .c(FE_OFN2207_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__Q), .o(n_10902) );
ao22f02 g56850_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__Q), .o(n_10901) );
ao22f02 g56851_u0 ( .a(FE_OFN2216_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__Q), .o(n_11730) );
ao22f02 g56853_u0 ( .a(FE_OFN2131_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__Q), .c(FE_OFN1528_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q), .o(n_10584) );
ao22f02 g56854_u0 ( .a(n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__Q), .o(n_9997) );
in01f02 g56856_u0 ( .a(n_10898), .o(n_11727) );
ao22f02 g56857_u0 ( .a(FE_OFN1493_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__Q), .o(n_10898) );
ao22f02 g56858_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__Q), .o(n_10579) );
ao22f02 g56860_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__Q), .c(FE_OFN2207_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__Q), .o(n_10895) );
ao22f02 g56862_u0 ( .a(n_9991), .b(n_337), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__Q), .o(n_9993) );
ao22f02 g56863_u0 ( .a(FE_OFN2137_n_15534), .b(n_354), .c(FE_OFN2145_n_16992), .d(n_393), .o(n_16844) );
ao22f02 g56864_u0 ( .a(FE_OFN2131_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__Q), .c(FE_OFN1528_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__Q), .o(n_10577) );
in01f02 g56865_u0 ( .a(n_11725), .o(n_11880) );
ao22f02 g56866_u0 ( .a(FE_OFN2216_n_10143), .b(n_251), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__Q), .o(n_11725) );
ao22f02 g56867_u0 ( .a(FE_OFN2150_n_10595), .b(n_317), .c(FE_OFN2207_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__Q), .o(n_10891) );
ao22f02 g56868_u0 ( .a(FE_OFN1493_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__Q), .o(n_10576) );
ao22f02 g56869_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__Q), .o(n_10890) );
ao22f02 g56870_u0 ( .a(FE_OCPN1882_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__Q), .c(FE_OFN1502_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q), .o(n_9992) );
ao22f02 g56871_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q), .o(n_10575) );
ao22f02 g56873_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__Q), .o(n_10572) );
in01f02 g56874_u0 ( .a(n_10889), .o(n_11724) );
ao22f02 g56875_u0 ( .a(FE_OFN1538_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__Q), .c(FE_OCPN1915_FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__Q), .o(n_10889) );
ao22f02 g56876_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__Q), .o(n_11723) );
ao22f02 g56877_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__Q), .c(FE_OFN1545_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__Q), .o(n_10569) );
ao22f02 g56878_u0 ( .a(FE_OCPN1892_FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__Q), .c(FE_OCP_RBN1934_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__Q), .o(n_10885) );
ao22f02 g56879_u0 ( .a(n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__Q), .o(n_16851) );
ao22f01 g56880_u0 ( .a(FE_OFN2131_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__Q), .c(n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__Q), .o(n_10564) );
ao22f02 g56881_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__Q), .c(FE_OFN2141_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__Q), .o(n_16850) );
in01f02 g56883_u0 ( .a(n_10561), .o(n_10882) );
ao22f02 g56884_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__Q), .o(n_10561) );
ao22f02 g56885_u0 ( .a(FE_OFN2216_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__Q), .o(n_11720) );
ao22f02 g56886_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__Q), .c(FE_OFN2207_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__Q), .o(n_10881) );
ao22f02 g56887_u0 ( .a(FE_OFN1490_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__Q), .o(n_10880) );
ao22f02 g56890_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__Q), .c(FE_OCP_RBN2006_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__Q), .o(n_9976) );
ao22f02 g56891_u0 ( .a(FE_OCP_RBN1968_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__Q), .c(n_10232), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__Q), .o(n_10560) );
in01f02 g56892_u0 ( .a(n_10559), .o(n_10876) );
ao22f02 g56893_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__Q), .c(FE_OFN1498_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q), .o(n_10559) );
ao22f02 g56894_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__Q), .o(n_10875) );
ao22f02 g56895_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__Q), .c(FE_OCPN1873_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__Q), .o(n_10873) );
ao22f02 g56896_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__Q), .o(n_10870) );
ao22f02 g56897_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__Q), .o(n_10556) );
ao22f02 g56898_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q), .c(FE_OFN1723_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q), .o(n_9971) );
ao22f01 g56899_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q), .c(n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q), .o(n_10554) );
ao22f02 g56900_u0 ( .a(n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__Q), .c(FE_OFN1501_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__Q), .o(n_9968) );
in01f02 g56901_u0 ( .a(n_10553), .o(n_10867) );
ao22f02 g56902_u0 ( .a(FE_OCPN1892_FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__Q), .c(FE_OCP_RBN1934_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__Q), .o(n_10553) );
ao22f02 g56903_u0 ( .a(FE_OFN1539_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__Q), .c(FE_OFN1521_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__Q), .o(n_10866) );
ao22f02 g56904_u0 ( .a(FE_OFN1535_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__Q), .o(n_11719) );
ao22f02 g56905_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__Q), .c(n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__Q), .o(n_10865) );
ao22f02 g56906_u0 ( .a(FE_OCPN1882_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__Q), .c(FE_OFN1500_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__Q), .o(n_16837) );
ao22f02 g56907_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__Q), .o(n_9962) );
ao22f01 g56908_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__Q), .o(n_16836) );
ao22f01 g56909_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__Q), .o(n_10547) );
in01f02 g56910_u0 ( .a(n_10864), .o(n_11718) );
ao22f02 g56911_u0 ( .a(FE_OFN1538_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__Q), .c(FE_OCPN1915_FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__Q), .o(n_10864) );
ao22f02 g56912_u0 ( .a(FE_OFN1491_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__Q), .c(n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__Q), .o(n_10544) );
ao22f02 g56913_u0 ( .a(FE_OCPN1892_FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__Q), .c(FE_OCP_RBN1934_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__Q), .o(n_10541) );
ao22f02 g56914_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__Q), .o(n_11717) );
ao22f02 g56915_u0 ( .a(n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__8__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__8__Q), .o(n_16839) );
ao22f02 g56916_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q), .o(n_9956) );
ao22f02 g56917_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q), .c(FE_OFN2142_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__8__Q), .o(n_16838) );
in01f02 g56919_u0 ( .a(n_10530), .o(n_10860) );
ao22f02 g56921_u0 ( .a(FE_OFN1493_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__Q), .o(n_10527) );
ao22f02 g56922_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__Q), .c(FE_OFN2206_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__Q), .o(n_10859) );
ao22f02 g56923_u0 ( .a(FE_OFN2216_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__Q), .o(n_11716) );
ao22f02 g56924_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__Q), .c(FE_OCP_RBN1932_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__Q), .o(n_9953) );
ao22f02 g56925_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__Q), .o(n_9950) );
ao22f02 g56927_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__Q), .c(FE_OCPN2015_n_10195), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__Q), .o(n_10521) );
in01f02 g56928_u0 ( .a(n_10518), .o(n_10856) );
ao22f02 g56929_u0 ( .a(FE_OCPN1882_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__Q), .c(FE_OFN1502_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__Q), .o(n_10518) );
ao22f02 g56930_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__Q), .c(FE_OCPN1888_FE_OFN473_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__Q), .o(n_11715) );
ao22f02 g56931_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__Q), .o(n_10855) );
ao22f02 g56932_u0 ( .a(FE_OCPN1886_FE_OFN1508_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__Q), .o(n_10851) );
in01s03 g56933_u0 ( .a(pci_target_unit_fifos_pcir_flush_in), .o(g56933_sb) );
na02f02 TIMEBOOST_cell_41550 ( .a(TIMEBOOST_net_13013), .b(g57586_sb), .o(n_10799) );
na02f08 TIMEBOOST_cell_4109 ( .a(TIMEBOOST_net_634), .b(n_16167), .o(n_16299) );
na02f02 TIMEBOOST_cell_4110 ( .a(n_7712), .b(n_8452), .o(TIMEBOOST_net_635) );
in01s02 g56934_u0 ( .a(FE_OFN276_n_9941), .o(g56934_sb) );
na02s01 TIMEBOOST_cell_44911 ( .a(TIMEBOOST_net_9513), .b(FE_OFN1044_n_2037), .o(TIMEBOOST_net_14694) );
na02f02 TIMEBOOST_cell_4061 ( .a(n_7695), .b(TIMEBOOST_net_610), .o(n_14485) );
in01s01 TIMEBOOST_cell_32831 ( .a(TIMEBOOST_net_10332), .o(TIMEBOOST_net_10331) );
in01f01 g56959_u0 ( .a(n_8934), .o(n_8875) );
no02m06 g56960_u0 ( .a(n_2878), .b(n_8800), .o(n_8934) );
na02f02 TIMEBOOST_cell_44260 ( .a(TIMEBOOST_net_14368), .b(FE_OFN1421_n_8567), .o(TIMEBOOST_net_12892) );
in01f02 g56975_u0 ( .a(n_8941), .o(n_10789) );
na02f02 g56976_u0 ( .a(n_9152), .b(n_8939), .o(n_8941) );
na02f06 g56978_u0 ( .a(n_16605), .b(n_9173), .o(n_9256) );
na02f02 g56980_u0 ( .a(n_9173), .b(n_8939), .o(n_8940) );
no02f02 g56985_u0 ( .a(n_9173), .b(n_8924), .o(n_9163) );
in01f02 g56991_u0 ( .a(n_9174), .o(n_11795) );
na02f02 g56992_u0 ( .a(n_9173), .b(n_9171), .o(n_9174) );
in01f02 g56999_u0 ( .a(n_9172), .o(n_11138) );
na02f02 g57000_u0 ( .a(n_9152), .b(n_9171), .o(n_9172) );
in01f03 g57003_u0 ( .a(n_9153), .o(n_11125) );
na02f02 g57009_u0 ( .a(n_9152), .b(n_15516), .o(n_9153) );
na02f02 g57011_u0 ( .a(n_9173), .b(n_15516), .o(n_9170) );
oa12s02 g57019_u0 ( .a(n_8871), .b(pci_target_unit_fifos_pcir_flush_in), .c(n_8876), .o(n_9168) );
oa12f01 g57020_u0 ( .a(n_9160), .b(FE_OFN276_n_9941), .c(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(n_9942) );
oa12m02 g57021_u0 ( .a(n_8950), .b(FE_OFN1394_n_8567), .c(n_9928), .o(n_11710) );
oa12m02 g57022_u0 ( .a(n_8949), .b(FE_OFN2184_n_8567), .c(n_9926), .o(n_11708) );
oa12m02 g57023_u0 ( .a(n_8890), .b(FE_OFN2184_n_8567), .c(n_9924), .o(n_11707) );
oa12m02 g57024_u0 ( .a(n_8889), .b(FE_OFN1403_n_8567), .c(n_9922), .o(n_11706) );
oa12m02 g57025_u0 ( .a(n_8888), .b(FE_OFN1403_n_8567), .c(n_9920), .o(n_11705) );
oa12m02 g57026_u0 ( .a(n_8947), .b(FE_OFN1402_n_8567), .c(n_9918), .o(n_11712) );
oa12m02 g57027_u0 ( .a(n_8946), .b(FE_OFN2184_n_8567), .c(n_9916), .o(n_11703) );
oa12m02 g57028_u0 ( .a(n_8945), .b(FE_OFN1402_n_8567), .c(n_9914), .o(n_11702) );
oa12m02 g57029_u0 ( .a(n_8944), .b(FE_OFN2184_n_8567), .c(n_9912), .o(n_11701) );
no02s02 g57030_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_reg_16__Q), .b(n_3463), .o(g57030_p) );
ao12s02 g57030_u1 ( .a(g57030_p), .b(pci_target_unit_del_sync_comp_cycle_count_reg_16__Q), .c(n_3463), .o(n_4697) );
oa12m02 g57031_u0 ( .a(n_8943), .b(FE_OFN1402_n_8567), .c(n_9910), .o(n_11700) );
oa12m02 g57032_u0 ( .a(n_8887), .b(FE_OFN2184_n_8567), .c(n_9908), .o(n_11699) );
no02m02 g57033_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q), .b(n_3462), .o(g57033_p) );
ao12m02 g57033_u1 ( .a(g57033_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q), .c(n_3462), .o(n_4800) );
in01f01 g57034_u0 ( .a(FE_OFN1420_n_8567), .o(g57034_sb) );
na02m02 TIMEBOOST_cell_30791 ( .a(TIMEBOOST_net_9306), .b(n_2883), .o(TIMEBOOST_net_544) );
na02f02 TIMEBOOST_cell_4177 ( .a(FE_OFN1602_n_13995), .b(TIMEBOOST_net_668), .o(n_14504) );
na02s01 TIMEBOOST_cell_42862 ( .a(TIMEBOOST_net_13669), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_11218) );
in01f02 g57035_u0 ( .a(FE_OFN2179_n_8567), .o(g57035_sb) );
na02s02 TIMEBOOST_cell_45303 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__Q), .b(n_3643), .o(TIMEBOOST_net_14890) );
na02s01 TIMEBOOST_cell_41853 ( .a(g61837_sb), .b(g61837_db), .o(TIMEBOOST_net_13165) );
na02s01 TIMEBOOST_cell_41854 ( .a(TIMEBOOST_net_13165), .b(n_4618), .o(n_6973) );
in01f01 g57036_u0 ( .a(FE_OFN1422_n_8567), .o(g57036_sb) );
na02s01 TIMEBOOST_cell_42863 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__Q), .b(FE_OFN542_n_9690), .o(TIMEBOOST_net_13670) );
na02s01 TIMEBOOST_cell_41855 ( .a(g62783_sb), .b(g62783_db), .o(TIMEBOOST_net_13166) );
na02m02 TIMEBOOST_cell_21982 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__Q), .o(TIMEBOOST_net_6248) );
in01f01 g57037_u0 ( .a(FE_OFN1397_n_8567), .o(g57037_sb) );
na03f02 TIMEBOOST_cell_35991 ( .a(g54489_sb), .b(n_13617), .c(TIMEBOOST_net_10119), .o(n_13607) );
na02f02 TIMEBOOST_cell_21983 ( .a(TIMEBOOST_net_6248), .b(n_13901), .o(TIMEBOOST_net_3019) );
na03f02 TIMEBOOST_cell_35993 ( .a(TIMEBOOST_net_10117), .b(n_13617), .c(g54492_sb), .o(n_13601) );
in01f01 g57038_u0 ( .a(FE_OFN1374_n_8567), .o(g57038_sb) );
na04f02 TIMEBOOST_cell_35987 ( .a(wbu_addr_in_255), .b(g52619_sb), .c(g52619_db), .d(TIMEBOOST_net_6387), .o(n_11851) );
na02s01 TIMEBOOST_cell_42860 ( .a(TIMEBOOST_net_13668), .b(FE_OFN1635_n_9531), .o(TIMEBOOST_net_11208) );
in01f02 g57039_u0 ( .a(FE_OFN2170_n_8567), .o(g57039_sb) );
na03f02 TIMEBOOST_cell_4230 ( .a(n_17050), .b(n_17051), .c(n_9301), .o(TIMEBOOST_net_695) );
na02s02 TIMEBOOST_cell_45304 ( .a(TIMEBOOST_net_14890), .b(FE_OFN1295_n_4098), .o(TIMEBOOST_net_12523) );
na02f02 TIMEBOOST_cell_44570 ( .a(TIMEBOOST_net_14523), .b(FE_OFN2180_n_8567), .o(TIMEBOOST_net_13002) );
in01f02 g57040_u0 ( .a(FE_OFN2170_n_8567), .o(g57040_sb) );
na03s02 TIMEBOOST_cell_33269 ( .a(FE_OFN229_n_9120), .b(g58230_sb), .c(g58246_db), .o(n_9044) );
na02m02 TIMEBOOST_cell_44131 ( .a(n_9033), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__Q), .o(TIMEBOOST_net_14304) );
na02s01 TIMEBOOST_cell_37311 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__Q), .b(n_8140), .o(TIMEBOOST_net_10894) );
in01f01 g57041_u0 ( .a(FE_OFN1385_n_8567), .o(g57041_sb) );
na02s01 TIMEBOOST_cell_9763 ( .a(TIMEBOOST_net_1448), .b(g65908_db), .o(n_1855) );
na02f02 TIMEBOOST_cell_4187 ( .a(TIMEBOOST_net_673), .b(n_10127), .o(n_12155) );
na03f02 TIMEBOOST_cell_35995 ( .a(TIMEBOOST_net_10115), .b(n_13617), .c(g54494_sb), .o(n_13597) );
in01f01 g57042_u0 ( .a(FE_OFN1423_n_8567), .o(g57042_sb) );
na02s01 TIMEBOOST_cell_41856 ( .a(TIMEBOOST_net_13166), .b(n_4737), .o(n_7132) );
na02m02 TIMEBOOST_cell_41857 ( .a(FE_OFN1148_n_13249), .b(TIMEBOOST_net_9660), .o(TIMEBOOST_net_13167) );
na02m02 TIMEBOOST_cell_21984 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__Q), .o(TIMEBOOST_net_6249) );
in01f01 g57043_u0 ( .a(FE_OFN1389_n_8567), .o(g57043_sb) );
na02s01 TIMEBOOST_cell_42864 ( .a(TIMEBOOST_net_13670), .b(FE_OFN262_n_9851), .o(TIMEBOOST_net_11213) );
na02f02 TIMEBOOST_cell_21985 ( .a(TIMEBOOST_net_6249), .b(n_13901), .o(TIMEBOOST_net_3016) );
na02m02 TIMEBOOST_cell_41858 ( .a(TIMEBOOST_net_13167), .b(g54234_sb), .o(n_13441) );
in01f01 g57044_u0 ( .a(FE_OFN1349_n_8567), .o(g57044_sb) );
na02s01 TIMEBOOST_cell_36382 ( .a(TIMEBOOST_net_10429), .b(g63590_sb), .o(n_2564) );
na02s02 TIMEBOOST_cell_42970 ( .a(TIMEBOOST_net_13723), .b(g54196_db), .o(n_13422) );
na02s01 TIMEBOOST_cell_45626 ( .a(TIMEBOOST_net_15051), .b(g58186_db), .o(n_9600) );
in01f01 g57045_u0 ( .a(FE_OFN1420_n_8567), .o(g57045_sb) );
na02s01 TIMEBOOST_cell_42932 ( .a(TIMEBOOST_net_13704), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_11152) );
na02f02 TIMEBOOST_cell_41859 ( .a(TIMEBOOST_net_9655), .b(FE_OFN1148_n_13249), .o(TIMEBOOST_net_13168) );
na02s02 TIMEBOOST_cell_31934 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_391), .b(g54200_sb), .o(TIMEBOOST_net_9878) );
in01f02 g57046_u0 ( .a(FE_OFN2177_n_8567), .o(g57046_sb) );
na02m02 TIMEBOOST_cell_44689 ( .a(n_9199), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__Q), .o(TIMEBOOST_net_14583) );
na02s02 TIMEBOOST_cell_37310 ( .a(TIMEBOOST_net_10893), .b(FE_OFN636_n_4669), .o(TIMEBOOST_net_10518) );
na02s01 TIMEBOOST_cell_37313 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__Q), .b(FE_OFN630_n_4454), .o(TIMEBOOST_net_10895) );
in01f01 g57047_u0 ( .a(FE_OFN1390_n_8567), .o(g57047_sb) );
na02s01 TIMEBOOST_cell_37312 ( .a(TIMEBOOST_net_10894), .b(n_2169), .o(TIMEBOOST_net_9983) );
na02f02 TIMEBOOST_cell_38447 ( .a(FE_OCPN1823_n_16560), .b(n_15376), .o(TIMEBOOST_net_11462) );
na02s02 TIMEBOOST_cell_37315 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__Q), .b(FE_OFN633_n_4454), .o(TIMEBOOST_net_10896) );
in01f01 g57048_u0 ( .a(FE_OFN1407_n_8567), .o(g57048_sb) );
na02s01 g65235_u1 ( .a(n_2651), .b(g65235_sb), .o(g65235_da) );
na02m02 TIMEBOOST_cell_44571 ( .a(n_9435), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q), .o(TIMEBOOST_net_14524) );
na02f02 TIMEBOOST_cell_44132 ( .a(TIMEBOOST_net_14304), .b(FE_OFN1404_n_8567), .o(TIMEBOOST_net_12746) );
in01f02 g57049_u0 ( .a(FE_OFN2190_n_8567), .o(g57049_sb) );
na02s01 TIMEBOOST_cell_42980 ( .a(TIMEBOOST_net_13728), .b(g58189_db), .o(n_9058) );
na02s01 TIMEBOOST_cell_37314 ( .a(TIMEBOOST_net_10895), .b(g65027_sb), .o(TIMEBOOST_net_230) );
na02s02 TIMEBOOST_cell_37317 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__Q), .b(FE_OFN629_n_4454), .o(TIMEBOOST_net_10897) );
in01f02 g57050_u0 ( .a(FE_OFN2190_n_8567), .o(g57050_sb) );
na02s02 TIMEBOOST_cell_31026 ( .a(n_4476), .b(g64846_sb), .o(TIMEBOOST_net_9424) );
na02s02 TIMEBOOST_cell_37316 ( .a(TIMEBOOST_net_10896), .b(g65038_sb), .o(TIMEBOOST_net_9452) );
na02s01 TIMEBOOST_cell_37319 ( .a(g58132_sb), .b(g58132_db), .o(TIMEBOOST_net_10898) );
in01f01 g57051_u0 ( .a(FE_OFN1397_n_8567), .o(g57051_sb) );
na02f02 TIMEBOOST_cell_13038 ( .a(FE_OFN1558_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__Q), .o(TIMEBOOST_net_3086) );
na02f02 TIMEBOOST_cell_4197 ( .a(FE_RN_26_0), .b(TIMEBOOST_net_678), .o(n_12817) );
na02s02 TIMEBOOST_cell_45732 ( .a(TIMEBOOST_net_15104), .b(FE_OFN1274_n_4096), .o(TIMEBOOST_net_13272) );
in01f01 g57052_u0 ( .a(FE_OFN1383_n_8567), .o(g57052_sb) );
na02f02 TIMEBOOST_cell_41860 ( .a(TIMEBOOST_net_13168), .b(g54154_sb), .o(n_13445) );
na02f02 TIMEBOOST_cell_4199 ( .a(n_12714), .b(TIMEBOOST_net_679), .o(n_15937) );
na02s01 TIMEBOOST_cell_19051 ( .a(TIMEBOOST_net_4782), .b(g65432_db), .o(n_4673) );
in01f01 g57053_u0 ( .a(FE_OFN1385_n_8567), .o(g57053_sb) );
na02m02 TIMEBOOST_cell_44133 ( .a(n_9549), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__Q), .o(TIMEBOOST_net_14305) );
na02s02 TIMEBOOST_cell_45704 ( .a(TIMEBOOST_net_15090), .b(FE_OFN1270_n_4095), .o(TIMEBOOST_net_12586) );
na02s01 TIMEBOOST_cell_42777 ( .a(FE_OFN213_n_9124), .b(g57982_sb), .o(TIMEBOOST_net_13627) );
na02f02 TIMEBOOST_cell_13044 ( .a(FE_OFN1742_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__26__Q), .o(TIMEBOOST_net_3089) );
na02s02 TIMEBOOST_cell_37318 ( .a(TIMEBOOST_net_10897), .b(g65033_sb), .o(TIMEBOOST_net_9450) );
na02s01 TIMEBOOST_cell_37321 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__Q), .b(n_3739), .o(TIMEBOOST_net_10899) );
in01f02 g57055_u0 ( .a(FE_OFN2179_n_8567), .o(g57055_sb) );
na02f02 TIMEBOOST_cell_41484 ( .a(TIMEBOOST_net_12980), .b(g57312_sb), .o(n_11438) );
na03f02 TIMEBOOST_cell_22354 ( .a(n_10930), .b(n_9277), .c(n_10078), .o(TIMEBOOST_net_6434) );
na02f02 TIMEBOOST_cell_22355 ( .a(TIMEBOOST_net_6434), .b(n_9276), .o(n_12439) );
in01f01 g57056_u0 ( .a(FE_OFN1368_n_8567), .o(g57056_sb) );
na02f02 TIMEBOOST_cell_44572 ( .a(TIMEBOOST_net_14524), .b(FE_OFN2184_n_8567), .o(TIMEBOOST_net_13003) );
na02m02 TIMEBOOST_cell_44573 ( .a(n_9491), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__Q), .o(TIMEBOOST_net_14525) );
na02s01 TIMEBOOST_cell_42778 ( .a(TIMEBOOST_net_13627), .b(g57982_db), .o(n_9110) );
in01f01 g57057_u0 ( .a(FE_OFN1392_n_8567), .o(g57057_sb) );
na02f02 TIMEBOOST_cell_44574 ( .a(TIMEBOOST_net_14525), .b(FE_OFN2187_n_8567), .o(TIMEBOOST_net_13471) );
na02f02 TIMEBOOST_cell_44134 ( .a(TIMEBOOST_net_14305), .b(FE_OFN1392_n_8567), .o(TIMEBOOST_net_12732) );
na02s02 TIMEBOOST_cell_43476 ( .a(TIMEBOOST_net_13976), .b(FE_OFN2064_n_6391), .o(TIMEBOOST_net_12197) );
in01f02 g57058_u0 ( .a(FE_OFN2174_n_8567), .o(g57058_sb) );
na02s01 TIMEBOOST_cell_43290 ( .a(TIMEBOOST_net_13883), .b(g62047_sb), .o(n_7764) );
na02f02 TIMEBOOST_cell_41240 ( .a(TIMEBOOST_net_12858), .b(g57162_sb), .o(n_11588) );
na02s02 TIMEBOOST_cell_45305 ( .a(n_4256), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__Q), .o(TIMEBOOST_net_14891) );
in01f02 g57059_u0 ( .a(FE_OFN2178_n_8567), .o(g57059_sb) );
na02f02 TIMEBOOST_cell_44690 ( .a(TIMEBOOST_net_14583), .b(FE_OFN1402_n_8567), .o(TIMEBOOST_net_13028) );
na03f02 TIMEBOOST_cell_22358 ( .a(n_9329), .b(n_17046), .c(n_9330), .o(TIMEBOOST_net_6436) );
na02s02 TIMEBOOST_cell_43188 ( .a(TIMEBOOST_net_13832), .b(FE_OFN1218_n_6886), .o(TIMEBOOST_net_11542) );
in01f02 g57060_u0 ( .a(FE_OFN2174_n_8567), .o(g57060_sb) );
na02m02 TIMEBOOST_cell_16012 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_3263) );
in01f01 g57061_u0 ( .a(FE_OFN1377_n_8567), .o(g57061_sb) );
na02s01 TIMEBOOST_cell_42779 ( .a(FE_OFN215_n_9856), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__Q), .o(TIMEBOOST_net_13628) );
na02f02 TIMEBOOST_cell_4207 ( .a(TIMEBOOST_net_683), .b(n_9962), .o(n_12130) );
na02f02 TIMEBOOST_cell_44362 ( .a(TIMEBOOST_net_14419), .b(FE_OFN1387_n_8567), .o(TIMEBOOST_net_12734) );
in01f01 g57062_u0 ( .a(FE_OFN1399_n_8567), .o(g57062_sb) );
na02s01 TIMEBOOST_cell_42780 ( .a(TIMEBOOST_net_13628), .b(FE_OFN1634_n_9531), .o(TIMEBOOST_net_11013) );
na02s02 TIMEBOOST_cell_45306 ( .a(TIMEBOOST_net_14891), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_12533) );
na02m02 TIMEBOOST_cell_43855 ( .a(n_9570), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__Q), .o(TIMEBOOST_net_14166) );
in01f01 g57063_u0 ( .a(FE_OFN1394_n_8567), .o(g57063_sb) );
na02s02 TIMEBOOST_cell_37320 ( .a(TIMEBOOST_net_10898), .b(FE_OFN243_n_9116), .o(n_9073) );
na03m02 TIMEBOOST_cell_35695 ( .a(TIMEBOOST_net_10018), .b(FE_OFN1305_n_13124), .c(g54367_sb), .o(n_13123) );
na02f02 TIMEBOOST_cell_43856 ( .a(TIMEBOOST_net_14166), .b(FE_OFN1385_n_8567), .o(TIMEBOOST_net_12938) );
in01f02 g57064_u0 ( .a(FE_OFN2167_n_8567), .o(g57064_sb) );
na02f02 TIMEBOOST_cell_44671 ( .a(TIMEBOOST_net_10053), .b(FE_OFN1407_n_8567), .o(TIMEBOOST_net_14574) );
na03f02 TIMEBOOST_cell_34806 ( .a(TIMEBOOST_net_5444), .b(n_3135), .c(TIMEBOOST_net_594), .o(n_14846) );
na02s01 TIMEBOOST_cell_41795 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__Q), .b(g58387_sb), .o(TIMEBOOST_net_13136) );
in01f01 g57065_u0 ( .a(FE_OFN1412_n_8567), .o(g57065_sb) );
na02s01 TIMEBOOST_cell_42781 ( .a(FE_OFN207_n_9865), .b(g57977_sb), .o(TIMEBOOST_net_13629) );
na02s01 TIMEBOOST_cell_30896 ( .a(pci_target_unit_pcit_if_strd_addr_in_688), .b(n_2499), .o(TIMEBOOST_net_9359) );
na03f02 TIMEBOOST_cell_4212 ( .a(n_10602), .b(n_10020), .c(n_10017), .o(TIMEBOOST_net_686) );
in01f01 g57066_u0 ( .a(FE_OFN1397_n_8567), .o(g57066_sb) );
na02s01 TIMEBOOST_cell_42782 ( .a(TIMEBOOST_net_13629), .b(g57977_db), .o(n_9824) );
na02f02 TIMEBOOST_cell_4213 ( .a(TIMEBOOST_net_686), .b(n_10605), .o(n_12143) );
na02s02 TIMEBOOST_cell_43189 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__Q), .b(n_3715), .o(TIMEBOOST_net_13833) );
in01f02 g57067_u0 ( .a(FE_OFN2173_n_8567), .o(g57067_sb) );
na02f02 TIMEBOOST_cell_42434 ( .a(TIMEBOOST_net_13455), .b(g57281_sb), .o(n_10412) );
na02s02 TIMEBOOST_cell_42370 ( .a(TIMEBOOST_net_13423), .b(g54358_sb), .o(n_13084) );
na02s01 TIMEBOOST_cell_45577 ( .a(FE_OFN638_n_4669), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__Q), .o(TIMEBOOST_net_15027) );
in01f01 g57068_u0 ( .a(FE_OFN1423_n_8567), .o(g57068_sb) );
na02f02 TIMEBOOST_cell_13058 ( .a(FE_OFN1738_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__Q), .o(TIMEBOOST_net_3096) );
na02s02 TIMEBOOST_cell_45307 ( .a(n_4290), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__Q), .o(TIMEBOOST_net_14892) );
na02s02 TIMEBOOST_cell_43190 ( .a(TIMEBOOST_net_13833), .b(FE_OFN1282_n_4097), .o(TIMEBOOST_net_12035) );
in01f01 g57069_u0 ( .a(FE_OFN1421_n_8567), .o(g57069_sb) );
na02s01 TIMEBOOST_cell_42783 ( .a(g60678_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__Q), .o(TIMEBOOST_net_13630) );
na02s02 TIMEBOOST_cell_45308 ( .a(TIMEBOOST_net_14892), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_12534) );
na02s02 TIMEBOOST_cell_42784 ( .a(TIMEBOOST_net_13630), .b(g60678_da), .o(TIMEBOOST_net_11353) );
in01f01 g57070_u0 ( .a(FE_OFN1404_n_8567), .o(g57070_sb) );
na02m02 TIMEBOOST_cell_44575 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__Q), .b(n_9222), .o(TIMEBOOST_net_14526) );
na02f02 TIMEBOOST_cell_44576 ( .a(TIMEBOOST_net_14526), .b(FE_OFN2170_n_8567), .o(TIMEBOOST_net_13428) );
na02s01 TIMEBOOST_cell_45026 ( .a(TIMEBOOST_net_14751), .b(FE_OFN2021_n_4778), .o(TIMEBOOST_net_13654) );
in01f01 g57071_u0 ( .a(FE_OFN1425_n_8567), .o(g57071_sb) );
na02f02 TIMEBOOST_cell_13064 ( .a(FE_OFN1748_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__Q), .o(TIMEBOOST_net_3099) );
na02s02 TIMEBOOST_cell_45309 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__Q), .b(n_3580), .o(TIMEBOOST_net_14893) );
na02s01 TIMEBOOST_cell_42785 ( .a(g61885_sb), .b(g61960_db), .o(TIMEBOOST_net_13631) );
in01f02 g57072_u0 ( .a(FE_OFN1370_n_8567), .o(g57072_sb) );
na02m02 TIMEBOOST_cell_44577 ( .a(n_9221), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__Q), .o(TIMEBOOST_net_14527) );
na02f02 TIMEBOOST_cell_44578 ( .a(TIMEBOOST_net_14527), .b(FE_OFN2178_n_8567), .o(TIMEBOOST_net_13472) );
na02s01 TIMEBOOST_cell_42786 ( .a(TIMEBOOST_net_13631), .b(g63619_db), .o(TIMEBOOST_net_12439) );
in01f01 g57073_u0 ( .a(FE_OFN1415_n_8567), .o(g57073_sb) );
na02m02 TIMEBOOST_cell_44579 ( .a(n_9804), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__Q), .o(TIMEBOOST_net_14528) );
na02f02 TIMEBOOST_cell_44580 ( .a(TIMEBOOST_net_14528), .b(FE_OFN2191_n_8567), .o(TIMEBOOST_net_13023) );
na02s01 TIMEBOOST_cell_42787 ( .a(g61885_sb), .b(g61885_db), .o(TIMEBOOST_net_13632) );
in01f02 g57074_u0 ( .a(FE_OFN2169_n_8567), .o(g57074_sb) );
na02s02 TIMEBOOST_cell_43061 ( .a(n_4305), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__Q), .o(TIMEBOOST_net_13769) );
na02s02 TIMEBOOST_cell_42372 ( .a(TIMEBOOST_net_13424), .b(g54359_sb), .o(n_13083) );
na02f02 TIMEBOOST_cell_42161 ( .a(n_9887), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__Q), .o(TIMEBOOST_net_13319) );
in01f01 g57075_u0 ( .a(FE_OFN1405_n_8567), .o(g57075_sb) );
na02m02 TIMEBOOST_cell_44135 ( .a(n_9540), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__Q), .o(TIMEBOOST_net_14306) );
na02f02 TIMEBOOST_cell_44136 ( .a(TIMEBOOST_net_14306), .b(FE_OFN1370_n_8567), .o(TIMEBOOST_net_12756) );
na02s01 TIMEBOOST_cell_42788 ( .a(TIMEBOOST_net_13632), .b(g63603_db), .o(TIMEBOOST_net_12440) );
in01f02 g57076_u0 ( .a(FE_OFN2182_n_8567), .o(g57076_sb) );
na02s01 TIMEBOOST_cell_42963 ( .a(TIMEBOOST_net_4369), .b(g54188_sb), .o(TIMEBOOST_net_13720) );
na02s01 TIMEBOOST_cell_31072 ( .a(n_4479), .b(g65006_sb), .o(TIMEBOOST_net_9447) );
na02f02 TIMEBOOST_cell_43748 ( .a(TIMEBOOST_net_14112), .b(FE_OFN1397_n_8567), .o(TIMEBOOST_net_12884) );
in01f01 g57077_u0 ( .a(FE_OFN1408_n_8567), .o(g57077_sb) );
na02m02 TIMEBOOST_cell_44581 ( .a(n_9231), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__Q), .o(TIMEBOOST_net_14529) );
na02m02 TIMEBOOST_cell_44137 ( .a(n_9673), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__Q), .o(TIMEBOOST_net_14307) );
na02s02 TIMEBOOST_cell_43402 ( .a(TIMEBOOST_net_13939), .b(n_6431), .o(TIMEBOOST_net_12166) );
in01f02 g57078_u0 ( .a(FE_OFN1389_n_8567), .o(g57078_sb) );
na02m02 TIMEBOOST_cell_43857 ( .a(n_9725), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__Q), .o(TIMEBOOST_net_14167) );
na02f01 g57078_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__Q), .b(FE_OFN1345_n_8567), .o(g57078_db) );
na02s01 TIMEBOOST_cell_37323 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__Q), .b(n_3792), .o(TIMEBOOST_net_10900) );
in01f01 g57079_u0 ( .a(FE_OFN1349_n_8567), .o(g57079_sb) );
na02m02 TIMEBOOST_cell_15932 ( .a(n_1414), .b(n_1413), .o(TIMEBOOST_net_3223) );
na02s02 TIMEBOOST_cell_40696 ( .a(TIMEBOOST_net_12586), .b(g62555_sb), .o(n_6453) );
na02s02 TIMEBOOST_cell_40714 ( .a(TIMEBOOST_net_12595), .b(g62426_sb), .o(n_6745) );
in01f01 g57080_u0 ( .a(FE_OFN1421_n_8567), .o(g57080_sb) );
na02s01 TIMEBOOST_cell_42789 ( .a(g61885_sb), .b(g61977_db), .o(TIMEBOOST_net_13633) );
na02s01 TIMEBOOST_cell_30910 ( .a(pci_target_unit_pcit_if_strd_addr_in_697), .b(pci_target_unit_del_sync_addr_in_215), .o(TIMEBOOST_net_9366) );
na02s01 TIMEBOOST_cell_42790 ( .a(TIMEBOOST_net_13633), .b(g63605_db), .o(TIMEBOOST_net_12441) );
in01f01 g57081_u0 ( .a(FE_OFN1392_n_8567), .o(g57081_sb) );
na02f02 TIMEBOOST_cell_44582 ( .a(TIMEBOOST_net_14529), .b(FE_OFN2184_n_8567), .o(TIMEBOOST_net_13473) );
na02m02 TIMEBOOST_cell_44583 ( .a(n_8997), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q), .o(TIMEBOOST_net_14530) );
na02s01 TIMEBOOST_cell_16787 ( .a(TIMEBOOST_net_3650), .b(g58022_sb), .o(n_9101) );
in01f01 g57082_u0 ( .a(FE_OFN1406_n_8567), .o(g57082_sb) );
na02f02 TIMEBOOST_cell_44138 ( .a(TIMEBOOST_net_14307), .b(FE_OFN1412_n_8567), .o(TIMEBOOST_net_12710) );
na02f02 TIMEBOOST_cell_44584 ( .a(TIMEBOOST_net_14530), .b(FE_OFN2168_n_8567), .o(TIMEBOOST_net_13474) );
na03m02 TIMEBOOST_cell_35891 ( .a(TIMEBOOST_net_4832), .b(g59123_sb), .c(TIMEBOOST_net_5432), .o(n_14813) );
in01f01 g57083_u0 ( .a(FE_OFN1406_n_8567), .o(g57083_sb) );
na02m02 TIMEBOOST_cell_44585 ( .a(n_9705), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__Q), .o(TIMEBOOST_net_14531) );
na02f02 TIMEBOOST_cell_44586 ( .a(TIMEBOOST_net_14531), .b(FE_OFN2174_n_8567), .o(TIMEBOOST_net_13431) );
na03f02 TIMEBOOST_cell_4238 ( .a(n_10942), .b(n_9286), .c(n_10099), .o(TIMEBOOST_net_699) );
in01f01 g57084_u0 ( .a(FE_OFN1424_n_8567), .o(g57084_sb) );
no02f02 TIMEBOOST_cell_13082 ( .a(FE_RN_726_0), .b(FE_RN_725_0), .o(TIMEBOOST_net_3108) );
na02f02 TIMEBOOST_cell_4239 ( .a(TIMEBOOST_net_699), .b(n_9287), .o(n_17041) );
na02s01 TIMEBOOST_cell_41826 ( .a(g63613_da), .b(TIMEBOOST_net_13151), .o(n_7143) );
in01f01 g57085_u0 ( .a(FE_OFN1422_n_8567), .o(g57085_sb) );
na02s01 TIMEBOOST_cell_43191 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__Q), .b(n_4340), .o(TIMEBOOST_net_13834) );
na02m02 TIMEBOOST_cell_44587 ( .a(n_9208), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q), .o(TIMEBOOST_net_14532) );
na03s02 TIMEBOOST_cell_34423 ( .a(n_14679), .b(n_8757), .c(g52442_sb), .o(TIMEBOOST_net_10002) );
in01f02 g57086_u0 ( .a(FE_OFN1370_n_8567), .o(g57086_sb) );
na02m02 TIMEBOOST_cell_13086 ( .a(FE_OFN1566_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q), .o(TIMEBOOST_net_3110) );
na02f02 TIMEBOOST_cell_37073 ( .a(n_13936), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__Q), .o(TIMEBOOST_net_10775) );
na02f02 TIMEBOOST_cell_44588 ( .a(TIMEBOOST_net_14532), .b(FE_OFN2175_n_8567), .o(TIMEBOOST_net_13475) );
in01f01 g57087_u0 ( .a(FE_OFN1414_n_8567), .o(g57087_sb) );
na02m02 TIMEBOOST_cell_44139 ( .a(n_9546), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__Q), .o(TIMEBOOST_net_14308) );
na02m02 TIMEBOOST_cell_44589 ( .a(n_9210), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__Q), .o(TIMEBOOST_net_14533) );
na02s01 TIMEBOOST_cell_37322 ( .a(TIMEBOOST_net_10899), .b(FE_OFN648_n_4497), .o(TIMEBOOST_net_9532) );
in01f01 g57088_u0 ( .a(FE_OFN1414_n_8567), .o(g57088_sb) );
na02s01 TIMEBOOST_cell_16783 ( .a(TIMEBOOST_net_3648), .b(g57991_sb), .o(n_9109) );
na02f02 TIMEBOOST_cell_45858 ( .a(TIMEBOOST_net_15167), .b(n_12061), .o(n_12483) );
na02s02 TIMEBOOST_cell_41966 ( .a(TIMEBOOST_net_13221), .b(g62583_sb), .o(n_6386) );
in01f01 g57089_u0 ( .a(FE_OFN1419_n_8567), .o(g57089_sb) );
na02f02 TIMEBOOST_cell_44590 ( .a(TIMEBOOST_net_14533), .b(FE_OFN2184_n_8567), .o(TIMEBOOST_net_13476) );
na03f03 TIMEBOOST_cell_44591 ( .a(n_337), .b(n_8551), .c(g58610_sb), .o(TIMEBOOST_net_14534) );
na02s01 TIMEBOOST_cell_37325 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__Q), .b(FE_OFN1626_n_4438), .o(TIMEBOOST_net_10901) );
in01f01 g57090_u0 ( .a(FE_OFN1415_n_8567), .o(g57090_sb) );
na02s01 TIMEBOOST_cell_41828 ( .a(g63607_da), .b(TIMEBOOST_net_13152), .o(n_7151) );
na02f02 TIMEBOOST_cell_4251 ( .a(TIMEBOOST_net_705), .b(n_13711), .o(n_14072) );
na03f02 TIMEBOOST_cell_4252 ( .a(n_10708), .b(n_10711), .c(n_10131), .o(TIMEBOOST_net_706) );
in01f01 g57091_u0 ( .a(FE_OFN1368_n_8567), .o(g57091_sb) );
na02f02 TIMEBOOST_cell_45859 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__Q), .b(n_11907), .o(TIMEBOOST_net_15168) );
na02f02 TIMEBOOST_cell_4253 ( .a(TIMEBOOST_net_706), .b(n_12581), .o(n_12843) );
no02f02 TIMEBOOST_cell_4254 ( .a(FE_RN_723_0), .b(FE_RN_722_0), .o(TIMEBOOST_net_707) );
in01f01 g57092_u0 ( .a(FE_OFN1401_n_8567), .o(g57092_sb) );
na02f02 TIMEBOOST_cell_41302 ( .a(TIMEBOOST_net_12889), .b(g57096_sb), .o(n_10487) );
no02f02 TIMEBOOST_cell_4255 ( .a(n_12290), .b(TIMEBOOST_net_707), .o(n_12725) );
na02s02 TIMEBOOST_cell_37534 ( .a(TIMEBOOST_net_11005), .b(FE_OFN2084_n_8407), .o(TIMEBOOST_net_4097) );
in01f02 g57093_u0 ( .a(FE_OFN2169_n_8567), .o(g57093_sb) );
na02s01 TIMEBOOST_cell_42964 ( .a(TIMEBOOST_net_13720), .b(g54188_db), .o(n_13427) );
na02s01 TIMEBOOST_cell_43291 ( .a(TIMEBOOST_net_4771), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_13884) );
na02s01 TIMEBOOST_cell_43292 ( .a(TIMEBOOST_net_13884), .b(g62040_sb), .o(n_7774) );
in01f02 g57094_u0 ( .a(FE_OFN2184_n_8567), .o(g57094_sb) );
na02s02 TIMEBOOST_cell_43501 ( .a(n_4391), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__Q), .o(TIMEBOOST_net_13989) );
na02f02 TIMEBOOST_cell_43749 ( .a(n_9006), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__Q), .o(TIMEBOOST_net_14113) );
na02f02 TIMEBOOST_cell_43293 ( .a(n_3152), .b(wbm_adr_o_16_), .o(TIMEBOOST_net_13885) );
in01f01 g57095_u0 ( .a(FE_OFN1417_n_8567), .o(g57095_sb) );
na02s01 TIMEBOOST_cell_41830 ( .a(g63599_da), .b(TIMEBOOST_net_13153), .o(n_7191) );
na02s01 TIMEBOOST_cell_31806 ( .a(configuration_wb_err_addr_559), .b(conf_wb_err_addr_in_968), .o(TIMEBOOST_net_9814) );
no02f02 TIMEBOOST_cell_4258 ( .a(FE_RN_729_0), .b(FE_RN_728_0), .o(TIMEBOOST_net_709) );
in01f01 g57096_u0 ( .a(FE_OFN1377_n_8567), .o(g57096_sb) );
na02f02 TIMEBOOST_cell_13102 ( .a(FE_OFN1753_n_12086), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__Q), .o(TIMEBOOST_net_3118) );
no02f02 TIMEBOOST_cell_4259 ( .a(n_12215), .b(TIMEBOOST_net_709), .o(n_12636) );
no02f02 TIMEBOOST_cell_4260 ( .a(FE_OCPN1895_FE_OFN1559_n_12042), .b(FE_RN_717_0), .o(TIMEBOOST_net_710) );
in01f01 g57097_u0 ( .a(FE_OFN1403_n_8567), .o(g57097_sb) );
na02f02 TIMEBOOST_cell_45860 ( .a(TIMEBOOST_net_15168), .b(FE_OFN1577_n_12028), .o(n_12626) );
no02f02 TIMEBOOST_cell_4261 ( .a(n_12277), .b(TIMEBOOST_net_710), .o(n_12709) );
na03s02 TIMEBOOST_cell_41799 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__Q), .b(FE_OFN699_n_7845), .c(n_1838), .o(TIMEBOOST_net_13138) );
in01f01 g57098_u0 ( .a(FE_OFN1405_n_8567), .o(g57098_sb) );
na02f02 TIMEBOOST_cell_41306 ( .a(TIMEBOOST_net_12891), .b(g57192_sb), .o(n_11561) );
na02s02 TIMEBOOST_cell_45310 ( .a(TIMEBOOST_net_14893), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_12129) );
na02s02 TIMEBOOST_cell_42965 ( .a(TIMEBOOST_net_9833), .b(g54201_sb), .o(TIMEBOOST_net_13721) );
in01f01 g57099_u0 ( .a(FE_OFN1380_n_8567), .o(g57099_sb) );
na02f02 TIMEBOOST_cell_13108 ( .a(FE_OFN1556_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__Q), .o(TIMEBOOST_net_3121) );
na02m02 TIMEBOOST_cell_38850 ( .a(TIMEBOOST_net_11663), .b(g58486_sb), .o(n_9348) );
na02s02 TIMEBOOST_cell_38150 ( .a(TIMEBOOST_net_11313), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_4537) );
in01f01 g57100_u0 ( .a(FE_OFN1400_n_8567), .o(g57100_sb) );
na02s01 TIMEBOOST_cell_42815 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__Q), .b(g65277_sb), .o(TIMEBOOST_net_13646) );
na02s02 TIMEBOOST_cell_41706 ( .a(TIMEBOOST_net_13091), .b(g58786_db), .o(n_9876) );
in01f01 g57101_u0 ( .a(FE_OFN1382_n_8567), .o(g57101_sb) );
na02s01 TIMEBOOST_cell_42816 ( .a(TIMEBOOST_net_13646), .b(g65277_db), .o(n_3586) );
na02f02 TIMEBOOST_cell_38930 ( .a(TIMEBOOST_net_11703), .b(g58601_sb), .o(n_9241) );
na02s02 TIMEBOOST_cell_38152 ( .a(TIMEBOOST_net_11314), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_4682) );
in01f01 g57102_u0 ( .a(FE_OFN1420_n_8567), .o(g57102_sb) );
na04f04 TIMEBOOST_cell_35909 ( .a(pci_target_unit_pci_target_sm_n_3), .b(n_9175), .c(n_9177), .d(g55853_sb), .o(n_9176) );
na02f02 TIMEBOOST_cell_44592 ( .a(TIMEBOOST_net_14534), .b(FE_OFN2185_n_8567), .o(n_9188) );
na02s01 TIMEBOOST_cell_45627 ( .a(FE_OFN221_n_9846), .b(g58180_sb), .o(TIMEBOOST_net_15052) );
in01f01 g57103_u0 ( .a(FE_OFN1425_n_8567), .o(g57103_sb) );
na02f02 TIMEBOOST_cell_42830 ( .a(TIMEBOOST_net_13653), .b(TIMEBOOST_net_467), .o(TIMEBOOST_net_541) );
na02s01 TIMEBOOST_cell_31087 ( .a(TIMEBOOST_net_9454), .b(g65046_db), .o(n_4325) );
na02m02 TIMEBOOST_cell_43345 ( .a(TIMEBOOST_net_9969), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_13911) );
in01f01 g57104_u0 ( .a(FE_OFN1411_n_8567), .o(g57104_sb) );
na03s02 TIMEBOOST_cell_35913 ( .a(n_3872), .b(g63086_sb), .c(g63086_db), .o(n_5082) );
in01f02 TIMEBOOST_cell_32820 ( .a(TIMEBOOST_net_10321), .o(n_3157) );
na02s01 TIMEBOOST_cell_4276 ( .a(n_16818), .b(n_1323), .o(TIMEBOOST_net_718) );
in01f01 g57105_u0 ( .a(FE_OFN1404_n_8567), .o(g57105_sb) );
na03f02 TIMEBOOST_cell_35915 ( .a(wbu_addr_in_252), .b(g52616_sb), .c(TIMEBOOST_net_10085), .o(n_11854) );
na02s03 TIMEBOOST_cell_45765 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__Q), .b(n_13166), .o(TIMEBOOST_net_15121) );
na02s01 TIMEBOOST_cell_4278 ( .a(wbm_rty_i), .b(n_1280), .o(TIMEBOOST_net_719) );
in01f01 g57106_u0 ( .a(FE_OFN1423_n_8567), .o(g57106_sb) );
na02f02 TIMEBOOST_cell_13122 ( .a(n_12313), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__Q), .o(TIMEBOOST_net_3128) );
na02s01 TIMEBOOST_cell_4279 ( .a(TIMEBOOST_net_719), .b(pci_target_unit_wishbone_master_reset_rty_cnt), .o(TIMEBOOST_net_154) );
in01f01 g57107_u0 ( .a(FE_OFN1381_n_8567), .o(g57107_sb) );
na02s02 TIMEBOOST_cell_45713 ( .a(n_4277), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__Q), .o(TIMEBOOST_net_15095) );
na02s01 TIMEBOOST_cell_45010 ( .a(TIMEBOOST_net_14743), .b(g64311_db), .o(n_3864) );
na02f08 TIMEBOOST_cell_4282 ( .a(n_657), .b(n_47), .o(TIMEBOOST_net_721) );
in01f01 g57108_u0 ( .a(FE_OFN1415_n_8567), .o(g57108_sb) );
na02f02 TIMEBOOST_cell_41184 ( .a(TIMEBOOST_net_12830), .b(g57346_sb), .o(n_11405) );
na02f06 TIMEBOOST_cell_4283 ( .a(TIMEBOOST_net_721), .b(n_15302), .o(n_1514) );
na02s01 TIMEBOOST_cell_4284 ( .a(pci_target_unit_wishbone_master_rty_counter_5_), .b(pci_target_unit_wishbone_master_rty_counter_6_), .o(TIMEBOOST_net_722) );
in01f02 g57109_u0 ( .a(FE_OFN2167_n_8567), .o(g57109_sb) );
na02f02 TIMEBOOST_cell_4231 ( .a(TIMEBOOST_net_695), .b(n_10134), .o(n_12156) );
na02s01 TIMEBOOST_cell_30814 ( .a(n_3747), .b(g64810_sb), .o(TIMEBOOST_net_9318) );
na02s01 TIMEBOOST_cell_30818 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__Q), .b(FE_OFN527_n_9899), .o(TIMEBOOST_net_9320) );
in01f01 g57110_u0 ( .a(FE_OFN1405_n_8567), .o(g57110_sb) );
na02f02 TIMEBOOST_cell_13128 ( .a(n_12313), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__Q), .o(TIMEBOOST_net_3131) );
na02s02 TIMEBOOST_cell_4285 ( .a(TIMEBOOST_net_722), .b(n_929), .o(TIMEBOOST_net_43) );
no02f04 TIMEBOOST_cell_4286 ( .a(n_1291), .b(FE_OCPN1849_n_15998), .o(TIMEBOOST_net_723) );
in01f02 g57111_u0 ( .a(FE_OFN2182_n_8567), .o(g57111_sb) );
na02s01 TIMEBOOST_cell_45628 ( .a(TIMEBOOST_net_15052), .b(g58180_db), .o(n_9607) );
na02s01 TIMEBOOST_cell_30820 ( .a(pci_target_unit_fifos_pcir_data_in), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__Q), .o(TIMEBOOST_net_9321) );
na02s01 TIMEBOOST_cell_30824 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__Q), .o(TIMEBOOST_net_9323) );
in01f01 g57112_u0 ( .a(FE_OFN1409_n_8567), .o(g57112_sb) );
na02f02 TIMEBOOST_cell_22568 ( .a(FE_OFN1742_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__8__Q), .o(TIMEBOOST_net_6541) );
na02s01 TIMEBOOST_cell_42085 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__Q), .b(n_4362), .o(TIMEBOOST_net_13281) );
na02s01 TIMEBOOST_cell_37324 ( .a(TIMEBOOST_net_10900), .b(FE_OFN648_n_4497), .o(TIMEBOOST_net_9540) );
in01f01 g57113_u0 ( .a(FE_OFN1388_n_8567), .o(g57113_sb) );
na03f02 TIMEBOOST_cell_35919 ( .a(TIMEBOOST_net_10079), .b(n_10155), .c(n_10792), .o(n_10793) );
no02f08 TIMEBOOST_cell_4287 ( .a(TIMEBOOST_net_723), .b(FE_OCPN1868_n_16289), .o(TIMEBOOST_net_49) );
na02s01 TIMEBOOST_cell_4288 ( .a(FE_OFN1778_parchk_pci_ad_reg_in_1222), .b(g67074_db), .o(TIMEBOOST_net_724) );
in01f01 g57114_u0 ( .a(FE_OFN1421_n_8567), .o(g57114_sb) );
no03f02 TIMEBOOST_cell_35921 ( .a(n_4647), .b(n_7552), .c(n_4881), .o(g59344_p) );
na02s01 TIMEBOOST_cell_4289 ( .a(TIMEBOOST_net_724), .b(g67049_sb), .o(n_1428) );
na02s01 TIMEBOOST_cell_4290 ( .a(n_8486), .b(n_653), .o(TIMEBOOST_net_725) );
in01f01 g57115_u0 ( .a(FE_OFN1345_n_8567), .o(g57115_sb) );
na03s02 TIMEBOOST_cell_40715 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__Q), .b(n_4272), .c(FE_OFN1244_n_4092), .o(TIMEBOOST_net_12596) );
na02f01 g57115_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__Q), .b(FE_OFN1345_n_8567), .o(g57115_db) );
na02s01 TIMEBOOST_cell_36383 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__Q), .b(g65866_sb), .o(TIMEBOOST_net_10430) );
in01f01 g57116_u0 ( .a(FE_OFN1406_n_8567), .o(g57116_sb) );
no03f02 TIMEBOOST_cell_35923 ( .a(n_4644), .b(n_7552), .c(n_4878), .o(g59346_p) );
na02s01 TIMEBOOST_cell_4291 ( .a(TIMEBOOST_net_725), .b(n_177), .o(TIMEBOOST_net_574) );
na02s01 TIMEBOOST_cell_4292 ( .a(n_13766), .b(configuration_sync_command_bit8), .o(TIMEBOOST_net_726) );
in01f02 g57117_u0 ( .a(FE_OFN1389_n_8567), .o(g57117_sb) );
na02f02 TIMEBOOST_cell_43858 ( .a(TIMEBOOST_net_14167), .b(FE_OFN1423_n_8567), .o(TIMEBOOST_net_12847) );
na02f01 g57117_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__Q), .b(FE_OFN1345_n_8567), .o(g57117_db) );
na02m02 TIMEBOOST_cell_43859 ( .a(n_9807), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__Q), .o(TIMEBOOST_net_14168) );
in01f01 g57118_u0 ( .a(FE_OFN1368_n_8567), .o(g57118_sb) );
na02s01 TIMEBOOST_cell_42832 ( .a(TIMEBOOST_net_13654), .b(g63612_da), .o(n_7187) );
na02s01 TIMEBOOST_cell_4293 ( .a(TIMEBOOST_net_726), .b(n_7396), .o(TIMEBOOST_net_112) );
na02s01 TIMEBOOST_cell_4294 ( .a(wbu_addr_in_254), .b(g58794_sb), .o(TIMEBOOST_net_727) );
in01f02 g57119_u0 ( .a(FE_OFN2191_n_8567), .o(g57119_sb) );
na02f02 g55711_u0 ( .a(FE_OFN2202_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__Q), .o(n_12183) );
na03m04 TIMEBOOST_cell_34872 ( .a(g52400_db), .b(g60679_da), .c(TIMEBOOST_net_9992), .o(n_14819) );
na02f02 TIMEBOOST_cell_43750 ( .a(TIMEBOOST_net_14113), .b(FE_OFN1400_n_8567), .o(TIMEBOOST_net_12693) );
in01f01 g57120_u0 ( .a(FE_OFN1424_n_8567), .o(g57120_sb) );
na02s01 TIMEBOOST_cell_41839 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__Q), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_13158) );
na02s01 TIMEBOOST_cell_4295 ( .a(TIMEBOOST_net_727), .b(g58794_db), .o(n_9114) );
na02s01 TIMEBOOST_cell_40289 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__Q), .b(n_8069), .o(TIMEBOOST_net_12383) );
in01f01 g57121_u0 ( .a(FE_OFN1380_n_8567), .o(g57121_sb) );
na02f02 TIMEBOOST_cell_41186 ( .a(TIMEBOOST_net_12831), .b(g57098_sb), .o(n_10483) );
na02s02 TIMEBOOST_cell_45224 ( .a(TIMEBOOST_net_14850), .b(FE_OFN1212_n_4151), .o(TIMEBOOST_net_12105) );
na04s02 TIMEBOOST_cell_34239 ( .a(g64307_da), .b(g64307_db), .c(g63091_sb), .d(g63091_db), .o(n_5071) );
in01f01 g57122_u0 ( .a(FE_OFN1383_n_8567), .o(g57122_sb) );
na02s02 TIMEBOOST_cell_45714 ( .a(TIMEBOOST_net_15095), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_13306) );
na02s01 TIMEBOOST_cell_45011 ( .a(n_1899), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__Q), .o(TIMEBOOST_net_14744) );
na02s01 TIMEBOOST_cell_15856 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_73), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3185) );
in01f01 g57123_u0 ( .a(FE_OFN1345_n_8567), .o(g57123_sb) );
na02s01 TIMEBOOST_cell_36384 ( .a(TIMEBOOST_net_10430), .b(g65866_db), .o(n_1709) );
na04f02 TIMEBOOST_cell_35931 ( .a(wbu_addr_in_257), .b(g52621_sb), .c(g52621_db), .d(TIMEBOOST_net_6287), .o(n_11848) );
na02f02 TIMEBOOST_cell_43860 ( .a(TIMEBOOST_net_14168), .b(FE_OFN1406_n_8567), .o(TIMEBOOST_net_12827) );
in01f01 g57124_u0 ( .a(FE_OFN1419_n_8567), .o(g57124_sb) );
na02f02 TIMEBOOST_cell_36934 ( .a(TIMEBOOST_net_10705), .b(g52603_sb), .o(n_10250) );
na02s01 TIMEBOOST_cell_31041 ( .a(TIMEBOOST_net_9431), .b(g64913_db), .o(n_4398) );
na02s01 TIMEBOOST_cell_31040 ( .a(n_4645), .b(g64913_sb), .o(TIMEBOOST_net_9431) );
in01f01 g57125_u0 ( .a(FE_OFN1415_n_8567), .o(g57125_sb) );
na02f02 TIMEBOOST_cell_44126 ( .a(TIMEBOOST_net_14301), .b(FE_OFN1382_n_8567), .o(TIMEBOOST_net_12708) );
na02s02 TIMEBOOST_cell_45311 ( .a(n_4353), .b(n_139), .o(TIMEBOOST_net_14894) );
na02s02 TIMEBOOST_cell_43106 ( .a(TIMEBOOST_net_13791), .b(FE_OFN1218_n_6886), .o(TIMEBOOST_net_12086) );
in01f01 g57126_u0 ( .a(FE_OFN1368_n_8567), .o(g57126_sb) );
na02f02 TIMEBOOST_cell_41194 ( .a(TIMEBOOST_net_12835), .b(g57520_sb), .o(n_11220) );
na02s02 TIMEBOOST_cell_45629 ( .a(FE_OFN1642_n_4671), .b(g65316_da), .o(TIMEBOOST_net_15053) );
na02s01 TIMEBOOST_cell_45573 ( .a(n_4444), .b(g64997_sb), .o(TIMEBOOST_net_15025) );
in01f01 g57127_u0 ( .a(FE_OFN1401_n_8567), .o(g57127_sb) );
na02f02 TIMEBOOST_cell_41196 ( .a(TIMEBOOST_net_12836), .b(g57097_sb), .o(n_10485) );
na03s02 TIMEBOOST_cell_33220 ( .a(FE_OFN245_n_9114), .b(g58063_sb), .c(g58063_db), .o(n_9089) );
na02s01 TIMEBOOST_cell_4308 ( .a(n_16690), .b(n_2078), .o(TIMEBOOST_net_734) );
in01f01 g57128_u0 ( .a(FE_OFN1417_n_8567), .o(g57128_sb) );
na02f02 TIMEBOOST_cell_44140 ( .a(TIMEBOOST_net_14308), .b(FE_OFN1383_n_8567), .o(TIMEBOOST_net_12788) );
na02s02 TIMEBOOST_cell_4309 ( .a(TIMEBOOST_net_734), .b(n_2316), .o(TIMEBOOST_net_192) );
na02s01 TIMEBOOST_cell_4310 ( .a(pci_target_unit_pci_target_if_target_rd_completed), .b(n_12595), .o(TIMEBOOST_net_735) );
in01f01 g57129_u0 ( .a(FE_OFN1402_n_8567), .o(g57129_sb) );
na02m02 TIMEBOOST_cell_44593 ( .a(n_9414), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q), .o(TIMEBOOST_net_14535) );
na02s01 TIMEBOOST_cell_4311 ( .a(TIMEBOOST_net_735), .b(n_2287), .o(n_2746) );
na02s02 TIMEBOOST_cell_38154 ( .a(TIMEBOOST_net_11315), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_4680) );
in01f01 g57130_u0 ( .a(FE_OFN1417_n_8567), .o(g57130_sb) );
na02f02 TIMEBOOST_cell_44594 ( .a(TIMEBOOST_net_14535), .b(FE_OFN2177_n_8567), .o(TIMEBOOST_net_13009) );
na02s01 TIMEBOOST_cell_4313 ( .a(TIMEBOOST_net_736), .b(g67057_sb), .o(n_1474) );
na02s02 TIMEBOOST_cell_38584 ( .a(TIMEBOOST_net_11530), .b(g60625_sb), .o(n_4828) );
in01f01 g57131_u0 ( .a(FE_OFN1377_n_8567), .o(g57131_sb) );
na02f02 TIMEBOOST_cell_44595 ( .a(n_9049), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__Q), .o(TIMEBOOST_net_14536) );
na02s01 TIMEBOOST_cell_4315 ( .a(TIMEBOOST_net_737), .b(g67057_sb), .o(n_1652) );
na03s02 TIMEBOOST_cell_38423 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__Q), .b(FE_OFN1133_g64577_p), .c(n_3207), .o(TIMEBOOST_net_11450) );
in01f01 g57132_u0 ( .a(FE_OFN1409_n_8567), .o(g57132_sb) );
na02s01 TIMEBOOST_cell_43192 ( .a(TIMEBOOST_net_13834), .b(FE_OFN1260_n_4143), .o(TIMEBOOST_net_12034) );
na02s01 TIMEBOOST_cell_4317 ( .a(TIMEBOOST_net_738), .b(g67057_sb), .o(n_1614) );
na02s01 TIMEBOOST_cell_42592 ( .a(TIMEBOOST_net_13534), .b(g58217_sb), .o(TIMEBOOST_net_11942) );
in01f01 g57133_u0 ( .a(FE_OFN1416_n_8567), .o(g57133_sb) );
na03s02 TIMEBOOST_cell_33534 ( .a(g65210_sb), .b(pci_target_unit_del_sync_addr_in_219), .c(TIMEBOOST_net_801), .o(n_2679) );
na02s01 TIMEBOOST_cell_4319 ( .a(TIMEBOOST_net_739), .b(g67057_sb), .o(n_1654) );
na02m02 TIMEBOOST_cell_41625 ( .a(wbu_sel_in_314), .b(wishbone_slave_unit_fifos_wbr_be_in_266), .o(TIMEBOOST_net_13051) );
in01f01 g57134_u0 ( .a(FE_OFN1396_n_8567), .o(g57134_sb) );
na02s02 TIMEBOOST_cell_43457 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__Q), .b(n_4275), .o(TIMEBOOST_net_13967) );
na02s01 TIMEBOOST_cell_4321 ( .a(TIMEBOOST_net_740), .b(g67057_sb), .o(n_1683) );
in01f01 g57135_u0 ( .a(FE_OFN1413_n_8567), .o(g57135_sb) );
na02m02 TIMEBOOST_cell_44363 ( .a(n_9854), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__Q), .o(TIMEBOOST_net_14420) );
na02s02 TIMEBOOST_cell_45705 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q), .b(n_4489), .o(TIMEBOOST_net_15091) );
na02m02 TIMEBOOST_cell_44317 ( .a(n_9890), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q), .o(TIMEBOOST_net_14397) );
in01f01 g57136_u0 ( .a(FE_OFN1400_n_8567), .o(g57136_sb) );
na02s02 TIMEBOOST_cell_43636 ( .a(TIMEBOOST_net_14056), .b(FE_OFN1225_n_6391), .o(TIMEBOOST_net_12557) );
na02s01 TIMEBOOST_cell_4325 ( .a(TIMEBOOST_net_742), .b(g67057_sb), .o(n_1685) );
na02s01 TIMEBOOST_cell_31037 ( .a(TIMEBOOST_net_9429), .b(g64909_db), .o(n_4404) );
in01f02 g57137_u0 ( .a(FE_OFN2174_n_8567), .o(g57137_sb) );
na02s02 TIMEBOOST_cell_45312 ( .a(TIMEBOOST_net_14894), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_12542) );
na02s01 TIMEBOOST_cell_15838 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_72), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3176) );
na02s01 TIMEBOOST_cell_15840 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_101), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3177) );
in01f01 g57138_u0 ( .a(FE_OFN1425_n_8567), .o(g57138_sb) );
no04m10 TIMEBOOST_cell_13170 ( .a(parchk_pci_ad_out_in_1174), .b(parchk_pci_ad_out_in_1173), .c(FE_RN_731_0), .d(FE_RN_732_0), .o(n_585) );
na02s02 TIMEBOOST_cell_31086 ( .a(n_4470), .b(g65046_sb), .o(TIMEBOOST_net_9454) );
na02s01 TIMEBOOST_cell_4328 ( .a(n_7044), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(TIMEBOOST_net_744) );
in01f01 g57139_u0 ( .a(FE_OFN1411_n_8567), .o(g57139_sb) );
na02s02 TIMEBOOST_cell_45313 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__Q), .b(n_3561), .o(TIMEBOOST_net_14895) );
na02s01 TIMEBOOST_cell_4329 ( .a(TIMEBOOST_net_744), .b(n_243), .o(TIMEBOOST_net_93) );
na04m02 TIMEBOOST_cell_34769 ( .a(TIMEBOOST_net_4828), .b(g63203_sb), .c(g52450_sb), .d(g52450_db), .o(n_14841) );
in01f02 g57140_u0 ( .a(FE_OFN1406_n_8567), .o(g57140_sb) );
na02s02 TIMEBOOST_cell_42040 ( .a(TIMEBOOST_net_13258), .b(g62645_sb), .o(n_6259) );
na02f01 g57140_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__Q), .b(FE_OFN1345_n_8567), .o(g57140_db) );
in01f01 g57141_u0 ( .a(FE_OFN1423_n_8567), .o(g57141_sb) );
na02s02 TIMEBOOST_cell_45314 ( .a(TIMEBOOST_net_14895), .b(FE_OFN1283_n_4097), .o(TIMEBOOST_net_12544) );
na02s01 TIMEBOOST_cell_31036 ( .a(n_4493), .b(g64909_sb), .o(TIMEBOOST_net_9429) );
na02s02 TIMEBOOST_cell_41713 ( .a(TIMEBOOST_net_3258), .b(n_16271), .o(TIMEBOOST_net_13095) );
in01f01 g57142_u0 ( .a(FE_OFN1381_n_8567), .o(g57142_sb) );
na02s02 TIMEBOOST_cell_43193 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__Q), .b(n_3554), .o(TIMEBOOST_net_13835) );
na02f02 TIMEBOOST_cell_42436 ( .a(TIMEBOOST_net_13456), .b(g57235_sb), .o(n_10832) );
na02f02 TIMEBOOST_cell_44596 ( .a(TIMEBOOST_net_14536), .b(FE_OFN2168_n_8567), .o(TIMEBOOST_net_13010) );
in01f01 g57143_u0 ( .a(FE_OFN1345_n_8567), .o(g57143_sb) );
na02f02 TIMEBOOST_cell_4133 ( .a(TIMEBOOST_net_646), .b(n_6978), .o(n_7338) );
na02s02 TIMEBOOST_cell_43458 ( .a(TIMEBOOST_net_13967), .b(FE_OFN1230_n_6391), .o(TIMEBOOST_net_12191) );
na02s01 TIMEBOOST_cell_42018 ( .a(TIMEBOOST_net_13247), .b(g62589_sb), .o(n_6373) );
in01f02 g57144_u0 ( .a(FE_OFN2167_n_8567), .o(g57144_sb) );
na02f02 TIMEBOOST_cell_41354 ( .a(TIMEBOOST_net_12915), .b(g57244_sb), .o(n_11513) );
na02f02 TIMEBOOST_cell_22569 ( .a(n_11925), .b(TIMEBOOST_net_6541), .o(n_12492) );
na02f02 TIMEBOOST_cell_22566 ( .a(FE_OFN1738_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__Q), .o(TIMEBOOST_net_6540) );
in01f01 g57145_u0 ( .a(FE_OFN1405_n_8567), .o(g57145_sb) );
na02s01 TIMEBOOST_cell_45315 ( .a(n_3551), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q), .o(TIMEBOOST_net_14896) );
na02m02 TIMEBOOST_cell_44141 ( .a(n_9642), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__Q), .o(TIMEBOOST_net_14309) );
na02f02 TIMEBOOST_cell_44597 ( .a(n_9072), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__Q), .o(TIMEBOOST_net_14537) );
in01f02 g57146_u0 ( .a(FE_OFN2182_n_8567), .o(g57146_sb) );
na02s02 TIMEBOOST_cell_45316 ( .a(TIMEBOOST_net_14896), .b(FE_OFN1194_n_6935), .o(TIMEBOOST_net_12547) );
na02f02 TIMEBOOST_cell_22567 ( .a(n_11930), .b(TIMEBOOST_net_6540), .o(n_12651) );
na02f02 TIMEBOOST_cell_22564 ( .a(FE_OFN1739_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__Q), .o(TIMEBOOST_net_6539) );
in01f01 g57147_u0 ( .a(FE_OFN1409_n_8567), .o(g57147_sb) );
na02m02 TIMEBOOST_cell_43680 ( .a(TIMEBOOST_net_14078), .b(g58630_db), .o(n_8851) );
na03m02 TIMEBOOST_cell_32916 ( .a(TIMEBOOST_net_544), .b(n_1615), .c(n_2415), .o(TIMEBOOST_net_2007) );
na02s01 TIMEBOOST_cell_17174 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__Q), .b(g65401_sb), .o(TIMEBOOST_net_3844) );
in01f01 g57148_u0 ( .a(FE_OFN1345_n_8567), .o(g57148_sb) );
na02s01 TIMEBOOST_cell_31068 ( .a(n_4452), .b(g65003_sb), .o(TIMEBOOST_net_9445) );
na02f01 g57148_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__Q), .b(FE_OFN1345_n_8567), .o(g57148_db) );
na03m02 TIMEBOOST_cell_4136 ( .a(n_2768), .b(n_2626), .c(n_2902), .o(TIMEBOOST_net_648) );
in01f01 g57149_u0 ( .a(FE_OFN1388_n_8567), .o(g57149_sb) );
na02s01 g58068_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__Q), .b(FE_OFN1793_n_9904), .o(g58068_db) );
na02s01 TIMEBOOST_cell_17175 ( .a(TIMEBOOST_net_3844), .b(g65401_db), .o(n_3519) );
na02m02 TIMEBOOST_cell_4340 ( .a(n_15923), .b(n_2016), .o(TIMEBOOST_net_750) );
in01f01 g57150_u0 ( .a(FE_OFN1421_n_8567), .o(g57150_sb) );
na02m02 TIMEBOOST_cell_44213 ( .a(n_9108), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__Q), .o(TIMEBOOST_net_14345) );
na02f03 TIMEBOOST_cell_4341 ( .a(TIMEBOOST_net_750), .b(n_2028), .o(TIMEBOOST_net_157) );
na02f01 TIMEBOOST_cell_4342 ( .a(n_16424), .b(pciu_pref_en_in_320), .o(TIMEBOOST_net_751) );
in01f01 g57151_u0 ( .a(FE_OFN1406_n_8567), .o(g57151_sb) );
na03s01 TIMEBOOST_cell_13186 ( .a(n_1117), .b(pci_target_unit_fifos_pcir_flush_in), .c(g57780_sb), .o(TIMEBOOST_net_623) );
na02f01 TIMEBOOST_cell_4343 ( .a(TIMEBOOST_net_751), .b(n_15755), .o(n_2388) );
na02s02 TIMEBOOST_cell_45706 ( .a(TIMEBOOST_net_15091), .b(FE_OFN1257_n_4143), .o(TIMEBOOST_net_12532) );
in01f01 g57152_u0 ( .a(FE_OFN1392_n_8567), .o(g57152_sb) );
na04f20 TIMEBOOST_cell_13188 ( .a(FE_OCP_RBN2290_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .b(n_16175), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_1_), .o(n_15824) );
na02f02 TIMEBOOST_cell_41462 ( .a(TIMEBOOST_net_12969), .b(g57557_sb), .o(n_10300) );
na02f02 TIMEBOOST_cell_44598 ( .a(TIMEBOOST_net_14537), .b(FE_OFN2170_n_8567), .o(TIMEBOOST_net_13477) );
in01f02 g57153_u0 ( .a(FE_OFN1389_n_8567), .o(g57153_sb) );
na02f02 TIMEBOOST_cell_22325 ( .a(TIMEBOOST_net_6419), .b(FE_OFN1748_n_12004), .o(n_12732) );
na02f01 g57153_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__Q), .b(FE_OFN1345_n_8567), .o(g57153_db) );
na02m02 TIMEBOOST_cell_44251 ( .a(n_9600), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__Q), .o(TIMEBOOST_net_14364) );
in01f02 g57154_u0 ( .a(FE_OFN2191_n_8567), .o(g57154_sb) );
na02f02 TIMEBOOST_cell_41232 ( .a(TIMEBOOST_net_12854), .b(g57466_sb), .o(n_10343) );
na02f02 TIMEBOOST_cell_22565 ( .a(TIMEBOOST_net_6539), .b(n_11951), .o(n_12671) );
na02f02 TIMEBOOST_cell_41372 ( .a(TIMEBOOST_net_12924), .b(g57069_sb), .o(n_11672) );
in01f01 g57155_u0 ( .a(FE_OFN1424_n_8567), .o(g57155_sb) );
na04f40 TIMEBOOST_cell_13190 ( .a(FE_RN_551_0), .b(FE_OCP_RBN2277_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_), .o(n_16462) );
na02m02 TIMEBOOST_cell_44599 ( .a(n_9134), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__Q), .o(TIMEBOOST_net_14538) );
na02s01 TIMEBOOST_cell_45317 ( .a(n_28), .b(n_4472), .o(TIMEBOOST_net_14897) );
in01f01 g57156_u0 ( .a(FE_OFN1380_n_8567), .o(g57156_sb) );
na02s02 TIMEBOOST_cell_43050 ( .a(TIMEBOOST_net_13763), .b(FE_OFN1258_n_4143), .o(TIMEBOOST_net_12210) );
na02s02 TIMEBOOST_cell_31029 ( .a(TIMEBOOST_net_9425), .b(n_4645), .o(n_4431) );
na02m02 TIMEBOOST_cell_43861 ( .a(n_9802), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__Q), .o(TIMEBOOST_net_14169) );
in01f02 g57157_u0 ( .a(FE_OFN2191_n_8567), .o(g57157_sb) );
na02s01 TIMEBOOST_cell_31027 ( .a(TIMEBOOST_net_9424), .b(g64846_db), .o(n_4436) );
na03s02 TIMEBOOST_cell_32915 ( .a(n_1387), .b(n_1351), .c(n_1486), .o(TIMEBOOST_net_146) );
in01f01 g57158_u0 ( .a(FE_OFN1345_n_8567), .o(g57158_sb) );
na02f02 TIMEBOOST_cell_4137 ( .a(TIMEBOOST_net_648), .b(n_7033), .o(n_7504) );
na02f02 TIMEBOOST_cell_44508 ( .a(TIMEBOOST_net_14492), .b(FE_OFN2167_n_8567), .o(TIMEBOOST_net_13489) );
na02s01 TIMEBOOST_cell_38020 ( .a(TIMEBOOST_net_11248), .b(g61701_sb), .o(n_8426) );
in01f01 g57159_u0 ( .a(FE_OFN1384_n_8567), .o(g57159_sb) );
na02s02 TIMEBOOST_cell_43194 ( .a(TIMEBOOST_net_13835), .b(FE_OFN1288_n_4098), .o(TIMEBOOST_net_12049) );
na02f02 TIMEBOOST_cell_44600 ( .a(TIMEBOOST_net_14538), .b(FE_OFN2168_n_8567), .o(TIMEBOOST_net_13024) );
na02s01 TIMEBOOST_cell_45318 ( .a(TIMEBOOST_net_14897), .b(FE_OFN1219_n_6886), .o(TIMEBOOST_net_12538) );
in01f01 g57160_u0 ( .a(FE_OFN1345_n_8567), .o(g57160_sb) );
no02f02 TIMEBOOST_cell_4139 ( .a(TIMEBOOST_net_649), .b(n_7091), .o(n_13568) );
na02f01 g57160_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__Q), .b(FE_OFN1345_n_8567), .o(g57160_db) );
na02s01 TIMEBOOST_cell_44912 ( .a(TIMEBOOST_net_14694), .b(g65830_sb), .o(TIMEBOOST_net_328) );
in01f01 g57161_u0 ( .a(FE_OFN1368_n_8567), .o(g57161_sb) );
na03s01 TIMEBOOST_cell_13196 ( .a(n_2629), .b(n_2311), .c(n_15407), .o(n_2616) );
na02f02 TIMEBOOST_cell_41466 ( .a(TIMEBOOST_net_12971), .b(g57551_sb), .o(n_11193) );
na02f02 TIMEBOOST_cell_41472 ( .a(TIMEBOOST_net_12974), .b(g57572_sb), .o(n_11179) );
in01f01 g57162_u0 ( .a(FE_OFN1401_n_8567), .o(g57162_sb) );
na02f02 TIMEBOOST_cell_44364 ( .a(TIMEBOOST_net_14420), .b(FE_OFN1408_n_8567), .o(TIMEBOOST_net_12731) );
na02s02 TIMEBOOST_cell_45319 ( .a(n_4374), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__Q), .o(TIMEBOOST_net_14898) );
na02f02 TIMEBOOST_cell_41482 ( .a(TIMEBOOST_net_12979), .b(g57539_sb), .o(n_11203) );
in01f02 g57163_u0 ( .a(FE_OFN2169_n_8567), .o(g57163_sb) );
na02s01 TIMEBOOST_cell_9060 ( .a(wishbone_slave_unit_del_sync_sync_req_comp_pending), .b(g66456_sb), .o(TIMEBOOST_net_1097) );
na02s02 TIMEBOOST_cell_45320 ( .a(TIMEBOOST_net_14898), .b(FE_OFN1250_n_4093), .o(TIMEBOOST_net_12571) );
na02f02 TIMEBOOST_cell_41464 ( .a(TIMEBOOST_net_12970), .b(g57161_sb), .o(n_10460) );
in01f01 g57164_u0 ( .a(FE_OFN1377_n_8567), .o(g57164_sb) );
na02s02 TIMEBOOST_cell_45321 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__Q), .b(n_4291), .o(TIMEBOOST_net_14899) );
na02s02 TIMEBOOST_cell_45322 ( .a(TIMEBOOST_net_14899), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_12076) );
na02s01 TIMEBOOST_cell_31085 ( .a(TIMEBOOST_net_9453), .b(g65039_db), .o(n_4329) );
in01f01 g57165_u0 ( .a(FE_OFN1416_n_8567), .o(g57165_sb) );
na02s01 TIMEBOOST_cell_43195 ( .a(n_4369), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__31__Q), .o(TIMEBOOST_net_13836) );
na02s02 TIMEBOOST_cell_45323 ( .a(wbm_adr_o_18_), .b(FE_OFN1700_n_5751), .o(TIMEBOOST_net_14900) );
na02f02 TIMEBOOST_cell_41476 ( .a(TIMEBOOST_net_12976), .b(g57569_sb), .o(n_11182) );
in01s02 g57166_u0 ( .a(FE_OFN1377_n_8567), .o(g57166_sb) );
na02f02 TIMEBOOST_cell_43862 ( .a(TIMEBOOST_net_14169), .b(FE_OFN1424_n_8567), .o(TIMEBOOST_net_12897) );
na02s02 TIMEBOOST_cell_45324 ( .a(TIMEBOOST_net_14900), .b(g58799_sb), .o(TIMEBOOST_net_587) );
na02f02 TIMEBOOST_cell_41470 ( .a(TIMEBOOST_net_12973), .b(g57303_sb), .o(n_10405) );
in01f01 g57167_u0 ( .a(FE_OFN1409_n_8567), .o(g57167_sb) );
na02m02 TIMEBOOST_cell_44365 ( .a(n_9003), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__Q), .o(TIMEBOOST_net_14421) );
na02m02 TIMEBOOST_cell_45325 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_), .b(n_2274), .o(TIMEBOOST_net_14901) );
na02f02 TIMEBOOST_cell_41454 ( .a(TIMEBOOST_net_12965), .b(g57374_sb), .o(n_11373) );
in01f01 g57168_u0 ( .a(FE_OFN1396_n_8567), .o(g57168_sb) );
na02m02 TIMEBOOST_cell_45326 ( .a(TIMEBOOST_net_14901), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_13274) );
na02f02 TIMEBOOST_cell_41474 ( .a(TIMEBOOST_net_12975), .b(g57317_sb), .o(n_11434) );
na03s02 TIMEBOOST_cell_45327 ( .a(n_3535), .b(FE_OFN1272_n_4096), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__Q), .o(TIMEBOOST_net_14902) );
in01f01 g57169_u0 ( .a(FE_OFN1416_n_8567), .o(g57169_sb) );
na02s01 TIMEBOOST_cell_15960 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__Q), .b(g65957_sb), .o(TIMEBOOST_net_3237) );
na02f02 TIMEBOOST_cell_41456 ( .a(TIMEBOOST_net_12966), .b(g57388_sb), .o(n_11355) );
na02m02 TIMEBOOST_cell_32558 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__Q), .o(TIMEBOOST_net_10190) );
in01f01 g57170_u0 ( .a(FE_OFN1413_n_8567), .o(g57170_sb) );
na02s01 TIMEBOOST_cell_43196 ( .a(TIMEBOOST_net_13836), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_12057) );
na03s01 TIMEBOOST_cell_34245 ( .a(TIMEBOOST_net_9801), .b(FE_OFN1164_n_5615), .c(g62102_sb), .o(n_5600) );
na02s02 TIMEBOOST_cell_45328 ( .a(TIMEBOOST_net_14902), .b(g63002_sb), .o(n_5878) );
in01f01 g57171_u0 ( .a(FE_OFN1370_n_8567), .o(g57171_sb) );
na02s01 TIMEBOOST_cell_45329 ( .a(TIMEBOOST_net_4801), .b(FE_OFN1203_n_4090), .o(TIMEBOOST_net_14903) );
na02s01 TIMEBOOST_cell_4375 ( .a(TIMEBOOST_net_767), .b(g63590_sb), .o(n_1411) );
na02s01 TIMEBOOST_cell_4376 ( .a(n_1816), .b(n_709), .o(TIMEBOOST_net_768) );
in01f02 g57172_u0 ( .a(FE_OFN2173_n_8567), .o(g57172_sb) );
na02m02 TIMEBOOST_cell_41598 ( .a(FE_OFN1438_n_9372), .b(TIMEBOOST_net_13037), .o(TIMEBOOST_net_11664) );
na02s01 TIMEBOOST_cell_45330 ( .a(TIMEBOOST_net_14903), .b(g63149_sb), .o(n_5842) );
na03s02 TIMEBOOST_cell_45331 ( .a(n_4458), .b(FE_OFN1278_n_4097), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__Q), .o(TIMEBOOST_net_14904) );
in01f01 g57173_u0 ( .a(FE_OFN1425_n_8567), .o(g57173_sb) );
na02s01 TIMEBOOST_cell_43197 ( .a(n_4466), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q), .o(TIMEBOOST_net_13837) );
na02s01 TIMEBOOST_cell_4377 ( .a(TIMEBOOST_net_768), .b(n_4686), .o(TIMEBOOST_net_135) );
na02s01 TIMEBOOST_cell_39222 ( .a(TIMEBOOST_net_11849), .b(g65744_db), .o(n_1927) );
in01f02 g57174_u0 ( .a(FE_OFN1427_n_8567), .o(g57174_sb) );
na02s01 TIMEBOOST_cell_31025 ( .a(TIMEBOOST_net_9423), .b(g64842_db), .o(n_4439) );
na02s02 TIMEBOOST_cell_43682 ( .a(TIMEBOOST_net_14079), .b(g58633_db), .o(n_8848) );
na02s02 TIMEBOOST_cell_45630 ( .a(TIMEBOOST_net_15053), .b(n_4450), .o(n_4271) );
in01f02 g57175_u0 ( .a(FE_OFN2177_n_8567), .o(g57175_sb) );
in01s01 TIMEBOOST_cell_32841 ( .a(TIMEBOOST_net_10342), .o(TIMEBOOST_net_10341) );
na03s01 TIMEBOOST_cell_5155 ( .a(g58208_sb), .b(g58208_db), .c(FE_OFN266_n_9884), .o(n_9578) );
na02s01 TIMEBOOST_cell_45332 ( .a(TIMEBOOST_net_14904), .b(g62440_sb), .o(n_6716) );
in01f01 g57176_u0 ( .a(FE_OFN1408_n_8567), .o(g57176_sb) );
na02s02 TIMEBOOST_cell_45333 ( .a(TIMEBOOST_net_4815), .b(FE_OFN1203_n_4090), .o(TIMEBOOST_net_14905) );
na02s02 TIMEBOOST_cell_40718 ( .a(TIMEBOOST_net_12597), .b(g62915_sb), .o(n_6049) );
na02s01 TIMEBOOST_cell_39224 ( .a(TIMEBOOST_net_11850), .b(g65800_db), .o(n_2004) );
in01f02 g57177_u0 ( .a(FE_OFN1370_n_8567), .o(g57177_sb) );
na02s01 TIMEBOOST_cell_44913 ( .a(TIMEBOOST_net_9515), .b(FE_OFN1043_n_2037), .o(TIMEBOOST_net_14695) );
na02s02 TIMEBOOST_cell_40720 ( .a(TIMEBOOST_net_12598), .b(g62384_sb), .o(n_6833) );
na02s01 TIMEBOOST_cell_39226 ( .a(TIMEBOOST_net_11851), .b(g65730_db), .o(n_1981) );
in01f01 g57178_u0 ( .a(FE_OFN1345_n_8567), .o(g57178_sb) );
na02f04 TIMEBOOST_cell_4141 ( .a(n_16970), .b(TIMEBOOST_net_650), .o(n_13703) );
na02f01 g57178_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__Q), .b(FE_OFN1345_n_8567), .o(g57178_db) );
na02s01 TIMEBOOST_cell_38638 ( .a(TIMEBOOST_net_11557), .b(g59113_sb), .o(n_8699) );
in01f02 g57179_u0 ( .a(FE_OFN2180_n_8567), .o(g57179_sb) );
na03s02 TIMEBOOST_cell_41993 ( .a(n_4422), .b(FE_OFN1284_n_4097), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__Q), .o(TIMEBOOST_net_13235) );
na02s02 TIMEBOOST_cell_41818 ( .a(TIMEBOOST_net_13147), .b(g58371_db), .o(n_9010) );
in01f01 g57180_u0 ( .a(FE_OFN1406_n_8567), .o(g57180_sb) );
na02s01 TIMEBOOST_cell_43198 ( .a(TIMEBOOST_net_13837), .b(FE_OFN1223_n_6391), .o(TIMEBOOST_net_12595) );
na02s02 TIMEBOOST_cell_40722 ( .a(TIMEBOOST_net_12599), .b(g62539_sb), .o(n_6490) );
na02f02 TIMEBOOST_cell_41458 ( .a(TIMEBOOST_net_12967), .b(g57366_sb), .o(n_10384) );
in01f01 g57181_u0 ( .a(FE_OFN1394_n_8567), .o(g57181_sb) );
na02s01 TIMEBOOST_cell_31280 ( .a(configuration_wb_err_cs_bit_570), .b(parchk_pci_cbe_out_in_1204), .o(TIMEBOOST_net_9551) );
na02s02 TIMEBOOST_cell_38022 ( .a(TIMEBOOST_net_11249), .b(g61827_sb), .o(n_8132) );
na02s01 TIMEBOOST_cell_31261 ( .a(TIMEBOOST_net_9541), .b(g65970_sb), .o(n_2154) );
in01f01 g57182_u0 ( .a(FE_OFN1408_n_8567), .o(g57182_sb) );
na02s02 TIMEBOOST_cell_45334 ( .a(TIMEBOOST_net_14905), .b(g63185_sb), .o(n_5782) );
na02s02 TIMEBOOST_cell_45335 ( .a(TIMEBOOST_net_4797), .b(FE_OFN1244_n_4092), .o(TIMEBOOST_net_14906) );
na02s01 TIMEBOOST_cell_4386 ( .a(g65994_sb), .b(wbu_pciif_devsel_reg_in), .o(TIMEBOOST_net_773) );
in01f01 g57183_u0 ( .a(FE_OFN1387_n_8567), .o(g57183_sb) );
na02s01 TIMEBOOST_cell_43199 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__Q), .b(n_4917), .o(TIMEBOOST_net_13838) );
na02f02 TIMEBOOST_cell_41452 ( .a(TIMEBOOST_net_12964), .b(g57554_sb), .o(n_10302) );
na02m02 TIMEBOOST_cell_42259 ( .a(n_9756), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__Q), .o(TIMEBOOST_net_13368) );
in01f01 g57184_u0 ( .a(FE_OFN1349_n_8567), .o(g57184_sb) );
na02m02 TIMEBOOST_cell_44403 ( .a(n_9582), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__Q), .o(TIMEBOOST_net_14440) );
in01s01 TIMEBOOST_cell_45925 ( .a(wbm_dat_i_21_), .o(TIMEBOOST_net_15232) );
na02f02 TIMEBOOST_cell_42957 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_413), .b(g54149_sb), .o(TIMEBOOST_net_13717) );
in01f01 g57185_u0 ( .a(FE_OFN1391_n_8567), .o(g57185_sb) );
na02s02 TIMEBOOST_cell_45336 ( .a(TIMEBOOST_net_14906), .b(g62710_sb), .o(n_6150) );
na02m02 TIMEBOOST_cell_41629 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_2__Q), .b(FE_OFN237_n_9118), .o(TIMEBOOST_net_13053) );
na02s02 TIMEBOOST_cell_4390 ( .a(n_188), .b(n_5757), .o(TIMEBOOST_net_775) );
in01f01 g57186_u0 ( .a(FE_OFN1406_n_8567), .o(g57186_sb) );
na02s01 TIMEBOOST_cell_31148 ( .a(n_3774), .b(g64886_sb), .o(TIMEBOOST_net_9485) );
na02s02 TIMEBOOST_cell_43200 ( .a(TIMEBOOST_net_13838), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_12041) );
na02s01 TIMEBOOST_cell_39485 ( .a(wbs_dat_i_1_), .b(g63601_db), .o(TIMEBOOST_net_11981) );
in01f01 g57187_u0 ( .a(FE_OFN1392_n_8567), .o(g57187_sb) );
na02s01 TIMEBOOST_cell_31147 ( .a(TIMEBOOST_net_9484), .b(g65066_db), .o(n_3609) );
na02m04 TIMEBOOST_cell_39023 ( .a(wbs_wbb3_2_wbb2_dat_o_i_118), .b(wbs_dat_o_19_), .o(TIMEBOOST_net_11750) );
na02s02 TIMEBOOST_cell_42813 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__Q), .b(g65284_sb), .o(TIMEBOOST_net_13645) );
in01f01 g57188_u0 ( .a(FE_OFN1389_n_8567), .o(g57188_sb) );
na02s01 TIMEBOOST_cell_42674 ( .a(TIMEBOOST_net_13575), .b(g65037_db), .o(n_4331) );
na02s01 TIMEBOOST_cell_45048 ( .a(TIMEBOOST_net_14762), .b(FE_OFN719_n_8060), .o(TIMEBOOST_net_11239) );
no02s01 TIMEBOOST_cell_4392 ( .a(wbu_pciif_frame_out_in), .b(wishbone_slave_unit_pci_initiator_sm_timeout), .o(TIMEBOOST_net_776) );
in01f01 g57189_u0 ( .a(FE_OFN1387_n_8567), .o(g57189_sb) );
na03m02 TIMEBOOST_cell_45337 ( .a(g52399_db), .b(n_3478), .c(g52399_sb), .o(TIMEBOOST_net_14907) );
no02s01 TIMEBOOST_cell_4393 ( .a(TIMEBOOST_net_776), .b(n_3126), .o(g63307_p) );
na02s01 TIMEBOOST_cell_4394 ( .a(pciu_cache_lsize_not_zero_in), .b(n_16818), .o(TIMEBOOST_net_777) );
in01f01 g57190_u0 ( .a(FE_OFN1387_n_8567), .o(g57190_sb) );
na02s01 TIMEBOOST_cell_43201 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__Q), .b(n_4456), .o(TIMEBOOST_net_13839) );
na02s01 TIMEBOOST_cell_4395 ( .a(TIMEBOOST_net_777), .b(FE_OCPN1832_n_16949), .o(TIMEBOOST_net_597) );
no02s01 TIMEBOOST_cell_4396 ( .a(wishbone_slave_unit_pcim_if_del_we_in), .b(n_1014), .o(TIMEBOOST_net_778) );
in01f01 g57191_u0 ( .a(FE_OFN1382_n_8567), .o(g57191_sb) );
na02m02 TIMEBOOST_cell_45338 ( .a(TIMEBOOST_net_14907), .b(TIMEBOOST_net_590), .o(n_14821) );
no02s01 TIMEBOOST_cell_4397 ( .a(TIMEBOOST_net_778), .b(FE_OCPN1832_n_16949), .o(g61618_BP) );
na03s02 TIMEBOOST_cell_42041 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__Q), .b(n_4356), .c(FE_OFN1214_n_4151), .o(TIMEBOOST_net_13259) );
in01f01 g57192_u0 ( .a(FE_OFN1387_n_8567), .o(g57192_sb) );
na02s02 TIMEBOOST_cell_43018 ( .a(TIMEBOOST_net_13747), .b(g63051_db), .o(n_5149) );
na02s01 TIMEBOOST_cell_42593 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__Q), .b(FE_OFN519_n_9697), .o(TIMEBOOST_net_13535) );
na02s01 TIMEBOOST_cell_4400 ( .a(n_1802), .b(n_3334), .o(TIMEBOOST_net_780) );
in01f01 g57193_u0 ( .a(FE_OFN1385_n_8567), .o(g57193_sb) );
na02f02 TIMEBOOST_cell_44216 ( .a(TIMEBOOST_net_14346), .b(FE_OFN1405_n_8567), .o(TIMEBOOST_net_12885) );
na02f01 TIMEBOOST_cell_4401 ( .a(TIMEBOOST_net_780), .b(n_2410), .o(TIMEBOOST_net_260) );
na02s01 TIMEBOOST_cell_4402 ( .a(n_188), .b(n_1459), .o(TIMEBOOST_net_781) );
in01f02 g57194_u0 ( .a(FE_OFN2177_n_8567), .o(g57194_sb) );
na02m02 TIMEBOOST_cell_44225 ( .a(n_9532), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__Q), .o(TIMEBOOST_net_14351) );
na02s01 TIMEBOOST_cell_31141 ( .a(TIMEBOOST_net_9481), .b(g65916_db), .o(n_1852) );
na03s02 TIMEBOOST_cell_5160 ( .a(g65020_sb), .b(g65020_db), .c(n_4447), .o(n_4340) );
in01f01 g57195_u0 ( .a(FE_OFN1385_n_8567), .o(g57195_sb) );
na02f02 TIMEBOOST_cell_42512 ( .a(TIMEBOOST_net_13494), .b(g57046_sb), .o(n_11688) );
na02m02 TIMEBOOST_cell_32488 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q), .o(TIMEBOOST_net_10155) );
na02s01 TIMEBOOST_cell_45339 ( .a(n_2170), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__Q), .o(TIMEBOOST_net_14908) );
in01f01 g57196_u0 ( .a(FE_OFN1412_n_8567), .o(g57196_sb) );
na02m02 TIMEBOOST_cell_43863 ( .a(n_9553), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__Q), .o(TIMEBOOST_net_14170) );
na02s02 TIMEBOOST_cell_45340 ( .a(TIMEBOOST_net_14908), .b(FE_OFN706_n_8119), .o(TIMEBOOST_net_11067) );
na02f02 TIMEBOOST_cell_42504 ( .a(TIMEBOOST_net_13490), .b(g57536_sb), .o(n_11206) );
in01f01 g57197_u0 ( .a(FE_OFN1401_n_8567), .o(g57197_sb) );
na02s01 TIMEBOOST_cell_15870 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_93), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3192) );
na03s02 TIMEBOOST_cell_34246 ( .a(TIMEBOOST_net_9800), .b(FE_OFN1171_n_5592), .c(g62131_sb), .o(n_5565) );
na02s01 TIMEBOOST_cell_4408 ( .a(n_3395), .b(n_188), .o(TIMEBOOST_net_784) );
in01f01 g57198_u0 ( .a(FE_OFN1373_n_8567), .o(g57198_sb) );
na02s01 TIMEBOOST_cell_31140 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__Q), .b(g65916_sb), .o(TIMEBOOST_net_9481) );
na02s02 TIMEBOOST_cell_42973 ( .a(g61842_sb), .b(g61842_db), .o(TIMEBOOST_net_13725) );
in01f02 g57199_u0 ( .a(FE_OFN1427_n_8567), .o(g57199_sb) );
na03s02 TIMEBOOST_cell_41975 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__Q), .b(n_3538), .c(FE_OFN1295_n_4098), .o(TIMEBOOST_net_13226) );
na02s02 TIMEBOOST_cell_45341 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__Q), .b(n_4507), .o(TIMEBOOST_net_14909) );
na03s01 TIMEBOOST_cell_5162 ( .a(n_3761), .b(g64759_sb), .c(g64759_db), .o(n_3787) );
in01f01 g57200_u0 ( .a(FE_OFN1405_n_8567), .o(g57200_sb) );
na02f02 TIMEBOOST_cell_44142 ( .a(TIMEBOOST_net_14309), .b(FE_OFN1407_n_8567), .o(TIMEBOOST_net_12719) );
na02f02 TIMEBOOST_cell_44669 ( .a(TIMEBOOST_net_10054), .b(FE_OFN1407_n_8567), .o(TIMEBOOST_net_14573) );
in01f01 g57201_u0 ( .a(FE_OFN1402_n_8567), .o(g57201_sb) );
na02s01 TIMEBOOST_cell_22246 ( .a(g52465_da), .b(FE_OFN1022_n_11877), .o(TIMEBOOST_net_6380) );
na02m01 TIMEBOOST_cell_4409 ( .a(TIMEBOOST_net_784), .b(FE_OFN2121_n_2687), .o(TIMEBOOST_net_309) );
na02s02 TIMEBOOST_cell_22063 ( .a(n_10247), .b(TIMEBOOST_net_6288), .o(n_11867) );
in01f01 g57202_u0 ( .a(FE_OFN1399_n_8567), .o(g57202_sb) );
na02m02 TIMEBOOST_cell_30802 ( .a(wbu_addr_in_257), .b(g58797_sb), .o(TIMEBOOST_net_9312) );
na02m02 TIMEBOOST_cell_38783 ( .a(TIMEBOOST_net_9654), .b(FE_OFN2093_n_2301), .o(TIMEBOOST_net_11630) );
na02f02 TIMEBOOST_cell_43864 ( .a(TIMEBOOST_net_14170), .b(FE_OFN1383_n_8567), .o(TIMEBOOST_net_12828) );
in01f01 g57203_u0 ( .a(FE_OFN1394_n_8567), .o(g57203_sb) );
na02s02 TIMEBOOST_cell_43615 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__Q), .b(n_3539), .o(TIMEBOOST_net_14046) );
in01f01 g57204_u0 ( .a(FE_OFN1384_n_8567), .o(g57204_sb) );
na02s01 TIMEBOOST_cell_22248 ( .a(g52470_da), .b(FE_OFN1025_n_11877), .o(TIMEBOOST_net_6381) );
na02m02 TIMEBOOST_cell_43865 ( .a(n_9866), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__Q), .o(TIMEBOOST_net_14171) );
na02s01 TIMEBOOST_cell_4414 ( .a(n_2503), .b(g66423_db), .o(TIMEBOOST_net_787) );
in01f01 g57205_u0 ( .a(FE_OFN1412_n_8567), .o(g57205_sb) );
na02s02 TIMEBOOST_cell_43202 ( .a(TIMEBOOST_net_13839), .b(FE_OFN1246_n_4093), .o(TIMEBOOST_net_12123) );
na02s01 TIMEBOOST_cell_4415 ( .a(TIMEBOOST_net_787), .b(g66398_sb), .o(n_2504) );
no02s02 TIMEBOOST_cell_4416 ( .a(n_1827), .b(n_7114), .o(TIMEBOOST_net_788) );
in01f01 g57206_u0 ( .a(FE_OFN1400_n_8567), .o(g57206_sb) );
na02s02 TIMEBOOST_cell_45712 ( .a(TIMEBOOST_net_15094), .b(FE_OFN1248_n_4093), .o(TIMEBOOST_net_13232) );
na02f04 TIMEBOOST_cell_45836 ( .a(TIMEBOOST_net_15156), .b(FE_OFN2134_n_13124), .o(TIMEBOOST_net_14998) );
na02f02 TIMEBOOST_cell_44247 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__8__Q), .b(n_9433), .o(TIMEBOOST_net_14362) );
in01f02 g57207_u0 ( .a(FE_OFN1427_n_8567), .o(g57207_sb) );
na02f02 TIMEBOOST_cell_42438 ( .a(TIMEBOOST_net_13457), .b(g57239_sb), .o(n_10428) );
na02s02 TIMEBOOST_cell_43203 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__Q), .b(n_3530), .o(TIMEBOOST_net_13840) );
na02s02 TIMEBOOST_cell_45342 ( .a(TIMEBOOST_net_14909), .b(n_6645), .o(TIMEBOOST_net_12621) );
in01f01 g57208_u0 ( .a(FE_OFN1425_n_8567), .o(g57208_sb) );
na03f06 TIMEBOOST_cell_33262 ( .a(n_16156), .b(pci_target_unit_wishbone_master_burst_chopped), .c(n_15388), .o(n_15389) );
na02s01 TIMEBOOST_cell_17657 ( .a(TIMEBOOST_net_4085), .b(g65404_db), .o(n_4234) );
na02s02 TIMEBOOST_cell_17255 ( .a(TIMEBOOST_net_3884), .b(g65403_da), .o(n_4235) );
in01f01 g57209_u0 ( .a(FE_OFN1420_n_8567), .o(g57209_sb) );
na02m02 TIMEBOOST_cell_43598 ( .a(TIMEBOOST_net_14037), .b(FE_OFN1317_n_6624), .o(TIMEBOOST_net_12238) );
na02s01 TIMEBOOST_cell_4421 ( .a(TIMEBOOST_net_790), .b(n_2301), .o(TIMEBOOST_net_540) );
na02m02 TIMEBOOST_cell_41587 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_31__Q), .b(FE_OFN241_n_9830), .o(TIMEBOOST_net_13032) );
in01f01 g57210_u0 ( .a(FE_OFN1407_n_8567), .o(g57210_sb) );
in01f01 g57211_u0 ( .a(FE_OFN1422_n_8567), .o(g57211_sb) );
na02s01 TIMEBOOST_cell_30876 ( .a(pci_target_unit_pcit_if_strd_addr_in_699), .b(pci_target_unit_del_sync_addr_in_217), .o(TIMEBOOST_net_9349) );
na02f02 TIMEBOOST_cell_41669 ( .a(FE_OFN1775_n_13800), .b(TIMEBOOST_net_10151), .o(TIMEBOOST_net_13073) );
na02f02 TIMEBOOST_cell_32555 ( .a(n_12313), .b(TIMEBOOST_net_10188), .o(TIMEBOOST_net_6560) );
in01f01 g57212_u0 ( .a(FE_OFN1397_n_8567), .o(g57212_sb) );
na02s02 TIMEBOOST_cell_43269 ( .a(n_4500), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__13__Q), .o(TIMEBOOST_net_13873) );
na02m02 TIMEBOOST_cell_32554 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__Q), .o(TIMEBOOST_net_10188) );
no02s01 TIMEBOOST_cell_4426 ( .a(n_1667), .b(n_1995), .o(TIMEBOOST_net_793) );
in01f01 g57213_u0 ( .a(FE_OFN1374_n_8567), .o(g57213_sb) );
na02f02 TIMEBOOST_cell_41510 ( .a(TIMEBOOST_net_12993), .b(g57112_sb), .o(TIMEBOOST_net_11641) );
no02s01 TIMEBOOST_cell_4427 ( .a(TIMEBOOST_net_793), .b(FE_OFN1024_n_11877), .o(n_3453) );
na02s01 TIMEBOOST_cell_17012 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(g65798_sb), .o(TIMEBOOST_net_3763) );
in01f02 g57214_u0 ( .a(FE_OFN2168_n_8567), .o(g57214_sb) );
na02f02 TIMEBOOST_cell_41588 ( .a(FE_OFN1436_n_9372), .b(TIMEBOOST_net_13032), .o(TIMEBOOST_net_11677) );
na02m02 TIMEBOOST_cell_43684 ( .a(TIMEBOOST_net_14080), .b(g58632_db), .o(n_8849) );
na02s02 TIMEBOOST_cell_45343 ( .a(n_4915), .b(n_395), .o(TIMEBOOST_net_14910) );
in01f02 g57215_u0 ( .a(FE_OFN2168_n_8567), .o(g57215_sb) );
na02f02 TIMEBOOST_cell_44206 ( .a(TIMEBOOST_net_14341), .b(FE_OFN1374_n_8567), .o(TIMEBOOST_net_12741) );
na02s01 TIMEBOOST_cell_17013 ( .a(TIMEBOOST_net_3763), .b(g65798_db), .o(n_1665) );
na02f02 TIMEBOOST_cell_44444 ( .a(TIMEBOOST_net_14460), .b(g58589_sb), .o(n_8912) );
in01f02 g57216_u0 ( .a(FE_OFN1376_n_8567), .o(g57216_sb) );
na02s02 TIMEBOOST_cell_45217 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__Q), .b(n_4367), .o(TIMEBOOST_net_14847) );
na02s02 TIMEBOOST_cell_39632 ( .a(TIMEBOOST_net_12054), .b(g62754_sb), .o(n_6129) );
in01s01 TIMEBOOST_cell_45954 ( .a(TIMEBOOST_net_15260), .o(TIMEBOOST_net_15261) );
in01f01 g57217_u0 ( .a(FE_OFN1423_n_8567), .o(g57217_sb) );
na02f02 TIMEBOOST_cell_41512 ( .a(TIMEBOOST_net_12994), .b(g57187_sb), .o(n_11565) );
na02s02 TIMEBOOST_cell_39634 ( .a(TIMEBOOST_net_12055), .b(g62761_sb), .o(n_6119) );
na02s01 TIMEBOOST_cell_45344 ( .a(TIMEBOOST_net_14910), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_12611) );
in01f01 g57218_u0 ( .a(FE_OFN1389_n_8567), .o(g57218_sb) );
na02s02 TIMEBOOST_cell_45749 ( .a(n_4408), .b(n_0), .o(TIMEBOOST_net_15113) );
na02s01 TIMEBOOST_cell_17955 ( .a(TIMEBOOST_net_4234), .b(g65392_da), .o(n_4240) );
na02s01 TIMEBOOST_cell_17224 ( .a(n_4452), .b(FE_OFN653_n_4508), .o(TIMEBOOST_net_3869) );
in01f01 g57219_u0 ( .a(FE_OFN1349_n_8567), .o(g57219_sb) );
na02f02 TIMEBOOST_cell_4145 ( .a(TIMEBOOST_net_652), .b(FE_RN_438_0), .o(FE_RN_439_0) );
na02f02 TIMEBOOST_cell_43866 ( .a(TIMEBOOST_net_14171), .b(FE_OFN1421_n_8567), .o(TIMEBOOST_net_12924) );
na02s02 TIMEBOOST_cell_42653 ( .a(n_3783), .b(g64992_sb), .o(TIMEBOOST_net_13565) );
in01f01 g57220_u0 ( .a(FE_OFN1421_n_8567), .o(g57220_sb) );
na02s02 TIMEBOOST_cell_42949 ( .a(TIMEBOOST_net_9643), .b(FE_OFN1670_n_9477), .o(TIMEBOOST_net_13713) );
na02s01 TIMEBOOST_cell_17225 ( .a(TIMEBOOST_net_3869), .b(g65375_da), .o(n_4249) );
na02f04 TIMEBOOST_cell_43685 ( .a(TIMEBOOST_net_5574), .b(FE_OFN1712_n_13563), .o(TIMEBOOST_net_14081) );
in01f02 g57221_u0 ( .a(FE_OFN2177_n_8567), .o(g57221_sb) );
na03s02 TIMEBOOST_cell_34243 ( .a(TIMEBOOST_net_9803), .b(FE_OFN1171_n_5592), .c(g62130_sb), .o(n_5566) );
na02s01 TIMEBOOST_cell_43340 ( .a(TIMEBOOST_net_13908), .b(g62995_sb), .o(n_5892) );
na02s01 TIMEBOOST_cell_45345 ( .a(n_4347), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__Q), .o(TIMEBOOST_net_14911) );
in01f01 g57222_u0 ( .a(FE_OFN1390_n_8567), .o(g57222_sb) );
na02s01 TIMEBOOST_cell_43467 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__Q), .b(n_2379), .o(TIMEBOOST_net_13972) );
na02s01 TIMEBOOST_cell_45087 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__Q), .b(FE_OFN535_n_9823), .o(TIMEBOOST_net_14782) );
in01f01 g57223_u0 ( .a(FE_OFN1407_n_8567), .o(g57223_sb) );
na02f02 TIMEBOOST_cell_43294 ( .a(TIMEBOOST_net_13885), .b(FE_OFN1699_n_5751), .o(TIMEBOOST_net_11525) );
na02s01 TIMEBOOST_cell_4439 ( .a(TIMEBOOST_net_799), .b(n_4177), .o(n_4711) );
na02f01 TIMEBOOST_cell_4440 ( .a(n_1805), .b(FE_OFN2121_n_2687), .o(TIMEBOOST_net_800) );
in01f02 g57224_u0 ( .a(FE_OFN2187_n_8567), .o(g57224_sb) );
na02f02 TIMEBOOST_cell_41564 ( .a(TIMEBOOST_net_13020), .b(g57229_sb), .o(n_11526) );
na02s02 TIMEBOOST_cell_43204 ( .a(TIMEBOOST_net_13840), .b(FE_OFN1242_n_4092), .o(TIMEBOOST_net_11543) );
na03s02 TIMEBOOST_cell_5170 ( .a(n_3752), .b(g64806_sb), .c(g64806_db), .o(n_3753) );
in01f02 g57225_u0 ( .a(FE_OFN2189_n_8567), .o(g57225_sb) );
na03m06 TIMEBOOST_cell_32932 ( .a(n_1629), .b(TIMEBOOST_net_3218), .c(n_1551), .o(TIMEBOOST_net_627) );
na02s01 TIMEBOOST_cell_45346 ( .a(TIMEBOOST_net_14911), .b(n_6287), .o(TIMEBOOST_net_12625) );
na02f02 TIMEBOOST_cell_22560 ( .a(FE_OFN1739_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__Q), .o(TIMEBOOST_net_6537) );
in01f01 g57226_u0 ( .a(FE_OFN1397_n_8567), .o(g57226_sb) );
na02f02 TIMEBOOST_cell_41540 ( .a(TIMEBOOST_net_13008), .b(g57464_sb), .o(n_11268) );
na02m04 TIMEBOOST_cell_4441 ( .a(TIMEBOOST_net_800), .b(FE_OFN2052_n_6965), .o(TIMEBOOST_net_472) );
na02s01 TIMEBOOST_cell_4442 ( .a(FE_OFN785_n_2678), .b(pci_target_unit_pcit_if_strd_addr_in_701), .o(TIMEBOOST_net_801) );
in01f01 g57227_u0 ( .a(FE_OFN1387_n_8567), .o(g57227_sb) );
na02f02 TIMEBOOST_cell_41508 ( .a(TIMEBOOST_net_12992), .b(g57362_sb), .o(n_10385) );
na02s01 TIMEBOOST_cell_17043 ( .a(TIMEBOOST_net_3778), .b(g64957_db), .o(n_3661) );
na02s02 TIMEBOOST_cell_38722 ( .a(TIMEBOOST_net_11599), .b(g62523_sb), .o(n_6530) );
in01f01 g57228_u0 ( .a(FE_OFN1385_n_8567), .o(g57228_sb) );
na02f02 TIMEBOOST_cell_44366 ( .a(TIMEBOOST_net_14421), .b(FE_OFN1396_n_8567), .o(TIMEBOOST_net_12715) );
na02m02 TIMEBOOST_cell_18063 ( .a(TIMEBOOST_net_4288), .b(g54235_sb), .o(n_13439) );
na02f02 TIMEBOOST_cell_42274 ( .a(TIMEBOOST_net_13375), .b(g57118_sb), .o(n_11628) );
in01f02 g57229_u0 ( .a(FE_OFN2177_n_8567), .o(g57229_sb) );
na03f08 TIMEBOOST_cell_32931 ( .a(n_7044), .b(n_2883), .c(FE_RN_533_0), .o(n_15402) );
na02s01 TIMEBOOST_cell_43205 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__Q), .b(n_4307), .o(TIMEBOOST_net_13841) );
na02s02 TIMEBOOST_cell_45347 ( .a(n_3767), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__Q), .o(TIMEBOOST_net_14912) );
in01f02 g57230_u0 ( .a(FE_OFN2179_n_8567), .o(g57230_sb) );
na02f02 TIMEBOOST_cell_44656 ( .a(TIMEBOOST_net_14566), .b(FE_OFN1377_n_8567), .o(TIMEBOOST_net_12786) );
in01f01 g57231_u0 ( .a(FE_OFN1413_n_8567), .o(g57231_sb) );
na02m02 TIMEBOOST_cell_43867 ( .a(n_9063), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__Q), .o(TIMEBOOST_net_14172) );
na02s01 TIMEBOOST_cell_37179 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_10828) );
na02s02 TIMEBOOST_cell_38156 ( .a(TIMEBOOST_net_11316), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_4536) );
in01f02 g57232_u0 ( .a(FE_OFN2174_n_8567), .o(g57232_sb) );
na02s02 TIMEBOOST_cell_45348 ( .a(TIMEBOOST_net_14912), .b(FE_OFN1250_n_4093), .o(TIMEBOOST_net_12521) );
na02s01 TIMEBOOST_cell_31129 ( .a(TIMEBOOST_net_9475), .b(g64767_db), .o(n_4487) );
na02s02 TIMEBOOST_cell_45349 ( .a(n_83), .b(n_3613), .o(TIMEBOOST_net_14913) );
in01f01 g57233_u0 ( .a(FE_OFN1401_n_8567), .o(g57233_sb) );
na02s01 TIMEBOOST_cell_18067 ( .a(TIMEBOOST_net_4290), .b(g61867_sb), .o(n_8102) );
na03s02 TIMEBOOST_cell_34033 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(g63544_sb), .c(g63544_db), .o(n_4612) );
in01f02 g57234_u0 ( .a(FE_OFN2178_n_8567), .o(g57234_sb) );
na02f02 TIMEBOOST_cell_41552 ( .a(TIMEBOOST_net_13014), .b(g57591_sb), .o(n_10288) );
na02s01 TIMEBOOST_cell_31128 ( .a(g64767_sb), .b(n_4498), .o(TIMEBOOST_net_9475) );
in01f02 g57235_u0 ( .a(FE_OFN2174_n_8567), .o(g57235_sb) );
na02f02 TIMEBOOST_cell_41480 ( .a(TIMEBOOST_net_12978), .b(g57545_sb), .o(n_11198) );
na02s02 TIMEBOOST_cell_44432 ( .a(TIMEBOOST_net_14454), .b(FE_OFN1305_n_13124), .o(TIMEBOOST_net_13419) );
in01f01 g57236_u0 ( .a(FE_OFN1377_n_8567), .o(g57236_sb) );
na02s02 TIMEBOOST_cell_45350 ( .a(TIMEBOOST_net_14913), .b(FE_OFN1232_n_6391), .o(TIMEBOOST_net_12640) );
na03s01 TIMEBOOST_cell_38127 ( .a(g64167_da), .b(g64167_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__Q), .o(TIMEBOOST_net_11302) );
na02s02 TIMEBOOST_cell_39163 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_26__Q), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_409), .o(TIMEBOOST_net_11820) );
in01f01 g57237_u0 ( .a(FE_OFN1399_n_8567), .o(g57237_sb) );
na02f02 TIMEBOOST_cell_22269 ( .a(TIMEBOOST_net_6391), .b(n_9265), .o(n_12145) );
na02s02 TIMEBOOST_cell_38158 ( .a(TIMEBOOST_net_11317), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_4527) );
na03s02 TIMEBOOST_cell_34034 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(g65680_sb), .c(g65680_db), .o(n_3215) );
in01f01 g57238_u0 ( .a(FE_OFN1396_n_8567), .o(g57238_sb) );
na02s01 TIMEBOOST_cell_31125 ( .a(TIMEBOOST_net_9473), .b(g64868_sb), .o(n_3712) );
na02m02 TIMEBOOST_cell_44545 ( .a(n_9430), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__Q), .o(TIMEBOOST_net_14511) );
na02f02 TIMEBOOST_cell_43868 ( .a(TIMEBOOST_net_14172), .b(FE_OFN1380_n_8567), .o(TIMEBOOST_net_12953) );
in01f02 g57239_u0 ( .a(FE_OFN2169_n_8567), .o(g57239_sb) );
na02s01 TIMEBOOST_cell_45578 ( .a(TIMEBOOST_net_15027), .b(n_4493), .o(TIMEBOOST_net_10913) );
na02s01 TIMEBOOST_cell_31123 ( .a(TIMEBOOST_net_9472), .b(g64876_db), .o(n_4420) );
na02s01 TIMEBOOST_cell_31122 ( .a(g64876_sb), .b(n_4498), .o(TIMEBOOST_net_9472) );
in01f01 g57240_u0 ( .a(FE_OFN1382_n_8567), .o(g57240_sb) );
na02m02 TIMEBOOST_cell_44367 ( .a(n_9525), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__Q), .o(TIMEBOOST_net_14422) );
na02f02 TIMEBOOST_cell_18071 ( .a(TIMEBOOST_net_4292), .b(g54239_sb), .o(n_13435) );
na02s02 TIMEBOOST_cell_45351 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__Q), .b(n_3684), .o(TIMEBOOST_net_14914) );
in01f01 g57241_u0 ( .a(FE_OFN1397_n_8567), .o(g57241_sb) );
in01s01 TIMEBOOST_cell_45955 ( .a(wbm_dat_i_6_), .o(TIMEBOOST_net_15262) );
na02s02 TIMEBOOST_cell_4457 ( .a(TIMEBOOST_net_808), .b(FE_OFN2245_n_4792), .o(n_7210) );
na02f02 TIMEBOOST_cell_4458 ( .a(n_1798), .b(n_3341), .o(TIMEBOOST_net_809) );
in01f02 g57242_u0 ( .a(FE_OFN2173_n_8567), .o(g57242_sb) );
na02s01 TIMEBOOST_cell_45631 ( .a(g64281_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__21__Q), .o(TIMEBOOST_net_15054) );
na02f02 TIMEBOOST_cell_22147 ( .a(TIMEBOOST_net_6330), .b(FE_OFN1600_n_13995), .o(n_16242) );
na04m04 TIMEBOOST_cell_35819 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_14__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_779), .c(FE_OFN2135_n_13124), .d(g54343_sb), .o(n_12970) );
in01f01 g57243_u0 ( .a(FE_OFN1408_n_8567), .o(g57243_sb) );
na03f02 TIMEBOOST_cell_22240 ( .a(n_10554), .b(n_10556), .c(n_9971), .o(TIMEBOOST_net_6377) );
na02f01 TIMEBOOST_cell_4459 ( .a(TIMEBOOST_net_809), .b(n_7321), .o(TIMEBOOST_net_322) );
na02m01 TIMEBOOST_cell_4460 ( .a(n_16451), .b(FE_OCPN1875_n_14526), .o(TIMEBOOST_net_810) );
in01f01 g57244_u0 ( .a(FE_OFN1420_n_8567), .o(g57244_sb) );
na02m02 TIMEBOOST_cell_43869 ( .a(n_9877), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__Q), .o(TIMEBOOST_net_14173) );
na02f01 TIMEBOOST_cell_4461 ( .a(n_16452), .b(TIMEBOOST_net_810), .o(TIMEBOOST_net_600) );
na02f01 TIMEBOOST_cell_4462 ( .a(n_16452), .b(n_7622), .o(TIMEBOOST_net_811) );
in01f02 g57245_u0 ( .a(FE_OFN2177_n_8567), .o(g57245_sb) );
na02s01 TIMEBOOST_cell_44868 ( .a(TIMEBOOST_net_14672), .b(g65274_sb), .o(TIMEBOOST_net_12403) );
na02s01 TIMEBOOST_cell_31119 ( .a(TIMEBOOST_net_9470), .b(g65054_db), .o(n_3617) );
in01f01 g57246_u0 ( .a(FE_OFN1423_n_8567), .o(g57246_sb) );
na02f02 TIMEBOOST_cell_41128 ( .a(TIMEBOOST_net_12802), .b(g57458_sb), .o(n_10346) );
na02f01 TIMEBOOST_cell_4463 ( .a(TIMEBOOST_net_811), .b(n_7725), .o(TIMEBOOST_net_582) );
na02s02 TIMEBOOST_cell_45352 ( .a(TIMEBOOST_net_14914), .b(FE_OFN1232_n_6391), .o(TIMEBOOST_net_12638) );
in01f01 g57247_u0 ( .a(FE_OFN1397_n_8567), .o(g57247_sb) );
na02m02 TIMEBOOST_cell_44143 ( .a(n_9037), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__Q), .o(TIMEBOOST_net_14310) );
na04m02 TIMEBOOST_cell_7759 ( .a(TIMEBOOST_net_595), .b(n_3134), .c(g52443_sb), .d(g52443_db), .o(n_14808) );
na02s01 TIMEBOOST_cell_9756 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__Q), .b(g65978_sb), .o(TIMEBOOST_net_1445) );
in01f01 g57248_u0 ( .a(FE_OFN1385_n_8567), .o(g57248_sb) );
na02s01 TIMEBOOST_cell_43403 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__Q), .b(n_3681), .o(TIMEBOOST_net_13940) );
na02s01 TIMEBOOST_cell_9757 ( .a(TIMEBOOST_net_1445), .b(g65978_db), .o(n_1836) );
na02s01 TIMEBOOST_cell_40391 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__Q), .b(g65366_sb), .o(TIMEBOOST_net_12434) );
in01f02 g57249_u0 ( .a(FE_OFN2180_n_8567), .o(g57249_sb) );
na02f02 TIMEBOOST_cell_41566 ( .a(TIMEBOOST_net_13021), .b(g57518_sb), .o(n_11222) );
na02s02 TIMEBOOST_cell_45353 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__Q), .b(n_3610), .o(TIMEBOOST_net_14915) );
na02s01 TIMEBOOST_cell_31118 ( .a(n_3752), .b(g65054_sb), .o(TIMEBOOST_net_9470) );
in01f01 g57250_u0 ( .a(FE_OFN1384_n_8567), .o(g57250_sb) );
na02s02 TIMEBOOST_cell_45354 ( .a(TIMEBOOST_net_14915), .b(FE_OFN1232_n_6391), .o(TIMEBOOST_net_12637) );
na02s01 TIMEBOOST_cell_42594 ( .a(TIMEBOOST_net_13535), .b(g58149_sb), .o(TIMEBOOST_net_11940) );
na02s01 TIMEBOOST_cell_9760 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__Q), .b(g65818_sb), .o(TIMEBOOST_net_1447) );
in01f01 g57251_u0 ( .a(FE_OFN1376_n_8567), .o(g57251_sb) );
na02s01 TIMEBOOST_cell_22250 ( .a(g52469_da), .b(FE_OFN1022_n_11877), .o(TIMEBOOST_net_6382) );
na02s01 TIMEBOOST_cell_9761 ( .a(TIMEBOOST_net_1447), .b(g65818_db), .o(n_1898) );
na02s01 TIMEBOOST_cell_39551 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__Q), .b(g58295_sb), .o(TIMEBOOST_net_12014) );
in01f01 g57252_u0 ( .a(FE_OFN1399_n_8567), .o(g57252_sb) );
na02f04 TIMEBOOST_cell_44780 ( .a(TIMEBOOST_net_14628), .b(n_16352), .o(TIMEBOOST_net_3293) );
na02s02 TIMEBOOST_cell_39636 ( .a(TIMEBOOST_net_12056), .b(g62419_sb), .o(n_6759) );
na02s01 TIMEBOOST_cell_40321 ( .a(n_4493), .b(g65031_sb), .o(TIMEBOOST_net_12399) );
in01f01 g57253_u0 ( .a(FE_OFN1387_n_8567), .o(g57253_sb) );
na03f02 TIMEBOOST_cell_22270 ( .a(n_16844), .b(n_9993), .c(n_16845), .o(TIMEBOOST_net_6392) );
na02s02 TIMEBOOST_cell_39638 ( .a(TIMEBOOST_net_12057), .b(g62675_sb), .o(n_6189) );
na02f02 TIMEBOOST_cell_36676 ( .a(TIMEBOOST_net_10576), .b(FE_OFN2128_n_16497), .o(n_13028) );
in01f01 g57254_u0 ( .a(FE_OFN1374_n_8567), .o(g57254_sb) );
na02s01 TIMEBOOST_cell_44914 ( .a(TIMEBOOST_net_14695), .b(g65837_sb), .o(TIMEBOOST_net_333) );
na02f02 TIMEBOOST_cell_36677 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_411), .b(TIMEBOOST_net_477), .o(TIMEBOOST_net_10577) );
na02f02 TIMEBOOST_cell_36678 ( .a(TIMEBOOST_net_10577), .b(g54146_sb), .o(n_13454) );
in01f01 g57255_u0 ( .a(FE_OFN1421_n_8567), .o(g57255_sb) );
na02s02 TIMEBOOST_cell_40848 ( .a(TIMEBOOST_net_12662), .b(FE_OFN1327_n_13547), .o(TIMEBOOST_net_11618) );
na02s01 TIMEBOOST_cell_36679 ( .a(parchk_pci_trdy_reg_in), .b(g66000_db), .o(TIMEBOOST_net_10578) );
na02s01 TIMEBOOST_cell_44915 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__Q), .b(g65363_sb), .o(TIMEBOOST_net_14696) );
in01f02 g57256_u0 ( .a(FE_OFN2177_n_8567), .o(g57256_sb) );
na03s02 TIMEBOOST_cell_41967 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__1__Q), .b(n_3759), .c(FE_OFN1219_n_6886), .o(TIMEBOOST_net_13222) );
na02s01 TIMEBOOST_cell_39640 ( .a(TIMEBOOST_net_12058), .b(g63171_sb), .o(n_5800) );
na02f02 TIMEBOOST_cell_36944 ( .a(TIMEBOOST_net_10710), .b(n_14971), .o(TIMEBOOST_net_6266) );
in01f01 g57257_u0 ( .a(FE_OFN1412_n_8567), .o(g57257_sb) );
na02s01 TIMEBOOST_cell_30848 ( .a(n_3783), .b(g65021_sb), .o(TIMEBOOST_net_9335) );
no02f02 TIMEBOOST_cell_36945 ( .a(TIMEBOOST_net_4765), .b(FE_RN_562_0), .o(TIMEBOOST_net_10711) );
na02f02 TIMEBOOST_cell_4484 ( .a(n_4814), .b(n_16914), .o(TIMEBOOST_net_822) );
in01f02 g57258_u0 ( .a(FE_OFN2179_n_8567), .o(g57258_sb) );
na02s02 TIMEBOOST_cell_45355 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__Q), .b(n_3622), .o(TIMEBOOST_net_14916) );
in01f02 g57259_u0 ( .a(FE_OFN2187_n_8567), .o(g57259_sb) );
na04m04 TIMEBOOST_cell_32974 ( .a(g58777_sb), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_19__Q), .c(n_8884), .d(wbu_addr_in_268), .o(n_9849) );
na02s01 TIMEBOOST_cell_31115 ( .a(TIMEBOOST_net_9468), .b(g64968_db), .o(n_4373) );
na02s01 TIMEBOOST_cell_31114 ( .a(n_4473), .b(g64968_sb), .o(TIMEBOOST_net_9468) );
in01f01 g57260_u0 ( .a(FE_OFN1422_n_8567), .o(g57260_sb) );
in01f01 g57261_u0 ( .a(FE_OFN1397_n_8567), .o(g57261_sb) );
na02s01 TIMEBOOST_cell_22278 ( .a(g52458_da), .b(FE_OFN1023_n_11877), .o(TIMEBOOST_net_6396) );
na02f02 TIMEBOOST_cell_4485 ( .a(TIMEBOOST_net_822), .b(n_7038), .o(TIMEBOOST_net_480) );
na02f02 TIMEBOOST_cell_43870 ( .a(TIMEBOOST_net_14173), .b(FE_OFN1385_n_8567), .o(TIMEBOOST_net_12770) );
in01f01 g57262_u0 ( .a(FE_OFN1386_n_8567), .o(g57262_sb) );
na02m02 TIMEBOOST_cell_43871 ( .a(n_9602), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__Q), .o(TIMEBOOST_net_14174) );
na02m02 TIMEBOOST_cell_43751 ( .a(n_9093), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__Q), .o(TIMEBOOST_net_14114) );
in01f01 g57263_u0 ( .a(FE_OFN1374_n_8567), .o(g57263_sb) );
na02s01 TIMEBOOST_cell_22280 ( .a(g52457_da), .b(FE_OFN1025_n_11877), .o(TIMEBOOST_net_6397) );
na02s01 TIMEBOOST_cell_9211 ( .a(TIMEBOOST_net_1172), .b(g65850_sb), .o(n_1585) );
na02s02 TIMEBOOST_cell_40461 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__Q), .b(g58288_sb), .o(TIMEBOOST_net_12469) );
in01f01 g57264_u0 ( .a(FE_OFN1384_n_8567), .o(g57264_sb) );
na02s01 TIMEBOOST_cell_30844 ( .a(n_3792), .b(g64903_sb), .o(TIMEBOOST_net_9333) );
na02s02 TIMEBOOST_cell_40450 ( .a(TIMEBOOST_net_12463), .b(g62117_sb), .o(TIMEBOOST_net_11380) );
na02f02 TIMEBOOST_cell_43872 ( .a(TIMEBOOST_net_14174), .b(FE_OFN1383_n_8567), .o(TIMEBOOST_net_12919) );
in01f01 g57265_u0 ( .a(FE_OFN1407_n_8567), .o(g57265_sb) );
na02m02 TIMEBOOST_cell_44509 ( .a(n_9008), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__Q), .o(TIMEBOOST_net_14493) );
na02s01 TIMEBOOST_cell_39267 ( .a(pci_target_unit_fifos_pciw_addr_data_in_123), .b(g64166_sb), .o(TIMEBOOST_net_11872) );
in01f01 g57266_u0 ( .a(FE_OFN1392_n_8567), .o(g57266_sb) );
na02m02 TIMEBOOST_cell_32536 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__Q), .o(TIMEBOOST_net_10179) );
na02s01 TIMEBOOST_cell_39228 ( .a(TIMEBOOST_net_11852), .b(g65804_db), .o(n_1906) );
na02m02 TIMEBOOST_cell_4496 ( .a(n_4822), .b(n_13732), .o(TIMEBOOST_net_828) );
in01f01 g57267_u0 ( .a(FE_OFN1392_n_8567), .o(g57267_sb) );
na02m02 TIMEBOOST_cell_43873 ( .a(n_9863), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__Q), .o(TIMEBOOST_net_14175) );
na02f04 TIMEBOOST_cell_37796 ( .a(TIMEBOOST_net_11136), .b(FE_RN_413_0), .o(TIMEBOOST_net_6209) );
in01f02 g57268_u0 ( .a(FE_OFN2170_n_8567), .o(g57268_sb) );
na02s02 TIMEBOOST_cell_41962 ( .a(TIMEBOOST_net_13219), .b(g62698_sb), .o(n_6158) );
na02s02 TIMEBOOST_cell_31111 ( .a(TIMEBOOST_net_9466), .b(g65058_db), .o(n_4318) );
na02s02 TIMEBOOST_cell_31110 ( .a(n_4493), .b(g65058_sb), .o(TIMEBOOST_net_9466) );
in01f01 g57269_u0 ( .a(FE_OFN1399_n_8567), .o(g57269_sb) );
na02f02 TIMEBOOST_cell_43874 ( .a(TIMEBOOST_net_14175), .b(FE_OFN1404_n_8567), .o(TIMEBOOST_net_12861) );
na02s02 TIMEBOOST_cell_4499 ( .a(TIMEBOOST_net_829), .b(n_3832), .o(n_4884) );
na02s01 TIMEBOOST_cell_39229 ( .a(pci_target_unit_fifos_pcir_control_in_192), .b(g64142_sb), .o(TIMEBOOST_net_11853) );
in01f01 g57270_u0 ( .a(FE_OFN1396_n_8567), .o(g57270_sb) );
na02s01 TIMEBOOST_cell_31109 ( .a(TIMEBOOST_net_9465), .b(g64979_db), .o(n_4366) );
na02s01 TIMEBOOST_cell_21976 ( .a(g52480_da), .b(FE_OFN9_n_11877), .o(TIMEBOOST_net_6245) );
na02s01 TIMEBOOST_cell_31108 ( .a(n_4476), .b(g64979_sb), .o(TIMEBOOST_net_9465) );
in01f02 g57271_u0 ( .a(FE_OFN2170_n_8567), .o(g57271_sb) );
na04m04 TIMEBOOST_cell_32972 ( .a(g58768_sb), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_10__Q), .c(n_8884), .d(wbu_addr_in_259), .o(n_9862) );
na03s02 TIMEBOOST_cell_43019 ( .a(n_4739), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__Q), .c(FE_OFN1119_g64577_p), .o(TIMEBOOST_net_13748) );
na02m02 TIMEBOOST_cell_22426 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__Q), .o(TIMEBOOST_net_6470) );
in01f02 g57272_u0 ( .a(FE_OFN1382_n_8567), .o(g57272_sb) );
na02m02 TIMEBOOST_cell_43875 ( .a(n_9793), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__Q), .o(TIMEBOOST_net_14176) );
na02s01 TIMEBOOST_cell_39230 ( .a(TIMEBOOST_net_11853), .b(g64142_db), .o(n_4523) );
na02s01 TIMEBOOST_cell_36680 ( .a(TIMEBOOST_net_10578), .b(g67051_sb), .o(n_2718) );
in01f01 g57273_u0 ( .a(FE_OFN1399_n_8567), .o(g57273_sb) );
na02f02 TIMEBOOST_cell_38923 ( .a(n_2719), .b(wbu_addr_in_261), .o(TIMEBOOST_net_11700) );
na02s02 TIMEBOOST_cell_43295 ( .a(n_7078), .b(n_9), .o(TIMEBOOST_net_13886) );
na02s01 TIMEBOOST_cell_36682 ( .a(TIMEBOOST_net_10579), .b(g62808_sb), .o(TIMEBOOST_net_4407) );
in01f01 g57274_u0 ( .a(FE_OFN1420_n_8567), .o(g57274_sb) );
na02s01 TIMEBOOST_cell_30886 ( .a(pci_target_unit_pcit_if_strd_addr_in_708), .b(pci_target_unit_del_sync_addr_in_226), .o(TIMEBOOST_net_9354) );
na04f02 TIMEBOOST_cell_34897 ( .a(TIMEBOOST_net_609), .b(g52402_sb), .c(g52445_db), .d(n_3357), .o(n_14847) );
na02s01 TIMEBOOST_cell_36684 ( .a(TIMEBOOST_net_10580), .b(g62757_sb), .o(TIMEBOOST_net_5293) );
in01f01 g57275_u0 ( .a(FE_OFN1423_n_8567), .o(g57275_sb) );
na02f02 TIMEBOOST_cell_44510 ( .a(TIMEBOOST_net_14493), .b(FE_OFN2168_n_8567), .o(TIMEBOOST_net_13453) );
na02s01 TIMEBOOST_cell_45027 ( .a(pci_target_unit_fifos_pciw_addr_data_in_125), .b(g64117_sb), .o(TIMEBOOST_net_14752) );
na02m02 TIMEBOOST_cell_4508 ( .a(n_13745), .b(n_15405), .o(TIMEBOOST_net_834) );
in01f01 g57276_u0 ( .a(FE_OFN1421_n_8567), .o(g57276_sb) );
na02s02 TIMEBOOST_cell_45707 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__Q), .b(n_3668), .o(TIMEBOOST_net_15092) );
na02m02 TIMEBOOST_cell_4509 ( .a(FE_OCPN1836_n_16798), .b(TIMEBOOST_net_834), .o(TIMEBOOST_net_583) );
na02f02 TIMEBOOST_cell_41450 ( .a(TIMEBOOST_net_12963), .b(g57460_sb), .o(n_10344) );
in01f01 g57277_u0 ( .a(FE_OFN1404_n_8567), .o(g57277_sb) );
na02s01 TIMEBOOST_cell_43404 ( .a(TIMEBOOST_net_13940), .b(n_6232), .o(TIMEBOOST_net_11571) );
na02s02 TIMEBOOST_cell_45356 ( .a(TIMEBOOST_net_14916), .b(FE_OFN1235_n_6391), .o(TIMEBOOST_net_12628) );
na02f02 TIMEBOOST_cell_22628 ( .a(FE_OFN1735_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__Q), .o(TIMEBOOST_net_6571) );
in01f01 g57278_u0 ( .a(FE_OFN1425_n_8567), .o(g57278_sb) );
na02f02 TIMEBOOST_cell_22359 ( .a(TIMEBOOST_net_6436), .b(n_17045), .o(n_12164) );
na02f02 TIMEBOOST_cell_41468 ( .a(TIMEBOOST_net_12972), .b(g57307_sb), .o(n_11443) );
na02f02 TIMEBOOST_cell_41430 ( .a(TIMEBOOST_net_12953), .b(g57304_sb), .o(n_10404) );
in01m01 g57279_u0 ( .a(FE_OFN1381_n_8567), .o(g57279_sb) );
na02f02 TIMEBOOST_cell_43876 ( .a(TIMEBOOST_net_14176), .b(FE_OFN1417_n_8567), .o(TIMEBOOST_net_12859) );
na02s02 TIMEBOOST_cell_45357 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__Q), .b(n_4271), .o(TIMEBOOST_net_14917) );
na02s02 TIMEBOOST_cell_42950 ( .a(TIMEBOOST_net_13713), .b(g58366_sb), .o(n_9013) );
in01f01 g57280_u0 ( .a(FE_OFN1415_n_8567), .o(g57280_sb) );
na02s02 TIMEBOOST_cell_42742 ( .a(TIMEBOOST_net_13609), .b(g65394_db), .o(n_3522) );
na02f02 TIMEBOOST_cell_41478 ( .a(TIMEBOOST_net_12977), .b(g57355_sb), .o(n_11393) );
no02f02 TIMEBOOST_cell_32803 ( .a(TIMEBOOST_net_10312), .b(n_12816), .o(FE_RN_23_0) );
in01f02 g57281_u0 ( .a(FE_OFN2169_n_8567), .o(g57281_sb) );
na02s02 TIMEBOOST_cell_41714 ( .a(TIMEBOOST_net_13095), .b(g56934_sb), .o(TIMEBOOST_net_10092) );
na02f02 TIMEBOOST_cell_22427 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_6470), .o(TIMEBOOST_net_3085) );
na02s01 TIMEBOOST_cell_43020 ( .a(TIMEBOOST_net_13748), .b(g62753_sb), .o(n_7134) );
in01f01 g57282_u0 ( .a(FE_OFN1405_n_8567), .o(g57282_sb) );
na02s02 TIMEBOOST_cell_30893 ( .a(TIMEBOOST_net_9357), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_3741) );
na02s02 TIMEBOOST_cell_45358 ( .a(TIMEBOOST_net_14917), .b(FE_OFN1235_n_6391), .o(TIMEBOOST_net_12635) );
no02f02 TIMEBOOST_cell_32802 ( .a(n_12920), .b(n_12707), .o(TIMEBOOST_net_10312) );
in01f02 g57283_u0 ( .a(FE_OFN2182_n_8567), .o(g57283_sb) );
na02m02 TIMEBOOST_cell_44649 ( .a(n_9484), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q), .o(TIMEBOOST_net_14563) );
na02f02 TIMEBOOST_cell_43752 ( .a(TIMEBOOST_net_14114), .b(FE_OFN1389_n_8567), .o(TIMEBOOST_net_12834) );
na02s01 TIMEBOOST_cell_31102 ( .a(n_3774), .b(g64815_sb), .o(TIMEBOOST_net_9462) );
in01f02 g57284_u0 ( .a(FE_OFN2188_n_8567), .o(g57284_sb) );
na02f02 TIMEBOOST_cell_41522 ( .a(TIMEBOOST_net_12999), .b(g57341_sb), .o(n_11410) );
na02f02 TIMEBOOST_cell_41610 ( .a(FE_OFN1436_n_9372), .b(TIMEBOOST_net_13043), .o(TIMEBOOST_net_11650) );
na02s02 TIMEBOOST_cell_31101 ( .a(TIMEBOOST_net_9461), .b(g64764_sb), .o(n_3784) );
in01f01 g57285_u0 ( .a(FE_OFN1345_n_8567), .o(g57285_sb) );
na02f02 TIMEBOOST_cell_4147 ( .a(TIMEBOOST_net_653), .b(n_5717), .o(n_7312) );
na02m02 TIMEBOOST_cell_43877 ( .a(n_9731), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__Q), .o(TIMEBOOST_net_14177) );
na02f02 TIMEBOOST_cell_4148 ( .a(n_2839), .b(n_2969), .o(TIMEBOOST_net_654) );
in01f01 g57286_u0 ( .a(FE_OFN1390_n_8567), .o(g57286_sb) );
na02m04 TIMEBOOST_cell_22312 ( .a(g52464_da), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_6413) );
na02s02 TIMEBOOST_cell_45359 ( .a(n_4257), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__18__Q), .o(TIMEBOOST_net_14918) );
na03f04 TIMEBOOST_cell_32800 ( .a(n_11805), .b(n_11903), .c(n_12203), .o(TIMEBOOST_net_10311) );
in01f01 g57287_u0 ( .a(FE_OFN1411_n_8567), .o(g57287_sb) );
na02s01 TIMEBOOST_cell_30894 ( .a(pci_target_unit_pcit_if_strd_addr_in_700), .b(pci_target_unit_del_sync_addr_in_218), .o(TIMEBOOST_net_9358) );
na02f02 TIMEBOOST_cell_41432 ( .a(TIMEBOOST_net_12954), .b(g57226_sb), .o(n_10434) );
na02s02 TIMEBOOST_cell_45360 ( .a(TIMEBOOST_net_14918), .b(FE_OFN1231_n_6391), .o(TIMEBOOST_net_13287) );
in01f01 g57288_u0 ( .a(FE_OFN1407_n_8567), .o(g57288_sb) );
na02f02 TIMEBOOST_cell_44412 ( .a(TIMEBOOST_net_14444), .b(FE_OFN1413_n_8567), .o(TIMEBOOST_net_12716) );
na02s02 TIMEBOOST_cell_45361 ( .a(n_36), .b(n_4320), .o(TIMEBOOST_net_14919) );
na03f04 TIMEBOOST_cell_32798 ( .a(n_11806), .b(n_11908), .c(n_12206), .o(TIMEBOOST_net_10310) );
in01f01 g57289_u0 ( .a(FE_OFN1368_n_8567), .o(g57289_sb) );
na02f02 TIMEBOOST_cell_22315 ( .a(TIMEBOOST_net_6414), .b(FE_OFN1749_n_12004), .o(n_12737) );
na02s02 TIMEBOOST_cell_45362 ( .a(TIMEBOOST_net_14919), .b(FE_OFN2063_n_6391), .o(TIMEBOOST_net_12619) );
na02f02 TIMEBOOST_cell_41288 ( .a(TIMEBOOST_net_12882), .b(g57456_sb), .o(n_11277) );
in01f01 g57290_u0 ( .a(FE_OFN1345_n_8567), .o(g57290_sb) );
na02f02 TIMEBOOST_cell_4149 ( .a(TIMEBOOST_net_654), .b(n_4125), .o(n_4855) );
na02f02 TIMEBOOST_cell_44546 ( .a(TIMEBOOST_net_14511), .b(FE_OFN1428_n_8567), .o(TIMEBOOST_net_13491) );
na02m02 TIMEBOOST_cell_4150 ( .a(n_3019), .b(n_3017), .o(TIMEBOOST_net_655) );
in01f01 g57291_u0 ( .a(FE_OFN1422_n_8567), .o(g57291_sb) );
na02m02 TIMEBOOST_cell_44601 ( .a(n_9488), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__Q), .o(TIMEBOOST_net_14539) );
na02s02 TIMEBOOST_cell_42743 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__Q), .b(g58278_sb), .o(TIMEBOOST_net_13610) );
na02s02 TIMEBOOST_cell_31627 ( .a(TIMEBOOST_net_9724), .b(g57948_sb), .o(n_9861) );
in01f01 g57292_u0 ( .a(FE_OFN1424_n_8567), .o(g57292_sb) );
na03f02 TIMEBOOST_cell_22326 ( .a(n_10116), .b(n_10112), .c(n_9294), .o(TIMEBOOST_net_6420) );
na02f02 TIMEBOOST_cell_41434 ( .a(TIMEBOOST_net_12955), .b(g57484_sb), .o(n_11252) );
na02s02 TIMEBOOST_cell_45363 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__Q), .b(n_3713), .o(TIMEBOOST_net_14920) );
in01f01 g57293_u0 ( .a(FE_OFN1380_n_8567), .o(g57293_sb) );
na02f02 TIMEBOOST_cell_22327 ( .a(TIMEBOOST_net_6420), .b(n_9295), .o(n_11847) );
na02f02 g55434_u0 ( .a(FE_OFN1577_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__Q), .o(n_12023) );
na02s02 TIMEBOOST_cell_45364 ( .a(TIMEBOOST_net_14920), .b(FE_OFN1233_n_6391), .o(TIMEBOOST_net_12634) );
in01f01 g57294_u0 ( .a(FE_OFN1383_n_8567), .o(g57294_sb) );
na02m02 TIMEBOOST_cell_32548 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__Q), .o(TIMEBOOST_net_10185) );
na02f02 TIMEBOOST_cell_41460 ( .a(TIMEBOOST_net_12968), .b(g57416_sb), .o(n_11326) );
na02s02 TIMEBOOST_cell_45365 ( .a(n_17), .b(n_3618), .o(TIMEBOOST_net_14921) );
in01f01 g57295_u0 ( .a(FE_OFN1414_n_8567), .o(g57295_sb) );
na03f02 TIMEBOOST_cell_22328 ( .a(n_16838), .b(n_9956), .c(n_16839), .o(TIMEBOOST_net_6421) );
na02f02 g54968_u0 ( .a(n_12023), .b(n_12022), .o(n_12527) );
na02f02 TIMEBOOST_cell_41436 ( .a(TIMEBOOST_net_12956), .b(g57403_sb), .o(n_11338) );
in01f01 g57296_u0 ( .a(FE_OFN1419_n_8567), .o(g57296_sb) );
na02f02 TIMEBOOST_cell_22329 ( .a(TIMEBOOST_net_6421), .b(n_10533), .o(n_12129) );
na02f02 TIMEBOOST_cell_41286 ( .a(TIMEBOOST_net_12881), .b(g57088_sb), .o(n_11653) );
na02s02 TIMEBOOST_cell_45366 ( .a(TIMEBOOST_net_14921), .b(FE_OFN2063_n_6391), .o(TIMEBOOST_net_12627) );
in01f01 g57297_u0 ( .a(FE_OFN1415_n_8567), .o(g57297_sb) );
na03f02 TIMEBOOST_cell_22330 ( .a(n_16850), .b(n_16851), .c(n_9982), .o(TIMEBOOST_net_6422) );
na02f02 TIMEBOOST_cell_22561 ( .a(n_11970), .b(TIMEBOOST_net_6537), .o(n_12680) );
na02s01 TIMEBOOST_cell_40309 ( .a(n_4493), .b(g64803_sb), .o(TIMEBOOST_net_12393) );
in01f01 g57298_u0 ( .a(FE_OFN1368_n_8567), .o(g57298_sb) );
na02f02 TIMEBOOST_cell_22331 ( .a(TIMEBOOST_net_6422), .b(n_10564), .o(n_12134) );
na02m02 TIMEBOOST_cell_43753 ( .a(n_9451), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__Q), .o(TIMEBOOST_net_14115) );
na02s01 TIMEBOOST_cell_39642 ( .a(TIMEBOOST_net_12059), .b(g62512_sb), .o(n_7381) );
in01f01 g57299_u0 ( .a(FE_OFN1417_n_8567), .o(g57299_sb) );
na03f02 TIMEBOOST_cell_22332 ( .a(n_16849), .b(n_16848), .c(n_9309), .o(TIMEBOOST_net_6423) );
na02s02 TIMEBOOST_cell_4543 ( .a(TIMEBOOST_net_851), .b(n_4202), .o(n_5748) );
na02m02 TIMEBOOST_cell_44547 ( .a(n_9752), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__Q), .o(TIMEBOOST_net_14512) );
in01f01 g57300_u0 ( .a(FE_OFN1344_n_8567), .o(g57300_sb) );
na02f02 TIMEBOOST_cell_4151 ( .a(TIMEBOOST_net_655), .b(n_6983), .o(n_7325) );
na02f01 g57300_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__Q), .b(FE_OFN1344_n_8567), .o(g57300_db) );
na02f04 TIMEBOOST_cell_4152 ( .a(n_16967), .b(n_16974), .o(TIMEBOOST_net_656) );
in01f01 g57301_u0 ( .a(FE_OFN1390_n_8567), .o(g57301_sb) );
na02f02 TIMEBOOST_cell_44276 ( .a(TIMEBOOST_net_14376), .b(FE_OFN1405_n_8567), .o(TIMEBOOST_net_12805) );
na02f02 TIMEBOOST_cell_43878 ( .a(TIMEBOOST_net_14177), .b(FE_OFN1401_n_8567), .o(TIMEBOOST_net_12775) );
na02m02 TIMEBOOST_cell_43879 ( .a(n_9847), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__Q), .o(TIMEBOOST_net_14178) );
in01f01 g57302_u0 ( .a(FE_OFN1401_n_8567), .o(g57302_sb) );
na02f02 TIMEBOOST_cell_43880 ( .a(TIMEBOOST_net_14178), .b(FE_OFN1406_n_8567), .o(TIMEBOOST_net_12774) );
na02s01 TIMEBOOST_cell_43405 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__Q), .b(n_3547), .o(TIMEBOOST_net_13941) );
na02f01 TIMEBOOST_cell_4548 ( .a(n_7622), .b(n_16914), .o(TIMEBOOST_net_854) );
in01f01 g57303_u0 ( .a(FE_OFN1416_n_8567), .o(g57303_sb) );
na02m02 TIMEBOOST_cell_44511 ( .a(n_9076), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__Q), .o(TIMEBOOST_net_14494) );
na02m06 TIMEBOOST_cell_4549 ( .a(TIMEBOOST_net_854), .b(n_7216), .o(TIMEBOOST_net_481) );
na02s02 TIMEBOOST_cell_39644 ( .a(TIMEBOOST_net_12060), .b(g62952_sb), .o(n_5977) );
in01f01 g57304_u0 ( .a(FE_OFN1380_n_8567), .o(g57304_sb) );
na02m02 TIMEBOOST_cell_43881 ( .a(n_9702), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__Q), .o(TIMEBOOST_net_14179) );
na02s02 TIMEBOOST_cell_4551 ( .a(TIMEBOOST_net_855), .b(n_4659), .o(n_6982) );
na02s02 TIMEBOOST_cell_39646 ( .a(TIMEBOOST_net_12061), .b(g62360_sb), .o(n_6878) );
in01f01 g57305_u0 ( .a(FE_OFN1398_n_8567), .o(g57305_sb) );
na02s02 TIMEBOOST_cell_43206 ( .a(TIMEBOOST_net_13841), .b(FE_OFN1241_n_4092), .o(TIMEBOOST_net_12124) );
na02s02 TIMEBOOST_cell_4553 ( .a(TIMEBOOST_net_856), .b(n_4664), .o(n_6984) );
na02s02 TIMEBOOST_cell_39648 ( .a(TIMEBOOST_net_12062), .b(g62886_sb), .o(n_6105) );
in01f01 g57306_u0 ( .a(FE_OFN1420_n_8567), .o(g57306_sb) );
na02s02 TIMEBOOST_cell_45367 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__Q), .b(n_4239), .o(TIMEBOOST_net_14922) );
na02m02 TIMEBOOST_cell_4555 ( .a(TIMEBOOST_net_857), .b(n_4663), .o(n_6987) );
na02s01 TIMEBOOST_cell_18643 ( .a(TIMEBOOST_net_4578), .b(g63131_sb), .o(n_4988) );
in01f01 g57307_u0 ( .a(FE_OFN1425_n_8567), .o(g57307_sb) );
na02s02 TIMEBOOST_cell_43207 ( .a(n_3782), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__25__Q), .o(TIMEBOOST_net_13842) );
na02s02 TIMEBOOST_cell_45632 ( .a(TIMEBOOST_net_15054), .b(g64281_da), .o(TIMEBOOST_net_11270) );
na02f02 TIMEBOOST_cell_10343 ( .a(TIMEBOOST_net_1738), .b(g54317_da), .o(n_13291) );
in01f01 g57308_u0 ( .a(FE_OFN1420_n_8567), .o(g57308_sb) );
na02s02 TIMEBOOST_cell_45368 ( .a(TIMEBOOST_net_14922), .b(FE_OFN1236_n_6391), .o(TIMEBOOST_net_12616) );
na02s01 TIMEBOOST_cell_41753 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__Q), .b(g58310_sb), .o(TIMEBOOST_net_13115) );
na02f02 TIMEBOOST_cell_38932 ( .a(TIMEBOOST_net_11704), .b(g58640_sb), .o(n_9238) );
in01f01 g57309_u0 ( .a(FE_OFN1404_n_8567), .o(g57309_sb) );
na02f02 TIMEBOOST_cell_43882 ( .a(TIMEBOOST_net_14179), .b(FE_OFN1423_n_8567), .o(TIMEBOOST_net_12773) );
in01s01 TIMEBOOST_cell_45922 ( .a(TIMEBOOST_net_15228), .o(TIMEBOOST_net_15229) );
na02s02 TIMEBOOST_cell_38160 ( .a(TIMEBOOST_net_11318), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_4579) );
in01f01 g57310_u0 ( .a(FE_OFN1425_n_8567), .o(g57310_sb) );
na02m02 TIMEBOOST_cell_43883 ( .a(n_9079), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__Q), .o(TIMEBOOST_net_14180) );
na02s01 TIMEBOOST_cell_44874 ( .a(TIMEBOOST_net_14675), .b(g64276_db), .o(n_3897) );
na02f02 TIMEBOOST_cell_38934 ( .a(TIMEBOOST_net_11705), .b(FE_OFN2157_n_16439), .o(TIMEBOOST_net_10727) );
in01f01 g57311_u0 ( .a(FE_OFN1381_n_8567), .o(g57311_sb) );
na02f02 TIMEBOOST_cell_44512 ( .a(TIMEBOOST_net_14494), .b(FE_OFN2179_n_8567), .o(TIMEBOOST_net_13454) );
na02m02 TIMEBOOST_cell_43809 ( .a(n_9055), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__Q), .o(TIMEBOOST_net_14143) );
na02s01 TIMEBOOST_cell_38162 ( .a(TIMEBOOST_net_11319), .b(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_4496) );
in01f01 g57312_u0 ( .a(FE_OFN1415_n_8567), .o(g57312_sb) );
na02f02 TIMEBOOST_cell_43884 ( .a(TIMEBOOST_net_14180), .b(FE_OFN1401_n_8567), .o(TIMEBOOST_net_12772) );
na02s01 TIMEBOOST_cell_45633 ( .a(g64277_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__18__Q), .o(TIMEBOOST_net_15055) );
na02s02 TIMEBOOST_cell_39650 ( .a(TIMEBOOST_net_12063), .b(g62497_sb), .o(n_6589) );
in01f02 g57313_u0 ( .a(FE_OFN2169_n_8567), .o(g57313_sb) );
na02s02 TIMEBOOST_cell_45369 ( .a(n_3627), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__Q), .o(TIMEBOOST_net_14923) );
na02f02 TIMEBOOST_cell_43885 ( .a(n_9119), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__Q), .o(TIMEBOOST_net_14181) );
na02s01 TIMEBOOST_cell_31099 ( .a(TIMEBOOST_net_9460), .b(g65032_db), .o(n_3626) );
in01f01 g57314_u0 ( .a(FE_OFN1405_n_8567), .o(g57314_sb) );
na02s02 TIMEBOOST_cell_43208 ( .a(TIMEBOOST_net_13842), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_12648) );
na02m02 TIMEBOOST_cell_4569 ( .a(TIMEBOOST_net_864), .b(n_4661), .o(n_6985) );
na02m02 TIMEBOOST_cell_4570 ( .a(n_1784), .b(n_13784), .o(TIMEBOOST_net_865) );
in01f02 g57315_u0 ( .a(FE_OFN2182_n_8567), .o(g57315_sb) );
na03m02 TIMEBOOST_cell_32893 ( .a(wbu_addr_in_261), .b(g58770_sb), .c(g58770_db), .o(n_9126) );
na02f02 TIMEBOOST_cell_4571 ( .a(TIMEBOOST_net_865), .b(n_13442), .o(FE_RN_213_0) );
na02f02 TIMEBOOST_cell_43886 ( .a(TIMEBOOST_net_14181), .b(FE_OFN1368_n_8567), .o(TIMEBOOST_net_12763) );
in01f02 g57316_u0 ( .a(FE_OFN2188_n_8567), .o(g57316_sb) );
na03m02 TIMEBOOST_cell_32892 ( .a(wbu_addr_in_266), .b(g58775_sb), .c(g58775_db), .o(n_9853) );
na02s01 TIMEBOOST_cell_31098 ( .a(n_3785), .b(g65032_sb), .o(TIMEBOOST_net_9460) );
na02s01 TIMEBOOST_cell_31097 ( .a(TIMEBOOST_net_9459), .b(g64751_db), .o(n_4502) );
in01f01 g57317_u0 ( .a(FE_OFN1388_n_8567), .o(g57317_sb) );
na02m02 TIMEBOOST_cell_43887 ( .a(n_9099), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__Q), .o(TIMEBOOST_net_14182) );
na02f02 TIMEBOOST_cell_43888 ( .a(TIMEBOOST_net_14182), .b(FE_OFN1368_n_8567), .o(TIMEBOOST_net_12970) );
no02f08 TIMEBOOST_cell_44761 ( .a(FE_RN_764_0), .b(FE_RN_821_0), .o(TIMEBOOST_net_14619) );
in01f01 g57318_u0 ( .a(FE_OFN1411_n_8567), .o(g57318_sb) );
na02m02 TIMEBOOST_cell_44513 ( .a(n_9069), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__Q), .o(TIMEBOOST_net_14495) );
na02s02 TIMEBOOST_cell_40380 ( .a(TIMEBOOST_net_12428), .b(FE_OFN231_n_9839), .o(n_9734) );
na02s02 TIMEBOOST_cell_4576 ( .a(n_9175), .b(n_1304), .o(TIMEBOOST_net_868) );
in01f01 g57319_u0 ( .a(FE_OFN1407_n_8567), .o(g57319_sb) );
na02f02 TIMEBOOST_cell_22065 ( .a(FE_OFN1602_n_13995), .b(TIMEBOOST_net_6289), .o(n_14481) );
na03f02 TIMEBOOST_cell_4578 ( .a(n_2849), .b(n_5230), .c(n_3370), .o(TIMEBOOST_net_869) );
in01f01 g57320_u0 ( .a(FE_OFN1389_n_8567), .o(g57320_sb) );
na02f02 TIMEBOOST_cell_22441 ( .a(FE_OFN1753_n_12086), .b(TIMEBOOST_net_6477), .o(n_12711) );
na03s02 TIMEBOOST_cell_37931 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__Q), .b(FE_OFN1668_n_9477), .c(FE_OFN272_n_9828), .o(TIMEBOOST_net_11204) );
na02m02 TIMEBOOST_cell_4580 ( .a(n_2111), .b(FE_OFN2059_n_13447), .o(TIMEBOOST_net_870) );
in01f01 g57321_u0 ( .a(FE_OFN1368_n_8567), .o(g57321_sb) );
na03s02 TIMEBOOST_cell_43341 ( .a(n_3678), .b(FE_OFN1223_n_6391), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__Q), .o(TIMEBOOST_net_13909) );
na02s02 TIMEBOOST_cell_43640 ( .a(TIMEBOOST_net_14058), .b(FE_OFN1235_n_6391), .o(TIMEBOOST_net_12160) );
na02s02 TIMEBOOST_cell_38164 ( .a(TIMEBOOST_net_11320), .b(FE_OFN1135_g64577_p), .o(TIMEBOOST_net_4719) );
in01f01 g57322_u0 ( .a(FE_OFN1345_n_8567), .o(g57322_sb) );
na02f08 TIMEBOOST_cell_4153 ( .a(TIMEBOOST_net_656), .b(FE_OCP_RBN2018_n_16970), .o(n_13743) );
na02m02 TIMEBOOST_cell_43889 ( .a(n_9770), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q), .o(TIMEBOOST_net_14183) );
na02f02 TIMEBOOST_cell_41098 ( .a(TIMEBOOST_net_12787), .b(g57386_sb), .o(n_10377) );
in01f01 g57323_u0 ( .a(FE_OFN1422_n_8567), .o(g57323_sb) );
na02s01 TIMEBOOST_cell_42042 ( .a(TIMEBOOST_net_13259), .b(g62397_sb), .o(n_6806) );
na02f02 TIMEBOOST_cell_43890 ( .a(TIMEBOOST_net_14183), .b(FE_OFN1406_n_8567), .o(TIMEBOOST_net_12887) );
na03s02 TIMEBOOST_cell_41805 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__Q), .b(FE_OFN699_n_7845), .c(n_1903), .o(TIMEBOOST_net_13141) );
in01f01 g57324_u0 ( .a(FE_OFN1424_n_8567), .o(g57324_sb) );
na02f02 TIMEBOOST_cell_22467 ( .a(TIMEBOOST_net_6490), .b(FE_OFN1513_n_14987), .o(n_12685) );
na02s01 TIMEBOOST_cell_18661 ( .a(TIMEBOOST_net_4587), .b(g62862_sb), .o(n_5242) );
na02f02 TIMEBOOST_cell_44632 ( .a(TIMEBOOST_net_14554), .b(FE_OFN2169_n_8567), .o(TIMEBOOST_net_13482) );
in01f01 g57325_u0 ( .a(FE_OFN1381_n_8567), .o(g57325_sb) );
na02s02 TIMEBOOST_cell_30911 ( .a(TIMEBOOST_net_9366), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_3739) );
na02s02 TIMEBOOST_cell_38166 ( .a(TIMEBOOST_net_11321), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_4654) );
na02f02 TIMEBOOST_cell_41356 ( .a(TIMEBOOST_net_12916), .b(g57530_sb), .o(n_10314) );
in01f01 g57326_u0 ( .a(FE_OFN1383_n_8567), .o(g57326_sb) );
na02s01 TIMEBOOST_cell_30912 ( .a(pci_target_unit_pcit_if_strd_addr_in_715), .b(pci_target_unit_del_sync_addr_in_233), .o(TIMEBOOST_net_9367) );
na02f02 g55198_u0 ( .a(n_12337), .b(n_12062), .o(n_12606) );
na02s02 TIMEBOOST_cell_19271 ( .a(TIMEBOOST_net_4892), .b(g60624_sb), .o(n_4830) );
in01f01 g57327_u0 ( .a(FE_OFN1415_n_8567), .o(g57327_sb) );
na02m02 TIMEBOOST_cell_43891 ( .a(n_9745), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__15__Q), .o(TIMEBOOST_net_14184) );
na02s01 TIMEBOOST_cell_44810 ( .a(TIMEBOOST_net_14643), .b(g65762_db), .o(TIMEBOOST_net_272) );
na02s02 TIMEBOOST_cell_19273 ( .a(TIMEBOOST_net_4893), .b(g60628_sb), .o(n_5709) );
in01f01 g57328_u0 ( .a(FE_OFN1419_n_8567), .o(g57328_sb) );
na02s01 TIMEBOOST_cell_30914 ( .a(pci_target_unit_pcit_if_strd_addr_in_714), .b(pci_target_unit_del_sync_addr_in_232), .o(TIMEBOOST_net_9368) );
na02f02 TIMEBOOST_cell_44368 ( .a(TIMEBOOST_net_14422), .b(FE_OFN1384_n_8567), .o(TIMEBOOST_net_12759) );
na02s02 TIMEBOOST_cell_19275 ( .a(TIMEBOOST_net_4894), .b(g60630_sb), .o(n_5707) );
in01f01 g57329_u0 ( .a(FE_OFN1415_n_8567), .o(g57329_sb) );
na02s02 TIMEBOOST_cell_45370 ( .a(TIMEBOOST_net_14923), .b(FE_OFN1222_n_6391), .o(TIMEBOOST_net_13255) );
na02s01 TIMEBOOST_cell_44811 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__Q), .b(FE_OFN539_n_9690), .o(TIMEBOOST_net_14644) );
na02s02 TIMEBOOST_cell_19277 ( .a(TIMEBOOST_net_4895), .b(g60632_sb), .o(n_5704) );
in01f01 g57330_u0 ( .a(FE_OFN1368_n_8567), .o(g57330_sb) );
na02f02 TIMEBOOST_cell_44548 ( .a(TIMEBOOST_net_14512), .b(FE_OFN2173_n_8567), .o(TIMEBOOST_net_13463) );
na02s01 TIMEBOOST_cell_44812 ( .a(TIMEBOOST_net_14644), .b(g58239_sb), .o(TIMEBOOST_net_13161) );
na02s02 TIMEBOOST_cell_19353 ( .a(TIMEBOOST_net_4933), .b(g60616_sb), .o(n_4838) );
in01f01 g57331_u0 ( .a(FE_OFN1344_n_8567), .o(g57331_sb) );
na02s01 TIMEBOOST_cell_41782 ( .a(TIMEBOOST_net_13129), .b(FE_OFN211_n_9858), .o(TIMEBOOST_net_10047) );
na02f01 g57331_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__Q), .b(FE_OFN1344_n_8567), .o(g57331_db) );
na02m02 TIMEBOOST_cell_32486 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__Q), .o(TIMEBOOST_net_10154) );
in01f01 g57332_u0 ( .a(FE_OFN1417_n_8567), .o(g57332_sb) );
na02f02 TIMEBOOST_cell_43892 ( .a(TIMEBOOST_net_14184), .b(FE_OFN1406_n_8567), .o(TIMEBOOST_net_12984) );
na02s02 TIMEBOOST_cell_44813 ( .a(n_3741), .b(g64930_sb), .o(TIMEBOOST_net_14645) );
na02s01 TIMEBOOST_cell_4598 ( .a(pci_target_unit_wbm_sm_pciw_fifo_cbe_in), .b(n_8757), .o(TIMEBOOST_net_879) );
in01f01 g57333_u0 ( .a(FE_OFN1390_n_8567), .o(g57333_sb) );
na02f02 TIMEBOOST_cell_44514 ( .a(TIMEBOOST_net_14495), .b(FE_OFN2169_n_8567), .o(TIMEBOOST_net_13455) );
na02m02 TIMEBOOST_cell_11469 ( .a(n_14387), .b(TIMEBOOST_net_2301), .o(n_14394) );
na02s01 TIMEBOOST_cell_4600 ( .a(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_81), .b(n_8757), .o(TIMEBOOST_net_880) );
in01f01 g57334_u0 ( .a(FE_OFN1401_n_8567), .o(g57334_sb) );
na02f02 TIMEBOOST_cell_42162 ( .a(TIMEBOOST_net_13319), .b(FE_OFN1389_n_8567), .o(TIMEBOOST_net_12272) );
na02s01 TIMEBOOST_cell_37184 ( .a(TIMEBOOST_net_10830), .b(wbu_addr_in_275), .o(n_9839) );
na02s01 TIMEBOOST_cell_4602 ( .a(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_82), .b(n_8757), .o(TIMEBOOST_net_881) );
in01f01 g57335_u0 ( .a(FE_OFN1416_n_8567), .o(g57335_sb) );
na02s02 TIMEBOOST_cell_43114 ( .a(TIMEBOOST_net_13795), .b(FE_OFN1268_n_4095), .o(TIMEBOOST_net_12094) );
na03s02 TIMEBOOST_cell_38147 ( .a(TIMEBOOST_net_3513), .b(g64254_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__Q), .o(TIMEBOOST_net_11312) );
na02s01 TIMEBOOST_cell_4604 ( .a(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_83), .b(n_8757), .o(TIMEBOOST_net_882) );
in01f01 g57336_u0 ( .a(FE_OFN1380_n_8567), .o(g57336_sb) );
na02f02 TIMEBOOST_cell_42531 ( .a(n_17044), .b(n_10069), .o(TIMEBOOST_net_13504) );
na02m02 TIMEBOOST_cell_19221 ( .a(g53897_db), .b(TIMEBOOST_net_4867), .o(n_13552) );
na02s02 TIMEBOOST_cell_43486 ( .a(TIMEBOOST_net_13981), .b(FE_OFN1232_n_6391), .o(TIMEBOOST_net_12615) );
in01f02 g57337_u0 ( .a(FE_OFN1370_n_8567), .o(g57337_sb) );
na02s01 TIMEBOOST_cell_44875 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__Q), .b(g65812_sb), .o(TIMEBOOST_net_14676) );
na02s02 g52444_u2 ( .a(n_14676), .b(n_14839), .o(g52444_db) );
na02f02 TIMEBOOST_cell_39100 ( .a(TIMEBOOST_net_6447), .b(TIMEBOOST_net_11788), .o(n_16220) );
in01f01 g57338_u0 ( .a(FE_OFN1420_n_8567), .o(g57338_sb) );
na02s01 TIMEBOOST_cell_42757 ( .a(FE_OFN207_n_9865), .b(g58169_sb), .o(TIMEBOOST_net_13617) );
na02s02 TIMEBOOST_cell_18479 ( .a(TIMEBOOST_net_4496), .b(g61835_sb), .o(n_6977) );
na02s02 TIMEBOOST_cell_38600 ( .a(TIMEBOOST_net_11538), .b(g60639_sb), .o(n_5691) );
in01f01 g57339_u0 ( .a(FE_OFN1425_n_8567), .o(g57339_sb) );
na02f02 TIMEBOOST_cell_42532 ( .a(TIMEBOOST_net_13504), .b(FE_RN_715_0), .o(n_12148) );
na02s02 TIMEBOOST_cell_18481 ( .a(TIMEBOOST_net_4497), .b(g62735_sb), .o(n_5509) );
na02s01 TIMEBOOST_cell_41889 ( .a(n_255), .b(n_4729), .o(TIMEBOOST_net_13183) );
in01f02 g57340_u0 ( .a(FE_OFN1428_n_8567), .o(g57340_sb) );
na02f02 TIMEBOOST_cell_41500 ( .a(TIMEBOOST_net_12988), .b(g57535_sb), .o(n_11207) );
na02m02 TIMEBOOST_cell_43893 ( .a(n_9698), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__Q), .o(TIMEBOOST_net_14185) );
na02s02 TIMEBOOST_cell_31096 ( .a(n_4672), .b(g64751_sb), .o(TIMEBOOST_net_9459) );
in01f02 g57341_u0 ( .a(FE_OFN2179_n_8567), .o(g57341_sb) );
na02s02 TIMEBOOST_cell_43489 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__Q), .b(n_4419), .o(TIMEBOOST_net_13983) );
na02s01 TIMEBOOST_cell_31104 ( .a(n_3770), .b(g64821_sb), .o(TIMEBOOST_net_9463) );
na02s01 TIMEBOOST_cell_31084 ( .a(n_4482), .b(g65039_sb), .o(TIMEBOOST_net_9453) );
in01f01 g57342_u0 ( .a(FE_OFN1423_n_8567), .o(g57342_sb) );
na02s02 TIMEBOOST_cell_45634 ( .a(TIMEBOOST_net_15055), .b(g64277_da), .o(TIMEBOOST_net_11261) );
na02s01 TIMEBOOST_cell_41890 ( .a(TIMEBOOST_net_13183), .b(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_4572) );
na02s02 TIMEBOOST_cell_19249 ( .a(TIMEBOOST_net_4881), .b(g60656_sb), .o(n_5666) );
in01f01 g57343_u0 ( .a(FE_OFN1376_n_8567), .o(g57343_sb) );
na02s02 TIMEBOOST_cell_43532 ( .a(TIMEBOOST_net_14004), .b(FE_OFN1249_n_4093), .o(TIMEBOOST_net_12063) );
na02m02 TIMEBOOST_cell_4615 ( .a(n_14387), .b(TIMEBOOST_net_887), .o(n_14388) );
na02s02 TIMEBOOST_cell_19247 ( .a(TIMEBOOST_net_4880), .b(g60606_sb), .o(n_4848) );
in01f01 g57344_u0 ( .a(FE_OFN1398_n_8567), .o(g57344_sb) );
na02s01 TIMEBOOST_cell_45371 ( .a(TIMEBOOST_net_4814), .b(FE_OFN1200_n_4090), .o(TIMEBOOST_net_14924) );
na02m02 TIMEBOOST_cell_4617 ( .a(n_14390), .b(TIMEBOOST_net_888), .o(n_14391) );
na02s02 TIMEBOOST_cell_19245 ( .a(TIMEBOOST_net_4879), .b(g60654_sb), .o(n_5669) );
in01f02 g57345_u0 ( .a(FE_OFN2180_n_8567), .o(g57345_sb) );
na03f08 TIMEBOOST_cell_32889 ( .a(n_16434), .b(n_16462), .c(n_16265), .o(n_16499) );
na03s02 TIMEBOOST_cell_34427 ( .a(TIMEBOOST_net_512), .b(g54180_da), .c(g53938_da), .o(n_13508) );
na02s01 TIMEBOOST_cell_30900 ( .a(pci_target_unit_pcit_if_strd_addr_in_698), .b(pci_target_unit_del_sync_addr_in_216), .o(TIMEBOOST_net_9361) );
in01f01 g57346_u0 ( .a(FE_OFN1384_n_8567), .o(g57346_sb) );
na02s01 TIMEBOOST_cell_43209 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__28__Q), .b(n_4300), .o(TIMEBOOST_net_13843) );
na02m02 TIMEBOOST_cell_4619 ( .a(n_14392), .b(TIMEBOOST_net_889), .o(n_14393) );
na02s02 TIMEBOOST_cell_38168 ( .a(TIMEBOOST_net_11322), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_4660) );
in01f01 g57347_u0 ( .a(FE_OFN1376_n_8567), .o(g57347_sb) );
na02s02 TIMEBOOST_cell_43555 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__Q), .b(n_3722), .o(TIMEBOOST_net_14016) );
na02f02 TIMEBOOST_cell_43894 ( .a(TIMEBOOST_net_14185), .b(FE_OFN1420_n_8567), .o(TIMEBOOST_net_12804) );
na02f02 TIMEBOOST_cell_44738 ( .a(TIMEBOOST_net_14607), .b(n_16629), .o(n_12628) );
in01f01 g57348_u0 ( .a(FE_OFN1399_n_8567), .o(g57348_sb) );
na02s02 TIMEBOOST_cell_40247 ( .a(n_2258), .b(n_2235), .o(TIMEBOOST_net_12362) );
na02m02 TIMEBOOST_cell_15933 ( .a(TIMEBOOST_net_3223), .b(n_2228), .o(TIMEBOOST_net_103) );
na03s02 TIMEBOOST_cell_38097 ( .a(TIMEBOOST_net_3469), .b(g64327_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__Q), .o(TIMEBOOST_net_11287) );
in01f01 g57349_u0 ( .a(FE_OFN1389_n_8567), .o(g57349_sb) );
na02s01 TIMEBOOST_cell_45372 ( .a(TIMEBOOST_net_14924), .b(g62617_sb), .o(n_6323) );
na02m02 TIMEBOOST_cell_4623 ( .a(n_8529), .b(TIMEBOOST_net_891), .o(n_8530) );
na03s02 TIMEBOOST_cell_38167 ( .a(TIMEBOOST_net_3546), .b(g64344_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__Q), .o(TIMEBOOST_net_11322) );
in01f01 g57350_u0 ( .a(FE_OFN1374_n_8567), .o(g57350_sb) );
na02m02 TIMEBOOST_cell_41646 ( .a(FE_OFN1438_n_9372), .b(TIMEBOOST_net_13061), .o(TIMEBOOST_net_11655) );
na02s01 TIMEBOOST_cell_39316 ( .a(TIMEBOOST_net_11896), .b(g65845_db), .o(n_1875) );
na02f06 TIMEBOOST_cell_4626 ( .a(n_16436), .b(n_4686), .o(TIMEBOOST_net_893) );
in01f01 g57351_u0 ( .a(FE_OFN1421_n_8567), .o(g57351_sb) );
na02s01 TIMEBOOST_cell_43210 ( .a(TIMEBOOST_net_13843), .b(FE_OFN1214_n_4151), .o(TIMEBOOST_net_12133) );
na02s01 TIMEBOOST_cell_39358 ( .a(TIMEBOOST_net_11917), .b(g61761_sb), .o(n_8291) );
na02s02 TIMEBOOST_cell_37902 ( .a(TIMEBOOST_net_11189), .b(g58282_sb), .o(n_9520) );
in01f01 g57352_u0 ( .a(FE_OFN1376_n_8567), .o(g57352_sb) );
na03f02 TIMEBOOST_cell_42533 ( .a(n_10524), .b(n_9953), .c(n_9950), .o(TIMEBOOST_net_13505) );
in01s01 TIMEBOOST_cell_45896 ( .a(TIMEBOOST_net_15202), .o(TIMEBOOST_net_15203) );
na02f02 TIMEBOOST_cell_42163 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__Q), .b(n_9645), .o(TIMEBOOST_net_13320) );
in01f01 g57353_u0 ( .a(FE_OFN1349_n_8567), .o(g57353_sb) );
na02f02 TIMEBOOST_cell_41100 ( .a(TIMEBOOST_net_12788), .b(g57390_sb), .o(n_11353) );
na03s02 TIMEBOOST_cell_38159 ( .a(TIMEBOOST_net_3512), .b(g64227_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__Q), .o(TIMEBOOST_net_11318) );
na02m02 TIMEBOOST_cell_32484 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__Q), .o(TIMEBOOST_net_10153) );
in01f02 g57354_u0 ( .a(FE_OFN2179_n_8567), .o(g57354_sb) );
na02s02 TIMEBOOST_cell_41953 ( .a(TIMEBOOST_net_4468), .b(FE_OFN1085_n_13221), .o(TIMEBOOST_net_13215) );
na02f02 TIMEBOOST_cell_12867 ( .a(TIMEBOOST_net_3000), .b(n_13960), .o(n_14256) );
na02f02 TIMEBOOST_cell_42440 ( .a(TIMEBOOST_net_13458), .b(g57179_sb), .o(n_10450) );
in01f01 g57355_u0 ( .a(FE_OFN1390_n_8567), .o(g57355_sb) );
na02s01 TIMEBOOST_cell_9338 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(g64135_sb), .o(TIMEBOOST_net_1236) );
na02f02 TIMEBOOST_cell_12869 ( .a(n_13958), .b(TIMEBOOST_net_3001), .o(n_14254) );
na02m02 TIMEBOOST_cell_41640 ( .a(FE_OFN1439_n_9372), .b(TIMEBOOST_net_13058), .o(TIMEBOOST_net_11648) );
in01f02 g57356_u0 ( .a(FE_OFN2190_n_8567), .o(g57356_sb) );
na03f20 TIMEBOOST_cell_32857 ( .a(n_16942), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .c(n_16635), .o(n_15417) );
na02s02 TIMEBOOST_cell_43211 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__Q), .b(n_4269), .o(TIMEBOOST_net_13844) );
na02s02 TIMEBOOST_cell_43212 ( .a(TIMEBOOST_net_13844), .b(FE_OFN1264_n_4095), .o(TIMEBOOST_net_12051) );
in01f01 g57357_u0 ( .a(FE_OFN1397_n_8567), .o(g57357_sb) );
na02s02 TIMEBOOST_cell_44433 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_789), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_24__Q), .o(TIMEBOOST_net_14455) );
na02m02 TIMEBOOST_cell_43895 ( .a(n_9624), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__Q), .o(TIMEBOOST_net_14186) );
na02s01 TIMEBOOST_cell_4636 ( .a(pci_target_unit_fifos_pcir_flush_in), .b(g57787_da), .o(TIMEBOOST_net_898) );
in01f01 g57358_u0 ( .a(FE_OFN1388_n_8567), .o(g57358_sb) );
na03s03 TIMEBOOST_cell_45373 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__Q), .b(n_3773), .c(FE_OFN2064_n_6391), .o(TIMEBOOST_net_14925) );
na02f02 TIMEBOOST_cell_43896 ( .a(TIMEBOOST_net_14186), .b(FE_OFN1370_n_8567), .o(TIMEBOOST_net_12806) );
na02s01 TIMEBOOST_cell_4638 ( .a(pci_target_unit_fifos_pcir_flush_in), .b(g57789_da), .o(TIMEBOOST_net_899) );
in01f01 g57359_u0 ( .a(FE_OFN1374_n_8567), .o(g57359_sb) );
na02m02 TIMEBOOST_cell_44369 ( .a(n_9062), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__Q), .o(TIMEBOOST_net_14423) );
na02s01 TIMEBOOST_cell_17268 ( .a(n_3739), .b(FE_OFN651_n_4508), .o(TIMEBOOST_net_3891) );
na02s01 TIMEBOOST_cell_4640 ( .a(pci_target_unit_fifos_pcir_flush_in), .b(g57788_da), .o(TIMEBOOST_net_900) );
in01f01 g57360_u0 ( .a(FE_OFN1384_n_8567), .o(g57360_sb) );
no03f06 TIMEBOOST_cell_35169 ( .a(TIMEBOOST_net_5430), .b(FE_RN_127_0), .c(TIMEBOOST_net_926), .o(TIMEBOOST_net_6291) );
na02m02 TIMEBOOST_cell_43897 ( .a(n_9605), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__Q), .o(TIMEBOOST_net_14187) );
na02s01 TIMEBOOST_cell_44814 ( .a(TIMEBOOST_net_14645), .b(g64930_db), .o(n_3678) );
in01f01 g57361_u0 ( .a(FE_OFN1406_n_8567), .o(g57361_sb) );
na02s02 TIMEBOOST_cell_43213 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__Q), .b(n_3771), .o(TIMEBOOST_net_13845) );
na02s02 TIMEBOOST_cell_43406 ( .a(TIMEBOOST_net_13941), .b(n_6645), .o(TIMEBOOST_net_12168) );
na02f04 TIMEBOOST_cell_4644 ( .a(n_3410), .b(FE_RN_158_0), .o(TIMEBOOST_net_902) );
in01f01 g57362_u0 ( .a(FE_OFN1392_n_8567), .o(g57362_sb) );
na02s02 TIMEBOOST_cell_40690 ( .a(TIMEBOOST_net_12583), .b(g62559_sb), .o(n_6443) );
na02f04 TIMEBOOST_cell_4645 ( .a(TIMEBOOST_net_902), .b(n_14967), .o(n_16161) );
na02s02 TIMEBOOST_cell_43641 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__Q), .b(n_3701), .o(TIMEBOOST_net_14059) );
in01f01 g57363_u0 ( .a(FE_OFN1392_n_8567), .o(g57363_sb) );
na02f02 TIMEBOOST_cell_43898 ( .a(TIMEBOOST_net_14187), .b(FE_OFN1368_n_8567), .o(TIMEBOOST_net_12857) );
na02s02 TIMEBOOST_cell_38449 ( .a(TIMEBOOST_net_9852), .b(FE_OFN1085_n_13221), .o(TIMEBOOST_net_11463) );
no02m02 TIMEBOOST_cell_4648 ( .a(n_1513), .b(FE_RN_281_0), .o(TIMEBOOST_net_904) );
in01f02 g57364_u0 ( .a(FE_OFN2170_n_8567), .o(g57364_sb) );
na02s01 TIMEBOOST_cell_42947 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__Q), .b(FE_OFN592_n_9694), .o(TIMEBOOST_net_13712) );
na02s02 TIMEBOOST_cell_30927 ( .a(TIMEBOOST_net_9374), .b(FE_OFN784_n_2678), .o(TIMEBOOST_net_3737) );
in01f01 g57365_u0 ( .a(FE_OFN1399_n_8567), .o(g57365_sb) );
na02s02 TIMEBOOST_cell_42744 ( .a(TIMEBOOST_net_13610), .b(g58278_db), .o(n_9524) );
no02f02 TIMEBOOST_cell_4649 ( .a(TIMEBOOST_net_904), .b(n_8819), .o(FE_RN_283_0) );
na02s02 TIMEBOOST_cell_39652 ( .a(TIMEBOOST_net_12064), .b(g62954_sb), .o(n_5973) );
in01f01 g57366_u0 ( .a(FE_OFN1396_n_8567), .o(g57366_sb) );
na02s02 TIMEBOOST_cell_43124 ( .a(TIMEBOOST_net_13800), .b(FE_OFN1288_n_4098), .o(TIMEBOOST_net_12108) );
na02s01 TIMEBOOST_cell_37602 ( .a(TIMEBOOST_net_11039), .b(g61806_sb), .o(n_8182) );
na02s04 TIMEBOOST_cell_45374 ( .a(TIMEBOOST_net_14925), .b(g62381_sb), .o(n_6840) );
in01f02 g57367_u0 ( .a(FE_OFN2170_n_8567), .o(g57367_sb) );
na02s02 TIMEBOOST_cell_41949 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__Q), .b(g58275_sb), .o(TIMEBOOST_net_13213) );
na02f02 TIMEBOOST_cell_44370 ( .a(TIMEBOOST_net_14423), .b(FE_OFN1381_n_8567), .o(TIMEBOOST_net_12717) );
na02s02 TIMEBOOST_cell_45375 ( .a(n_3757), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__Q), .o(TIMEBOOST_net_14926) );
in01f01 g57368_u0 ( .a(FE_OFN1382_n_8567), .o(g57368_sb) );
na02s01 TIMEBOOST_cell_30928 ( .a(pci_target_unit_pcit_if_strd_addr_in_694), .b(n_2503), .o(TIMEBOOST_net_9375) );
na02m02 TIMEBOOST_cell_44371 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__Q), .b(n_9906), .o(TIMEBOOST_net_14424) );
na02f02 TIMEBOOST_cell_44288 ( .a(TIMEBOOST_net_14382), .b(FE_OFN1402_n_8567), .o(TIMEBOOST_net_12793) );
in01f01 g57369_u0 ( .a(FE_OFN1399_n_8567), .o(g57369_sb) );
na02s01 TIMEBOOST_cell_42675 ( .a(n_4498), .b(g64914_sb), .o(TIMEBOOST_net_13576) );
na02f04 TIMEBOOST_cell_4655 ( .a(TIMEBOOST_net_907), .b(n_16331), .o(n_8820) );
na02s02 TIMEBOOST_cell_45376 ( .a(TIMEBOOST_net_14926), .b(FE_OFN1224_n_6391), .o(TIMEBOOST_net_13273) );
in01f01 g57370_u0 ( .a(FE_OFN1420_n_8567), .o(g57370_sb) );
na02m02 TIMEBOOST_cell_43899 ( .a(n_9623), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__Q), .o(TIMEBOOST_net_14188) );
na03s02 TIMEBOOST_cell_35101 ( .a(TIMEBOOST_net_10003), .b(n_5732), .c(n_7326), .o(n_7721) );
na03f02 TIMEBOOST_cell_22348 ( .a(n_9321), .b(n_10985), .c(n_9322), .o(TIMEBOOST_net_6431) );
in01f01 g57371_u0 ( .a(FE_OFN1423_n_8567), .o(g57371_sb) );
na02m02 TIMEBOOST_cell_42072 ( .a(TIMEBOOST_net_13274), .b(g59090_sb), .o(n_8714) );
na02f02 TIMEBOOST_cell_41202 ( .a(TIMEBOOST_net_12839), .b(g57492_sb), .o(n_11244) );
na02f02 TIMEBOOST_cell_42270 ( .a(TIMEBOOST_net_13373), .b(g57908_sb), .o(n_8920) );
in01f01 g57372_u0 ( .a(FE_OFN1411_n_8567), .o(g57372_sb) );
na02f04 TIMEBOOST_cell_43686 ( .a(TIMEBOOST_net_14081), .b(TIMEBOOST_net_5590), .o(n_13731) );
na02s01 TIMEBOOST_cell_37177 ( .a(n_8831), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_25__Q), .o(TIMEBOOST_net_10827) );
na02s01 TIMEBOOST_cell_38024 ( .a(TIMEBOOST_net_11250), .b(g61716_sb), .o(n_8393) );
in01f01 g57373_u0 ( .a(FE_OFN1419_n_8567), .o(g57373_sb) );
na02f02 TIMEBOOST_cell_44723 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__Q), .b(FE_OCP_RBN1980_n_10273), .o(TIMEBOOST_net_14600) );
no02f02 TIMEBOOST_cell_4661 ( .a(TIMEBOOST_net_910), .b(n_7709), .o(n_13566) );
na02s02 TIMEBOOST_cell_45377 ( .a(n_3695), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__Q), .o(TIMEBOOST_net_14927) );
in01f01 g57374_u0 ( .a(FE_OFN1422_n_8567), .o(g57374_sb) );
na02f02 TIMEBOOST_cell_22433 ( .a(TIMEBOOST_net_6473), .b(FE_OFN1752_n_12086), .o(n_12596) );
na02s01 TIMEBOOST_cell_37175 ( .a(FE_OFN2054_n_8831), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_32__Q), .o(TIMEBOOST_net_10826) );
na02f02 TIMEBOOST_cell_42272 ( .a(TIMEBOOST_net_13374), .b(g57393_sb), .o(n_11349) );
in01f01 g57375_u0 ( .a(FE_OFN1381_n_8567), .o(g57375_sb) );
na02m02 TIMEBOOST_cell_43346 ( .a(TIMEBOOST_net_13911), .b(g59098_sb), .o(n_8713) );
no02f04 TIMEBOOST_cell_37173 ( .a(FE_RN_315_0), .b(FE_RN_317_0), .o(TIMEBOOST_net_10825) );
na02s01 TIMEBOOST_cell_43270 ( .a(TIMEBOOST_net_13873), .b(FE_OFN1284_n_4097), .o(TIMEBOOST_net_12643) );
in01f01 g57376_u0 ( .a(FE_OFN1414_n_8567), .o(g57376_sb) );
na02s02 TIMEBOOST_cell_43347 ( .a(TIMEBOOST_net_338), .b(n_2770), .o(TIMEBOOST_net_13912) );
na02s01 TIMEBOOST_cell_39317 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__Q), .b(g65843_sb), .o(TIMEBOOST_net_11897) );
na02s02 TIMEBOOST_cell_43616 ( .a(TIMEBOOST_net_14046), .b(FE_OFN1314_n_6624), .o(TIMEBOOST_net_12245) );
in01f02 g57377_u0 ( .a(FE_OFN2169_n_8567), .o(g57377_sb) );
na02f02 TIMEBOOST_cell_44640 ( .a(TIMEBOOST_net_14558), .b(FE_OFN2189_n_8567), .o(TIMEBOOST_net_13432) );
na02s02 TIMEBOOST_cell_39654 ( .a(TIMEBOOST_net_12065), .b(g62445_sb), .o(n_6705) );
na02f02 TIMEBOOST_cell_39102 ( .a(TIMEBOOST_net_11789), .b(n_12772), .o(n_12951) );
in01f01 g57378_u0 ( .a(FE_OFN1384_n_8567), .o(g57378_sb) );
na02s02 TIMEBOOST_cell_42745 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__Q), .b(g58304_sb), .o(TIMEBOOST_net_13611) );
na02m02 TIMEBOOST_cell_19145 ( .a(TIMEBOOST_net_4829), .b(g63576_sb), .o(n_3427) );
na02s01 TIMEBOOST_cell_38026 ( .a(TIMEBOOST_net_11251), .b(g62026_sb), .o(n_7844) );
in01f02 g57379_u0 ( .a(FE_OFN2185_n_8567), .o(g57379_sb) );
na02s01 TIMEBOOST_cell_42946 ( .a(TIMEBOOST_net_13711), .b(FE_OFN262_n_9851), .o(TIMEBOOST_net_11147) );
na02s02 TIMEBOOST_cell_21943 ( .a(TIMEBOOST_net_6228), .b(g62746_sb), .o(n_5489) );
na02s01 TIMEBOOST_cell_30850 ( .a(n_3764), .b(g65024_sb), .o(TIMEBOOST_net_9336) );
in01f01 g57380_u0 ( .a(FE_OFN1409_n_8567), .o(g57380_sb) );
na02f02 TIMEBOOST_cell_43807 ( .a(n_9530), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__Q), .o(TIMEBOOST_net_14142) );
no02f02 TIMEBOOST_cell_4671 ( .a(TIMEBOOST_net_915), .b(n_7702), .o(n_13571) );
na03f02 g63279_u0 ( .a(n_2826), .b(n_3287), .c(n_3040), .o(n_4652) );
in01f01 g57381_u0 ( .a(FE_OFN1383_n_8567), .o(g57381_sb) );
na02s02 TIMEBOOST_cell_43407 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__Q), .b(n_4463), .o(TIMEBOOST_net_13942) );
na02s02 TIMEBOOST_cell_38586 ( .a(TIMEBOOST_net_11531), .b(g60664_sb), .o(n_5655) );
na02f02 TIMEBOOST_cell_42534 ( .a(TIMEBOOST_net_13505), .b(n_10521), .o(n_12128) );
in01f01 g57382_u0 ( .a(FE_OFN1390_n_8567), .o(g57382_sb) );
na02f02 TIMEBOOST_cell_43900 ( .a(TIMEBOOST_net_14188), .b(FE_OFN1425_n_8567), .o(TIMEBOOST_net_12972) );
na02f02 TIMEBOOST_cell_41102 ( .a(TIMEBOOST_net_12789), .b(g57555_sb), .o(n_10806) );
na02m02 TIMEBOOST_cell_36893 ( .a(n_9413), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__29__Q), .o(TIMEBOOST_net_10685) );
in01f01 g57383_u0 ( .a(FE_OFN1411_n_8567), .o(g57383_sb) );
na02m02 TIMEBOOST_cell_43901 ( .a(n_9885), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__Q), .o(TIMEBOOST_net_14189) );
na02f02 TIMEBOOST_cell_36894 ( .a(TIMEBOOST_net_10685), .b(FE_OFN1385_n_8567), .o(TIMEBOOST_net_6059) );
na02s01 TIMEBOOST_cell_44916 ( .a(TIMEBOOST_net_14696), .b(g65363_db), .o(n_3535) );
in01f01 g57384_u0 ( .a(FE_OFN1419_n_8567), .o(g57384_sb) );
na02s01 TIMEBOOST_cell_30982 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(g65921_sb), .o(TIMEBOOST_net_9402) );
na02s02 TIMEBOOST_cell_38724 ( .a(TIMEBOOST_net_11600), .b(g62498_sb), .o(n_6587) );
na02s01 TIMEBOOST_cell_39656 ( .a(TIMEBOOST_net_12066), .b(g63007_sb), .o(n_5868) );
in01f01 g57385_u0 ( .a(FE_OFN1392_n_8567), .o(g57385_sb) );
na02f02 TIMEBOOST_cell_43902 ( .a(TIMEBOOST_net_14189), .b(FE_OFN1421_n_8567), .o(TIMEBOOST_net_12981) );
na03m02 TIMEBOOST_cell_1790 ( .a(n_3427), .b(g52449_sb), .c(g52449_db), .o(n_14842) );
na02s02 TIMEBOOST_cell_45378 ( .a(TIMEBOOST_net_14927), .b(FE_OFN1224_n_6391), .o(TIMEBOOST_net_13221) );
in01f01 g57386_u0 ( .a(FE_OFN1406_n_8567), .o(g57386_sb) );
na02s02 TIMEBOOST_cell_43214 ( .a(TIMEBOOST_net_13845), .b(FE_OFN1213_n_4151), .o(TIMEBOOST_net_12131) );
na02f02 TIMEBOOST_cell_40926 ( .a(TIMEBOOST_net_12701), .b(g57289_sb), .o(n_11463) );
na02s01 TIMEBOOST_cell_32024 ( .a(configuration_pci_err_data_524), .b(wbm_dat_o_23_), .o(TIMEBOOST_net_9923) );
in01f02 g57387_u0 ( .a(FE_OFN2191_n_8567), .o(g57387_sb) );
na03s02 TIMEBOOST_cell_32856 ( .a(pci_target_unit_del_sync_comp_cycle_count_5_), .b(pci_target_unit_del_sync_comp_cycle_count_2_), .c(n_948), .o(TIMEBOOST_net_31) );
na02s01 TIMEBOOST_cell_15862 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_84), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3188) );
na02m02 TIMEBOOST_cell_43903 ( .a(n_9617), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__Q), .o(TIMEBOOST_net_14190) );
in01f01 g57388_u0 ( .a(FE_OFN1424_n_8567), .o(g57388_sb) );
na02s01 TIMEBOOST_cell_43215 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__Q), .b(n_3550), .o(TIMEBOOST_net_13846) );
na02s01 TIMEBOOST_cell_45379 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_14928) );
na02f02 TIMEBOOST_cell_41366 ( .a(TIMEBOOST_net_12921), .b(g57263_sb), .o(n_11490) );
in01f01 g57389_u0 ( .a(FE_OFN1381_n_8567), .o(g57389_sb) );
na02f02 TIMEBOOST_cell_43904 ( .a(TIMEBOOST_net_14190), .b(FE_OFN1415_n_8567), .o(TIMEBOOST_net_12980) );
na02f02 TIMEBOOST_cell_40928 ( .a(TIMEBOOST_net_12702), .b(g57527_sb), .o(n_11214) );
na02f02 TIMEBOOST_cell_41438 ( .a(TIMEBOOST_net_12957), .b(g57037_sb), .o(n_10515) );
in01f01 g57390_u0 ( .a(FE_OFN1414_n_8567), .o(g57390_sb) );
na02s01 TIMEBOOST_cell_30980 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__Q), .b(pci_target_unit_fifos_pcir_data_in_167), .o(TIMEBOOST_net_9401) );
na02s02 TIMEBOOST_cell_39658 ( .a(TIMEBOOST_net_12067), .b(g62760_sb), .o(n_6121) );
na03f02 TIMEBOOST_cell_4210 ( .a(n_16986), .b(n_9334), .c(n_9335), .o(TIMEBOOST_net_685) );
in01f01 g57391_u0 ( .a(FE_OFN1414_n_8567), .o(g57391_sb) );
na02s01 TIMEBOOST_cell_30983 ( .a(TIMEBOOST_net_9402), .b(g65921_db), .o(n_1850) );
na02m02 TIMEBOOST_cell_32282 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__Q), .b(n_9693), .o(TIMEBOOST_net_10052) );
na02s01 TIMEBOOST_cell_38028 ( .a(TIMEBOOST_net_11252), .b(g61762_sb), .o(n_8288) );
in01f01 g57392_u0 ( .a(FE_OFN1406_n_8567), .o(g57392_sb) );
na02s02 TIMEBOOST_cell_43408 ( .a(TIMEBOOST_net_13942), .b(n_6554), .o(TIMEBOOST_net_12196) );
na02s02 TIMEBOOST_cell_39660 ( .a(TIMEBOOST_net_12068), .b(g62342_sb), .o(n_6915) );
na02s01 TIMEBOOST_cell_32038 ( .a(configuration_pci_err_data_509), .b(wbm_dat_o_8_), .o(TIMEBOOST_net_9930) );
in01f01 g57393_u0 ( .a(FE_OFN1404_n_8567), .o(g57393_sb) );
in01s01 TIMEBOOST_cell_22638 ( .a(TIMEBOOST_net_6576), .o(wbs_dat_i_9_) );
na02s02 TIMEBOOST_cell_32037 ( .a(TIMEBOOST_net_9929), .b(FE_OFN1179_n_3476), .o(TIMEBOOST_net_4911) );
na03s02 TIMEBOOST_cell_37799 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__Q), .b(FE_OFN2257_n_8060), .c(n_1582), .o(TIMEBOOST_net_11138) );
in01f02 g57394_u0 ( .a(FE_OFN1368_n_8567), .o(g57394_sb) );
na03s02 TIMEBOOST_cell_5057 ( .a(g64814_sb), .b(g64814_db), .c(n_4473), .o(n_4459) );
na02f01 g57394_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__Q), .b(FE_OFN1344_n_8567), .o(g57394_db) );
na02f02 TIMEBOOST_cell_41672 ( .a(TIMEBOOST_net_13074), .b(FE_OFN1773_n_13800), .o(g53254_p) );
in01f01 g57395_u0 ( .a(FE_OFN1344_n_8567), .o(g57395_sb) );
na02s01 TIMEBOOST_cell_42698 ( .a(TIMEBOOST_net_13587), .b(g65337_sb), .o(TIMEBOOST_net_10929) );
na02f01 g57395_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__Q), .b(FE_OFN1344_n_8567), .o(g57395_db) );
na02f02 TIMEBOOST_cell_43754 ( .a(TIMEBOOST_net_14115), .b(FE_OFN1374_n_8567), .o(TIMEBOOST_net_12835) );
in01f01 g57396_u0 ( .a(FE_OFN1417_n_8567), .o(g57396_sb) );
in01s01 TIMEBOOST_cell_22639 ( .a(TIMEBOOST_net_6577), .o(TIMEBOOST_net_6576) );
na02s01 TIMEBOOST_cell_38546 ( .a(TIMEBOOST_net_11511), .b(g62059_sb), .o(n_7751) );
na02m02 TIMEBOOST_cell_21978 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__Q), .o(TIMEBOOST_net_6246) );
in01f01 g57397_u0 ( .a(FE_OFN1390_n_8567), .o(g57397_sb) );
in01s01 TIMEBOOST_cell_22640 ( .a(TIMEBOOST_net_6578), .o(wbs_dat_i_20_) );
na02f02 TIMEBOOST_cell_37035 ( .a(FE_OFN1771_n_14054), .b(TIMEBOOST_net_10142), .o(TIMEBOOST_net_10756) );
na03s02 TIMEBOOST_cell_36769 ( .a(g64343_da), .b(g64343_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__Q), .o(TIMEBOOST_net_10623) );
in01f01 g57398_u0 ( .a(FE_OFN1401_n_8567), .o(g57398_sb) );
na02s02 TIMEBOOST_cell_41754 ( .a(TIMEBOOST_net_13115), .b(g58310_db), .o(n_9026) );
na02s01 TIMEBOOST_cell_39662 ( .a(TIMEBOOST_net_12069), .b(g62596_sb), .o(n_6361) );
na02s02 TIMEBOOST_cell_43617 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__Q), .b(n_4457), .o(TIMEBOOST_net_14047) );
in01f01 g57399_u0 ( .a(FE_OFN1405_n_8567), .o(g57399_sb) );
na02s02 TIMEBOOST_cell_43062 ( .a(TIMEBOOST_net_13769), .b(FE_OFN1224_n_6391), .o(TIMEBOOST_net_12585) );
na02m02 TIMEBOOST_cell_11476 ( .a(FE_OFN1699_n_5751), .b(n_3168), .o(TIMEBOOST_net_2305) );
no02f08 TIMEBOOST_cell_36318 ( .a(TIMEBOOST_net_10397), .b(n_16030), .o(n_1279) );
in01f01 g57400_u0 ( .a(FE_OFN1413_n_8567), .o(g57400_sb) );
na02s02 TIMEBOOST_cell_45635 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__Q), .b(g63569_sb), .o(TIMEBOOST_net_15056) );
na02m02 TIMEBOOST_cell_32278 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_1_), .o(TIMEBOOST_net_10050) );
na02s01 TIMEBOOST_cell_38030 ( .a(TIMEBOOST_net_11253), .b(g61744_sb), .o(n_8329) );
in01f01 g57401_u0 ( .a(FE_OFN1380_n_8567), .o(g57401_sb) );
na02f02 TIMEBOOST_cell_42442 ( .a(TIMEBOOST_net_13459), .b(g57316_sb), .o(n_11435) );
no02f02 TIMEBOOST_cell_4707 ( .a(TIMEBOOST_net_933), .b(n_7708), .o(n_13565) );
na02s01 TIMEBOOST_cell_18086 ( .a(FE_OFN252_n_9868), .b(FE_OFN1635_n_9531), .o(TIMEBOOST_net_4300) );
in01f02 g57402_u0 ( .a(FE_OFN2173_n_8567), .o(g57402_sb) );
na02f02 TIMEBOOST_cell_21817 ( .a(TIMEBOOST_net_6165), .b(FE_OFN2260_n_2775), .o(n_4170) );
na02s01 TIMEBOOST_cell_15841 ( .a(TIMEBOOST_net_3177), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_414), .o(TIMEBOOST_net_75) );
na02s01 TIMEBOOST_cell_17853 ( .a(TIMEBOOST_net_4183), .b(g65349_db), .o(n_3542) );
in01f01 g57403_u0 ( .a(FE_OFN1422_n_8567), .o(g57403_sb) );
na02s01 TIMEBOOST_cell_45636 ( .a(TIMEBOOST_net_15056), .b(g63569_db), .o(n_4593) );
na02s02 TIMEBOOST_cell_18087 ( .a(TIMEBOOST_net_4300), .b(TIMEBOOST_net_1537), .o(n_9433) );
na02s01 TIMEBOOST_cell_39664 ( .a(TIMEBOOST_net_12070), .b(g62680_sb), .o(n_6179) );
in01f02 g57404_u0 ( .a(FE_OFN2175_n_8567), .o(g57404_sb) );
na02s01 TIMEBOOST_cell_45380 ( .a(TIMEBOOST_net_14928), .b(FE_OFN1801_n_9690), .o(TIMEBOOST_net_11219) );
na02m02 TIMEBOOST_cell_43905 ( .a(n_9432), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__Q), .o(TIMEBOOST_net_14191) );
na02s02 TIMEBOOST_cell_45695 ( .a(n_4480), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__Q), .o(TIMEBOOST_net_15086) );
in01f02 g57405_u0 ( .a(FE_OFN2184_n_8567), .o(g57405_sb) );
na02m02 TIMEBOOST_cell_44641 ( .a(n_9869), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__8__Q), .o(TIMEBOOST_net_14559) );
na02f02 TIMEBOOST_cell_44274 ( .a(TIMEBOOST_net_14375), .b(FE_OFN1404_n_8567), .o(TIMEBOOST_net_13404) );
in01f02 g57406_u0 ( .a(FE_OFN2175_n_8567), .o(g57406_sb) );
na02s02 TIMEBOOST_cell_45752 ( .a(TIMEBOOST_net_15114), .b(FE_OFN1284_n_4097), .o(TIMEBOOST_net_13267) );
na02s02 TIMEBOOST_cell_43125 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__Q), .b(n_3723), .o(TIMEBOOST_net_13801) );
na02s01 TIMEBOOST_cell_42595 ( .a(FE_OFN205_n_9140), .b(g58417_sb), .o(TIMEBOOST_net_13536) );
in01f01 g57407_u0 ( .a(FE_OFN1391_n_8567), .o(g57407_sb) );
na02f02 TIMEBOOST_cell_42444 ( .a(TIMEBOOST_net_13460), .b(g57340_sb), .o(n_11411) );
na02m02 TIMEBOOST_cell_43739 ( .a(n_9892), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__Q), .o(TIMEBOOST_net_14108) );
na02s01 TIMEBOOST_cell_17952 ( .a(n_4447), .b(FE_OFN1677_n_4655), .o(TIMEBOOST_net_4233) );
in01f01 g57408_u0 ( .a(FE_OFN1411_n_8567), .o(g57408_sb) );
na02m02 TIMEBOOST_cell_45637 ( .a(pci_target_unit_pcit_if_strd_addr_in_687), .b(g52644_sb), .o(TIMEBOOST_net_15057) );
na02s02 TIMEBOOST_cell_17953 ( .a(TIMEBOOST_net_4233), .b(g65387_da), .o(n_4244) );
na02s02 TIMEBOOST_cell_32005 ( .a(TIMEBOOST_net_9913), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_4895) );
in01f01 g57409_u0 ( .a(FE_OFN1419_n_8567), .o(g57409_sb) );
na03s02 TIMEBOOST_cell_33571 ( .a(TIMEBOOST_net_9551), .b(n_5633), .c(g62078_sb), .o(n_5632) );
na02f02 TIMEBOOST_cell_4715 ( .a(FE_OCP_RBN1983_FE_OFN1591_n_13741), .b(TIMEBOOST_net_937), .o(g53182_p) );
na02m02 TIMEBOOST_cell_32452 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__Q), .o(TIMEBOOST_net_10137) );
in01f01 g57410_u0 ( .a(FE_OFN1422_n_8567), .o(g57410_sb) );
na02f02 TIMEBOOST_cell_42446 ( .a(TIMEBOOST_net_13461), .b(g57174_sb), .o(n_11582) );
na02f02 TIMEBOOST_cell_4717 ( .a(FE_OCP_RBN1981_FE_OFN1591_n_13741), .b(TIMEBOOST_net_938), .o(g53170_p) );
na02f02 TIMEBOOST_cell_40930 ( .a(TIMEBOOST_net_12703), .b(g57310_sb), .o(n_11440) );
in01f01 g57411_u0 ( .a(FE_OFN1381_n_8567), .o(g57411_sb) );
na02f02 TIMEBOOST_cell_4719 ( .a(FE_OCP_RBN1984_FE_OFN1591_n_13741), .b(TIMEBOOST_net_939), .o(g53211_p) );
na02m02 TIMEBOOST_cell_37791 ( .a(n_662), .b(g63195_sb), .o(TIMEBOOST_net_11134) );
in01f01 g57412_u0 ( .a(FE_OFN1414_n_8567), .o(g57412_sb) );
na03s02 TIMEBOOST_cell_33568 ( .a(TIMEBOOST_net_9550), .b(n_5633), .c(g62072_sb), .o(n_5639) );
na03m02 TIMEBOOST_cell_32276 ( .a(TIMEBOOST_net_585), .b(g52405_sb), .c(n_4688), .o(TIMEBOOST_net_10049) );
na02s01 TIMEBOOST_cell_39666 ( .a(TIMEBOOST_net_12071), .b(g62459_sb), .o(n_6678) );
in01f02 g57413_u0 ( .a(FE_OFN2169_n_8567), .o(g57413_sb) );
na02s02 TIMEBOOST_cell_43487 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__Q), .b(n_4317), .o(TIMEBOOST_net_13982) );
na02m02 TIMEBOOST_cell_44289 ( .a(n_9029), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__Q), .o(TIMEBOOST_net_14383) );
na02f02 TIMEBOOST_cell_42278 ( .a(TIMEBOOST_net_13377), .b(g57496_sb), .o(n_11241) );
in01f01 g57414_u0 ( .a(FE_OFN1384_n_8567), .o(g57414_sb) );
na02m02 TIMEBOOST_cell_45638 ( .a(TIMEBOOST_net_15057), .b(g52644_db), .o(n_14746) );
na02s02 TIMEBOOST_cell_38465 ( .a(g58437_da), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__31__Q), .o(TIMEBOOST_net_11471) );
na02m02 TIMEBOOST_cell_32482 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__Q), .o(TIMEBOOST_net_10152) );
in01f02 g57415_u0 ( .a(FE_OFN2185_n_8567), .o(g57415_sb) );
na02m02 TIMEBOOST_cell_44215 ( .a(n_9857), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__Q), .o(TIMEBOOST_net_14346) );
na02m02 TIMEBOOST_cell_43572 ( .a(TIMEBOOST_net_14024), .b(FE_OFN1311_n_6624), .o(TIMEBOOST_net_12217) );
na02f02 TIMEBOOST_cell_22443 ( .a(TIMEBOOST_net_6478), .b(FE_OFN1752_n_12086), .o(n_12706) );
in01f01 g57416_u0 ( .a(FE_OFN1383_n_8567), .o(g57416_sb) );
na03f02 TIMEBOOST_cell_33624 ( .a(TIMEBOOST_net_3823), .b(FE_OFN1063_n_15808), .c(TIMEBOOST_net_4360), .o(n_15732) );
na02f02 TIMEBOOST_cell_42535 ( .a(FE_OFN1554_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q), .o(TIMEBOOST_net_13506) );
na02s01 TIMEBOOST_cell_38032 ( .a(TIMEBOOST_net_11254), .b(g61699_sb), .o(n_8430) );
in01f01 g57417_u0 ( .a(FE_OFN1409_n_8567), .o(g57417_sb) );
na02s01 TIMEBOOST_cell_43063 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__Q), .b(n_3748), .o(TIMEBOOST_net_13770) );
in01s01 TIMEBOOST_cell_45897 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_), .o(TIMEBOOST_net_15204) );
na02s01 TIMEBOOST_cell_38170 ( .a(TIMEBOOST_net_11323), .b(FE_OFN877_g64577_p), .o(TIMEBOOST_net_4543) );
in01f01 g57418_u0 ( .a(FE_OFN1390_n_8567), .o(g57418_sb) );
na02s02 TIMEBOOST_cell_42106 ( .a(TIMEBOOST_net_13291), .b(FE_OFN1315_n_6624), .o(TIMEBOOST_net_11588) );
na02s01 TIMEBOOST_cell_37932 ( .a(TIMEBOOST_net_11204), .b(g58368_sb), .o(n_9458) );
na02s01 TIMEBOOST_cell_39481 ( .a(wbs_dat_i_9_), .b(g63616_db), .o(TIMEBOOST_net_11979) );
in01f01 g57419_u0 ( .a(FE_OFN1411_n_8567), .o(g57419_sb) );
na02f02 TIMEBOOST_cell_22547 ( .a(TIMEBOOST_net_6530), .b(FE_OFN1736_n_16317), .o(n_12523) );
na02s02 TIMEBOOST_cell_38172 ( .a(TIMEBOOST_net_11324), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_4605) );
na03s01 TIMEBOOST_cell_38173 ( .a(TIMEBOOST_net_3354), .b(g64128_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__Q), .o(TIMEBOOST_net_11325) );
in01f01 g57420_u0 ( .a(FE_OFN1419_n_8567), .o(g57420_sb) );
na02s02 TIMEBOOST_cell_43216 ( .a(TIMEBOOST_net_13846), .b(FE_OFN1242_n_4092), .o(TIMEBOOST_net_12046) );
na02s01 TIMEBOOST_cell_38174 ( .a(TIMEBOOST_net_11325), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_4566) );
na02s02 TIMEBOOST_cell_38662 ( .a(TIMEBOOST_net_11569), .b(g62404_sb), .o(n_6791) );
in01f01 g57421_u0 ( .a(FE_OFN1349_n_8567), .o(g57421_sb) );
na02m06 TIMEBOOST_cell_15922 ( .a(n_1196), .b(n_1383), .o(TIMEBOOST_net_3218) );
na03s02 TIMEBOOST_cell_38181 ( .a(TIMEBOOST_net_4076), .b(g64258_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__Q), .o(TIMEBOOST_net_11329) );
na02s01 TIMEBOOST_cell_42608 ( .a(TIMEBOOST_net_13542), .b(g58095_db), .o(n_9081) );
in01f01 g57422_u0 ( .a(FE_OFN1404_n_8567), .o(g57422_sb) );
na02f02 TIMEBOOST_cell_22549 ( .a(TIMEBOOST_net_6531), .b(FE_OFN1736_n_16317), .o(n_12701) );
na02s02 TIMEBOOST_cell_18097 ( .a(TIMEBOOST_net_4305), .b(g63058_sb), .o(n_5134) );
na02s01 TIMEBOOST_cell_37326 ( .a(TIMEBOOST_net_10901), .b(g64854_sb), .o(TIMEBOOST_net_9425) );
in01f01 g57423_u0 ( .a(FE_OFN1424_n_8567), .o(g57423_sb) );
na02s02 TIMEBOOST_cell_43217 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__Q), .b(n_3657), .o(TIMEBOOST_net_13847) );
na02s01 TIMEBOOST_cell_37327 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__Q), .b(FE_OFN584_n_9692), .o(TIMEBOOST_net_10902) );
na02s01 TIMEBOOST_cell_37328 ( .a(TIMEBOOST_net_10902), .b(g58260_sb), .o(TIMEBOOST_net_408) );
in01f01 g57424_u0 ( .a(FE_OFN1424_n_8567), .o(g57424_sb) );
na02f02 TIMEBOOST_cell_22551 ( .a(TIMEBOOST_net_6532), .b(FE_OFN1735_n_16317), .o(n_12683) );
na02s01 TIMEBOOST_cell_37329 ( .a(n_4479), .b(g64779_sb), .o(TIMEBOOST_net_10903) );
na02s01 TIMEBOOST_cell_37330 ( .a(TIMEBOOST_net_10903), .b(g64779_db), .o(n_4481) );
in01f01 g57425_u0 ( .a(FE_OFN1381_n_8567), .o(g57425_sb) );
na02s02 TIMEBOOST_cell_43544 ( .a(TIMEBOOST_net_14010), .b(FE_OFN1315_n_6624), .o(TIMEBOOST_net_12220) );
na02s01 TIMEBOOST_cell_37331 ( .a(n_4488), .b(g64761_sb), .o(TIMEBOOST_net_10904) );
no02f08 TIMEBOOST_cell_17974 ( .a(FE_RN_66_0), .b(n_15402), .o(TIMEBOOST_net_4244) );
in01f02 g57426_u0 ( .a(FE_OFN2191_n_8567), .o(g57426_sb) );
na02f02 TIMEBOOST_cell_44647 ( .a(n_9061), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__Q), .o(TIMEBOOST_net_14562) );
no02f08 TIMEBOOST_cell_17975 ( .a(TIMEBOOST_net_4244), .b(FE_RN_67_0), .o(n_15403) );
na02s02 TIMEBOOST_cell_36736 ( .a(TIMEBOOST_net_10606), .b(g63620_sb), .o(n_4748) );
in01f01 g57427_u0 ( .a(FE_OFN1414_n_8567), .o(g57427_sb) );
in01s01 TIMEBOOST_cell_22641 ( .a(TIMEBOOST_net_6579), .o(TIMEBOOST_net_6578) );
na02s02 TIMEBOOST_cell_37904 ( .a(TIMEBOOST_net_11190), .b(g58286_sb), .o(n_9517) );
na02s01 TIMEBOOST_cell_18104 ( .a(FE_OFN264_n_9849), .b(g58048_sb), .o(TIMEBOOST_net_4309) );
in01f01 g57428_u0 ( .a(FE_OFN1384_n_8567), .o(g57428_sb) );
na02s01 TIMEBOOST_cell_39668 ( .a(TIMEBOOST_net_12072), .b(g62333_sb), .o(n_6934) );
na02s01 TIMEBOOST_cell_18105 ( .a(TIMEBOOST_net_4309), .b(g58048_db), .o(n_9741) );
na02m02 TIMEBOOST_cell_43348 ( .a(TIMEBOOST_net_13912), .b(TIMEBOOST_net_4813), .o(n_13504) );
in01f01 g57429_u0 ( .a(FE_OFN1404_n_8567), .o(g57429_sb) );
in01s01 TIMEBOOST_cell_22642 ( .a(TIMEBOOST_net_6580), .o(wbs_dat_i_1_) );
na02s02 TIMEBOOST_cell_18187 ( .a(TIMEBOOST_net_4350), .b(g58373_sb), .o(n_9456) );
na02f02 TIMEBOOST_cell_42536 ( .a(n_12427), .b(TIMEBOOST_net_13506), .o(n_12661) );
in01f01 g57430_u0 ( .a(FE_OFN1368_n_8567), .o(g57430_sb) );
in01s01 TIMEBOOST_cell_22643 ( .a(TIMEBOOST_net_6581), .o(TIMEBOOST_net_6580) );
na02s01 TIMEBOOST_cell_18195 ( .a(TIMEBOOST_net_4354), .b(g61901_sb), .o(n_8021) );
na02s01 TIMEBOOST_cell_45028 ( .a(TIMEBOOST_net_14752), .b(g64117_db), .o(n_4043) );
in01f01 g57431_u0 ( .a(FE_OFN1401_n_8567), .o(g57431_sb) );
na02f02 TIMEBOOST_cell_41662 ( .a(TIMEBOOST_net_13069), .b(FE_OFN2158_n_16439), .o(TIMEBOOST_net_11737) );
na02s02 TIMEBOOST_cell_18191 ( .a(TIMEBOOST_net_4352), .b(g58351_sb), .o(n_9470) );
na03s02 TIMEBOOST_cell_38175 ( .a(TIMEBOOST_net_4042), .b(g65915_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__Q), .o(TIMEBOOST_net_11326) );
in01f01 g57432_u0 ( .a(FE_OFN1417_n_8567), .o(g57432_sb) );
na02f04 TIMEBOOST_cell_44767 ( .a(FE_RN_269_0), .b(FE_RN_271_0), .o(TIMEBOOST_net_14622) );
na02s02 TIMEBOOST_cell_38176 ( .a(TIMEBOOST_net_11326), .b(FE_OFN1125_g64577_p), .o(TIMEBOOST_net_4595) );
na02f02 TIMEBOOST_cell_42537 ( .a(FE_OFN1553_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__Q), .o(TIMEBOOST_net_13507) );
in01f01 g57433_u0 ( .a(FE_OFN1377_n_8567), .o(g57433_sb) );
no02f02 TIMEBOOST_cell_44764 ( .a(TIMEBOOST_net_14620), .b(FE_RN_353_0), .o(FE_RN_354_0) );
na02s02 TIMEBOOST_cell_38178 ( .a(TIMEBOOST_net_11327), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_4547) );
na02f02 TIMEBOOST_cell_38824 ( .a(TIMEBOOST_net_11650), .b(g58456_sb), .o(n_9400) );
in01f02 g57434_u0 ( .a(FE_OFN1416_n_8567), .o(g57434_sb) );
na03s02 TIMEBOOST_cell_33880 ( .a(g64302_da), .b(g64302_db), .c(g63085_sb), .o(TIMEBOOST_net_9714) );
na02s01 TIMEBOOST_cell_18509 ( .a(TIMEBOOST_net_4511), .b(g62815_sb), .o(n_5347) );
na03f02 TIMEBOOST_cell_44445 ( .a(n_8557), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__Q), .c(FE_OFN1403_n_8567), .o(TIMEBOOST_net_14461) );
in01f01 g57435_u0 ( .a(FE_OFN1377_n_8567), .o(g57435_sb) );
na02s02 TIMEBOOST_cell_42128 ( .a(TIMEBOOST_net_13302), .b(g62957_sb), .o(n_5967) );
na02f02 TIMEBOOST_cell_4761 ( .a(TIMEBOOST_net_960), .b(n_10281), .o(n_12169) );
na02m02 TIMEBOOST_cell_38852 ( .a(TIMEBOOST_net_11664), .b(g58838_sb), .o(n_8676) );
in01f01 g57436_u0 ( .a(FE_OFN1402_n_8567), .o(g57436_sb) );
na02f02 TIMEBOOST_cell_44252 ( .a(TIMEBOOST_net_14364), .b(FE_OFN1414_n_8567), .o(TIMEBOOST_net_12865) );
na02s02 TIMEBOOST_cell_18511 ( .a(TIMEBOOST_net_4512), .b(g62816_sb), .o(n_5345) );
na02f02 TIMEBOOST_cell_38936 ( .a(TIMEBOOST_net_11706), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10728) );
in01f01 g57437_u0 ( .a(FE_OFN1382_n_8567), .o(g57437_sb) );
na02s01 TIMEBOOST_cell_43141 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__Q), .b(n_4384), .o(TIMEBOOST_net_13809) );
na02s01 TIMEBOOST_cell_18513 ( .a(TIMEBOOST_net_4513), .b(g62818_sb), .o(n_5339) );
na02f02 TIMEBOOST_cell_4766 ( .a(FE_OFN1581_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__Q), .o(TIMEBOOST_net_963) );
in01f01 g57438_u0 ( .a(FE_OFN1403_n_8567), .o(g57438_sb) );
in01s01 TIMEBOOST_cell_45866 ( .a(TIMEBOOST_net_15173), .o(TIMEBOOST_net_15172) );
na02s02 TIMEBOOST_cell_45381 ( .a(n_3721), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__Q), .o(TIMEBOOST_net_14929) );
na02f02 TIMEBOOST_cell_41400 ( .a(TIMEBOOST_net_12938), .b(g57359_sb), .o(n_11388) );
in01f02 g57439_u0 ( .a(FE_OFN2170_n_8567), .o(g57439_sb) );
na02s02 TIMEBOOST_cell_41950 ( .a(TIMEBOOST_net_13213), .b(g58275_db), .o(n_9526) );
na02s02 TIMEBOOST_cell_37536 ( .a(TIMEBOOST_net_11006), .b(FE_OFN712_n_8140), .o(TIMEBOOST_net_4170) );
na02m01 TIMEBOOST_cell_37443 ( .a(wbs_adr_i_2_), .b(FE_OFN1023_n_11877), .o(TIMEBOOST_net_10960) );
in01f01 g57440_u0 ( .a(FE_OFN1380_n_8567), .o(g57440_sb) );
na02f02 TIMEBOOST_cell_44322 ( .a(TIMEBOOST_net_14399), .b(FE_OFN1376_n_8567), .o(TIMEBOOST_net_12318) );
na02s01 TIMEBOOST_cell_37442 ( .a(TIMEBOOST_net_10959), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(n_14741) );
na02f02 TIMEBOOST_cell_43906 ( .a(TIMEBOOST_net_14191), .b(FE_OFN1408_n_8567), .o(TIMEBOOST_net_12971) );
in01f01 g57441_u0 ( .a(FE_OFN1380_n_8567), .o(g57441_sb) );
na02f02 TIMEBOOST_cell_41682 ( .a(TIMEBOOST_net_13079), .b(FE_OFN1586_n_13736), .o(g53222_p) );
na02m02 TIMEBOOST_cell_43907 ( .a(n_9408), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__Q), .o(TIMEBOOST_net_14192) );
na02s01 TIMEBOOST_cell_44815 ( .a(FE_OFN209_n_9126), .b(g58230_sb), .o(TIMEBOOST_net_14646) );
in01f02 g57442_u0 ( .a(FE_OFN2173_n_8567), .o(g57442_sb) );
na02s02 TIMEBOOST_cell_45382 ( .a(TIMEBOOST_net_14929), .b(FE_OFN1222_n_6391), .o(TIMEBOOST_net_13262) );
na02m02 TIMEBOOST_cell_43687 ( .a(n_7698), .b(TIMEBOOST_net_868), .o(TIMEBOOST_net_14082) );
na02f02 TIMEBOOST_cell_22445 ( .a(TIMEBOOST_net_6479), .b(FE_OFN1752_n_12086), .o(n_12697) );
in01f01 g57443_u0 ( .a(FE_OFN1422_n_8567), .o(g57443_sb) );
na02s01 TIMEBOOST_cell_45383 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__Q), .o(TIMEBOOST_net_14930) );
na02f02 TIMEBOOST_cell_4776 ( .a(FE_OFN1735_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__Q), .o(TIMEBOOST_net_968) );
in01f01 g57444_u0 ( .a(FE_OFN1391_n_8567), .o(g57444_sb) );
na02f02 TIMEBOOST_cell_43908 ( .a(TIMEBOOST_net_14192), .b(FE_OFN1423_n_8567), .o(TIMEBOOST_net_12989) );
na02f02 TIMEBOOST_cell_44670 ( .a(TIMEBOOST_net_14573), .b(g57354_sb), .o(n_10388) );
na02s02 TIMEBOOST_cell_31095 ( .a(TIMEBOOST_net_9458), .b(g65415_db), .o(n_3513) );
in01f01 g57445_u0 ( .a(FE_OFN1407_n_8567), .o(g57445_sb) );
na02s01 TIMEBOOST_cell_31094 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__Q), .b(g65415_sb), .o(TIMEBOOST_net_9458) );
na02f02 TIMEBOOST_cell_44228 ( .a(TIMEBOOST_net_14352), .b(FE_OFN1383_n_8567), .o(TIMEBOOST_net_12803) );
na02s01 TIMEBOOST_cell_31093 ( .a(TIMEBOOST_net_9457), .b(g65053_db), .o(n_3618) );
in01f02 g57446_u0 ( .a(FE_OFN2187_n_8567), .o(g57446_sb) );
na02s02 TIMEBOOST_cell_41957 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__Q), .b(g58347_sb), .o(TIMEBOOST_net_13217) );
na02f02 TIMEBOOST_cell_43688 ( .a(TIMEBOOST_net_14082), .b(n_13919), .o(n_14308) );
na02s01 TIMEBOOST_cell_45384 ( .a(TIMEBOOST_net_14930), .b(FE_OFN569_n_9528), .o(TIMEBOOST_net_11189) );
in01f02 g57447_u0 ( .a(FE_OFN1370_n_8567), .o(g57447_sb) );
na02s02 TIMEBOOST_cell_43573 ( .a(n_4410), .b(n_4411), .o(TIMEBOOST_net_14025) );
na02f02 TIMEBOOST_cell_4777 ( .a(n_12334), .b(TIMEBOOST_net_968), .o(n_12768) );
na02s01 TIMEBOOST_cell_37333 ( .a(n_4465), .b(g65089_sb), .o(TIMEBOOST_net_10905) );
in01f01 g57448_u0 ( .a(FE_OFN1374_n_8567), .o(g57448_sb) );
na02s01 TIMEBOOST_cell_31092 ( .a(n_3777), .b(g65053_sb), .o(TIMEBOOST_net_9457) );
na02m02 TIMEBOOST_cell_43909 ( .a(n_9573), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__Q), .o(TIMEBOOST_net_14193) );
na02s02 TIMEBOOST_cell_31091 ( .a(TIMEBOOST_net_9456), .b(g65067_db), .o(n_4314) );
in01f02 g57449_u0 ( .a(FE_OFN2168_n_8567), .o(g57449_sb) );
na02s01 TIMEBOOST_cell_45029 ( .a(pci_target_unit_fifos_pciw_addr_data_in_150), .b(g64157_sb), .o(TIMEBOOST_net_14753) );
na02s02 TIMEBOOST_cell_43218 ( .a(TIMEBOOST_net_13847), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_12045) );
na02s01 TIMEBOOST_cell_42618 ( .a(TIMEBOOST_net_13547), .b(g58251_sb), .o(TIMEBOOST_net_11951) );
in01f02 g57450_u0 ( .a(FE_OFN2180_n_8567), .o(g57450_sb) );
na02f02 TIMEBOOST_cell_41524 ( .a(TIMEBOOST_net_13000), .b(g57439_sb), .o(n_10353) );
na02f02 TIMEBOOST_cell_22449 ( .a(TIMEBOOST_net_6481), .b(FE_OFN1753_n_12086), .o(n_12621) );
na02s02 TIMEBOOST_cell_43219 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__Q), .b(n_4911), .o(TIMEBOOST_net_13848) );
in01f01 g57451_u0 ( .a(FE_OFN1394_n_8567), .o(g57451_sb) );
na02s02 TIMEBOOST_cell_31090 ( .a(n_4470), .b(g65067_sb), .o(TIMEBOOST_net_9456) );
na03s02 TIMEBOOST_cell_38163 ( .a(g64331_da), .b(g64331_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__Q), .o(TIMEBOOST_net_11320) );
na02f02 TIMEBOOST_cell_22459 ( .a(TIMEBOOST_net_6486), .b(FE_OFN1752_n_12086), .o(n_12679) );
in01f01 g57452_u0 ( .a(FE_OFN1408_n_8567), .o(g57452_sb) );
na03s01 TIMEBOOST_cell_33488 ( .a(g61866_sb), .b(g61866_db), .c(n_2032), .o(n_8105) );
na02s01 TIMEBOOST_cell_37332 ( .a(TIMEBOOST_net_10904), .b(g64761_db), .o(n_4492) );
na02f02 TIMEBOOST_cell_43910 ( .a(TIMEBOOST_net_14193), .b(FE_OFN1390_n_8567), .o(TIMEBOOST_net_12977) );
in01f01 g57453_u0 ( .a(FE_OFN1374_n_8567), .o(g57453_sb) );
na03s01 TIMEBOOST_cell_34280 ( .a(TIMEBOOST_net_9812), .b(FE_OFN1174_n_5592), .c(g62113_sb), .o(n_5583) );
na02s01 TIMEBOOST_cell_45385 ( .a(n_3724), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__Q), .o(TIMEBOOST_net_14931) );
na02s02 TIMEBOOST_cell_39670 ( .a(TIMEBOOST_net_12073), .b(g62577_sb), .o(n_6400) );
in01f01 g57454_u0 ( .a(FE_OFN1386_n_8567), .o(g57454_sb) );
na02m02 TIMEBOOST_cell_32570 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__22__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__22__Q), .o(TIMEBOOST_net_10196) );
na02m02 TIMEBOOST_cell_44515 ( .a(n_9439), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__Q), .o(TIMEBOOST_net_14496) );
na03f20 TIMEBOOST_cell_4784 ( .a(n_279), .b(wishbone_slave_unit_wishbone_slave_c_state), .c(wishbone_slave_unit_wishbone_slave_c_state_2), .o(n_15370) );
in01f01 g57455_u0 ( .a(FE_OFN1391_n_8567), .o(g57455_sb) );
na02s02 TIMEBOOST_cell_43220 ( .a(TIMEBOOST_net_13848), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_12081) );
na02s01 TIMEBOOST_cell_43142 ( .a(TIMEBOOST_net_13809), .b(FE_OFN1241_n_4092), .o(TIMEBOOST_net_12040) );
na02m02 TIMEBOOST_cell_43911 ( .a(n_9610), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__Q), .o(TIMEBOOST_net_14194) );
in01f01 g57456_u0 ( .a(FE_OFN1376_n_8567), .o(g57456_sb) );
na02s01 TIMEBOOST_cell_45579 ( .a(FE_OFN639_n_4669), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__Q), .o(TIMEBOOST_net_15028) );
na02f02 TIMEBOOST_cell_43912 ( .a(TIMEBOOST_net_14194), .b(FE_OFN1388_n_8567), .o(TIMEBOOST_net_12975) );
na02m02 TIMEBOOST_cell_43913 ( .a(n_9423), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q), .o(TIMEBOOST_net_14195) );
in01f01 g57457_u0 ( .a(FE_OFN1349_n_8567), .o(g57457_sb) );
na03s02 TIMEBOOST_cell_38103 ( .a(TIMEBOOST_net_4248), .b(g64222_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__Q), .o(TIMEBOOST_net_11290) );
na02s02 TIMEBOOST_cell_43409 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__Q), .b(n_4293), .o(TIMEBOOST_net_13943) );
na02f02 TIMEBOOST_cell_4164 ( .a(n_15434), .b(n_3032), .o(TIMEBOOST_net_662) );
in01f01 g57458_u0 ( .a(FE_OFN1385_n_8567), .o(g57458_sb) );
na02s02 TIMEBOOST_cell_42358 ( .a(TIMEBOOST_net_13417), .b(g54361_sb), .o(n_13081) );
na02s01 TIMEBOOST_cell_37335 ( .a(g64841_sb), .b(n_4465), .o(TIMEBOOST_net_10906) );
na02s01 TIMEBOOST_cell_37334 ( .a(TIMEBOOST_net_10905), .b(g65089_db), .o(n_4301) );
in01f01 g57459_u0 ( .a(FE_OFN1390_n_8567), .o(g57459_sb) );
na02s02 TIMEBOOST_cell_41709 ( .a(g58790_sb), .b(wbu_addr_in_279), .o(TIMEBOOST_net_13093) );
na02s02 TIMEBOOST_cell_45784 ( .a(TIMEBOOST_net_15130), .b(FE_OFN1812_n_7845), .o(TIMEBOOST_net_11383) );
na02s01 TIMEBOOST_cell_37336 ( .a(TIMEBOOST_net_10906), .b(g64841_db), .o(n_4440) );
in01f01 g57460_u0 ( .a(FE_OFN1400_n_8567), .o(g57460_sb) );
na03s02 TIMEBOOST_cell_43021 ( .a(n_3965), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__Q), .c(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_13749) );
na02s02 TIMEBOOST_cell_37338 ( .a(TIMEBOOST_net_10907), .b(g65388_sb), .o(n_4243) );
na04f06 TIMEBOOST_cell_4794 ( .a(g75024_sb), .b(conf_w_addr_in_931), .c(n_16027), .d(conf_w_addr_in), .o(n_16393) );
in01f02 g57461_u0 ( .a(FE_OFN2187_n_8567), .o(g57461_sb) );
na02s02 TIMEBOOST_cell_45639 ( .a(g52642_sb), .b(pci_target_unit_pcit_if_strd_addr_in_713), .o(TIMEBOOST_net_15058) );
na02s01 TIMEBOOST_cell_45386 ( .a(TIMEBOOST_net_14931), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_12587) );
na02s01 TIMEBOOST_cell_42619 ( .a(n_3761), .b(g64788_sb), .o(TIMEBOOST_net_13548) );
in01f01 g57462_u0 ( .a(FE_OFN1388_n_8567), .o(g57462_sb) );
na02s01 TIMEBOOST_cell_44869 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__Q), .b(FE_OFN572_n_9502), .o(TIMEBOOST_net_14673) );
na02f02 TIMEBOOST_cell_44144 ( .a(TIMEBOOST_net_14310), .b(FE_OFN1391_n_8567), .o(TIMEBOOST_net_12808) );
na02s02 TIMEBOOST_cell_39672 ( .a(TIMEBOOST_net_12074), .b(g62889_sb), .o(n_6099) );
in01f01 g57463_u0 ( .a(FE_OFN1386_n_8567), .o(g57463_sb) );
na03s02 TIMEBOOST_cell_33367 ( .a(n_4672), .b(g64839_sb), .c(g64839_db), .o(n_4441) );
na02s02 TIMEBOOST_cell_43051 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__Q), .b(n_3600), .o(TIMEBOOST_net_13764) );
na02f02 TIMEBOOST_cell_44602 ( .a(TIMEBOOST_net_14539), .b(FE_OFN2177_n_8567), .o(TIMEBOOST_net_13008) );
in01f02 g57464_u0 ( .a(FE_OFN2177_n_8567), .o(g57464_sb) );
na02s02 TIMEBOOST_cell_38664 ( .a(TIMEBOOST_net_11570), .b(g62905_sb), .o(n_6067) );
na02f02 TIMEBOOST_cell_44446 ( .a(TIMEBOOST_net_14461), .b(g58591_sb), .o(n_8908) );
na02s01 TIMEBOOST_cell_43221 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__Q), .b(n_4459), .o(TIMEBOOST_net_13849) );
in01f01 g57465_u0 ( .a(FE_OFN1376_n_8567), .o(g57465_sb) );
na02f02 TIMEBOOST_cell_44739 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q), .b(FE_OFN1579_n_12306), .o(TIMEBOOST_net_14608) );
na02f02 TIMEBOOST_cell_43914 ( .a(TIMEBOOST_net_14195), .b(FE_OFN1408_n_8567), .o(TIMEBOOST_net_12976) );
na02m02 TIMEBOOST_cell_43915 ( .a(n_9345), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__Q), .o(TIMEBOOST_net_14196) );
in01f01 g57466_u0 ( .a(FE_OFN1413_n_8567), .o(g57466_sb) );
na02m02 TIMEBOOST_cell_44253 ( .a(n_9007), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__22__Q), .o(TIMEBOOST_net_14365) );
na02s02 TIMEBOOST_cell_39674 ( .a(TIMEBOOST_net_12075), .b(g62652_sb), .o(n_6240) );
no04f10 TIMEBOOST_cell_4802 ( .a(FE_RN_60_0), .b(FE_RN_61_0), .c(wishbone_slave_unit_fifos_pci_clk_inGreyCount_1_), .d(wishbone_slave_unit_fifos_outGreyCount_1_), .o(n_1829) );
in01f01 g57467_u0 ( .a(FE_OFN1396_n_8567), .o(g57467_sb) );
na02f02 TIMEBOOST_cell_42164 ( .a(TIMEBOOST_net_13320), .b(FE_OFN1390_n_8567), .o(TIMEBOOST_net_12326) );
no04f10 TIMEBOOST_cell_4803 ( .a(FE_RN_63_0), .b(FE_RN_64_0), .c(wishbone_slave_unit_fifos_pci_clk_inGreyCount_0_), .d(wishbone_slave_unit_fifos_outGreyCount_0_), .o(n_1828) );
na02f02 TIMEBOOST_cell_43755 ( .a(n_9015), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__Q), .o(TIMEBOOST_net_14116) );
in01f02 g57468_u0 ( .a(FE_OFN2175_n_8567), .o(g57468_sb) );
na02f02 TIMEBOOST_cell_21819 ( .a(TIMEBOOST_net_6166), .b(n_2819), .o(n_4167) );
na02s02 TIMEBOOST_cell_43556 ( .a(TIMEBOOST_net_14016), .b(FE_OFN1322_n_6436), .o(TIMEBOOST_net_12218) );
na02s01 TIMEBOOST_cell_43091 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__Q), .b(g58305_sb), .o(TIMEBOOST_net_13784) );
in01f02 g57469_u0 ( .a(FE_OFN2177_n_8567), .o(g57469_sb) );
na02s02 TIMEBOOST_cell_43689 ( .a(pci_target_unit_fifos_pcir_flush_in), .b(g57781_da), .o(TIMEBOOST_net_14083) );
na03f04 TIMEBOOST_cell_45837 ( .a(n_9219), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__Q), .c(FE_OFN2182_n_8567), .o(TIMEBOOST_net_15157) );
na02f02 TIMEBOOST_cell_22453 ( .a(TIMEBOOST_net_6483), .b(FE_OFN1753_n_12086), .o(n_12611) );
in01f01 g57470_u0 ( .a(FE_OFN1373_n_8567), .o(g57470_sb) );
na02s01 TIMEBOOST_cell_37341 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__Q), .b(FE_OFN580_n_9531), .o(TIMEBOOST_net_10909) );
in01s01 TIMEBOOST_cell_45956 ( .a(TIMEBOOST_net_15262), .o(TIMEBOOST_net_15263) );
na02s02 TIMEBOOST_cell_43222 ( .a(TIMEBOOST_net_13849), .b(FE_OFN1270_n_4095), .o(TIMEBOOST_net_12082) );
in01f02 g57471_u0 ( .a(FE_OFN2184_n_8567), .o(g57471_sb) );
na02s02 TIMEBOOST_cell_41968 ( .a(TIMEBOOST_net_13222), .b(g62347_sb), .o(n_6905) );
na02s02 TIMEBOOST_cell_37340 ( .a(TIMEBOOST_net_10908), .b(g65301_sb), .o(n_4277) );
na02s02 TIMEBOOST_cell_45785 ( .a(n_1875), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__Q), .o(TIMEBOOST_net_15131) );
in01f02 g57472_u0 ( .a(FE_OFN2184_n_8567), .o(g57472_sb) );
na03m02 TIMEBOOST_cell_32926 ( .a(n_2722), .b(TIMEBOOST_net_9304), .c(n_1359), .o(n_2723) );
na02f02 TIMEBOOST_cell_42448 ( .a(TIMEBOOST_net_13462), .b(g57450_sb), .o(n_11284) );
na02s02 TIMEBOOST_cell_43503 ( .a(n_3775), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__1__Q), .o(TIMEBOOST_net_13990) );
in01f01 g57473_u0 ( .a(FE_OFN1409_n_8567), .o(g57473_sb) );
na02m02 TIMEBOOST_cell_42165 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__Q), .b(n_9420), .o(TIMEBOOST_net_13321) );
na02s01 TIMEBOOST_cell_37342 ( .a(TIMEBOOST_net_10909), .b(g58395_sb), .o(TIMEBOOST_net_3937) );
na02s02 TIMEBOOST_cell_42835 ( .a(FE_OFN1145_n_15261), .b(conf_wb_err_addr_in_956), .o(TIMEBOOST_net_13656) );
in01f01 g57474_u0 ( .a(FE_OFN1396_n_8567), .o(g57474_sb) );
na02s01 TIMEBOOST_cell_43223 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__Q), .b(n_4379), .o(TIMEBOOST_net_13850) );
na03s02 TIMEBOOST_cell_36773 ( .a(TIMEBOOST_net_3547), .b(g64353_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q), .o(TIMEBOOST_net_10625) );
na02s01 TIMEBOOST_cell_44864 ( .a(TIMEBOOST_net_14670), .b(g65406_sb), .o(TIMEBOOST_net_11871) );
in01f02 g57475_u0 ( .a(FE_OFN2167_n_8567), .o(g57475_sb) );
na02m02 TIMEBOOST_cell_32788 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__Q), .o(TIMEBOOST_net_10305) );
na02s01 TIMEBOOST_cell_43224 ( .a(TIMEBOOST_net_13850), .b(FE_OFN1247_n_4093), .o(TIMEBOOST_net_11551) );
na02s01 TIMEBOOST_cell_45387 ( .a(TIMEBOOST_net_5307), .b(FE_OFN1232_n_6391), .o(TIMEBOOST_net_14932) );
in01f01 g57476_u0 ( .a(FE_OFN1382_n_8567), .o(g57476_sb) );
na02f02 TIMEBOOST_cell_44372 ( .a(TIMEBOOST_net_14424), .b(FE_OFN1394_n_8567), .o(TIMEBOOST_net_12718) );
na02s02 TIMEBOOST_cell_45640 ( .a(TIMEBOOST_net_15058), .b(g52642_db), .o(TIMEBOOST_net_11369) );
na02m02 TIMEBOOST_cell_44219 ( .a(n_9629), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__29__Q), .o(TIMEBOOST_net_14348) );
in01f01 g57477_u0 ( .a(FE_OFN1400_n_8567), .o(g57477_sb) );
na02f02 TIMEBOOST_cell_42166 ( .a(TIMEBOOST_net_13321), .b(FE_OFN1396_n_8567), .o(TIMEBOOST_net_12265) );
na02s02 TIMEBOOST_cell_31605 ( .a(TIMEBOOST_net_9713), .b(g58300_sb), .o(n_9508) );
na02s02 TIMEBOOST_cell_41710 ( .a(TIMEBOOST_net_13093), .b(g58790_db), .o(n_9832) );
in01f01 g57478_u0 ( .a(FE_OFN1373_n_8567), .o(g57478_sb) );
na02s02 TIMEBOOST_cell_16650 ( .a(n_3744), .b(g64963_sb), .o(TIMEBOOST_net_3582) );
na02s02 TIMEBOOST_cell_45049 ( .a(n_1851), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__Q), .o(TIMEBOOST_net_14763) );
na02s02 TIMEBOOST_cell_16797 ( .a(TIMEBOOST_net_3655), .b(g65343_db), .o(n_3545) );
in01f01 g57479_u0 ( .a(FE_OFN1408_n_8567), .o(g57479_sb) );
na02m02 TIMEBOOST_cell_42167 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__Q), .b(n_9715), .o(TIMEBOOST_net_13322) );
na02s02 TIMEBOOST_cell_37345 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__Q), .b(g58392_sb), .o(TIMEBOOST_net_10911) );
na02s02 TIMEBOOST_cell_37344 ( .a(TIMEBOOST_net_10910), .b(g65346_sb), .o(n_4260) );
in01f01 g57480_u0 ( .a(FE_OFN1421_n_8567), .o(g57480_sb) );
na02m02 TIMEBOOST_cell_43690 ( .a(TIMEBOOST_net_14083), .b(g58622_da), .o(TIMEBOOST_net_12259) );
na02s02 TIMEBOOST_cell_37346 ( .a(TIMEBOOST_net_10911), .b(g58392_db), .o(n_9006) );
in01f01 g57481_u0 ( .a(FE_OFN1419_n_8567), .o(g57481_sb) );
na02s02 TIMEBOOST_cell_42101 ( .a(n_2092), .b(n_3361), .o(TIMEBOOST_net_13289) );
na02f02 TIMEBOOST_cell_22349 ( .a(TIMEBOOST_net_6431), .b(n_10198), .o(n_12162) );
na03s02 TIMEBOOST_cell_34475 ( .a(wbm_adr_o_20_), .b(FE_OFN1699_n_5751), .c(g61855_sb), .o(TIMEBOOST_net_592) );
in01f01 g57482_u0 ( .a(FE_OFN1422_n_8567), .o(g57482_sb) );
na02s02 TIMEBOOST_cell_45641 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__Q), .b(FE_OFN1666_n_9477), .o(TIMEBOOST_net_15059) );
na02s02 TIMEBOOST_cell_31599 ( .a(TIMEBOOST_net_9710), .b(g58342_sb), .o(n_9478) );
na02s02 TIMEBOOST_cell_45388 ( .a(TIMEBOOST_net_14932), .b(g62570_sb), .o(n_6415) );
in01f01 g57483_u0 ( .a(FE_OFN1370_n_8567), .o(g57483_sb) );
na02m02 TIMEBOOST_cell_42265 ( .a(n_9442), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__Q), .o(TIMEBOOST_net_13371) );
na02s02 TIMEBOOST_cell_37348 ( .a(TIMEBOOST_net_10912), .b(g65299_sb), .o(n_4278) );
in01f01 g57484_u0 ( .a(FE_OFN1415_n_8567), .o(g57484_sb) );
na02s02 TIMEBOOST_cell_41755 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__Q), .b(g58378_sb), .o(TIMEBOOST_net_13116) );
na02s02 TIMEBOOST_cell_31595 ( .a(TIMEBOOST_net_9708), .b(g58487_sb), .o(n_9346) );
na02s01 TIMEBOOST_cell_41711 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_14__Q), .b(FE_OFN2054_n_8831), .o(TIMEBOOST_net_13094) );
in01f02 g57485_u0 ( .a(FE_OFN2167_n_8567), .o(g57485_sb) );
na02f02 TIMEBOOST_cell_41440 ( .a(TIMEBOOST_net_12958), .b(g57344_sb), .o(n_10391) );
na02f02 TIMEBOOST_cell_44256 ( .a(TIMEBOOST_net_14366), .b(FE_OFN1398_n_8567), .o(TIMEBOOST_net_12939) );
in01f01 g57486_u0 ( .a(FE_OFN1405_n_8567), .o(g57486_sb) );
na02s02 TIMEBOOST_cell_41756 ( .a(TIMEBOOST_net_13116), .b(g58378_db), .o(n_9009) );
na02s02 TIMEBOOST_cell_37351 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_28__Q), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_411), .o(TIMEBOOST_net_10914) );
na02s02 TIMEBOOST_cell_37350 ( .a(TIMEBOOST_net_10913), .b(g65418_sb), .o(n_4228) );
in01f02 g57487_u0 ( .a(FE_OFN2178_n_8567), .o(g57487_sb) );
na02m02 TIMEBOOST_cell_32786 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__26__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__26__Q), .o(TIMEBOOST_net_10304) );
na03s02 TIMEBOOST_cell_5259 ( .a(n_4473), .b(g65081_sb), .c(g65081_db), .o(n_4306) );
na02s01 TIMEBOOST_cell_41729 ( .a(FE_OFN205_n_9140), .b(g57896_sb), .o(TIMEBOOST_net_13103) );
in01f01 g57488_u0 ( .a(FE_OFN1408_n_8567), .o(g57488_sb) );
in01s01 TIMEBOOST_cell_45878 ( .a(TIMEBOOST_net_15184), .o(TIMEBOOST_net_15185) );
na02s01 TIMEBOOST_cell_37353 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__Q), .b(FE_OFN618_n_4490), .o(TIMEBOOST_net_10915) );
na02s02 TIMEBOOST_cell_37352 ( .a(TIMEBOOST_net_10914), .b(FE_OFN2072_n_15978), .o(TIMEBOOST_net_9853) );
in01f01 g57489_u0 ( .a(FE_OFN1345_n_8567), .o(g57489_sb) );
na02f02 TIMEBOOST_cell_4165 ( .a(TIMEBOOST_net_662), .b(n_15699), .o(n_4857) );
na02f01 g57489_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__Q), .b(FE_OFN1345_n_8567), .o(g57489_db) );
na02f02 TIMEBOOST_cell_4166 ( .a(n_16852), .b(n_3049), .o(TIMEBOOST_net_663) );
in01f01 g57490_u0 ( .a(FE_OFN1388_n_8567), .o(g57490_sb) );
na03s02 TIMEBOOST_cell_43691 ( .a(n_4427), .b(FE_OFN1219_n_6886), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__Q), .o(TIMEBOOST_net_14084) );
na02m02 TIMEBOOST_cell_44557 ( .a(n_9202), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__Q), .o(TIMEBOOST_net_14517) );
na02m02 TIMEBOOST_cell_44145 ( .a(n_9123), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__Q), .o(TIMEBOOST_net_14311) );
in01f01 g57491_u0 ( .a(FE_OFN1421_n_8567), .o(g57491_sb) );
na02s01 TIMEBOOST_cell_37355 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__10__Q), .b(FE_OFN572_n_9502), .o(TIMEBOOST_net_10916) );
na02s01 TIMEBOOST_cell_37354 ( .a(TIMEBOOST_net_10915), .b(g65092_sb), .o(TIMEBOOST_net_239) );
in01f01 g57492_u0 ( .a(FE_OFN1406_n_8567), .o(g57492_sb) );
na02m02 TIMEBOOST_cell_43349 ( .a(TIMEBOOST_net_9972), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_13913) );
na02s01 TIMEBOOST_cell_37357 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__Q), .b(FE_OFN612_n_4501), .o(TIMEBOOST_net_10917) );
na02s01 TIMEBOOST_cell_37356 ( .a(TIMEBOOST_net_10916), .b(g58308_sb), .o(TIMEBOOST_net_409) );
in01f01 g57493_u0 ( .a(FE_OFN1392_n_8567), .o(g57493_sb) );
na02s01 TIMEBOOST_cell_42716 ( .a(TIMEBOOST_net_13596), .b(g65009_db), .o(TIMEBOOST_net_10953) );
na02f02 TIMEBOOST_cell_43916 ( .a(TIMEBOOST_net_14196), .b(FE_OFN1391_n_8567), .o(TIMEBOOST_net_12974) );
na02f02 TIMEBOOST_cell_43917 ( .a(n_9751), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__Q), .o(TIMEBOOST_net_14197) );
in01f01 g57494_u0 ( .a(FE_OFN1407_n_8567), .o(g57494_sb) );
na02s01 TIMEBOOST_cell_37359 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q), .b(FE_OFN1660_n_4490), .o(TIMEBOOST_net_10918) );
na02s01 TIMEBOOST_cell_37358 ( .a(TIMEBOOST_net_10917), .b(g64877_sb), .o(TIMEBOOST_net_235) );
in01f01 g57495_u0 ( .a(FE_OFN1424_n_8567), .o(g57495_sb) );
in01s01 TIMEBOOST_cell_45881 ( .a(n_14388), .o(TIMEBOOST_net_15188) );
na02s01 TIMEBOOST_cell_43459 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__22__Q), .b(n_3712), .o(TIMEBOOST_net_13968) );
na02f02 TIMEBOOST_cell_43918 ( .a(TIMEBOOST_net_14197), .b(FE_OFN1425_n_8567), .o(TIMEBOOST_net_12797) );
in01f01 g57496_u0 ( .a(FE_OFN1424_n_8567), .o(g57496_sb) );
na02f02 TIMEBOOST_cell_42450 ( .a(TIMEBOOST_net_13463), .b(g57172_sb), .o(n_11584) );
na02m02 TIMEBOOST_cell_43919 ( .a(n_9547), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__Q), .o(TIMEBOOST_net_14198) );
na02f02 TIMEBOOST_cell_43920 ( .a(TIMEBOOST_net_14198), .b(FE_OFN1424_n_8567), .o(TIMEBOOST_net_12966) );
in01f01 g57497_u0 ( .a(FE_OFN1413_n_8567), .o(g57497_sb) );
na02s02 TIMEBOOST_cell_45642 ( .a(TIMEBOOST_net_15059), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_11207) );
na02m02 TIMEBOOST_cell_43921 ( .a(n_9050), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__Q), .o(TIMEBOOST_net_14199) );
na02f02 TIMEBOOST_cell_43922 ( .a(TIMEBOOST_net_14199), .b(FE_OFN1396_n_8567), .o(TIMEBOOST_net_12967) );
in01f01 g57498_u0 ( .a(FE_OFN1383_n_8567), .o(g57498_sb) );
na02s02 TIMEBOOST_cell_43557 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__Q), .b(n_4461), .o(TIMEBOOST_net_14017) );
na02s02 TIMEBOOST_cell_31259 ( .a(TIMEBOOST_net_9540), .b(g64943_sb), .o(n_3671) );
na02m02 TIMEBOOST_cell_43923 ( .a(n_9544), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__Q), .o(TIMEBOOST_net_14200) );
in01f01 g57499_u0 ( .a(FE_OFN1414_n_8567), .o(g57499_sb) );
no02f04 TIMEBOOST_cell_44765 ( .a(n_2866), .b(FE_RN_637_0), .o(TIMEBOOST_net_14621) );
na03m04 TIMEBOOST_cell_35837 ( .a(FE_OFN2088_n_13124), .b(TIMEBOOST_net_10023), .c(g54346_sb), .o(n_12966) );
na02f02 TIMEBOOST_cell_44516 ( .a(TIMEBOOST_net_14496), .b(FE_OFN2177_n_8567), .o(TIMEBOOST_net_13490) );
in01f01 g57500_u0 ( .a(FE_OFN1419_n_8567), .o(g57500_sb) );
na02s01 TIMEBOOST_cell_43037 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_), .b(FE_OFN1117_g64577_p), .o(TIMEBOOST_net_13757) );
na02s02 TIMEBOOST_cell_41954 ( .a(TIMEBOOST_net_13215), .b(g54181_da), .o(g53897_db) );
na02s02 TIMEBOOST_cell_45389 ( .a(TIMEBOOST_net_4812), .b(FE_OFN1203_n_4090), .o(TIMEBOOST_net_14933) );
in01f01 g57501_u0 ( .a(FE_OFN1415_n_8567), .o(g57501_sb) );
na02s02 TIMEBOOST_cell_42107 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__Q), .b(n_3717), .o(TIMEBOOST_net_13292) );
na02s01 TIMEBOOST_cell_31257 ( .a(TIMEBOOST_net_9539), .b(g65670_db), .o(n_1959) );
no04f10 TIMEBOOST_cell_4854 ( .a(FE_RN_57_0), .b(FE_RN_58_0), .c(wishbone_slave_unit_fifos_pci_clk_inGreyCount_2_), .d(wishbone_slave_unit_fifos_outGreyCount_2_), .o(n_15735) );
in01f01 g57502_u0 ( .a(FE_OFN1368_n_8567), .o(g57502_sb) );
na02s01 TIMEBOOST_cell_43022 ( .a(TIMEBOOST_net_13749), .b(g62802_sb), .o(n_5378) );
na02s01 TIMEBOOST_cell_39676 ( .a(TIMEBOOST_net_12076), .b(g62897_sb), .o(n_6083) );
na02m02 TIMEBOOST_cell_15911 ( .a(n_1549), .b(TIMEBOOST_net_3212), .o(TIMEBOOST_net_138) );
in01f01 g57503_u0 ( .a(FE_OFN1401_n_8567), .o(g57503_sb) );
na02f02 TIMEBOOST_cell_42452 ( .a(TIMEBOOST_net_13464), .b(g57475_sb), .o(n_10338) );
na02s01 TIMEBOOST_cell_31256 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(g65670_sb), .o(TIMEBOOST_net_9539) );
na02f02 TIMEBOOST_cell_44146 ( .a(TIMEBOOST_net_14311), .b(FE_OFN1404_n_8567), .o(TIMEBOOST_net_13387) );
in01f01 g57504_u0 ( .a(FE_OFN1417_n_8567), .o(g57504_sb) );
na02s03 TIMEBOOST_cell_45774 ( .a(TIMEBOOST_net_15125), .b(FE_OFN1326_n_13547), .o(TIMEBOOST_net_14960) );
na02s02 TIMEBOOST_cell_43225 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__Q), .b(n_3685), .o(TIMEBOOST_net_13851) );
na02s02 TIMEBOOST_cell_43226 ( .a(TIMEBOOST_net_13851), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_11547) );
in01f02 g57505_u0 ( .a(FE_OFN2184_n_8567), .o(g57505_sb) );
na02f02 TIMEBOOST_cell_41442 ( .a(TIMEBOOST_net_12959), .b(g57408_sb), .o(n_11336) );
na02s02 TIMEBOOST_cell_41784 ( .a(TIMEBOOST_net_13130), .b(n_4450), .o(n_4298) );
na02s02 TIMEBOOST_cell_41785 ( .a(n_4447), .b(g64832_db), .o(TIMEBOOST_net_13131) );
in01f01 g57506_u0 ( .a(FE_OFN1416_n_8567), .o(g57506_sb) );
na02s03 TIMEBOOST_cell_45775 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__Q), .b(n_13104), .o(TIMEBOOST_net_15126) );
na02s02 TIMEBOOST_cell_43692 ( .a(TIMEBOOST_net_14084), .b(g62528_sb), .o(n_6518) );
na02s01 TIMEBOOST_cell_45030 ( .a(TIMEBOOST_net_14753), .b(g64157_db), .o(n_4008) );
in01f01 g57507_u0 ( .a(FE_OFN1411_n_8567), .o(g57507_sb) );
na02s02 TIMEBOOST_cell_45031 ( .a(conf_wb_err_addr_in_951), .b(FE_OFN1144_n_15261), .o(TIMEBOOST_net_14754) );
na02m02 TIMEBOOST_cell_43350 ( .a(TIMEBOOST_net_13913), .b(g59118_sb), .o(n_8694) );
na02m02 TIMEBOOST_cell_44373 ( .a(n_9489), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__Q), .o(TIMEBOOST_net_14425) );
in01f01 g57508_u0 ( .a(FE_OFN1402_n_8567), .o(g57508_sb) );
na02s02 TIMEBOOST_cell_43081 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__Q), .b(n_4420), .o(TIMEBOOST_net_13779) );
na02s02 TIMEBOOST_cell_43227 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__Q), .b(n_3545), .o(TIMEBOOST_net_13852) );
na02s02 TIMEBOOST_cell_41819 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__Q), .b(g58406_sb), .o(TIMEBOOST_net_13148) );
in01f01 g57509_u0 ( .a(FE_OFN1400_n_8567), .o(g57509_sb) );
na02s01 TIMEBOOST_cell_42583 ( .a(TIMEBOOST_net_9315), .b(FE_OFN959_n_2299), .o(TIMEBOOST_net_13530) );
no03f02 TIMEBOOST_cell_35838 ( .a(n_4652), .b(n_12595), .c(n_4879), .o(g59345_p) );
na02m02 TIMEBOOST_cell_44603 ( .a(n_9215), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__Q), .o(TIMEBOOST_net_14540) );
in01f01 g57510_u0 ( .a(FE_OFN1403_n_8567), .o(g57510_sb) );
na02m02 TIMEBOOST_cell_44147 ( .a(n_9051), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__Q), .o(TIMEBOOST_net_14312) );
na02m02 TIMEBOOST_cell_44231 ( .a(n_9767), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__Q), .o(TIMEBOOST_net_14354) );
na02s02 TIMEBOOST_cell_43463 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__Q), .b(n_3687), .o(TIMEBOOST_net_13970) );
in01f01 g57511_u0 ( .a(FE_OFN1405_n_8567), .o(g57511_sb) );
na02s02 TIMEBOOST_cell_43128 ( .a(TIMEBOOST_net_13802), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_11552) );
na02s01 TIMEBOOST_cell_42913 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__Q), .b(FE_OFN608_n_9904), .o(TIMEBOOST_net_13695) );
in01f01 g57512_u0 ( .a(FE_OFN1380_n_8567), .o(g57512_sb) );
na02s02 TIMEBOOST_cell_43129 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__Q), .b(n_4475), .o(TIMEBOOST_net_13803) );
na02m02 TIMEBOOST_cell_44157 ( .a(n_9709), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__Q), .o(TIMEBOOST_net_14317) );
na02f02 TIMEBOOST_cell_44158 ( .a(TIMEBOOST_net_14317), .b(FE_OFN1385_n_8567), .o(TIMEBOOST_net_12769) );
in01f01 g57513_u0 ( .a(FE_OFN1409_n_8567), .o(g57513_sb) );
na02s02 TIMEBOOST_cell_43130 ( .a(TIMEBOOST_net_13803), .b(FE_OFN1285_n_4097), .o(TIMEBOOST_net_12115) );
na02m02 TIMEBOOST_cell_43351 ( .a(TIMEBOOST_net_9970), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_13914) );
na02s01 TIMEBOOST_cell_42717 ( .a(FE_OFN225_n_9122), .b(g58052_sb), .o(TIMEBOOST_net_13597) );
in01f01 g57514_u0 ( .a(FE_OFN1420_n_8567), .o(g57514_sb) );
na02s01 TIMEBOOST_cell_43131 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__Q), .b(n_1576), .o(TIMEBOOST_net_13804) );
na02s02 TIMEBOOST_cell_37361 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN615_n_4501), .o(TIMEBOOST_net_10919) );
na02f02 TIMEBOOST_cell_41502 ( .a(TIMEBOOST_net_12989), .b(g57595_sb), .o(n_11158) );
in01f01 g57515_u0 ( .a(FE_OFN1425_n_8567), .o(g57515_sb) );
na02m04 TIMEBOOST_cell_45823 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_16__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_781), .o(TIMEBOOST_net_15150) );
na03f08 TIMEBOOST_cell_4877 ( .a(n_15981), .b(n_16940), .c(FE_RN_56_0), .o(n_15982) );
na03s01 TIMEBOOST_cell_33498 ( .a(n_2165), .b(g61994_sb), .c(g61994_db), .o(n_7907) );
na02f01 g57516_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__Q), .b(FE_OFN1379_n_8567), .o(g57516_db) );
na02f02 TIMEBOOST_cell_44290 ( .a(TIMEBOOST_net_14383), .b(FE_OFN1403_n_8567), .o(TIMEBOOST_net_13406) );
in01f01 g57517_u0 ( .a(FE_OFN1407_n_8567), .o(g57517_sb) );
na02f04 TIMEBOOST_cell_45824 ( .a(TIMEBOOST_net_15150), .b(FE_OFN2134_n_13124), .o(TIMEBOOST_net_14992) );
na02s01 TIMEBOOST_cell_37360 ( .a(TIMEBOOST_net_10918), .b(g64765_sb), .o(TIMEBOOST_net_232) );
na02s01 TIMEBOOST_cell_31555 ( .a(TIMEBOOST_net_9688), .b(g57929_sb), .o(n_9881) );
in01f02 g57518_u0 ( .a(FE_OFN2188_n_8567), .o(g57518_sb) );
na02m02 TIMEBOOST_cell_32784 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__Q), .o(TIMEBOOST_net_10303) );
na02f02 TIMEBOOST_cell_44148 ( .a(TIMEBOOST_net_14312), .b(FE_OFN1413_n_8567), .o(TIMEBOOST_net_12992) );
na02s01 TIMEBOOST_cell_31069 ( .a(TIMEBOOST_net_9445), .b(g65003_db), .o(n_4352) );
in01f01 g57519_u0 ( .a(FE_OFN1370_n_8567), .o(g57519_sb) );
na03s01 TIMEBOOST_cell_33496 ( .a(n_1577), .b(g61929_sb), .c(g61929_db), .o(n_7965) );
na02f02 TIMEBOOST_cell_42280 ( .a(TIMEBOOST_net_13378), .b(g57293_sb), .o(n_10410) );
na02s01 TIMEBOOST_cell_31255 ( .a(TIMEBOOST_net_9538), .b(g64805_db), .o(n_3754) );
in01f01 g57520_u0 ( .a(FE_OFN1374_n_8567), .o(g57520_sb) );
na03s01 TIMEBOOST_cell_33495 ( .a(n_2204), .b(g61707_sb), .c(g61707_db), .o(n_8413) );
na02m02 TIMEBOOST_cell_15910 ( .a(n_1409), .b(n_3007), .o(TIMEBOOST_net_3212) );
na04m02 TIMEBOOST_cell_34765 ( .a(TIMEBOOST_net_4827), .b(g63202_sb), .c(g52454_sb), .d(g52454_db), .o(n_14836) );
in01f02 g57521_u0 ( .a(FE_OFN2168_n_8567), .o(g57521_sb) );
na02f02 TIMEBOOST_cell_41444 ( .a(TIMEBOOST_net_12960), .b(g57057_sb), .o(n_11680) );
na02f06 TIMEBOOST_cell_43693 ( .a(n_13289), .b(FE_RN_578_0), .o(TIMEBOOST_net_14085) );
na02f02 TIMEBOOST_cell_22469 ( .a(TIMEBOOST_net_6491), .b(FE_OFN1513_n_14987), .o(n_12629) );
in01f02 g57522_u0 ( .a(FE_OFN2180_n_8567), .o(g57522_sb) );
na02m02 TIMEBOOST_cell_32782 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__Q), .b(n_351), .o(TIMEBOOST_net_10302) );
na02f02 TIMEBOOST_cell_42144 ( .a(TIMEBOOST_net_13310), .b(g57457_sb), .o(n_11276) );
na02f06 TIMEBOOST_cell_43694 ( .a(TIMEBOOST_net_14085), .b(n_7821), .o(FE_RN_176_0) );
in01f01 g57523_u0 ( .a(FE_OFN1394_n_8567), .o(g57523_sb) );
na02s02 TIMEBOOST_cell_41952 ( .a(TIMEBOOST_net_13214), .b(FE_OFN1258_n_4143), .o(TIMEBOOST_net_11544) );
na02f02 TIMEBOOST_cell_43924 ( .a(TIMEBOOST_net_14200), .b(FE_OFN1406_n_8567), .o(TIMEBOOST_net_12820) );
in01f01 g57524_u0 ( .a(FE_OFN1399_n_8567), .o(g57524_sb) );
na02f02 TIMEBOOST_cell_44678 ( .a(TIMEBOOST_net_14577), .b(g57415_sb), .o(n_11327) );
na02f02 TIMEBOOST_cell_43925 ( .a(n_9105), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__Q), .o(TIMEBOOST_net_14201) );
na02s01 TIMEBOOST_cell_37363 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__Q), .b(FE_OFN579_n_9531), .o(TIMEBOOST_net_10920) );
in01f01 g57525_u0 ( .a(FE_OFN1374_n_8567), .o(g57525_sb) );
na02s01 TIMEBOOST_cell_39318 ( .a(TIMEBOOST_net_11897), .b(g65843_db), .o(n_1877) );
na02s02 TIMEBOOST_cell_41757 ( .a(n_3774), .b(g64946_sb), .o(TIMEBOOST_net_13117) );
in01f01 g57526_u0 ( .a(FE_OFN1388_n_8567), .o(g57526_sb) );
na02s01 TIMEBOOST_cell_45643 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__Q), .b(FE_OFN588_n_9692), .o(TIMEBOOST_net_15060) );
na02m02 TIMEBOOST_cell_42253 ( .a(n_9843), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__Q), .o(TIMEBOOST_net_13365) );
na02f02 TIMEBOOST_cell_42454 ( .a(TIMEBOOST_net_13465), .b(g57146_sb), .o(n_11604) );
in01f01 g57527_u0 ( .a(FE_OFN1391_n_8567), .o(g57527_sb) );
na02s02 TIMEBOOST_cell_43228 ( .a(TIMEBOOST_net_13852), .b(FE_OFN1257_n_4143), .o(TIMEBOOST_net_12111) );
na02s02 TIMEBOOST_cell_45390 ( .a(TIMEBOOST_net_14933), .b(g62594_sb), .o(n_6364) );
na02s01 TIMEBOOST_cell_45644 ( .a(TIMEBOOST_net_15060), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_11184) );
in01f02 g57528_u0 ( .a(FE_OFN2182_n_8567), .o(g57528_sb) );
na02f02 TIMEBOOST_cell_41446 ( .a(TIMEBOOST_net_12961), .b(g57101_sb), .o(n_11645) );
na02f02 TIMEBOOST_cell_22471 ( .a(TIMEBOOST_net_6492), .b(FE_OCPN1827_n_14995), .o(n_12746) );
na02f02 TIMEBOOST_cell_43926 ( .a(TIMEBOOST_net_14201), .b(FE_OFN1416_n_8567), .o(TIMEBOOST_net_12925) );
in01f01 g57529_u0 ( .a(FE_OFN1349_n_8567), .o(g57529_sb) );
na02f02 TIMEBOOST_cell_4167 ( .a(TIMEBOOST_net_663), .b(n_16853), .o(n_4858) );
na02f02 TIMEBOOST_cell_44549 ( .a(n_9020), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__Q), .o(TIMEBOOST_net_14513) );
na02m02 TIMEBOOST_cell_40197 ( .a(wbs_wbb3_2_wbb2_dat_o_i_103), .b(wbs_dat_o_4_), .o(TIMEBOOST_net_12337) );
in01m01 g57530_u0 ( .a(FE_OFN1385_n_8567), .o(g57530_sb) );
na02s04 TIMEBOOST_cell_45764 ( .a(TIMEBOOST_net_15120), .b(FE_OFN1332_n_13547), .o(TIMEBOOST_net_14955) );
na02f02 TIMEBOOST_cell_42456 ( .a(TIMEBOOST_net_13466), .b(g57111_sb), .o(n_11635) );
na02s01 TIMEBOOST_cell_45645 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__Q), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_15061) );
in01f01 g57531_u0 ( .a(FE_OFN1390_n_8567), .o(g57531_sb) );
no03f06 TIMEBOOST_cell_33212 ( .a(n_15142), .b(TIMEBOOST_net_3443), .c(g74749_p), .o(n_15458) );
na02f02 TIMEBOOST_cell_41652 ( .a(FE_OFN1440_n_9372), .b(TIMEBOOST_net_13064), .o(TIMEBOOST_net_11680) );
na02f02 TIMEBOOST_cell_42458 ( .a(TIMEBOOST_net_13467), .b(g57487_sb), .o(n_11250) );
in01f02 g57532_u0 ( .a(FE_OFN2187_n_8567), .o(g57532_sb) );
na02m02 TIMEBOOST_cell_32780 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__Q), .o(TIMEBOOST_net_10301) );
na02s01 TIMEBOOST_cell_30926 ( .a(pci_target_unit_pcit_if_strd_addr_in_709), .b(pci_target_unit_del_sync_addr_in_227), .o(TIMEBOOST_net_9374) );
na02s01 TIMEBOOST_cell_45646 ( .a(TIMEBOOST_net_15061), .b(FE_OFN526_n_9899), .o(TIMEBOOST_net_11167) );
in01f01 g57533_u0 ( .a(FE_OFN1400_n_8567), .o(g57533_sb) );
na02f02 TIMEBOOST_cell_41622 ( .a(FE_OFN1441_n_9372), .b(TIMEBOOST_net_13049), .o(TIMEBOOST_net_11661) );
na02f02 TIMEBOOST_cell_42460 ( .a(TIMEBOOST_net_13468), .b(g57559_sb), .o(n_10802) );
na02s02 TIMEBOOST_cell_42374 ( .a(TIMEBOOST_net_13425), .b(g54362_sb), .o(n_13080) );
in01f01 g57534_u0 ( .a(FE_OFN1388_n_8567), .o(g57534_sb) );
na02s02 TIMEBOOST_cell_43080 ( .a(TIMEBOOST_net_13778), .b(FE_OFN1293_n_4098), .o(TIMEBOOST_net_12077) );
na02m02 TIMEBOOST_cell_41653 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_28__Q), .b(FE_OFN270_n_9836), .o(TIMEBOOST_net_13065) );
in01f01 g57535_u0 ( .a(FE_OFN1387_n_8567), .o(g57535_sb) );
na02s01 TIMEBOOST_cell_42992 ( .a(TIMEBOOST_net_13734), .b(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_11439) );
na02f02 TIMEBOOST_cell_44720 ( .a(TIMEBOOST_net_14598), .b(FE_OFN1586_n_13736), .o(n_14419) );
na02s04 TIMEBOOST_cell_45808 ( .a(TIMEBOOST_net_15142), .b(FE_OFN2135_n_13124), .o(TIMEBOOST_net_14984) );
in01f02 g57536_u0 ( .a(FE_OFN2177_n_8567), .o(g57536_sb) );
na02s01 TIMEBOOST_cell_45391 ( .a(n_4227), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__Q), .o(TIMEBOOST_net_14934) );
na02f04 TIMEBOOST_cell_45838 ( .a(TIMEBOOST_net_15157), .b(g57405_sb), .o(n_10829) );
na02f02 TIMEBOOST_cell_44672 ( .a(TIMEBOOST_net_14574), .b(g57035_sb), .o(n_11697) );
in01f01 g57537_u0 ( .a(FE_OFN1376_n_8567), .o(g57537_sb) );
na02s02 TIMEBOOST_cell_37362 ( .a(TIMEBOOST_net_10919), .b(g64962_sb), .o(TIMEBOOST_net_236) );
na02f02 TIMEBOOST_cell_44691 ( .a(wbu_addr_in_258), .b(g52622_sb), .o(TIMEBOOST_net_14584) );
na02s02 TIMEBOOST_cell_31079 ( .a(TIMEBOOST_net_9450), .b(n_4493), .o(n_4334) );
in01f01 g57538_u0 ( .a(FE_OFN1412_n_8567), .o(g57538_sb) );
na03s02 TIMEBOOST_cell_42019 ( .a(n_4323), .b(n_4324), .c(FE_OFN1208_n_6356), .o(TIMEBOOST_net_13248) );
na02f02 TIMEBOOST_cell_40894 ( .a(TIMEBOOST_net_12685), .b(g57491_sb), .o(n_11245) );
na02s01 TIMEBOOST_cell_31254 ( .a(n_3752), .b(g64805_sb), .o(TIMEBOOST_net_9538) );
in01f01 g57539_u0 ( .a(FE_OFN1396_n_8567), .o(g57539_sb) );
na02s01 TIMEBOOST_cell_42020 ( .a(TIMEBOOST_net_13248), .b(g62682_sb), .o(n_6175) );
na02m02 TIMEBOOST_cell_15925 ( .a(TIMEBOOST_net_3219), .b(n_2982), .o(TIMEBOOST_net_180) );
na03f02 TIMEBOOST_cell_36112 ( .a(n_10744), .b(FE_RN_95_0), .c(n_12585), .o(n_12847) );
in01f02 g57540_u0 ( .a(FE_OFN2167_n_8567), .o(g57540_sb) );
na02f02 TIMEBOOST_cell_41402 ( .a(TIMEBOOST_net_12939), .b(g57177_sb), .o(n_10451) );
na02s03 TIMEBOOST_cell_45766 ( .a(TIMEBOOST_net_15121), .b(FE_OFN1327_n_13547), .o(TIMEBOOST_net_14956) );
in01f02 g57541_u0 ( .a(FE_OFN2177_n_8567), .o(g57541_sb) );
na02s02 TIMEBOOST_cell_45392 ( .a(TIMEBOOST_net_14934), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_12580) );
na02s02 TIMEBOOST_cell_45218 ( .a(TIMEBOOST_net_14847), .b(FE_OFN1241_n_4092), .o(TIMEBOOST_net_12122) );
in01f02 g57542_u0 ( .a(FE_OFN2175_n_8567), .o(g57542_sb) );
na02f02 TIMEBOOST_cell_41404 ( .a(TIMEBOOST_net_12940), .b(g57189_sb), .o(n_11564) );
in01s01 TIMEBOOST_cell_45957 ( .a(wbm_dat_i_7_), .o(TIMEBOOST_net_15264) );
na03s02 TIMEBOOST_cell_45393 ( .a(n_4010), .b(FE_OFN1138_g64577_p), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q), .o(TIMEBOOST_net_14935) );
in01f01 g57543_u0 ( .a(FE_OFN1391_n_8567), .o(g57543_sb) );
na02s01 TIMEBOOST_cell_31075 ( .a(TIMEBOOST_net_9448), .b(g65012_db), .o(n_4346) );
na02f01 g57543_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__Q), .b(FE_OFN1379_n_8567), .o(g57543_db) );
na03f02 TIMEBOOST_cell_34491 ( .a(n_2768), .b(n_3593), .c(n_3454), .o(TIMEBOOST_net_653) );
in01f02 g57544_u0 ( .a(FE_OFN2185_n_8567), .o(g57544_sb) );
na02f02 TIMEBOOST_cell_41406 ( .a(TIMEBOOST_net_12941), .b(g57480_sb), .o(n_11256) );
na02m02 TIMEBOOST_cell_41626 ( .a(FE_OFN1438_n_9372), .b(TIMEBOOST_net_13051), .o(TIMEBOOST_net_11662) );
na02f02 TIMEBOOST_cell_44374 ( .a(TIMEBOOST_net_14425), .b(FE_OFN1389_n_8567), .o(TIMEBOOST_net_12720) );
in01f01 g57545_u0 ( .a(FE_OFN1409_n_8567), .o(g57545_sb) );
na02s02 TIMEBOOST_cell_42993 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__Q), .b(g58293_sb), .o(TIMEBOOST_net_13735) );
na02f02 TIMEBOOST_cell_44604 ( .a(TIMEBOOST_net_14540), .b(FE_OFN2177_n_8567), .o(TIMEBOOST_net_13026) );
na02s01 TIMEBOOST_cell_45088 ( .a(TIMEBOOST_net_14782), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_11163) );
in01f01 g57546_u0 ( .a(FE_OFN1396_n_8567), .o(g57546_sb) );
na02s02 TIMEBOOST_cell_42044 ( .a(TIMEBOOST_net_13260), .b(g62530_sb), .o(n_6514) );
na02f04 TIMEBOOST_cell_41515 ( .a(TIMEBOOST_net_10074), .b(n_7095), .o(TIMEBOOST_net_12996) );
na02s02 TIMEBOOST_cell_39678 ( .a(TIMEBOOST_net_12077), .b(g62962_sb), .o(n_5958) );
in01f02 g57547_u0 ( .a(FE_OFN2167_n_8567), .o(g57547_sb) );
na02m02 TIMEBOOST_cell_32774 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__Q), .o(TIMEBOOST_net_10298) );
na02f02 TIMEBOOST_cell_39104 ( .a(TIMEBOOST_net_11790), .b(FE_OFN1554_n_12104), .o(FE_RN_908_0) );
na02s03 TIMEBOOST_cell_45776 ( .a(TIMEBOOST_net_15126), .b(FE_OFN1327_n_13547), .o(TIMEBOOST_net_14961) );
in01f01 g57548_u0 ( .a(FE_OFN1382_n_8567), .o(g57548_sb) );
na03s02 TIMEBOOST_cell_33204 ( .a(n_4312), .b(FE_OFN618_n_4490), .c(g65068_sb), .o(TIMEBOOST_net_238) );
na02f04 TIMEBOOST_cell_41516 ( .a(n_7724), .b(TIMEBOOST_net_12996), .o(n_8576) );
na02s02 TIMEBOOST_cell_41958 ( .a(TIMEBOOST_net_13217), .b(g58347_db), .o(n_9474) );
in01f01 g57549_u0 ( .a(FE_OFN1400_n_8567), .o(g57549_sb) );
na02s02 TIMEBOOST_cell_43533 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__Q), .b(n_3581), .o(TIMEBOOST_net_14005) );
na03s02 TIMEBOOST_cell_45647 ( .a(g63543_da), .b(g63543_db), .c(g61836_sb), .o(TIMEBOOST_net_15062) );
na02s02 TIMEBOOST_cell_43229 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__Q), .b(n_4377), .o(TIMEBOOST_net_13853) );
in01f01 g57550_u0 ( .a(FE_OFN1373_n_8567), .o(g57550_sb) );
na02s02 TIMEBOOST_cell_43296 ( .a(TIMEBOOST_net_13886), .b(g60409_sb), .o(TIMEBOOST_net_11535) );
na02s01 TIMEBOOST_cell_44917 ( .a(TIMEBOOST_net_9505), .b(FE_OFN1044_n_2037), .o(TIMEBOOST_net_14697) );
na02s02 TIMEBOOST_cell_45032 ( .a(TIMEBOOST_net_14754), .b(g59121_sb), .o(TIMEBOOST_net_338) );
in01f01 g57551_u0 ( .a(FE_OFN1408_n_8567), .o(g57551_sb) );
na03s02 TIMEBOOST_cell_42045 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__Q), .b(n_4502), .c(FE_OFN1219_n_6886), .o(TIMEBOOST_net_13261) );
na02m02 TIMEBOOST_cell_44605 ( .a(n_9901), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__Q), .o(TIMEBOOST_net_14541) );
na02s01 TIMEBOOST_cell_41955 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__Q), .b(g58271_sb), .o(TIMEBOOST_net_13216) );
in01f01 g57552_u0 ( .a(FE_OFN1402_n_8567), .o(g57552_sb) );
na02m02 TIMEBOOST_cell_43352 ( .a(TIMEBOOST_net_13914), .b(g59110_sb), .o(n_8693) );
na02f02 TIMEBOOST_cell_44218 ( .a(TIMEBOOST_net_14347), .b(FE_OFN1387_n_8567), .o(TIMEBOOST_net_12988) );
na02s01 TIMEBOOST_cell_37365 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(g64155_sb), .o(TIMEBOOST_net_10921) );
in01f01 g57553_u0 ( .a(FE_OFN1416_n_8567), .o(g57553_sb) );
na02m02 TIMEBOOST_cell_43927 ( .a(n_9779), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__Q), .o(TIMEBOOST_net_14202) );
na02s01 TIMEBOOST_cell_37364 ( .a(TIMEBOOST_net_10920), .b(g58408_sb), .o(TIMEBOOST_net_3899) );
na02f02 TIMEBOOST_cell_41526 ( .a(TIMEBOOST_net_13001), .b(g57040_sb), .o(n_11694) );
in01f01 g57554_u0 ( .a(FE_OFN1411_n_8567), .o(g57554_sb) );
na02s01 TIMEBOOST_cell_42718 ( .a(TIMEBOOST_net_13597), .b(g58052_db), .o(n_9093) );
na02s01 TIMEBOOST_cell_37367 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__Q), .b(g58323_sb), .o(TIMEBOOST_net_10922) );
na02s01 TIMEBOOST_cell_37366 ( .a(TIMEBOOST_net_10921), .b(g64155_db), .o(n_4010) );
in01f01 g57555_u0 ( .a(FE_OFN1402_n_8567), .o(g57555_sb) );
na03s02 TIMEBOOST_cell_33201 ( .a(n_4394), .b(FE_OFN618_n_4490), .c(g64920_sb), .o(TIMEBOOST_net_3943) );
na02s01 TIMEBOOST_cell_41823 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__Q), .b(g58298_sb), .o(TIMEBOOST_net_13150) );
na02s02 TIMEBOOST_cell_41824 ( .a(TIMEBOOST_net_13150), .b(g58298_db), .o(n_9030) );
in01f01 g57556_u0 ( .a(FE_OFN1416_n_8567), .o(g57556_sb) );
na02s02 TIMEBOOST_cell_42046 ( .a(TIMEBOOST_net_13261), .b(g62541_sb), .o(n_6485) );
na02s01 TIMEBOOST_cell_37369 ( .a(n_3774), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__Q), .o(TIMEBOOST_net_10923) );
na02s02 TIMEBOOST_cell_37368 ( .a(TIMEBOOST_net_10922), .b(g58323_db), .o(n_9023) );
in01f01 g57557_u0 ( .a(FE_OFN1377_n_8567), .o(g57557_sb) );
na02s02 TIMEBOOST_cell_41976 ( .a(TIMEBOOST_net_13226), .b(g62989_sb), .o(n_5904) );
na02s01 TIMEBOOST_cell_37371 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__Q), .b(g58322_sb), .o(TIMEBOOST_net_10924) );
na02s01 TIMEBOOST_cell_37370 ( .a(TIMEBOOST_net_10923), .b(FE_OFN640_n_4669), .o(TIMEBOOST_net_9653) );
in01f02 g57558_u0 ( .a(FE_OFN2182_n_8567), .o(g57558_sb) );
na02f02 TIMEBOOST_cell_41408 ( .a(TIMEBOOST_net_12942), .b(g57262_sb), .o(n_11492) );
na03s01 TIMEBOOST_cell_34797 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__Q), .b(g63198_sb), .c(g63198_db), .o(n_5768) );
na02f02 TIMEBOOST_cell_44606 ( .a(TIMEBOOST_net_14541), .b(FE_OFN2189_n_8567), .o(TIMEBOOST_net_13011) );
in01f02 g57559_u0 ( .a(FE_OFN2175_n_8567), .o(g57559_sb) );
na02m02 TIMEBOOST_cell_32772 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__Q), .o(TIMEBOOST_net_10297) );
na02f02 TIMEBOOST_cell_22473 ( .a(FE_OCPN1827_n_14995), .b(TIMEBOOST_net_6493), .o(n_12710) );
na03s02 TIMEBOOST_cell_5288 ( .a(n_4473), .b(g64791_sb), .c(g64791_db), .o(n_4474) );
in01f01 g57560_u0 ( .a(FE_OFN1391_n_8567), .o(g57560_sb) );
na02s02 TIMEBOOST_cell_41988 ( .a(TIMEBOOST_net_13232), .b(g62556_sb), .o(n_6451) );
na02s02 TIMEBOOST_cell_37172 ( .a(TIMEBOOST_net_10824), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_9831) );
na02m02 TIMEBOOST_cell_31536 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_779), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_14__Q), .o(TIMEBOOST_net_9679) );
in01f02 g57561_u0 ( .a(FE_OFN1428_n_8567), .o(g57561_sb) );
na02f02 TIMEBOOST_cell_41410 ( .a(TIMEBOOST_net_12943), .b(g57126_sb), .o(n_10474) );
na02f02 TIMEBOOST_cell_44745 ( .a(FE_OFN1753_n_12086), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__Q), .o(TIMEBOOST_net_14611) );
na02s02 TIMEBOOST_cell_43230 ( .a(TIMEBOOST_net_13853), .b(FE_OFN1283_n_4097), .o(TIMEBOOST_net_12084) );
in01f02 g57562_u0 ( .a(FE_OFN2180_n_8567), .o(g57562_sb) );
na02m02 TIMEBOOST_cell_32770 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__Q), .o(TIMEBOOST_net_10296) );
na02f02 TIMEBOOST_cell_22475 ( .a(TIMEBOOST_net_6494), .b(FE_OCPN1827_n_14995), .o(n_12511) );
na02s01 TIMEBOOST_cell_43231 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__Q), .b(n_3552), .o(TIMEBOOST_net_13854) );
in01f02 g57563_u0 ( .a(FE_OFN2188_n_8567), .o(g57563_sb) );
na02f02 TIMEBOOST_cell_41412 ( .a(TIMEBOOST_net_12944), .b(g57432_sb), .o(n_11302) );
na02f02 TIMEBOOST_cell_44746 ( .a(TIMEBOOST_net_14611), .b(n_12406), .o(n_12729) );
na02f02 TIMEBOOST_cell_22477 ( .a(TIMEBOOST_net_6495), .b(FE_OCPN1827_n_14995), .o(n_12654) );
in01f02 g57564_u0 ( .a(FE_OFN1370_n_8567), .o(g57564_sb) );
na03s02 TIMEBOOST_cell_41989 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__Q), .b(n_3519), .c(FE_OFN1214_n_4151), .o(TIMEBOOST_net_13233) );
no02f04 TIMEBOOST_cell_37174 ( .a(TIMEBOOST_net_10825), .b(FE_RN_322_0), .o(FE_RN_323_0) );
na02m02 TIMEBOOST_cell_31534 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_778), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_13__Q), .o(TIMEBOOST_net_9678) );
in01f01 g57565_u0 ( .a(FE_OFN1345_n_8567), .o(g57565_sb) );
na02m02 TIMEBOOST_cell_16013 ( .a(TIMEBOOST_net_3263), .b(g56934_sb), .o(TIMEBOOST_net_2540) );
na02f01 g57565_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__Q), .b(FE_OFN1345_n_8567), .o(g57565_db) );
na02s01 TIMEBOOST_cell_36738 ( .a(TIMEBOOST_net_10607), .b(n_4743), .o(TIMEBOOST_net_206) );
in01f02 g57566_u0 ( .a(FE_OFN2177_n_8567), .o(g57566_sb) );
na02m02 TIMEBOOST_cell_32768 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__Q), .o(TIMEBOOST_net_10295) );
na02f02 TIMEBOOST_cell_45839 ( .a(n_9299), .b(n_9298), .o(TIMEBOOST_net_15158) );
na02f02 TIMEBOOST_cell_45840 ( .a(TIMEBOOST_net_15158), .b(n_10124), .o(TIMEBOOST_net_673) );
in01f01 g57567_u0 ( .a(FE_OFN1384_n_8567), .o(g57567_sb) );
na02s01 TIMEBOOST_cell_17666 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__Q), .b(g65285_sb), .o(TIMEBOOST_net_4090) );
na03s02 TIMEBOOST_cell_33199 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__Q), .b(FE_OFN653_n_4508), .c(g65433_sb), .o(TIMEBOOST_net_305) );
na02m02 TIMEBOOST_cell_45033 ( .a(g59383_sb), .b(n_3345), .o(TIMEBOOST_net_14755) );
in01f01 g57568_u0 ( .a(FE_OFN1394_n_8567), .o(g57568_sb) );
na02m02 TIMEBOOST_cell_44291 ( .a(n_9455), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__Q), .o(TIMEBOOST_net_14384) );
na02s01 TIMEBOOST_cell_37176 ( .a(TIMEBOOST_net_10826), .b(n_8832), .o(n_9230) );
na02s01 TIMEBOOST_cell_40381 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__Q), .b(g65391_sb), .o(TIMEBOOST_net_12429) );
in01f01 g57569_u0 ( .a(FE_OFN1408_n_8567), .o(g57569_sb) );
na02m02 TIMEBOOST_cell_31532 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_774), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_9__Q), .o(TIMEBOOST_net_9677) );
na02s02 TIMEBOOST_cell_43232 ( .a(TIMEBOOST_net_13854), .b(FE_OFN1212_n_4151), .o(TIMEBOOST_net_12083) );
in01f01 g57570_u0 ( .a(FE_OFN1387_n_8567), .o(g57570_sb) );
na02s01 TIMEBOOST_cell_42719 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__Q), .b(FE_OFN1793_n_9904), .o(TIMEBOOST_net_13598) );
na02s02 TIMEBOOST_cell_43143 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__Q), .b(n_3615), .o(TIMEBOOST_net_13810) );
na02s01 TIMEBOOST_cell_37178 ( .a(TIMEBOOST_net_10827), .b(TIMEBOOST_net_1065), .o(n_9120) );
in01f01 g57571_u0 ( .a(FE_OFN1349_n_8567), .o(g57571_sb) );
na02s02 TIMEBOOST_cell_45593 ( .a(TIMEBOOST_net_9347), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_15035) );
na02f02 TIMEBOOST_cell_43928 ( .a(TIMEBOOST_net_14202), .b(FE_OFN1405_n_8567), .o(TIMEBOOST_net_12880) );
na03f02 TIMEBOOST_cell_4172 ( .a(n_16842), .b(n_9328), .c(n_16843), .o(TIMEBOOST_net_666) );
in01f01 g57572_u0 ( .a(FE_OFN1391_n_8567), .o(g57572_sb) );
na02m02 TIMEBOOST_cell_43695 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__Q), .b(n_9850), .o(TIMEBOOST_net_14086) );
na02m02 TIMEBOOST_cell_31530 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_776), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_11__Q), .o(TIMEBOOST_net_9676) );
no02f08 TIMEBOOST_cell_37162 ( .a(TIMEBOOST_net_10819), .b(n_15744), .o(n_15755) );
in01f02 g57573_u0 ( .a(FE_OFN2180_n_8567), .o(g57573_sb) );
na02f02 TIMEBOOST_cell_41414 ( .a(TIMEBOOST_net_12945), .b(g57332_sb), .o(n_11418) );
na02f02 TIMEBOOST_cell_45841 ( .a(FE_RN_185_0), .b(n_10895), .o(TIMEBOOST_net_15159) );
in01f01 g57574_u0 ( .a(FE_OFN1412_n_8567), .o(g57574_sb) );
na02m02 TIMEBOOST_cell_43353 ( .a(TIMEBOOST_net_9968), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_13915) );
na02s02 TIMEBOOST_cell_43490 ( .a(TIMEBOOST_net_13983), .b(FE_OFN2063_n_6391), .o(TIMEBOOST_net_12617) );
na02s02 TIMEBOOST_cell_31528 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_65), .b(pci_target_unit_pcit_if_strd_addr_in_701), .o(TIMEBOOST_net_9675) );
in01f01 g57575_u0 ( .a(FE_OFN1389_n_8567), .o(g57575_sb) );
na02s02 TIMEBOOST_cell_42048 ( .a(TIMEBOOST_net_13262), .b(g62513_sb), .o(n_6553) );
na02s01 TIMEBOOST_cell_36687 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__Q), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_10582) );
na02s01 TIMEBOOST_cell_36686 ( .a(TIMEBOOST_net_10581), .b(FE_OFN1689_n_9528), .o(TIMEBOOST_net_9713) );
in01f01 g57576_u0 ( .a(FE_OFN1387_n_8567), .o(g57576_sb) );
na02s02 TIMEBOOST_cell_36689 ( .a(n_3970), .b(g62844_sb), .o(TIMEBOOST_net_10583) );
na02s01 TIMEBOOST_cell_36688 ( .a(TIMEBOOST_net_10582), .b(FE_OFN1668_n_9477), .o(TIMEBOOST_net_9708) );
in01f01 g57577_u0 ( .a(FE_OFN1387_n_8567), .o(g57577_sb) );
na03s02 TIMEBOOST_cell_42015 ( .a(n_3691), .b(n_3692), .c(FE_OFN1206_n_6356), .o(TIMEBOOST_net_13246) );
na02f02 TIMEBOOST_cell_36691 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_401), .b(TIMEBOOST_net_494), .o(TIMEBOOST_net_10584) );
na02s01 TIMEBOOST_cell_36690 ( .a(TIMEBOOST_net_10583), .b(g62844_db), .o(n_5283) );
in01f01 g57578_u0 ( .a(FE_OFN1382_n_8567), .o(g57578_sb) );
na02s01 TIMEBOOST_cell_30826 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__Q), .o(TIMEBOOST_net_9324) );
na02f02 TIMEBOOST_cell_44550 ( .a(TIMEBOOST_net_14513), .b(FE_OFN2167_n_8567), .o(TIMEBOOST_net_13464) );
na02s02 TIMEBOOST_cell_31024 ( .a(n_4488), .b(g64842_sb), .o(TIMEBOOST_net_9423) );
in01f01 g57579_u0 ( .a(FE_OFN1387_n_8567), .o(g57579_sb) );
na02m02 TIMEBOOST_cell_41611 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_15__Q), .b(n_9856), .o(TIMEBOOST_net_13044) );
na02f02 TIMEBOOST_cell_36693 ( .a(TIMEBOOST_net_1725), .b(g54147_db), .o(TIMEBOOST_net_10585) );
na02f02 TIMEBOOST_cell_36692 ( .a(TIMEBOOST_net_10584), .b(g54135_sb), .o(n_13463) );
in01f01 g57580_u0 ( .a(FE_OFN1389_n_8567), .o(g57580_sb) );
na02f02 TIMEBOOST_cell_41612 ( .a(FE_OFN1436_n_9372), .b(TIMEBOOST_net_13044), .o(TIMEBOOST_net_11665) );
na02s01 TIMEBOOST_cell_37676 ( .a(TIMEBOOST_net_11076), .b(g62066_sb), .o(n_7833) );
na02f02 TIMEBOOST_cell_22271 ( .a(TIMEBOOST_net_6392), .b(n_10577), .o(n_12137) );
in01f02 g57581_u0 ( .a(FE_OFN2177_n_8567), .o(g57581_sb) );
na02m02 TIMEBOOST_cell_32766 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__Q), .o(TIMEBOOST_net_10294) );
na02f02 TIMEBOOST_cell_43696 ( .a(TIMEBOOST_net_14086), .b(FE_OFN1349_n_8567), .o(TIMEBOOST_net_13309) );
na02f02 g55392_u0 ( .a(FE_OFN1577_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__Q), .o(n_12328) );
in01f02 g57582_u0 ( .a(FE_OFN2179_n_8567), .o(g57582_sb) );
na02f02 TIMEBOOST_cell_41416 ( .a(TIMEBOOST_net_12946), .b(g57081_sb), .o(n_11661) );
na03s02 TIMEBOOST_cell_4955 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .b(g57797_sb), .c(FE_OFN276_n_9941), .o(TIMEBOOST_net_618) );
na02s01 TIMEBOOST_cell_42620 ( .a(TIMEBOOST_net_13548), .b(g64788_db), .o(n_3762) );
in01f01 g57583_u0 ( .a(FE_OFN1412_n_8567), .o(g57583_sb) );
na02m02 TIMEBOOST_cell_41613 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_12__Q), .b(FE_OFN209_n_9126), .o(TIMEBOOST_net_13045) );
na02s01 TIMEBOOST_cell_39680 ( .a(TIMEBOOST_net_12078), .b(g62591_sb), .o(n_6371) );
na02m02 TIMEBOOST_cell_31518 ( .a(n_2261), .b(g63196_sb), .o(TIMEBOOST_net_9670) );
in01f01 g57584_u0 ( .a(FE_OFN1396_n_8567), .o(g57584_sb) );
na02f02 TIMEBOOST_cell_41614 ( .a(FE_OFN1441_n_9372), .b(TIMEBOOST_net_13045), .o(TIMEBOOST_net_11683) );
na02s02 TIMEBOOST_cell_43578 ( .a(TIMEBOOST_net_14027), .b(FE_OFN1323_n_6436), .o(TIMEBOOST_net_12229) );
na03f08 TIMEBOOST_cell_4960 ( .a(n_15735), .b(n_15736), .c(n_15739), .o(n_16486) );
na02m02 TIMEBOOST_cell_41615 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_21__Q), .b(FE_OFN223_n_9844), .o(TIMEBOOST_net_13046) );
na02f01 g57585_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q), .b(FE_OFN1379_n_8567), .o(g57585_db) );
na02s02 TIMEBOOST_cell_42077 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__Q), .b(n_4333), .o(TIMEBOOST_net_13277) );
in01f02 g57586_u0 ( .a(FE_OFN2170_n_8567), .o(g57586_sb) );
na02m02 TIMEBOOST_cell_32764 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__Q), .o(TIMEBOOST_net_10293) );
na02f02 TIMEBOOST_cell_41358 ( .a(TIMEBOOST_net_12917), .b(g57099_sb), .o(n_10481) );
na02s01 TIMEBOOST_cell_45394 ( .a(TIMEBOOST_net_14935), .b(FE_OFN1135_g64577_p), .o(n_5388) );
in01f01 g57587_u0 ( .a(FE_OFN1391_n_8567), .o(g57587_sb) );
na02s02 TIMEBOOST_cell_42078 ( .a(TIMEBOOST_net_13277), .b(n_6232), .o(TIMEBOOST_net_11577) );
na02f02 TIMEBOOST_cell_36694 ( .a(TIMEBOOST_net_10585), .b(g54147_sb), .o(n_13453) );
na02f02 TIMEBOOST_cell_36697 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_410), .b(TIMEBOOST_net_490), .o(TIMEBOOST_net_10587) );
in01f02 g57588_u0 ( .a(FE_OFN2184_n_8567), .o(g57588_sb) );
na02f02 TIMEBOOST_cell_32763 ( .a(FE_OFN1742_n_11019), .b(TIMEBOOST_net_10292), .o(TIMEBOOST_net_6536) );
na02s02 TIMEBOOST_cell_45395 ( .a(n_3563), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__Q), .o(TIMEBOOST_net_14936) );
na02s01 TIMEBOOST_cell_43548 ( .a(TIMEBOOST_net_14012), .b(g62387_sb), .o(n_6826) );
in01f01 g57589_u0 ( .a(FE_OFN1409_n_8567), .o(g57589_sb) );
na02s02 TIMEBOOST_cell_42079 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q), .b(n_4462), .o(TIMEBOOST_net_13278) );
na02f02 TIMEBOOST_cell_36696 ( .a(TIMEBOOST_net_10586), .b(TIMEBOOST_net_503), .o(FE_RN_367_0) );
na02s02 TIMEBOOST_cell_36699 ( .a(TIMEBOOST_net_326), .b(g61891_sb), .o(TIMEBOOST_net_10588) );
in01f01 g57590_u0 ( .a(FE_OFN1374_n_8567), .o(g57590_sb) );
na02s02 TIMEBOOST_cell_42080 ( .a(TIMEBOOST_net_13278), .b(n_6645), .o(TIMEBOOST_net_11576) );
na02f02 TIMEBOOST_cell_36698 ( .a(TIMEBOOST_net_10587), .b(g54145_sb), .o(n_13455) );
na02s02 TIMEBOOST_cell_36701 ( .a(TIMEBOOST_net_328), .b(g61895_sb), .o(TIMEBOOST_net_10589) );
in01f02 g57591_u0 ( .a(FE_OFN2170_n_8567), .o(g57591_sb) );
na02m02 TIMEBOOST_cell_32762 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__14__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__14__Q), .o(TIMEBOOST_net_10292) );
no04f04 TIMEBOOST_cell_4967 ( .a(FE_RN_669_0), .b(FE_RN_671_0), .c(FE_RN_674_0), .d(FE_RN_670_0), .o(FE_RN_675_0) );
na02s01 TIMEBOOST_cell_36700 ( .a(TIMEBOOST_net_10588), .b(g61891_db), .o(n_8047) );
in01f01 g57592_u0 ( .a(FE_OFN1412_n_8567), .o(g57592_sb) );
na02s02 TIMEBOOST_cell_36703 ( .a(TIMEBOOST_net_330), .b(g61897_sb), .o(TIMEBOOST_net_10590) );
na02s01 TIMEBOOST_cell_36702 ( .a(TIMEBOOST_net_10589), .b(g61895_db), .o(n_8036) );
in01f01 g57593_u0 ( .a(FE_OFN1399_n_8567), .o(g57593_sb) );
na02f02 TIMEBOOST_cell_43756 ( .a(TIMEBOOST_net_14116), .b(FE_OFN1413_n_8567), .o(TIMEBOOST_net_12810) );
na02f02 TIMEBOOST_cell_37100 ( .a(TIMEBOOST_net_10788), .b(n_12588), .o(n_12850) );
na03m02 TIMEBOOST_cell_4972 ( .a(n_15065), .b(wbu_map_in_131), .c(n_2341), .o(n_3017) );
in01f02 g57594_u0 ( .a(FE_OFN1427_n_8567), .o(g57594_sb) );
na02f02 TIMEBOOST_cell_41374 ( .a(TIMEBOOST_net_12925), .b(g57133_sb), .o(n_10470) );
na02m02 TIMEBOOST_cell_43779 ( .a(n_9001), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__Q), .o(TIMEBOOST_net_14128) );
na02f02 TIMEBOOST_cell_41338 ( .a(TIMEBOOST_net_12907), .b(g57103_sb), .o(n_11642) );
in01f01 g57595_u0 ( .a(FE_OFN1425_n_8567), .o(g57595_sb) );
na02s02 TIMEBOOST_cell_43386 ( .a(TIMEBOOST_net_13931), .b(n_6319), .o(TIMEBOOST_net_12209) );
na02s01 TIMEBOOST_cell_15822 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_80), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3168) );
na02s01 TIMEBOOST_cell_15826 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_85), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3170) );
in01f01 g57596_u0 ( .a(FE_OFN1402_n_8567), .o(g57596_sb) );
na02f02 TIMEBOOST_cell_41568 ( .a(TIMEBOOST_net_13022), .b(g57215_sb), .o(n_11543) );
na02m02 TIMEBOOST_cell_31506 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_772), .b(g54040_sb), .o(TIMEBOOST_net_9664) );
na02f02 TIMEBOOST_cell_37079 ( .a(FE_OCP_RBN1996_n_13971), .b(TIMEBOOST_net_10235), .o(TIMEBOOST_net_10778) );
in01f01 g57597_u0 ( .a(FE_OFN1416_n_8567), .o(g57597_sb) );
na02s02 TIMEBOOST_cell_45396 ( .a(TIMEBOOST_net_14936), .b(FE_OFN1194_n_6935), .o(TIMEBOOST_net_12576) );
na02f02 TIMEBOOST_cell_37078 ( .a(TIMEBOOST_net_10777), .b(FE_OFN1587_n_13736), .o(g53267_p) );
na02f02 TIMEBOOST_cell_37081 ( .a(FE_OCP_RBN1998_n_13971), .b(TIMEBOOST_net_10240), .o(TIMEBOOST_net_10779) );
in01f01 g57598_u0 ( .a(FE_OFN1377_n_8567), .o(g57598_sb) );
na02f02 TIMEBOOST_cell_42538 ( .a(n_12124), .b(TIMEBOOST_net_13507), .o(n_12715) );
na02s01 TIMEBOOST_cell_30884 ( .a(pci_target_unit_pcit_if_strd_addr_in_706), .b(pci_target_unit_del_sync_addr_in_224), .o(TIMEBOOST_net_9353) );
na03s02 TIMEBOOST_cell_4980 ( .a(g58115_sb), .b(g58115_db), .c(FE_OFN262_n_9851), .o(n_9678) );
na02f02 g57641_u0 ( .a(n_8842), .b(FE_OFN276_n_9941), .o(n_9160) );
na02f02 TIMEBOOST_cell_4065 ( .a(TIMEBOOST_net_612), .b(n_17040), .o(n_4878) );
in01f04 g57644_u0 ( .a(n_8800), .o(n_8801) );
no02s01 g57646_u0 ( .a(n_3330), .b(FE_OFN778_n_4152), .o(n_4153) );
na02f02 g57648_u0 ( .a(n_8794), .b(pci_target_unit_fifos_pcir_flush_in), .o(n_8871) );
no02s02 g57649_u0 ( .a(n_3329), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8662) );
na02f02 g57654_u0 ( .a(n_16535), .b(n_8866), .o(n_16888) );
in01f04 g57667_u0 ( .a(n_8932), .o(n_10588) );
na02f02 g57668_u0 ( .a(n_16535), .b(n_16105), .o(n_8932) );
in01f08 g57671_u0 ( .a(n_15589), .o(n_10680) );
in01f03 g57676_u0 ( .a(n_16572), .o(n_9991) );
in01f06 g57698_u0 ( .a(n_8864), .o(n_10566) );
na02f04 g57699_u0 ( .a(n_8863), .b(n_8866), .o(n_8864) );
in01f02 g57700_u0 ( .a(n_8928), .o(n_9320) );
na02f02 g57710_u0 ( .a(n_16579), .b(n_16535), .o(n_8928) );
in01f02 g57725_u0 ( .a(n_8861), .o(n_9975) );
na02f02 g57726_u0 ( .a(n_16566), .b(n_8866), .o(n_8861) );
in01f10 g57734_u0 ( .a(FE_OCPN1905_n_8927), .o(n_11728) );
in01f04 g57735_u0 ( .a(FE_OCPN1905_n_8927), .o(n_10185) );
in01f02 g57736_u0 ( .a(FE_OCPN1905_n_8927), .o(n_10141) );
in01f02 g57737_u0 ( .a(FE_OCPN1905_n_8927), .o(n_10232) );
in01f01 g57738_u0 ( .a(n_8927), .o(n_10195) );
na02f02 g57739_u0 ( .a(n_8860), .b(n_16535), .o(n_8927) );
in01f04 g57747_u0 ( .a(n_9155), .o(n_10143) );
na02f03 g57751_u0 ( .a(n_8863), .b(n_15453), .o(n_9155) );
in01f03 g57755_u0 ( .a(n_8859), .o(n_10853) );
na02f02 g57756_u0 ( .a(n_8863), .b(n_8860), .o(n_8859) );
in01f02 g57759_u0 ( .a(n_15560), .o(n_10693) );
in01f02 g57770_u0 ( .a(n_8857), .o(n_10892) );
na02f02 g57771_u0 ( .a(n_8867), .b(n_8860), .o(n_8857) );
na02m02 g57779_u1 ( .a(n_6136), .b(g56934_sb), .o(g57779_da) );
na02s02 TIMEBOOST_cell_19299 ( .a(TIMEBOOST_net_4906), .b(g60657_sb), .o(n_5664) );
na02s01 TIMEBOOST_cell_32036 ( .a(configuration_pci_err_addr_484), .b(wbm_adr_o_14_), .o(TIMEBOOST_net_9929) );
in01s03 g57780_u0 ( .a(pci_target_unit_fifos_pcir_flush_in), .o(g57780_sb) );
na02s01 g57780_u1 ( .a(n_7835), .b(g57780_sb), .o(g57780_da) );
na02f02 TIMEBOOST_cell_4116 ( .a(n_2904), .b(n_3034), .o(TIMEBOOST_net_638) );
na02s02 TIMEBOOST_cell_38180 ( .a(TIMEBOOST_net_11328), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_4658) );
na02s01 g57781_u1 ( .a(n_7569), .b(g57780_sb), .o(g57781_da) );
na02s02 TIMEBOOST_cell_37878 ( .a(TIMEBOOST_net_11177), .b(g57925_sb), .o(n_9885) );
na02m02 TIMEBOOST_cell_44517 ( .a(n_9200), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__Q), .o(TIMEBOOST_net_14497) );
na02s02 TIMEBOOST_cell_42952 ( .a(TIMEBOOST_net_13714), .b(g58348_sb), .o(n_9473) );
na02f02 TIMEBOOST_cell_4063 ( .a(TIMEBOOST_net_611), .b(n_17049), .o(n_4881) );
na02f02 TIMEBOOST_cell_41084 ( .a(TIMEBOOST_net_12780), .b(g57276_sb), .o(n_11478) );
na02s02 TIMEBOOST_cell_32023 ( .a(TIMEBOOST_net_9922), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_4904) );
na02s01 TIMEBOOST_cell_36386 ( .a(TIMEBOOST_net_10431), .b(g65719_db), .o(n_2066) );
na03s02 TIMEBOOST_cell_42699 ( .a(g58152_sb), .b(g58152_db), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__Q), .o(TIMEBOOST_net_13588) );
na02s01 TIMEBOOST_cell_45648 ( .a(TIMEBOOST_net_15062), .b(g61836_db), .o(n_6975) );
na02f02 TIMEBOOST_cell_12788 ( .a(FE_OFN1599_n_13995), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__Q), .o(TIMEBOOST_net_2961) );
na02s02 TIMEBOOST_cell_43092 ( .a(TIMEBOOST_net_13784), .b(g58305_db), .o(n_9506) );
na02s02 TIMEBOOST_cell_44853 ( .a(n_4473), .b(g64969_sb), .o(TIMEBOOST_net_14665) );
na02s01 TIMEBOOST_cell_36369 ( .a(FE_OFN945_n_2248), .b(g65849_sb), .o(TIMEBOOST_net_10423) );
na02f02 TIMEBOOST_cell_44747 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__28__Q), .b(FE_OFN1753_n_12086), .o(TIMEBOOST_net_14612) );
na02s01 TIMEBOOST_cell_45580 ( .a(TIMEBOOST_net_15028), .b(n_4452), .o(TIMEBOOST_net_10935) );
na02s02 TIMEBOOST_cell_37538 ( .a(TIMEBOOST_net_11007), .b(FE_OFN712_n_8140), .o(TIMEBOOST_net_4171) );
na02m02 TIMEBOOST_cell_43775 ( .a(n_9107), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__Q), .o(TIMEBOOST_net_14126) );
na02s01 g57787_u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_), .b(g56933_sb), .o(g57787_da) );
na03s02 TIMEBOOST_cell_39359 ( .a(n_1923), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__Q), .c(FE_OFN2081_n_8176), .o(TIMEBOOST_net_11918) );
na03s02 TIMEBOOST_cell_34260 ( .a(TIMEBOOST_net_9815), .b(FE_OFN1168_n_5592), .c(g62098_sb), .o(n_5606) );
na02s01 g57788_u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_), .b(g56933_sb), .o(g57788_da) );
na02s02 TIMEBOOST_cell_43410 ( .a(TIMEBOOST_net_13943), .b(n_6287), .o(TIMEBOOST_net_12207) );
na02f02 TIMEBOOST_cell_41086 ( .a(TIMEBOOST_net_12781), .b(g57427_sb), .o(n_11307) );
na02s01 g57789_u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_), .b(g56933_sb), .o(g57789_da) );
na02f02 TIMEBOOST_cell_4075 ( .a(TIMEBOOST_net_617), .b(n_4619), .o(n_7214) );
na02f02 TIMEBOOST_cell_4211 ( .a(TIMEBOOST_net_685), .b(n_16987), .o(n_12166) );
in01s40 g57790_u0 ( .a(parchk_pci_cbe_en_in), .o(g57790_sb) );
na02s02 TIMEBOOST_cell_42087 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__Q), .b(n_3709), .o(TIMEBOOST_net_13282) );
na02f02 TIMEBOOST_cell_4117 ( .a(TIMEBOOST_net_638), .b(n_4119), .o(n_4856) );
na02s01 TIMEBOOST_cell_16576 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__28__Q), .b(g64336_sb), .o(TIMEBOOST_net_3545) );
na02f02 TIMEBOOST_cell_41188 ( .a(TIMEBOOST_net_12832), .b(g57275_sb), .o(n_11479) );
na02m02 TIMEBOOST_cell_3989 ( .a(TIMEBOOST_net_574), .b(n_7626), .o(n_8487) );
na02f04 TIMEBOOST_cell_3990 ( .a(n_16163), .b(n_3422), .o(TIMEBOOST_net_575) );
in01f04 g57792_u0 ( .a(n_9173), .o(n_9152) );
in01f06 g57794_u0 ( .a(n_8747), .o(g57794_sb) );
na02f10 g57794_u1 ( .a(g57794_sb), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(g57794_da) );
na02f10 g57794_u2 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__Q), .b(n_8747), .o(g57794_db) );
na02f10 g57794_u3 ( .a(g57794_da), .b(g57794_db), .o(n_9173) );
in01s02 g57795_u0 ( .a(FE_OFN276_n_9941), .o(g57795_sb) );
na02s01 g57795_u1 ( .a(n_4939), .b(g57795_sb), .o(g57795_da) );
na02m02 TIMEBOOST_cell_3982 ( .a(n_2753), .b(n_1355), .o(TIMEBOOST_net_571) );
na02s02 TIMEBOOST_cell_32035 ( .a(TIMEBOOST_net_9928), .b(FE_OFN1180_n_3476), .o(TIMEBOOST_net_4910) );
na02s02 TIMEBOOST_cell_40375 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__Q), .b(g58353_sb), .o(TIMEBOOST_net_12426) );
na02m02 TIMEBOOST_cell_12622 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__Q), .o(TIMEBOOST_net_2878) );
na02s02 TIMEBOOST_cell_39456 ( .a(TIMEBOOST_net_11966), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_4650) );
in01s04 g57797_u0 ( .a(FE_OFN276_n_9941), .o(g57797_sb) );
na03s02 TIMEBOOST_cell_40601 ( .a(n_74), .b(n_4378), .c(FE_OFN1261_n_4143), .o(TIMEBOOST_net_12539) );
na02s01 TIMEBOOST_cell_38182 ( .a(TIMEBOOST_net_11329), .b(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_4489) );
na02s02 TIMEBOOST_cell_38666 ( .a(TIMEBOOST_net_11571), .b(g62630_sb), .o(n_6295) );
na02s02 TIMEBOOST_cell_45397 ( .a(n_3559), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__Q), .o(TIMEBOOST_net_14937) );
na02f04 TIMEBOOST_cell_3991 ( .a(TIMEBOOST_net_575), .b(n_5722), .o(n_8452) );
na02s01 TIMEBOOST_cell_44816 ( .a(TIMEBOOST_net_14646), .b(g58230_db), .o(n_9047) );
na02f02 TIMEBOOST_cell_41180 ( .a(TIMEBOOST_net_12828), .b(g57381_sb), .o(n_11365) );
na02s01 TIMEBOOST_cell_44817 ( .a(n_3780), .b(g64977_sb), .o(TIMEBOOST_net_14647) );
na02m01 TIMEBOOST_cell_3994 ( .a(n_1299), .b(n_15370), .o(TIMEBOOST_net_577) );
na02m02 TIMEBOOST_cell_32760 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__Q), .o(TIMEBOOST_net_10291) );
na02m01 TIMEBOOST_cell_3995 ( .a(n_16520), .b(TIMEBOOST_net_577), .o(n_8660) );
na02s01 TIMEBOOST_cell_44918 ( .a(TIMEBOOST_net_14697), .b(g65832_sb), .o(TIMEBOOST_net_330) );
na02s02 TIMEBOOST_cell_45398 ( .a(TIMEBOOST_net_14937), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_12572) );
na02s01 TIMEBOOST_cell_18529 ( .a(TIMEBOOST_net_4521), .b(g62845_sb), .o(n_5281) );
na02s01 TIMEBOOST_cell_39682 ( .a(TIMEBOOST_net_12079), .b(g62585_sb), .o(n_6382) );
na02f02 TIMEBOOST_cell_32759 ( .a(FE_OFN1738_n_11019), .b(TIMEBOOST_net_10290), .o(TIMEBOOST_net_6534) );
na02s02 TIMEBOOST_cell_40794 ( .a(TIMEBOOST_net_12635), .b(g62931_sb), .o(n_6019) );
na02s01 TIMEBOOST_cell_4000 ( .a(n_16818), .b(wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q), .o(TIMEBOOST_net_580) );
in01f01 g57803_u0 ( .a(n_16368), .o(n_8926) );
na03s01 TIMEBOOST_cell_6011 ( .a(n_2048), .b(g61734_sb), .c(g61734_db), .o(n_8351) );
na02m02 g57850_u0 ( .a(n_3363), .b(n_8571), .o(n_8688) );
na03s02 TIMEBOOST_cell_43297 ( .a(n_4304), .b(FE_OFN1206_n_6356), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__Q), .o(TIMEBOOST_net_13887) );
na02s02 TIMEBOOST_cell_43549 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__20__Q), .b(n_3754), .o(TIMEBOOST_net_14013) );
na02f02 g57856_u0 ( .a(n_15515), .b(n_15517), .o(g57856_p) );
in01f02 g57856_u1 ( .a(g57856_p), .o(n_8939) );
in01f02 g57857_u0 ( .a(n_8924), .o(n_16605) );
na02f04 g57858_u0 ( .a(n_8790), .b(n_8792), .o(n_8924) );
na02f04 g57863_u0 ( .a(n_16537), .b(n_16534), .o(g57863_p) );
in01f04 g57863_u1 ( .a(g57863_p), .o(n_8863) );
na02f02 g57864_u0 ( .a(n_8686), .b(n_16533), .o(g57864_p) );
in01f02 g57864_u1 ( .a(g57864_p), .o(n_8867) );
no02f04 g57865_u0 ( .a(n_8790), .b(n_15517), .o(n_9171) );
in01f02 g57867_u0 ( .a(n_15581), .o(n_10258) );
oa12f01 g57871_u0 ( .a(n_9143), .b(wishbone_slave_unit_fifos_wbw_inTransactionCount_1_), .c(n_9144), .o(n_9146) );
oa12s02 g57872_u0 ( .a(n_8575), .b(pci_target_unit_pci_target_sm_rd_request), .c(FE_OFN2093_n_2301), .o(n_8687) );
oa12f01 g57874_u0 ( .a(n_9143), .b(wishbone_slave_unit_fifos_inGreyCount_0_), .c(n_9144), .o(n_9145) );
in01f01 g57875_u0 ( .a(n_9144), .o(g57875_sb) );
na02f02 TIMEBOOST_cell_37080 ( .a(TIMEBOOST_net_10778), .b(FE_OFN1588_n_13736), .o(g53250_p) );
na03s02 TIMEBOOST_cell_38361 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__Q), .b(FE_OFN1130_g64577_p), .c(n_3881), .o(TIMEBOOST_net_11419) );
na02s02 TIMEBOOST_cell_36705 ( .a(TIMEBOOST_net_335), .b(g61889_sb), .o(TIMEBOOST_net_10591) );
no02s01 g57876_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_12_), .b(n_3024), .o(g57876_p) );
ao12s01 g57876_u1 ( .a(g57876_p), .b(pci_target_unit_del_sync_comp_cycle_count_12_), .c(n_3024), .o(n_3330) );
ao12m02 g57877_u0 ( .a(n_5754), .b(conf_wb_err_addr_in_971), .c(FE_OFN1145_n_15261), .o(n_7362) );
no02s02 g57878_u0 ( .a(n_206), .b(n_3073), .o(g57878_p) );
ao12s02 g57878_u1 ( .a(g57878_p), .b(n_206), .c(n_3073), .o(n_3329) );
ao12s01 g57879_u0 ( .a(n_8971), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__Q), .c(FE_OFN601_n_9687), .o(n_9928) );
ao12s01 g57880_u0 ( .a(n_8970), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__Q), .c(FE_OFN562_n_9895), .o(n_9926) );
ao12s01 g57881_u0 ( .a(n_8968), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__Q), .c(FE_OFN554_n_9864), .o(n_9924) );
ao12s01 g57882_u0 ( .a(n_8967), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__Q), .c(FE_OFN519_n_9697), .o(n_9922) );
ao12s01 g57883_u0 ( .a(n_8966), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__Q), .c(FE_OFN587_n_9692), .o(n_9920) );
ao12s01 g57884_u0 ( .a(n_8965), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__Q), .c(FE_OFN532_n_9823), .o(n_9918) );
ao12s01 g57885_u0 ( .a(n_8964), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__Q), .c(FE_OFN595_n_9694), .o(n_9916) );
ao12s01 g57886_u0 ( .a(n_8963), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__Q), .c(FE_OFN529_n_9899), .o(n_9914) );
ao12s01 g57887_u0 ( .a(n_8962), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__Q), .c(FE_OFN606_n_9904), .o(n_9912) );
ao12s01 g57888_u0 ( .a(n_8961), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__Q), .c(FE_OFN1803_n_9690), .o(n_9910) );
ao12s01 g57889_u0 ( .a(n_8960), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q), .c(FE_OFN577_n_9902), .o(n_9908) );
in01s01 g57890_u0 ( .a(FE_OFN576_n_9902), .o(g57890_sb) );
na02s01 g57890_u1 ( .a(FE_OFN205_n_9140), .b(g57890_sb), .o(g57890_da) );
na02s01 g57890_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__Q), .b(FE_OFN576_n_9902), .o(g57890_db) );
na02s01 g57890_u3 ( .a(g57890_da), .b(g57890_db), .o(n_9142) );
in01s01 g57891_u0 ( .a(FE_OFN562_n_9895), .o(g57891_sb) );
na04s02 TIMEBOOST_cell_34337 ( .a(n_2692), .b(g63193_sb), .c(g53942_db), .d(TIMEBOOST_net_890), .o(n_13503) );
na02s01 g57891_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__Q), .b(FE_OFN562_n_9895), .o(g57891_db) );
na02s02 TIMEBOOST_cell_19319 ( .a(TIMEBOOST_net_4916), .b(g60611_sb), .o(n_4843) );
in01s01 g57892_u0 ( .a(FE_OFN564_n_9895), .o(g57892_sb) );
na02s01 g57892_u1 ( .a(FE_OFN203_n_9228), .b(g57892_sb), .o(g57892_da) );
na02s01 g57892_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__Q), .b(FE_OFN564_n_9895), .o(g57892_db) );
na02s01 g57892_u3 ( .a(g57892_da), .b(g57892_db), .o(n_9232) );
in01s01 g57893_u0 ( .a(FE_OFN562_n_9895), .o(g57893_sb) );
na02s02 TIMEBOOST_cell_40408 ( .a(TIMEBOOST_net_12442), .b(FE_OFN2212_n_8407), .o(TIMEBOOST_net_1751) );
na02s01 g57893_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__Q), .b(FE_OFN562_n_9895), .o(g57893_db) );
na02s01 TIMEBOOST_cell_44919 ( .a(TIMEBOOST_net_9508), .b(FE_OFN1044_n_2037), .o(TIMEBOOST_net_14698) );
in01s01 g57894_u0 ( .a(FE_OFN554_n_9864), .o(g57894_sb) );
na02f02 TIMEBOOST_cell_42539 ( .a(FE_OFN1759_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__Q), .o(TIMEBOOST_net_13508) );
na02s01 g57894_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__Q), .b(FE_OFN554_n_9864), .o(g57894_db) );
na02s02 TIMEBOOST_cell_19321 ( .a(TIMEBOOST_net_4917), .b(g60613_sb), .o(n_4841) );
in01s01 g57895_u0 ( .a(FE_OFN556_n_9864), .o(g57895_sb) );
na02f02 TIMEBOOST_cell_42540 ( .a(n_11923), .b(TIMEBOOST_net_13508), .o(n_12491) );
na02s01 g57895_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__Q), .b(FE_OFN556_n_9864), .o(g57895_db) );
na02s02 TIMEBOOST_cell_19323 ( .a(TIMEBOOST_net_4918), .b(g60615_sb), .o(n_4839) );
in01s01 g57896_u0 ( .a(FE_OFN554_n_9864), .o(g57896_sb) );
na02s01 TIMEBOOST_cell_40452 ( .a(TIMEBOOST_net_12464), .b(g62125_sb), .o(n_5571) );
na02s01 g57896_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__Q), .b(FE_OFN554_n_9864), .o(g57896_db) );
na02s01 TIMEBOOST_cell_16188 ( .a(pci_target_unit_fifos_pciw_addr_data_in_124), .b(g64085_sb), .o(TIMEBOOST_net_3351) );
in01s01 g57897_u0 ( .a(FE_OFN532_n_9823), .o(g57897_sb) );
na02f06 TIMEBOOST_cell_42541 ( .a(FE_OCP_RBN1976_n_12381), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__Q), .o(TIMEBOOST_net_13509) );
na02s01 g57897_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__Q), .b(FE_OFN532_n_9823), .o(g57897_db) );
na02s02 TIMEBOOST_cell_19325 ( .a(TIMEBOOST_net_4919), .b(g60617_sb), .o(n_4837) );
in01s01 g57898_u0 ( .a(FE_OFN534_n_9823), .o(g57898_sb) );
na02s02 TIMEBOOST_cell_38622 ( .a(TIMEBOOST_net_11549), .b(g62554_sb), .o(n_6456) );
na02s01 g57898_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__Q), .b(FE_OFN534_n_9823), .o(g57898_db) );
na02s01 TIMEBOOST_cell_38184 ( .a(TIMEBOOST_net_11330), .b(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_4518) );
in01s01 g57899_u0 ( .a(FE_OFN532_n_9823), .o(g57899_sb) );
in01s01 TIMEBOOST_cell_45958 ( .a(TIMEBOOST_net_15264), .o(TIMEBOOST_net_15265) );
na02s01 g57899_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__Q), .b(FE_OFN532_n_9823), .o(g57899_db) );
na02s01 TIMEBOOST_cell_32034 ( .a(configuration_pci_err_data_505), .b(wbm_dat_o_4_), .o(TIMEBOOST_net_9928) );
in01s01 g57900_u0 ( .a(FE_OFN529_n_9899), .o(g57900_sb) );
na02f06 TIMEBOOST_cell_42542 ( .a(n_16402), .b(TIMEBOOST_net_13509), .o(n_16403) );
na02s01 g57900_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__Q), .b(FE_OFN529_n_9899), .o(g57900_db) );
na03s02 TIMEBOOST_cell_38101 ( .a(TIMEBOOST_net_4252), .b(g64086_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__Q), .o(TIMEBOOST_net_11289) );
in01s01 g57901_u0 ( .a(FE_OFN528_n_9899), .o(g57901_sb) );
na02s01 g57901_u1 ( .a(FE_OFN203_n_9228), .b(g57901_sb), .o(g57901_da) );
na02s01 g57901_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__Q), .b(FE_OFN528_n_9899), .o(g57901_db) );
na02s01 g57901_u3 ( .a(g57901_da), .b(g57901_db), .o(n_9224) );
in01s01 g57902_u0 ( .a(FE_OFN529_n_9899), .o(g57902_sb) );
na02f04 TIMEBOOST_cell_39520 ( .a(TIMEBOOST_net_11998), .b(g54148_sb), .o(n_13452) );
na02s01 g57902_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__Q), .b(FE_OFN529_n_9899), .o(g57902_db) );
na02m02 TIMEBOOST_cell_44149 ( .a(n_9035), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__Q), .o(TIMEBOOST_net_14313) );
in01s01 g57903_u0 ( .a(FE_OFN606_n_9904), .o(g57903_sb) );
na02m08 TIMEBOOST_cell_42543 ( .a(pci_trdy_i), .b(parchk_pci_trdy_en_in), .o(TIMEBOOST_net_13510) );
na02s01 g57903_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__Q), .b(FE_OFN606_n_9904), .o(g57903_db) );
na02s02 TIMEBOOST_cell_19331 ( .a(TIMEBOOST_net_4922), .b(g60638_sb), .o(n_5694) );
in01s01 g57904_u0 ( .a(FE_OFN606_n_9904), .o(g57904_sb) );
in01s01 TIMEBOOST_cell_45891 ( .a(n_9168), .o(TIMEBOOST_net_15198) );
na02s01 g57904_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__Q), .b(FE_OFN606_n_9904), .o(g57904_db) );
na02s02 TIMEBOOST_cell_38034 ( .a(TIMEBOOST_net_11255), .b(g61756_sb), .o(n_8302) );
in01s01 g57905_u0 ( .a(FE_OFN606_n_9904), .o(g57905_sb) );
na02s01 g57905_u1 ( .a(FE_OFN205_n_9140), .b(g57905_sb), .o(g57905_da) );
na02s01 g57905_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__Q), .b(FE_OFN606_n_9904), .o(g57905_db) );
na02s01 g57905_u3 ( .a(g57905_da), .b(g57905_db), .o(n_9136) );
in01s01 g57906_u0 ( .a(FE_OFN576_n_9902), .o(g57906_sb) );
na02s02 TIMEBOOST_cell_43115 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__Q), .b(n_3533), .o(TIMEBOOST_net_13796) );
na02s01 g57906_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__Q), .b(FE_OFN576_n_9902), .o(g57906_db) );
na02s02 TIMEBOOST_cell_19335 ( .a(TIMEBOOST_net_4924), .b(g60604_sb), .o(n_4851) );
in01s01 g57907_u0 ( .a(FE_OFN576_n_9902), .o(g57907_sb) );
na02s01 g57907_u1 ( .a(FE_OFN203_n_9228), .b(g57907_sb), .o(g57907_da) );
na02s01 g57907_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__Q), .b(FE_OFN576_n_9902), .o(g57907_db) );
na02s01 g57907_u3 ( .a(g57907_da), .b(g57907_db), .o(n_9220) );
in01f01 g57908_u0 ( .a(n_9144), .o(g57908_sb) );
na02s01 TIMEBOOST_cell_36704 ( .a(TIMEBOOST_net_10590), .b(g61897_db), .o(n_8032) );
no02f06 TIMEBOOST_cell_20068 ( .a(FE_RN_396_0), .b(FE_OFN1707_n_4868), .o(TIMEBOOST_net_5291) );
na02f04 TIMEBOOST_cell_37026 ( .a(TIMEBOOST_net_10751), .b(g52523_sb), .o(n_13697) );
in01s01 g57909_u0 ( .a(FE_OFN1795_n_9904), .o(g57909_sb) );
na02s01 TIMEBOOST_cell_9066 ( .a(pci_target_unit_fifos_pcir_data_in_188), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__Q), .o(TIMEBOOST_net_1100) );
na02s02 TIMEBOOST_cell_45050 ( .a(TIMEBOOST_net_14763), .b(FE_OFN719_n_8060), .o(TIMEBOOST_net_11256) );
na02s01 TIMEBOOST_cell_9067 ( .a(TIMEBOOST_net_1100), .b(FE_OFN945_n_2248), .o(TIMEBOOST_net_140) );
in01s01 g57910_u0 ( .a(FE_OFN576_n_9902), .o(g57910_sb) );
na02s02 TIMEBOOST_cell_45130 ( .a(TIMEBOOST_net_14803), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_11433) );
na03s02 TIMEBOOST_cell_41969 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__Q), .b(n_4342), .c(FE_OFN1293_n_4098), .o(TIMEBOOST_net_13223) );
na02f02 TIMEBOOST_cell_38938 ( .a(TIMEBOOST_net_11707), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10712) );
in01s01 g57911_u0 ( .a(FE_OFN527_n_9899), .o(g57911_sb) );
na02s02 TIMEBOOST_cell_38668 ( .a(TIMEBOOST_net_11572), .b(g62491_sb), .o(n_6603) );
in01s01 TIMEBOOST_cell_45959 ( .a(wbm_dat_i_8_), .o(TIMEBOOST_net_15266) );
na02f02 TIMEBOOST_cell_38854 ( .a(TIMEBOOST_net_11665), .b(g58461_sb), .o(n_9393) );
in01s01 g57912_u0 ( .a(FE_OFN576_n_9902), .o(g57912_sb) );
na02s01 g57912_u1 ( .a(FE_OFN252_n_9868), .b(g57912_sb), .o(g57912_da) );
na02s01 g57912_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__8__Q), .b(FE_OFN576_n_9902), .o(g57912_db) );
na02s01 g57912_u3 ( .a(g57912_da), .b(g57912_db), .o(n_9898) );
in01s01 g57913_u0 ( .a(FE_OFN1794_n_9904), .o(g57913_sb) );
na02s01 TIMEBOOST_cell_17470 ( .a(pci_target_unit_fifos_pciw_addr_data_in_150), .b(g64127_sb), .o(TIMEBOOST_net_3992) );
na02s01 g57913_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q), .b(FE_OFN1794_n_9904), .o(g57913_db) );
na02s02 TIMEBOOST_cell_45051 ( .a(n_1663), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__Q), .o(TIMEBOOST_net_14764) );
in01s01 g57914_u0 ( .a(FE_OFN562_n_9895), .o(g57914_sb) );
in01s01 TIMEBOOST_cell_45937 ( .a(wbm_dat_i_27_), .o(TIMEBOOST_net_15244) );
na02s01 g57914_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__Q), .b(FE_OFN562_n_9895), .o(g57914_db) );
na02m02 TIMEBOOST_cell_44637 ( .a(n_9232), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__Q), .o(TIMEBOOST_net_14557) );
in01s01 g57915_u0 ( .a(FE_OFN563_n_9895), .o(g57915_sb) );
na03s01 TIMEBOOST_cell_1017 ( .a(n_3928), .b(g63027_sb), .c(g63027_db), .o(n_5192) );
na02s01 TIMEBOOST_cell_39522 ( .a(TIMEBOOST_net_11999), .b(g61702_sb), .o(n_8423) );
na02s02 TIMEBOOST_cell_39684 ( .a(TIMEBOOST_net_12080), .b(g62959_sb), .o(n_5964) );
in01s01 g57916_u0 ( .a(FE_OFN561_n_9895), .o(g57916_sb) );
na02s01 TIMEBOOST_cell_44818 ( .a(TIMEBOOST_net_14647), .b(g64977_db), .o(n_3650) );
na02s01 TIMEBOOST_cell_36527 ( .a(pci_target_unit_fifos_pcir_data_in_173), .b(g65705_sb), .o(TIMEBOOST_net_10502) );
na03s02 TIMEBOOST_cell_1020 ( .a(n_3926), .b(g63031_sb), .c(g63031_db), .o(n_5185) );
in01s01 g57917_u0 ( .a(FE_OFN560_n_9895), .o(g57917_sb) );
na02s01 g57917_u1 ( .a(FE_OFN209_n_9126), .b(g57917_sb), .o(g57917_da) );
na02s01 g57917_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__Q), .b(FE_OFN560_n_9895), .o(g57917_db) );
na02s01 g57917_u3 ( .a(g57917_da), .b(g57917_db), .o(n_9135) );
in01s01 g57918_u0 ( .a(FE_OFN562_n_9895), .o(g57918_sb) );
na02s01 g57918_u1 ( .a(FE_OFN211_n_9858), .b(g57918_sb), .o(g57918_da) );
na02s01 g57918_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__Q), .b(FE_OFN563_n_9895), .o(g57918_db) );
na02s01 g57918_u3 ( .a(g57918_da), .b(g57918_db), .o(n_9892) );
in01s01 g57919_u0 ( .a(FE_OFN564_n_9895), .o(g57919_sb) );
na02s01 TIMEBOOST_cell_17474 ( .a(pci_target_unit_fifos_pciw_cbe_in_152), .b(g64110_sb), .o(TIMEBOOST_net_3994) );
na02s01 g57919_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__Q), .b(FE_OFN564_n_9895), .o(g57919_db) );
na02f02 TIMEBOOST_cell_44162 ( .a(TIMEBOOST_net_14319), .b(FE_OFN1415_n_8567), .o(TIMEBOOST_net_13390) );
in01s01 g57920_u0 ( .a(FE_OFN564_n_9895), .o(g57920_sb) );
na02s01 TIMEBOOST_cell_17476 ( .a(pci_target_unit_fifos_pciw_addr_data_in_145), .b(g64133_sb), .o(TIMEBOOST_net_3995) );
na02s01 g57920_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__Q), .b(FE_OFN564_n_9895), .o(g57920_db) );
na02f02 TIMEBOOST_cell_44404 ( .a(TIMEBOOST_net_14440), .b(FE_OFN1399_n_8567), .o(TIMEBOOST_net_12777) );
in01s01 g57921_u0 ( .a(FE_OFN562_n_9895), .o(g57921_sb) );
na02s01 g57921_u1 ( .a(FE_OFN217_n_9889), .b(g57921_sb), .o(g57921_da) );
na02s01 g57921_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q), .b(FE_OFN563_n_9895), .o(g57921_db) );
na02s01 g57921_u3 ( .a(g57921_da), .b(g57921_db), .o(n_9890) );
in01s01 g57922_u0 ( .a(FE_OFN561_n_9895), .o(g57922_sb) );
na02m02 TIMEBOOST_cell_43929 ( .a(n_9682), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__Q), .o(TIMEBOOST_net_14203) );
na02s01 g57922_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__Q), .b(FE_OFN561_n_9895), .o(g57922_db) );
na02s01 TIMEBOOST_cell_16190 ( .a(pci_target_unit_fifos_pciw_addr_data_in_144), .b(g64087_sb), .o(TIMEBOOST_net_3352) );
in01s01 g57923_u0 ( .a(FE_OFN563_n_9895), .o(g57923_sb) );
na02s01 TIMEBOOST_cell_44791 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__Q), .b(FE_OFN517_n_9697), .o(TIMEBOOST_net_14634) );
na03s02 TIMEBOOST_cell_38189 ( .a(g64309_da), .b(g64309_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__Q), .o(TIMEBOOST_net_11333) );
na02s01 TIMEBOOST_cell_37853 ( .a(FE_OFN264_n_9849), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__Q), .o(TIMEBOOST_net_11165) );
in01s01 g57924_u0 ( .a(FE_OFN562_n_9895), .o(g57924_sb) );
na02s02 TIMEBOOST_cell_39686 ( .a(TIMEBOOST_net_12081), .b(g62643_sb), .o(n_7371) );
na02f02 TIMEBOOST_cell_38788 ( .a(TIMEBOOST_net_11632), .b(g57331_db), .o(n_11419) );
na02s01 TIMEBOOST_cell_39320 ( .a(TIMEBOOST_net_11898), .b(g65874_db), .o(n_1869) );
in01s01 g57925_u0 ( .a(FE_OFN562_n_9895), .o(g57925_sb) );
na02s02 TIMEBOOST_cell_41773 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__Q), .b(g58349_sb), .o(TIMEBOOST_net_13125) );
na02s02 TIMEBOOST_cell_39688 ( .a(TIMEBOOST_net_12082), .b(g62693_sb), .o(n_6162) );
na03s02 TIMEBOOST_cell_37609 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__Q), .b(FE_OFN2256_n_8060), .c(n_1585), .o(TIMEBOOST_net_11043) );
in01s01 g57926_u0 ( .a(FE_OFN563_n_9895), .o(g57926_sb) );
na02s02 TIMEBOOST_cell_17478 ( .a(pci_target_unit_fifos_pciw_addr_data_in_151), .b(g64107_sb), .o(TIMEBOOST_net_3996) );
na02s01 g57926_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__Q), .b(FE_OFN563_n_9895), .o(g57926_db) );
na02s02 TIMEBOOST_cell_38687 ( .a(n_2093), .b(wishbone_slave_unit_pci_initiator_sm_rdata_selector), .o(TIMEBOOST_net_11582) );
in01s01 g57927_u0 ( .a(FE_OFN562_n_9895), .o(g57927_sb) );
na02s01 TIMEBOOST_cell_16191 ( .a(TIMEBOOST_net_3352), .b(g64087_db), .o(n_4068) );
na02s01 g57927_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__Q), .b(FE_OFN562_n_9895), .o(g57927_db) );
na02s01 TIMEBOOST_cell_16192 ( .a(pci_target_unit_fifos_pciw_addr_data_in_140), .b(g64095_sb), .o(TIMEBOOST_net_3353) );
in01s01 g57928_u0 ( .a(FE_OFN563_n_9895), .o(g57928_sb) );
na02m02 TIMEBOOST_cell_31498 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in), .b(TIMEBOOST_net_1637), .o(TIMEBOOST_net_9660) );
na02s01 g57928_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__Q), .b(FE_OFN563_n_9895), .o(g57928_db) );
na02s01 TIMEBOOST_cell_45052 ( .a(TIMEBOOST_net_14764), .b(FE_OFN2212_n_8407), .o(TIMEBOOST_net_11241) );
in01s01 g57929_u0 ( .a(FE_OFN561_n_9895), .o(g57929_sb) );
na03s01 TIMEBOOST_cell_38131 ( .a(g64201_da), .b(g64201_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__Q), .o(TIMEBOOST_net_11304) );
na03m02 TIMEBOOST_cell_7356 ( .a(TIMEBOOST_net_878), .b(g59799_da), .c(g59239_da), .o(n_7714) );
na02s01 TIMEBOOST_cell_38457 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__Q), .b(g58340_sb), .o(TIMEBOOST_net_11467) );
in01s01 g57930_u0 ( .a(FE_OFN561_n_9895), .o(g57930_sb) );
na02s01 TIMEBOOST_cell_16193 ( .a(TIMEBOOST_net_3353), .b(g64095_db), .o(n_4060) );
na02s01 g57930_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__Q), .b(FE_OFN561_n_9895), .o(g57930_db) );
na02s01 TIMEBOOST_cell_16194 ( .a(pci_target_unit_fifos_pciw_addr_data_in_147), .b(g64128_sb), .o(TIMEBOOST_net_3354) );
in01s01 g57931_u0 ( .a(FE_OFN560_n_9895), .o(g57931_sb) );
na02s01 g57931_u1 ( .a(FE_OFN229_n_9120), .b(g57931_sb), .o(g57931_da) );
na02s01 g57931_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__Q), .b(FE_OFN560_n_9895), .o(g57931_db) );
na02s02 g57931_u3 ( .a(g57931_da), .b(g57931_db), .o(n_9132) );
in01s01 g57932_u0 ( .a(FE_OFN561_n_9895), .o(g57932_sb) );
na02s01 TIMEBOOST_cell_43495 ( .a(n_4429), .b(n_4430), .o(TIMEBOOST_net_13986) );
na02s01 g57932_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q), .b(FE_OFN561_n_9895), .o(g57932_db) );
na02s01 TIMEBOOST_cell_39422 ( .a(TIMEBOOST_net_11949), .b(g54184_sb), .o(TIMEBOOST_net_11228) );
in01s01 g57933_u0 ( .a(FE_OFN563_n_9895), .o(g57933_sb) );
na02s01 TIMEBOOST_cell_43496 ( .a(TIMEBOOST_net_13986), .b(FE_OFN1235_n_6391), .o(TIMEBOOST_net_12144) );
na02s01 g57933_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__Q), .b(FE_OFN563_n_9895), .o(g57933_db) );
na02m02 TIMEBOOST_cell_38856 ( .a(TIMEBOOST_net_11666), .b(g58839_sb), .o(n_8675) );
in01s01 g57934_u0 ( .a(FE_OFN564_n_9895), .o(g57934_sb) );
na02f02 TIMEBOOST_cell_37965 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_403), .b(g54138_sb), .o(TIMEBOOST_net_11221) );
na02s01 g57934_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__Q), .b(FE_OFN564_n_9895), .o(g57934_db) );
na02s01 TIMEBOOST_cell_18929 ( .a(TIMEBOOST_net_4721), .b(g63551_sb), .o(n_4926) );
in01s01 g57935_u0 ( .a(FE_OFN563_n_9895), .o(g57935_sb) );
na02s01 TIMEBOOST_cell_17484 ( .a(pci_target_unit_fifos_pciw_addr_data_in_124), .b(g64098_sb), .o(TIMEBOOST_net_3999) );
na02s01 g57935_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__Q), .b(FE_OFN563_n_9895), .o(g57935_db) );
na02m02 TIMEBOOST_cell_44405 ( .a(n_9684), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__Q), .o(TIMEBOOST_net_14441) );
in01s01 g57936_u0 ( .a(FE_OFN562_n_9895), .o(g57936_sb) );
na02f02 TIMEBOOST_cell_43930 ( .a(TIMEBOOST_net_14203), .b(FE_OFN1376_n_8567), .o(TIMEBOOST_net_12879) );
na02s01 g57936_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__Q), .b(FE_OFN562_n_9895), .o(g57936_db) );
na02s01 TIMEBOOST_cell_16196 ( .a(pci_target_unit_fifos_pciw_addr_data_in_130), .b(g64202_sb), .o(TIMEBOOST_net_3355) );
in01s01 g57937_u0 ( .a(FE_OFN562_n_9895), .o(g57937_sb) );
na02s01 TIMEBOOST_cell_17486 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(g63549_sb), .o(TIMEBOOST_net_4000) );
na02s01 g57937_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__Q), .b(FE_OFN562_n_9895), .o(g57937_db) );
na02s01 TIMEBOOST_cell_17487 ( .a(TIMEBOOST_net_4000), .b(g63549_db), .o(n_4608) );
in01s01 g57938_u0 ( .a(FE_OFN564_n_9895), .o(g57938_sb) );
na02s02 TIMEBOOST_cell_36778 ( .a(TIMEBOOST_net_10627), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_4675) );
na02s01 g57938_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__Q), .b(FE_OFN564_n_9895), .o(g57938_db) );
na03s02 TIMEBOOST_cell_36779 ( .a(g65431_da), .b(g65431_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__Q), .o(TIMEBOOST_net_10628) );
in01s01 g57939_u0 ( .a(FE_OFN560_n_9895), .o(g57939_sb) );
na02m02 TIMEBOOST_cell_10981 ( .a(TIMEBOOST_net_2057), .b(g58636_sb), .o(TIMEBOOST_net_608) );
na02f02 TIMEBOOST_cell_44692 ( .a(TIMEBOOST_net_14584), .b(TIMEBOOST_net_10083), .o(n_11849) );
na02s01 TIMEBOOST_cell_39323 ( .a(TIMEBOOST_net_3893), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__Q), .o(TIMEBOOST_net_11900) );
in01s01 g57940_u0 ( .a(FE_OFN562_n_9895), .o(g57940_sb) );
na02m02 TIMEBOOST_cell_43931 ( .a(n_9653), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__Q), .o(TIMEBOOST_net_14204) );
na02s01 g57940_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__Q), .b(FE_OFN562_n_9895), .o(g57940_db) );
na02s01 TIMEBOOST_cell_16198 ( .a(pci_target_unit_fifos_pciw_addr_data_in_151), .b(g64216_sb), .o(TIMEBOOST_net_3356) );
in01s01 g57941_u0 ( .a(FE_OFN564_n_9895), .o(g57941_sb) );
na02s01 TIMEBOOST_cell_16199 ( .a(TIMEBOOST_net_3356), .b(g64216_db), .o(n_3953) );
na02s01 g57941_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__Q), .b(FE_OFN564_n_9895), .o(g57941_db) );
na02m02 TIMEBOOST_cell_43697 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__Q), .b(n_9493), .o(TIMEBOOST_net_14087) );
in01s01 g57942_u0 ( .a(FE_OFN559_n_9895), .o(g57942_sb) );
na02s01 TIMEBOOST_cell_36643 ( .a(parchk_pci_ad_reg_in_1216), .b(g65813_sb), .o(TIMEBOOST_net_10560) );
na02s01 g57942_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q), .b(FE_OFN559_n_9895), .o(g57942_db) );
na02s01 TIMEBOOST_cell_44819 ( .a(pci_target_unit_fifos_pcir_data_in_172), .b(g65725_sb), .o(TIMEBOOST_net_14648) );
na02f02 TIMEBOOST_cell_42514 ( .a(TIMEBOOST_net_13495), .b(g57221_sb), .o(n_11534) );
na02s01 g57943_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__Q), .b(FE_OFN560_n_9895), .o(g57943_db) );
na02s01 TIMEBOOST_cell_45649 ( .a(g58207_sb), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_15063) );
in01s01 g57944_u0 ( .a(FE_OFN564_n_9895), .o(g57944_sb) );
na02s01 TIMEBOOST_cell_17490 ( .a(n_4473), .b(FE_OFN643_n_4677), .o(TIMEBOOST_net_4002) );
na02s01 g57944_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__8__Q), .b(FE_OFN564_n_9895), .o(g57944_db) );
na02s01 TIMEBOOST_cell_17491 ( .a(TIMEBOOST_net_4002), .b(g65280_da), .o(n_4287) );
in01s01 g57945_u0 ( .a(FE_OFN561_n_9895), .o(g57945_sb) );
na02s01 TIMEBOOST_cell_17492 ( .a(pci_target_unit_fifos_pciw_addr_data_in_139), .b(g64223_sb), .o(TIMEBOOST_net_4003) );
na02s01 g57945_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__Q), .b(FE_OFN561_n_9895), .o(g57945_db) );
na03s01 TIMEBOOST_cell_39459 ( .a(TIMEBOOST_net_3957), .b(g64252_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__Q), .o(TIMEBOOST_net_11968) );
in01s01 g57946_u0 ( .a(FE_OFN554_n_9864), .o(g57946_sb) );
na02s01 TIMEBOOST_cell_17562 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__Q), .b(g64314_sb), .o(TIMEBOOST_net_4038) );
na02s01 g57946_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__Q), .b(FE_OFN554_n_9864), .o(g57946_db) );
na03s02 TIMEBOOST_cell_38357 ( .a(n_3938), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q), .c(FE_OFN2104_g64577_p), .o(TIMEBOOST_net_11417) );
in01s01 g57947_u0 ( .a(FE_OFN555_n_9864), .o(g57947_sb) );
na02s02 TIMEBOOST_cell_38602 ( .a(TIMEBOOST_net_11539), .b(g62334_sb), .o(n_6932) );
na02s01 g57947_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__Q), .b(FE_OFN555_n_9864), .o(g57947_db) );
na02s01 TIMEBOOST_cell_18483 ( .a(TIMEBOOST_net_4498), .b(g62737_sb), .o(n_5505) );
in01s01 g57948_u0 ( .a(FE_OFN553_n_9864), .o(g57948_sb) );
na02f02 TIMEBOOST_cell_38940 ( .a(TIMEBOOST_net_11708), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10723) );
na02s02 TIMEBOOST_cell_40662 ( .a(TIMEBOOST_net_12569), .b(g62364_sb), .o(n_6872) );
na02s01 TIMEBOOST_cell_44876 ( .a(TIMEBOOST_net_14676), .b(g65812_db), .o(n_1902) );
in01s01 g57949_u0 ( .a(FE_OFN551_n_9864), .o(g57949_sb) );
na02s01 g57949_u1 ( .a(FE_OFN209_n_9126), .b(g57949_sb), .o(g57949_da) );
na02s01 g57949_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__Q), .b(FE_OFN551_n_9864), .o(g57949_db) );
na02s01 g57949_u3 ( .a(g57949_da), .b(g57949_db), .o(n_9127) );
na02s01 g57950_u1 ( .a(FE_OFN211_n_9858), .b(g57965_sb), .o(g57950_da) );
na02s01 g57950_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__Q), .b(FE_OFN555_n_9864), .o(g57950_db) );
na02s01 g57950_u3 ( .a(g57950_da), .b(g57950_db), .o(n_9859) );
in01s01 g57951_u0 ( .a(FE_OFN556_n_9864), .o(g57951_sb) );
na02f02 TIMEBOOST_cell_44406 ( .a(TIMEBOOST_net_14441), .b(FE_OFN1385_n_8567), .o(TIMEBOOST_net_12776) );
na02s01 g57951_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__Q), .b(FE_OFN556_n_9864), .o(g57951_db) );
na02s02 TIMEBOOST_cell_39690 ( .a(TIMEBOOST_net_12083), .b(g63184_sb), .o(n_5784) );
in01s01 g57952_u0 ( .a(FE_OFN556_n_9864), .o(g57952_sb) );
na02s01 TIMEBOOST_cell_17280 ( .a(n_3780), .b(FE_OFN652_n_4508), .o(TIMEBOOST_net_3897) );
na02s01 g57952_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__Q), .b(FE_OFN556_n_9864), .o(g57952_db) );
na02s01 TIMEBOOST_cell_17281 ( .a(TIMEBOOST_net_3897), .b(g65428_da), .o(n_3507) );
in01s01 g57953_u0 ( .a(FE_OFN554_n_9864), .o(g57953_sb) );
na02s01 g57953_u1 ( .a(FE_OFN217_n_9889), .b(g57953_sb), .o(g57953_da) );
na02s01 g57953_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__Q), .b(FE_OFN554_n_9864), .o(g57953_db) );
na02s01 g57953_u3 ( .a(g57953_da), .b(g57953_db), .o(n_9855) );
in01s01 g57954_u0 ( .a(FE_OFN553_n_9864), .o(g57954_sb) );
na02s01 g57954_u1 ( .a(FE_OFN219_n_9853), .b(g57954_sb), .o(g57954_da) );
na02s01 g57954_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__Q), .b(FE_OFN553_n_9864), .o(g57954_db) );
na02s01 g57954_u3 ( .a(g57954_da), .b(g57954_db), .o(n_9854) );
na02s01 TIMEBOOST_cell_38036 ( .a(TIMEBOOST_net_11256), .b(g61860_sb), .o(n_8118) );
no02f04 TIMEBOOST_cell_19039 ( .a(TIMEBOOST_net_4776), .b(FE_RN_711_0), .o(TIMEBOOST_net_933) );
in01s01 g57956_u0 ( .a(FE_OFN554_n_9864), .o(g57956_sb) );
na02s01 TIMEBOOST_cell_38186 ( .a(TIMEBOOST_net_11331), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_4544) );
na02s01 TIMEBOOST_cell_40454 ( .a(TIMEBOOST_net_12465), .b(g62136_sb), .o(n_5557) );
na02s01 TIMEBOOST_cell_44820 ( .a(TIMEBOOST_net_14648), .b(g65725_db), .o(TIMEBOOST_net_268) );
in01s01 g57957_u0 ( .a(FE_OFN554_n_9864), .o(g57957_sb) );
na03s01 TIMEBOOST_cell_1039 ( .a(n_3897), .b(g63060_sb), .c(g63060_db), .o(n_5130) );
na02s01 TIMEBOOST_cell_40455 ( .a(parchk_pci_ad_out_in_1182), .b(configuration_wb_err_data_585), .o(TIMEBOOST_net_12466) );
na03s02 TIMEBOOST_cell_37893 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__Q), .b(FE_OFN539_n_9690), .c(FE_OFN264_n_9849), .o(TIMEBOOST_net_11185) );
in01s01 g57958_u0 ( .a(FE_OFN555_n_9864), .o(g57958_sb) );
na02m04 TIMEBOOST_cell_9604 ( .a(FE_RN_72_0), .b(FE_OCPN1854_n_2071), .o(TIMEBOOST_net_1369) );
na02s01 g57958_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__Q), .b(FE_OFN555_n_9864), .o(g57958_db) );
na02m04 TIMEBOOST_cell_9605 ( .a(FE_RN_73_0), .b(TIMEBOOST_net_1369), .o(TIMEBOOST_net_907) );
in01s01 g57959_u0 ( .a(FE_OFN554_n_9864), .o(g57959_sb) );
na02s01 g57959_u1 ( .a(FE_OFN223_n_9844), .b(g57959_sb), .o(g57959_da) );
na02s01 g57959_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__Q), .b(FE_OFN554_n_9864), .o(g57959_db) );
na02s01 g57959_u3 ( .a(g57959_da), .b(g57959_db), .o(n_9845) );
na02s01 g57960_u1 ( .a(FE_OFN225_n_9122), .b(g57958_sb), .o(g57960_da) );
na02s01 g57960_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__Q), .b(FE_OFN555_n_9864), .o(g57960_db) );
na02s01 g57960_u3 ( .a(g57960_da), .b(g57960_db), .o(n_9123) );
in01s01 g57961_u0 ( .a(FE_OFN553_n_9864), .o(g57961_sb) );
na02s01 TIMEBOOST_cell_39232 ( .a(TIMEBOOST_net_11854), .b(g58190_sb), .o(TIMEBOOST_net_10989) );
na02s02 TIMEBOOST_cell_40456 ( .a(TIMEBOOST_net_12466), .b(g62085_sb), .o(TIMEBOOST_net_11371) );
na02m02 TIMEBOOST_cell_32758 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__Q), .o(TIMEBOOST_net_10290) );
na02s01 g57962_u1 ( .a(FE_OFN227_n_9841), .b(g57961_sb), .o(g57962_da) );
na02s01 g57962_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__Q), .b(FE_OFN553_n_9864), .o(g57962_db) );
na02s02 g57962_u3 ( .a(g57962_da), .b(g57962_db), .o(n_9842) );
na02s01 g57963_u1 ( .a(FE_OFN229_n_9120), .b(g57949_sb), .o(g57963_da) );
na02s01 g57963_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__Q), .b(FE_OFN551_n_9864), .o(g57963_db) );
na02s02 g57963_u3 ( .a(g57963_da), .b(g57963_db), .o(n_9121) );
in01s01 g57964_u0 ( .a(FE_OFN555_n_9864), .o(g57964_sb) );
na02s01 g57964_u1 ( .a(FE_OFN231_n_9839), .b(g57964_sb), .o(g57964_da) );
na02s01 g57964_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__Q), .b(FE_OFN555_n_9864), .o(g57964_db) );
na02s02 g57964_u3 ( .a(g57964_da), .b(g57964_db), .o(n_9840) );
in01s01 g57965_u0 ( .a(FE_OFN555_n_9864), .o(g57965_sb) );
na02s01 g57965_u1 ( .a(FE_OFN233_n_9876), .b(g57965_sb), .o(g57965_da) );
na02s01 g57965_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__Q), .b(FE_OFN555_n_9864), .o(g57965_db) );
na02s01 g57965_u3 ( .a(g57965_da), .b(g57965_db), .o(n_9838) );
na02s02 TIMEBOOST_cell_38038 ( .a(TIMEBOOST_net_11257), .b(g61778_sb), .o(n_8251) );
na02m02 TIMEBOOST_cell_44303 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__Q), .b(n_9499), .o(TIMEBOOST_net_14390) );
na02s01 TIMEBOOST_cell_39234 ( .a(TIMEBOOST_net_11855), .b(g65682_db), .o(n_1955) );
na02s01 g57967_u1 ( .a(FE_OFN235_n_9834), .b(g57947_sb), .o(g57967_da) );
na02s01 g57967_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__Q), .b(FE_OFN555_n_9864), .o(g57967_db) );
na02s02 g57967_u3 ( .a(g57967_da), .b(g57967_db), .o(n_9835) );
in01s01 g57968_u0 ( .a(FE_OFN552_n_9864), .o(g57968_sb) );
na02s01 g57968_u1 ( .a(FE_OFN237_n_9118), .b(g57968_sb), .o(g57968_da) );
na02s01 g57968_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__Q), .b(FE_OFN552_n_9864), .o(g57968_db) );
na02s01 g57968_u3 ( .a(g57968_da), .b(g57968_db), .o(n_9119) );
in01s01 g57969_u0 ( .a(FE_OFN554_n_9864), .o(g57969_sb) );
na02s02 TIMEBOOST_cell_17588 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_11__Q), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_4051) );
na02s01 g57969_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__Q), .b(FE_OFN554_n_9864), .o(g57969_db) );
na02s02 TIMEBOOST_cell_17589 ( .a(TIMEBOOST_net_4051), .b(n_13221), .o(TIMEBOOST_net_522) );
in01s01 g57970_u0 ( .a(FE_OFN556_n_9864), .o(g57970_sb) );
na02s01 g57970_u1 ( .a(FE_OFN241_n_9830), .b(g57970_sb), .o(g57970_da) );
na02s01 g57970_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__Q), .b(FE_OFN556_n_9864), .o(g57970_db) );
na02s01 g57970_u3 ( .a(g57970_da), .b(g57970_db), .o(n_9831) );
in01s01 g57971_u0 ( .a(FE_OFN551_n_9864), .o(g57971_sb) );
na02s01 TIMEBOOST_cell_39236 ( .a(TIMEBOOST_net_11856), .b(g65728_db), .o(n_1937) );
na02s01 TIMEBOOST_cell_40458 ( .a(TIMEBOOST_net_12467), .b(g62118_sb), .o(n_5578) );
in01s01 g57972_u0 ( .a(FE_OFN554_n_9864), .o(g57972_sb) );
na02s01 g57972_u1 ( .a(FE_OFN243_n_9116), .b(g57972_sb), .o(g57972_da) );
na02s01 g57972_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__Q), .b(FE_OFN554_n_9864), .o(g57972_db) );
na02s01 g57972_u3 ( .a(g57972_da), .b(g57972_db), .o(n_9117) );
in01s01 g57973_u0 ( .a(FE_OFN556_n_9864), .o(g57973_sb) );
na02s01 TIMEBOOST_cell_44858 ( .a(TIMEBOOST_net_14667), .b(g58317_sb), .o(TIMEBOOST_net_12445) );
na02s01 g57973_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__Q), .b(FE_OFN556_n_9864), .o(g57973_db) );
na02f02 TIMEBOOST_cell_44304 ( .a(TIMEBOOST_net_14390), .b(FE_OFN1394_n_8567), .o(TIMEBOOST_net_12952) );
na02s02 TIMEBOOST_cell_39692 ( .a(TIMEBOOST_net_12084), .b(g62437_sb), .o(n_6722) );
na02m02 TIMEBOOST_cell_17494 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_4__Q), .b(n_12595), .o(TIMEBOOST_net_4004) );
na02s01 TIMEBOOST_cell_16925 ( .a(TIMEBOOST_net_3719), .b(g65410_db), .o(n_3516) );
in01s01 g57975_u0 ( .a(FE_OFN554_n_9864), .o(g57975_sb) );
na02s01 g57975_u1 ( .a(FE_OFN252_n_9868), .b(g57975_sb), .o(g57975_da) );
na02s01 g57975_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__Q), .b(FE_OFN554_n_9864), .o(g57975_db) );
na02s01 g57975_u3 ( .a(g57975_da), .b(g57975_db), .o(n_9827) );
na02s01 TIMEBOOST_cell_45140 ( .a(TIMEBOOST_net_14808), .b(n_5546), .o(TIMEBOOST_net_13761) );
na02s01 g57976_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__Q), .b(FE_OFN553_n_9864), .o(g57976_db) );
na02s02 TIMEBOOST_cell_39694 ( .a(TIMEBOOST_net_12085), .b(g62354_sb), .o(n_6892) );
in01s01 g57977_u0 ( .a(FE_OFN532_n_9823), .o(g57977_sb) );
na02s01 TIMEBOOST_cell_17590 ( .a(wbu_addr_in_250), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_4052) );
na02s01 g57977_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__Q), .b(FE_OFN532_n_9823), .o(g57977_db) );
na02s01 TIMEBOOST_cell_39696 ( .a(TIMEBOOST_net_12086), .b(g62383_sb), .o(n_6835) );
in01s01 g57978_u0 ( .a(FE_OFN535_n_9823), .o(g57978_sb) );
na02s01 TIMEBOOST_cell_39238 ( .a(TIMEBOOST_net_11857), .b(g64931_db), .o(n_4388) );
na02s01 TIMEBOOST_cell_39524 ( .a(TIMEBOOST_net_12000), .b(g61709_sb), .o(n_8409) );
na02s02 TIMEBOOST_cell_39240 ( .a(TIMEBOOST_net_11858), .b(g65409_sb), .o(n_4231) );
in01s01 g57979_u0 ( .a(FE_OFN533_n_9823), .o(g57979_sb) );
na02s01 TIMEBOOST_cell_38040 ( .a(TIMEBOOST_net_11258), .b(g61996_db), .o(n_7903) );
na02m02 TIMEBOOST_cell_44607 ( .a(n_9125), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__Q), .o(TIMEBOOST_net_14542) );
na02s02 TIMEBOOST_cell_39242 ( .a(TIMEBOOST_net_11859), .b(g58314_db), .o(n_9498) );
in01s01 g57980_u0 ( .a(FE_OFN1789_n_9823), .o(g57980_sb) );
na02s01 TIMEBOOST_cell_16668 ( .a(pci_target_unit_fifos_pciw_addr_data_in_145), .b(g64168_sb), .o(TIMEBOOST_net_3591) );
na02s01 g57980_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__Q), .b(FE_OFN1789_n_9823), .o(g57980_db) );
na02s01 TIMEBOOST_cell_45089 ( .a(FE_OFN258_n_9862), .b(g57947_sb), .o(TIMEBOOST_net_14783) );
in01s01 g57981_u0 ( .a(FE_OFN535_n_9823), .o(g57981_sb) );
na02s01 TIMEBOOST_cell_9612 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__Q), .b(g58319_sb), .o(TIMEBOOST_net_1373) );
na02s01 g57981_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__Q), .b(FE_OFN535_n_9823), .o(g57981_db) );
na02s01 TIMEBOOST_cell_9613 ( .a(TIMEBOOST_net_1373), .b(g58319_db), .o(n_9493) );
in01s01 g57982_u0 ( .a(FE_OFN534_n_9823), .o(g57982_sb) );
na02s01 TIMEBOOST_cell_36502 ( .a(TIMEBOOST_net_10489), .b(g66415_sb), .o(n_2502) );
na02s01 g57982_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__Q), .b(FE_OFN534_n_9823), .o(g57982_db) );
na02s01 TIMEBOOST_cell_36503 ( .a(pci_target_unit_del_sync_addr_in_221), .b(g66408_db), .o(TIMEBOOST_net_10490) );
in01s01 g57983_u0 ( .a(FE_OFN534_n_9823), .o(g57983_sb) );
na02s01 TIMEBOOST_cell_44920 ( .a(TIMEBOOST_net_14698), .b(g65943_sb), .o(TIMEBOOST_net_335) );
na02s01 g57983_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__Q), .b(FE_OFN534_n_9823), .o(g57983_db) );
na02s01 TIMEBOOST_cell_39698 ( .a(TIMEBOOST_net_12087), .b(g62940_sb), .o(n_6001) );
in01s01 g57984_u0 ( .a(FE_OFN531_n_9823), .o(g57984_sb) );
na02s01 TIMEBOOST_cell_40525 ( .a(wishbone_slave_unit_pcim_sm_data_in_658), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__Q), .o(TIMEBOOST_net_12501) );
na02s01 g57984_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__Q), .b(FE_OFN531_n_9823), .o(g57984_db) );
na02s01 TIMEBOOST_cell_40460 ( .a(TIMEBOOST_net_12468), .b(g62126_sb), .o(n_5570) );
in01s01 g57985_u0 ( .a(FE_OFN535_n_9823), .o(g57985_sb) );
na02s01 TIMEBOOST_cell_39322 ( .a(TIMEBOOST_net_11899), .b(FE_OFN211_n_9858), .o(TIMEBOOST_net_3898) );
na02s01 TIMEBOOST_cell_39526 ( .a(TIMEBOOST_net_12001), .b(g61710_sb), .o(n_8406) );
na02s02 TIMEBOOST_cell_38042 ( .a(TIMEBOOST_net_11259), .b(FE_OFN1128_g64577_p), .o(TIMEBOOST_net_4721) );
in01s01 g57986_u0 ( .a(FE_OFN533_n_9823), .o(g57986_sb) );
na02s02 TIMEBOOST_cell_40462 ( .a(TIMEBOOST_net_12469), .b(g58288_db), .o(n_9032) );
na02s01 g57986_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__Q), .b(FE_OFN533_n_9823), .o(g57986_db) );
na02s01 TIMEBOOST_cell_16661 ( .a(TIMEBOOST_net_3587), .b(g64198_db), .o(n_3971) );
in01s01 g57987_u0 ( .a(FE_OFN531_n_9823), .o(g57987_sb) );
na02s01 TIMEBOOST_cell_39244 ( .a(TIMEBOOST_net_11860), .b(g58425_db), .o(n_9423) );
na02s01 TIMEBOOST_cell_36489 ( .a(n_2541), .b(g66400_db), .o(TIMEBOOST_net_10483) );
na02s02 TIMEBOOST_cell_39246 ( .a(TIMEBOOST_net_11861), .b(g58338_db), .o(n_9482) );
in01s01 g57988_u0 ( .a(FE_OFN532_n_9823), .o(g57988_sb) );
in01s01 TIMEBOOST_cell_45898 ( .a(TIMEBOOST_net_15204), .o(TIMEBOOST_net_15205) );
na02s01 TIMEBOOST_cell_39528 ( .a(TIMEBOOST_net_12002), .b(g61703_sb), .o(n_8421) );
na02s02 TIMEBOOST_cell_38188 ( .a(TIMEBOOST_net_11332), .b(FE_OFN1134_g64577_p), .o(TIMEBOOST_net_4548) );
in01s01 g57989_u0 ( .a(FE_OFN535_n_9823), .o(g57989_sb) );
in01s01 TIMEBOOST_cell_45960 ( .a(TIMEBOOST_net_15266), .o(TIMEBOOST_net_15267) );
na02s01 g57989_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__Q), .b(FE_OFN535_n_9823), .o(g57989_db) );
na02s02 TIMEBOOST_cell_39700 ( .a(TIMEBOOST_net_12088), .b(g62676_sb), .o(n_7368) );
in01s01 g57990_u0 ( .a(FE_OFN531_n_9823), .o(g57990_sb) );
na02s01 g57990_u1 ( .a(FE_OFN223_n_9844), .b(g57990_sb), .o(g57990_da) );
na02s01 g57990_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__Q), .b(FE_OFN531_n_9823), .o(g57990_db) );
na02s01 g57990_u3 ( .a(g57990_da), .b(g57990_db), .o(n_9805) );
in01s01 g57991_u0 ( .a(FE_OFN535_n_9823), .o(g57991_sb) );
na02s02 TIMEBOOST_cell_42836 ( .a(TIMEBOOST_net_13656), .b(g62031_sb), .o(TIMEBOOST_net_579) );
na02f02 TIMEBOOST_cell_39095 ( .a(FE_OCP_RBN1995_n_13971), .b(TIMEBOOST_net_10233), .o(TIMEBOOST_net_11786) );
na02s02 TIMEBOOST_cell_39702 ( .a(TIMEBOOST_net_12089), .b(g62631_sb), .o(n_6292) );
in01s01 g57992_u0 ( .a(FE_OFN533_n_9823), .o(g57992_sb) );
na02s02 TIMEBOOST_cell_38044 ( .a(TIMEBOOST_net_11260), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_4585) );
na02s01 TIMEBOOST_cell_36517 ( .a(g58210_sb), .b(g58210_db), .o(TIMEBOOST_net_10497) );
na02s02 TIMEBOOST_cell_38190 ( .a(TIMEBOOST_net_11333), .b(FE_OFN1134_g64577_p), .o(TIMEBOOST_net_4581) );
in01s01 g57993_u0 ( .a(FE_OFN533_n_9823), .o(g57993_sb) );
na02s01 TIMEBOOST_cell_32016 ( .a(configuration_pci_err_data_519), .b(wbm_dat_o_18_), .o(TIMEBOOST_net_9919) );
na02s01 g57993_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__Q), .b(FE_OFN533_n_9823), .o(g57993_db) );
na02s01 TIMEBOOST_cell_32014 ( .a(configuration_pci_err_data_517), .b(wbm_dat_o_16_), .o(TIMEBOOST_net_9918) );
in01s01 g57994_u0 ( .a(FE_OFN1789_n_9823), .o(g57994_sb) );
na02s02 TIMEBOOST_cell_39704 ( .a(TIMEBOOST_net_12090), .b(g62958_sb), .o(n_5966) );
na02s01 g57994_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__Q), .b(FE_OFN1789_n_9823), .o(g57994_db) );
na02s01 TIMEBOOST_cell_44921 ( .a(FE_OFN241_n_9830), .b(g58191_sb), .o(TIMEBOOST_net_14699) );
in01s01 g57995_u0 ( .a(FE_OFN533_n_9823), .o(g57995_sb) );
na03f02 TIMEBOOST_cell_36228 ( .a(n_16397), .b(TIMEBOOST_net_6571), .c(n_16395), .o(n_16398) );
na02s01 g57995_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__Q), .b(FE_OFN533_n_9823), .o(g57995_db) );
na03f02 TIMEBOOST_cell_36229 ( .a(FE_RN_110_0), .b(n_12809), .c(n_12964), .o(n_13144) );
in01s01 g57996_u0 ( .a(FE_OFN535_n_9823), .o(g57996_sb) );
na02s01 TIMEBOOST_cell_18967 ( .a(TIMEBOOST_net_4740), .b(g58339_db), .o(n_9481) );
na02s01 TIMEBOOST_cell_39512 ( .a(TIMEBOOST_net_11994), .b(TIMEBOOST_net_9838), .o(n_5062) );
na02s02 TIMEBOOST_cell_18931 ( .a(TIMEBOOST_net_4722), .b(g58296_sb), .o(n_9217) );
in01s01 g57997_u0 ( .a(FE_OFN535_n_9823), .o(g57997_sb) );
na02s01 g57997_u1 ( .a(FE_OFN235_n_9834), .b(g57997_sb), .o(g57997_da) );
na02s01 g57997_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__Q), .b(FE_OFN535_n_9823), .o(g57997_db) );
na02s02 g57997_u3 ( .a(g57997_da), .b(g57997_db), .o(n_9796) );
in01s01 TIMEBOOST_cell_45961 ( .a(wbm_dat_i_9_), .o(TIMEBOOST_net_15268) );
na02s01 g57998_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__Q), .b(FE_OFN1789_n_9823), .o(g57998_db) );
na02s01 TIMEBOOST_cell_39706 ( .a(TIMEBOOST_net_12091), .b(g62487_sb), .o(n_6613) );
in01s01 g57999_u0 ( .a(FE_OFN531_n_9823), .o(g57999_sb) );
na02s01 TIMEBOOST_cell_36504 ( .a(TIMEBOOST_net_10490), .b(g66403_sb), .o(n_2530) );
na02s01 g57999_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__Q), .b(FE_OFN531_n_9823), .o(g57999_db) );
no02f02 g57_u0 ( .a(n_15585), .b(n_15562), .o(n_15586) );
in01s01 g58000_u0 ( .a(FE_OFN534_n_9823), .o(g58000_sb) );
na02s01 g58000_u1 ( .a(FE_OFN241_n_9830), .b(g58000_sb), .o(g58000_da) );
na02s01 g58000_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__Q), .b(FE_OFN534_n_9823), .o(g58000_db) );
na02s01 g58000_u3 ( .a(g58000_da), .b(g58000_db), .o(n_9793) );
in01s01 g58001_u0 ( .a(FE_OFN533_n_9823), .o(g58001_sb) );
na02m02 TIMEBOOST_cell_32264 ( .a(wishbone_slave_unit_fifos_inGreyCount_reg_2__Q), .b(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q), .o(TIMEBOOST_net_10043) );
na02f02 TIMEBOOST_cell_39106 ( .a(TIMEBOOST_net_11791), .b(FE_OFN1599_n_13995), .o(n_14457) );
in01s01 g58002_u0 ( .a(FE_OFN531_n_9823), .o(g58002_sb) );
na02s01 g58002_u1 ( .a(FE_OFN243_n_9116), .b(g58002_sb), .o(g58002_da) );
na02s01 g58002_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__Q), .b(FE_OFN531_n_9823), .o(g58002_db) );
na02s02 g58002_u3 ( .a(g58002_da), .b(g58002_db), .o(n_9106) );
in01s01 g58003_u0 ( .a(FE_OFN534_n_9823), .o(g58003_sb) );
na02s01 TIMEBOOST_cell_41780 ( .a(TIMEBOOST_net_13128), .b(g58004_db), .o(n_9104) );
na02s01 g58003_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__Q), .b(FE_OFN534_n_9823), .o(g58003_db) );
na02s01 TIMEBOOST_cell_44821 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(g65694_sb), .o(TIMEBOOST_net_14649) );
in01s01 g58004_u0 ( .a(FE_OFN1789_n_9823), .o(g58004_sb) );
na02m02 TIMEBOOST_cell_42235 ( .a(n_9476), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__Q), .o(TIMEBOOST_net_13356) );
na02s01 g58004_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__Q), .b(FE_OFN1789_n_9823), .o(g58004_db) );
na02s01 TIMEBOOST_cell_17599 ( .a(TIMEBOOST_net_4056), .b(g58405_sb), .o(n_9002) );
in01s01 g58005_u0 ( .a(FE_OFN1789_n_9823), .o(g58005_sb) );
na02s02 TIMEBOOST_cell_43052 ( .a(TIMEBOOST_net_13764), .b(FE_OFN1242_n_4092), .o(TIMEBOOST_net_12078) );
na02s01 g58005_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__Q), .b(FE_OFN1789_n_9823), .o(g58005_db) );
na02s02 TIMEBOOST_cell_16737 ( .a(TIMEBOOST_net_3625), .b(g65298_sb), .o(n_3575) );
in01s01 g58006_u0 ( .a(FE_OFN533_n_9823), .o(g58006_sb) );
na02s02 TIMEBOOST_cell_44922 ( .a(TIMEBOOST_net_14699), .b(g58191_db), .o(n_9593) );
na02s01 g58006_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__Q), .b(FE_OFN533_n_9823), .o(g58006_db) );
na02s01 TIMEBOOST_cell_39708 ( .a(TIMEBOOST_net_12092), .b(g63006_sb), .o(n_5870) );
na02s01 g58007_u1 ( .a(FE_OFN250_n_9789), .b(g57971_sb), .o(g58007_da) );
na02s01 g58007_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__Q), .b(FE_OFN551_n_9864), .o(g58007_db) );
na02s02 g58007_u3 ( .a(g58007_da), .b(g58007_db), .o(n_9787) );
in01s01 g58008_u0 ( .a(FE_OFN529_n_9899), .o(g58008_sb) );
na02s01 g58008_u1 ( .a(FE_OFN207_n_9865), .b(g58008_sb), .o(g58008_da) );
na02s01 g58008_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__Q), .b(FE_OFN529_n_9899), .o(g58008_db) );
na02s01 g58008_u3 ( .a(g58008_da), .b(g58008_db), .o(n_9786) );
in01s01 g58009_u0 ( .a(FE_OFN527_n_9899), .o(g58009_sb) );
na02s01 TIMEBOOST_cell_18613 ( .a(TIMEBOOST_net_4563), .b(g63118_sb), .o(n_5021) );
in01s01 TIMEBOOST_cell_45962 ( .a(TIMEBOOST_net_15268), .o(TIMEBOOST_net_15269) );
na02s02 TIMEBOOST_cell_38192 ( .a(TIMEBOOST_net_11334), .b(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_4598) );
in01s01 g58010_u0 ( .a(FE_OFN527_n_9899), .o(g58010_sb) );
na02s02 TIMEBOOST_cell_19223 ( .a(TIMEBOOST_net_4868), .b(g60620_sb), .o(n_4834) );
na02s02 TIMEBOOST_cell_22297 ( .a(n_10274), .b(TIMEBOOST_net_6405), .o(n_11873) );
na02f02 TIMEBOOST_cell_41050 ( .a(TIMEBOOST_net_12763), .b(g57091_sb), .o(n_10489) );
in01s01 g58011_u0 ( .a(FE_OFN525_n_9899), .o(g58011_sb) );
na02s01 g58011_u1 ( .a(FE_OFN209_n_9126), .b(g58011_sb), .o(g58011_da) );
na02s01 g58011_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__Q), .b(FE_OFN525_n_9899), .o(g58011_db) );
na02s01 g58011_u3 ( .a(g58011_da), .b(g58011_db), .o(n_9103) );
in01s01 g58012_u0 ( .a(FE_OFN527_n_9899), .o(g58012_sb) );
na02s02 TIMEBOOST_cell_45183 ( .a(n_4301), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__Q), .o(TIMEBOOST_net_14830) );
na02s01 g58012_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__Q), .b(FE_OFN527_n_9899), .o(g58012_db) );
na02s02 TIMEBOOST_cell_39710 ( .a(TIMEBOOST_net_12093), .b(g62353_sb), .o(n_6895) );
in01s01 g58013_u0 ( .a(FE_OFN528_n_9899), .o(g58013_sb) );
na03s02 TIMEBOOST_cell_33967 ( .a(n_1597), .b(g61807_sb), .c(g61807_db), .o(n_8180) );
na02s01 g58013_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__Q), .b(FE_OFN528_n_9899), .o(g58013_db) );
na02s01 TIMEBOOST_cell_36239 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_1_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_2_), .o(TIMEBOOST_net_10358) );
in01s01 g58014_u0 ( .a(FE_OFN528_n_9899), .o(g58014_sb) );
na03s02 TIMEBOOST_cell_39371 ( .a(g65844_da), .b(g65844_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__Q), .o(TIMEBOOST_net_11924) );
na02s01 g58014_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__Q), .b(FE_OFN528_n_9899), .o(g58014_db) );
na02s01 TIMEBOOST_cell_39372 ( .a(TIMEBOOST_net_11924), .b(FE_OFN704_n_8069), .o(TIMEBOOST_net_4355) );
in01s01 g58015_u0 ( .a(FE_OFN529_n_9899), .o(g58015_sb) );
na02s01 g58015_u1 ( .a(FE_OFN217_n_9889), .b(g58015_sb), .o(g58015_da) );
na02s01 g58015_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__Q), .b(FE_OFN529_n_9899), .o(g58015_db) );
na02s01 g58015_u3 ( .a(g58015_da), .b(g58015_db), .o(n_9777) );
in01s01 g58016_u0 ( .a(FE_OFN526_n_9899), .o(g58016_sb) );
na02s01 g58016_u1 ( .a(FE_OFN219_n_9853), .b(g58016_sb), .o(g58016_da) );
na02s01 g58016_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__Q), .b(FE_OFN526_n_9899), .o(g58016_db) );
na02s01 g58016_u3 ( .a(g58016_da), .b(g58016_db), .o(n_9776) );
in01s01 g58017_u0 ( .a(FE_OFN527_n_9899), .o(g58017_sb) );
na02s02 TIMEBOOST_cell_38046 ( .a(TIMEBOOST_net_11261), .b(FE_OFN1140_g64577_p), .o(TIMEBOOST_net_4659) );
na02f02 TIMEBOOST_cell_32589 ( .a(TIMEBOOST_net_10205), .b(n_11988), .o(n_12704) );
na02s02 TIMEBOOST_cell_19225 ( .a(TIMEBOOST_net_4869), .b(g60623_sb), .o(n_4831) );
in01s01 g58018_u0 ( .a(FE_OFN526_n_9899), .o(g58018_sb) );
na02s02 TIMEBOOST_cell_19227 ( .a(TIMEBOOST_net_4870), .b(g60626_sb), .o(n_5712) );
na02f02 TIMEBOOST_cell_37807 ( .a(TIMEBOOST_net_9678), .b(g54334_sb), .o(TIMEBOOST_net_11142) );
na02s02 TIMEBOOST_cell_19229 ( .a(TIMEBOOST_net_4871), .b(g60629_sb), .o(n_5708) );
in01s01 g58019_u0 ( .a(FE_OFN529_n_9899), .o(g58019_sb) );
na02s02 TIMEBOOST_cell_19231 ( .a(TIMEBOOST_net_4872), .b(g60631_sb), .o(n_5705) );
na02f02 TIMEBOOST_cell_32561 ( .a(n_12313), .b(TIMEBOOST_net_10191), .o(TIMEBOOST_net_6565) );
na02s02 TIMEBOOST_cell_19233 ( .a(TIMEBOOST_net_4873), .b(g60635_sb), .o(n_5701) );
in01s01 g58020_u0 ( .a(FE_OFN527_n_9899), .o(g58020_sb) );
na02s01 g58020_u1 ( .a(FE_OFN221_n_9846), .b(g58020_sb), .o(g58020_da) );
na02s01 g58020_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q), .b(FE_OFN527_n_9899), .o(g58020_db) );
na02s01 g58020_u3 ( .a(g58020_da), .b(g58020_db), .o(n_9770) );
in01s01 g58021_u0 ( .a(FE_OFN525_n_9899), .o(g58021_sb) );
na02s01 g58021_u1 ( .a(FE_OFN223_n_9844), .b(g58021_sb), .o(g58021_da) );
na02s01 g58021_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__Q), .b(FE_OFN525_n_9899), .o(g58021_db) );
na02s01 g58021_u3 ( .a(g58021_da), .b(g58021_db), .o(n_9768) );
in01s01 g58022_u0 ( .a(FE_OFN527_n_9899), .o(g58022_sb) );
na02s01 TIMEBOOST_cell_44923 ( .a(FE_OFN239_n_9832), .b(g57969_sb), .o(TIMEBOOST_net_14700) );
na02s01 TIMEBOOST_cell_39231 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__Q), .b(FE_OFN585_n_9692), .o(TIMEBOOST_net_11854) );
na02s02 TIMEBOOST_cell_39712 ( .a(TIMEBOOST_net_12094), .b(g62410_sb), .o(n_6778) );
in01s01 g58023_u0 ( .a(FE_OFN527_n_9899), .o(g58023_sb) );
na02s01 g58023_u1 ( .a(FE_OFN227_n_9841), .b(g58023_sb), .o(g58023_da) );
na02s01 g58023_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__Q), .b(FE_OFN527_n_9899), .o(g58023_db) );
na02s02 g58023_u3 ( .a(g58023_da), .b(g58023_db), .o(n_9767) );
in01s01 g58024_u0 ( .a(FE_OFN525_n_9899), .o(g58024_sb) );
na02s01 g58024_u1 ( .a(FE_OFN229_n_9120), .b(g58024_sb), .o(g58024_da) );
na02s01 g58024_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__Q), .b(FE_OFN525_n_9899), .o(g58024_db) );
na02s02 g58024_u3 ( .a(g58024_da), .b(g58024_db), .o(n_9100) );
in01s01 g58025_u0 ( .a(FE_OFN527_n_9899), .o(g58025_sb) );
na02s01 TIMEBOOST_cell_9634 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__Q), .b(g58388_sb), .o(TIMEBOOST_net_1384) );
na02s01 g58025_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__Q), .b(FE_OFN527_n_9899), .o(g58025_db) );
na02s01 TIMEBOOST_cell_9635 ( .a(TIMEBOOST_net_1384), .b(g58388_db), .o(n_9443) );
in01s01 g58026_u0 ( .a(FE_OFN527_n_9899), .o(g58026_sb) );
na03s02 TIMEBOOST_cell_39373 ( .a(g65872_da), .b(g65872_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__Q), .o(TIMEBOOST_net_11925) );
na02s01 g58026_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__Q), .b(FE_OFN527_n_9899), .o(g58026_db) );
na02f02 TIMEBOOST_cell_39108 ( .a(TIMEBOOST_net_11792), .b(FE_OFN1599_n_13995), .o(n_14469) );
in01s01 g58027_u0 ( .a(FE_OFN528_n_9899), .o(g58027_sb) );
na03s02 TIMEBOOST_cell_38095 ( .a(TIMEBOOST_net_3472), .b(g64335_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__Q), .o(TIMEBOOST_net_11286) );
na02f02 TIMEBOOST_cell_38942 ( .a(TIMEBOOST_net_11709), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10715) );
na03s02 TIMEBOOST_cell_38093 ( .a(TIMEBOOST_net_4253), .b(g64115_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__Q), .o(TIMEBOOST_net_11285) );
in01s01 g58028_u0 ( .a(FE_OFN527_n_9899), .o(g58028_sb) );
na02s01 TIMEBOOST_cell_44924 ( .a(TIMEBOOST_net_14700), .b(g57969_db), .o(n_9833) );
na02s01 TIMEBOOST_cell_36506 ( .a(TIMEBOOST_net_10491), .b(g66402_sb), .o(n_2539) );
na02s02 TIMEBOOST_cell_39714 ( .a(TIMEBOOST_net_12095), .b(g62422_sb), .o(n_6752) );
in01s01 g58029_u0 ( .a(FE_OFN525_n_9899), .o(g58029_sb) );
na02s01 g58029_u1 ( .a(FE_OFN237_n_9118), .b(g58029_sb), .o(g58029_da) );
na02s01 g58029_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__Q), .b(FE_OFN525_n_9899), .o(g58029_db) );
na02s01 g58029_u3 ( .a(g58029_da), .b(g58029_db), .o(n_9099) );
in01s01 g58030_u0 ( .a(FE_OFN526_n_9899), .o(g58030_sb) );
na02s01 g58030_u1 ( .a(FE_OFN239_n_9832), .b(g58030_sb), .o(g58030_da) );
na02s01 g58030_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__Q), .b(FE_OFN526_n_9899), .o(g58030_db) );
na02s01 g58030_u3 ( .a(g58030_da), .b(g58030_db), .o(n_9757) );
in01s01 g58031_u0 ( .a(FE_OFN528_n_9899), .o(g58031_sb) );
na02s01 g58031_u1 ( .a(FE_OFN241_n_9830), .b(g58031_sb), .o(g58031_da) );
na02s01 g58031_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__Q), .b(FE_OFN528_n_9899), .o(g58031_db) );
na02s01 g58031_u3 ( .a(g58031_da), .b(g58031_db), .o(n_9756) );
in01s01 g58032_u0 ( .a(FE_OFN526_n_9899), .o(g58032_sb) );
na02s02 TIMEBOOST_cell_19239 ( .a(TIMEBOOST_net_4876), .b(g60648_sb), .o(n_5678) );
na02f02 TIMEBOOST_cell_32569 ( .a(FE_OCPN1825_n_12030), .b(TIMEBOOST_net_10195), .o(TIMEBOOST_net_6557) );
na02s02 TIMEBOOST_cell_19241 ( .a(TIMEBOOST_net_4877), .b(g60650_sb), .o(n_5675) );
in01s01 g58033_u0 ( .a(FE_OFN526_n_9899), .o(g58033_sb) );
na02s01 g58033_u1 ( .a(FE_OFN243_n_9116), .b(g58033_sb), .o(g58033_da) );
na02s01 g58033_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__Q), .b(FE_OFN526_n_9899), .o(g58033_db) );
na02s01 g58033_u3 ( .a(g58033_da), .b(g58033_db), .o(n_9098) );
in01s01 g58034_u0 ( .a(FE_OFN528_n_9899), .o(g58034_sb) );
na02m02 TIMEBOOST_cell_44305 ( .a(n_9480), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__Q), .o(TIMEBOOST_net_14391) );
na02s01 g58034_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__Q), .b(FE_OFN528_n_9899), .o(g58034_db) );
na02s02 TIMEBOOST_cell_40464 ( .a(TIMEBOOST_net_12470), .b(g61843_sb), .o(n_7212) );
in01s01 g58035_u0 ( .a(FE_OFN525_n_9899), .o(g58035_sb) );
na02m02 TIMEBOOST_cell_38969 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_7__Q), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__Q), .o(TIMEBOOST_net_11723) );
na02s01 g58035_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__Q), .b(FE_OFN526_n_9899), .o(g58035_db) );
na02f02 TIMEBOOST_cell_38944 ( .a(TIMEBOOST_net_11710), .b(FE_OFN2157_n_16439), .o(TIMEBOOST_net_10736) );
in01s01 g58036_u0 ( .a(FE_OFN525_n_9899), .o(g58036_sb) );
na02s01 g58036_u1 ( .a(FE_OFN250_n_9789), .b(g58036_sb), .o(g58036_da) );
na02s01 g58036_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__Q), .b(FE_OFN525_n_9899), .o(g58036_db) );
na02s02 g58036_u3 ( .a(g58036_da), .b(g58036_db), .o(n_9753) );
in01s01 g58037_u0 ( .a(FE_OFN528_n_9899), .o(g58037_sb) );
na02s01 g58037_u1 ( .a(FE_OFN252_n_9868), .b(g58037_sb), .o(g58037_da) );
na02s01 g58037_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__Q), .b(FE_OFN528_n_9899), .o(g58037_db) );
na02s01 g58037_u3 ( .a(g58037_da), .b(g58037_db), .o(n_9752) );
na02s01 TIMEBOOST_cell_17606 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_3__Q), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_4060) );
na02s01 g58038_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__Q), .b(FE_OFN527_n_9899), .o(g58038_db) );
na02m01 TIMEBOOST_cell_17607 ( .a(TIMEBOOST_net_4060), .b(n_13221), .o(TIMEBOOST_net_515) );
in01s01 g58039_u0 ( .a(FE_OFN606_n_9904), .o(g58039_sb) );
na02s01 g58039_u1 ( .a(FE_OFN207_n_9865), .b(g58039_sb), .o(g58039_da) );
na02s01 g58039_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q), .b(FE_OFN606_n_9904), .o(g58039_db) );
na02s01 g58039_u3 ( .a(g58039_da), .b(g58039_db), .o(n_9750) );
in01s01 g58040_u0 ( .a(FE_OFN606_n_9904), .o(g58040_sb) );
na02s01 TIMEBOOST_cell_38048 ( .a(TIMEBOOST_net_11262), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_4546) );
na02s01 g58040_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__10__Q), .b(FE_OFN606_n_9904), .o(g58040_db) );
na02m01 TIMEBOOST_cell_37444 ( .a(TIMEBOOST_net_10960), .b(g52470_sb), .o(TIMEBOOST_net_6232) );
in01s01 g58041_u0 ( .a(FE_OFN608_n_9904), .o(g58041_sb) );
na02s01 TIMEBOOST_cell_37460 ( .a(TIMEBOOST_net_10968), .b(FE_OFN775_n_15366), .o(TIMEBOOST_net_10568) );
na02s02 TIMEBOOST_cell_42376 ( .a(TIMEBOOST_net_13426), .b(g54338_sb), .o(n_12980) );
na02s01 TIMEBOOST_cell_37462 ( .a(TIMEBOOST_net_10969), .b(FE_OFN775_n_15366), .o(TIMEBOOST_net_10569) );
in01s01 g58042_u0 ( .a(n_9904), .o(g58042_sb) );
na02s01 TIMEBOOST_cell_9243 ( .a(TIMEBOOST_net_1188), .b(g65706_db), .o(n_2200) );
na02s01 g58042_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__Q), .b(n_9904), .o(g58042_db) );
na02f02 TIMEBOOST_cell_40466 ( .a(TIMEBOOST_net_12471), .b(n_17034), .o(TIMEBOOST_net_611) );
in01s01 g58043_u0 ( .a(FE_OFN1794_n_9904), .o(g58043_sb) );
na02s01 TIMEBOOST_cell_36508 ( .a(TIMEBOOST_net_10492), .b(FE_OFN1631_n_9531), .o(TIMEBOOST_net_3610) );
na02m02 TIMEBOOST_cell_44163 ( .a(n_9511), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__Q), .o(TIMEBOOST_net_14320) );
na02s01 TIMEBOOST_cell_36509 ( .a(TIMEBOOST_net_1207), .b(FE_OFN992_n_2373), .o(TIMEBOOST_net_10493) );
in01s01 g58044_u0 ( .a(FE_OFN606_n_9904), .o(g58044_sb) );
na02s01 g58044_u1 ( .a(FE_OFN213_n_9124), .b(g58044_sb), .o(g58044_da) );
na02s01 g58044_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__Q), .b(FE_OFN606_n_9904), .o(g58044_db) );
na02s01 g58044_u3 ( .a(g58044_da), .b(g58044_db), .o(n_9094) );
in01s01 g58045_u0 ( .a(FE_OFN606_n_9904), .o(g58045_sb) );
na02s01 TIMEBOOST_cell_44842 ( .a(TIMEBOOST_net_14659), .b(g64774_db), .o(n_3775) );
na02s01 g58045_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__15__Q), .b(FE_OFN606_n_9904), .o(g58045_db) );
na02s02 TIMEBOOST_cell_17611 ( .a(TIMEBOOST_net_4062), .b(g58235_sb), .o(n_9556) );
in01s01 g58046_u0 ( .a(FE_OFN608_n_9904), .o(g58046_sb) );
na03s02 TIMEBOOST_cell_41781 ( .a(g58012_sb), .b(g58012_db), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__Q), .o(TIMEBOOST_net_13129) );
na02s01 g58046_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q), .b(FE_OFN608_n_9904), .o(g58046_db) );
na02s02 TIMEBOOST_cell_41822 ( .a(TIMEBOOST_net_13149), .b(g58346_db), .o(n_9017) );
in01s01 g58047_u0 ( .a(FE_OFN1793_n_9904), .o(g58047_sb) );
in01s01 TIMEBOOST_cell_45916 ( .a(TIMEBOOST_net_15222), .o(TIMEBOOST_net_15223) );
na02s01 g58047_u2 ( .a(n_15569), .b(FE_OFN1793_n_9904), .o(g58047_db) );
na02s01 TIMEBOOST_cell_38194 ( .a(TIMEBOOST_net_11335), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_4619) );
in01s01 g58048_u0 ( .a(FE_OFN1795_n_9904), .o(g58048_sb) );
na02m02 TIMEBOOST_cell_38858 ( .a(TIMEBOOST_net_11667), .b(g58474_sb), .o(n_9368) );
na02s01 g58048_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__Q), .b(FE_OFN1795_n_9904), .o(g58048_db) );
na02s02 TIMEBOOST_cell_18555 ( .a(TIMEBOOST_net_4534), .b(g62857_sb), .o(n_5253) );
in01s01 g58049_u0 ( .a(FE_OFN606_n_9904), .o(g58049_sb) );
na02s02 TIMEBOOST_cell_37464 ( .a(TIMEBOOST_net_10970), .b(n_8892), .o(n_9484) );
na02s01 g58049_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__Q), .b(FE_OFN606_n_9904), .o(g58049_db) );
na02s02 TIMEBOOST_cell_37466 ( .a(TIMEBOOST_net_10971), .b(n_8892), .o(n_9411) );
in01s01 g58050_u0 ( .a(FE_OFN606_n_9904), .o(g58050_sb) );
na03f02 TIMEBOOST_cell_36230 ( .a(FE_RN_20_0), .b(n_12632), .c(n_12957), .o(n_13131) );
na02s01 g58050_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__Q), .b(FE_OFN606_n_9904), .o(g58050_db) );
na04f04 TIMEBOOST_cell_36231 ( .a(n_12897), .b(n_12959), .c(n_12789), .d(n_12896), .o(n_13135) );
in01s01 g58051_u0 ( .a(FE_OFN607_n_9904), .o(g58051_sb) );
na03f04 TIMEBOOST_cell_45861 ( .a(n_11912), .b(n_11915), .c(n_11914), .o(TIMEBOOST_net_15169) );
na02m02 TIMEBOOST_cell_43354 ( .a(TIMEBOOST_net_13915), .b(g59098_sb), .o(n_8695) );
na02s02 TIMEBOOST_cell_43465 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__Q), .b(n_4266), .o(TIMEBOOST_net_13971) );
in01s01 g58052_u0 ( .a(FE_OFN1794_n_9904), .o(g58052_sb) );
na02s01 TIMEBOOST_cell_9068 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__Q), .o(TIMEBOOST_net_1101) );
na02s01 g58052_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__Q), .b(FE_OFN1794_n_9904), .o(g58052_db) );
na02s01 TIMEBOOST_cell_9069 ( .a(TIMEBOOST_net_1101), .b(FE_OFN945_n_2248), .o(TIMEBOOST_net_141) );
in01s01 g58053_u0 ( .a(FE_OFN1793_n_9904), .o(g58053_sb) );
na02s01 TIMEBOOST_cell_9070 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__Q), .o(TIMEBOOST_net_1102) );
na02s01 TIMEBOOST_cell_43355 ( .a(n_4515), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__Q), .o(TIMEBOOST_net_13916) );
na02s01 TIMEBOOST_cell_41920 ( .a(TIMEBOOST_net_13198), .b(g57898_db), .o(n_9226) );
na02s01 g58054_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__Q), .b(n_9904), .o(g58054_db) );
na02s01 TIMEBOOST_cell_41918 ( .a(TIMEBOOST_net_13197), .b(g57891_db), .o(n_9233) );
in01s01 g58055_u0 ( .a(FE_OFN1793_n_9904), .o(g58055_sb) );
na02s02 TIMEBOOST_cell_38726 ( .a(TIMEBOOST_net_11601), .b(g61864_db), .o(n_8109) );
na02f02 TIMEBOOST_cell_43698 ( .a(TIMEBOOST_net_14087), .b(FE_OFN1349_n_8567), .o(TIMEBOOST_net_13310) );
na02s02 TIMEBOOST_cell_17785 ( .a(TIMEBOOST_net_4149), .b(g62011_sb), .o(n_7873) );
in01s01 g58056_u0 ( .a(FE_OFN606_n_9904), .o(g58056_sb) );
na02s02 TIMEBOOST_cell_37468 ( .a(TIMEBOOST_net_10972), .b(FE_OFN2257_n_8060), .o(TIMEBOOST_net_4099) );
na02s01 g58056_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q), .b(FE_OFN606_n_9904), .o(g58056_db) );
na02s02 TIMEBOOST_cell_37470 ( .a(TIMEBOOST_net_10973), .b(FE_OFN716_n_8176), .o(TIMEBOOST_net_4129) );
in01s01 g58057_u0 ( .a(FE_OFN1794_n_9904), .o(g58057_sb) );
na02s01 TIMEBOOST_cell_44843 ( .a(n_3792), .b(g64862_sb), .o(TIMEBOOST_net_14660) );
na02s01 g58057_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q), .b(FE_OFN1794_n_9904), .o(g58057_db) );
na02s01 TIMEBOOST_cell_36237 ( .a(pci_target_unit_del_sync_comp_cycle_count_1_), .b(pci_target_unit_del_sync_comp_cycle_count_0_), .o(TIMEBOOST_net_10357) );
in01s01 g58058_u0 ( .a(FE_OFN607_n_9904), .o(g58058_sb) );
na02s01 g58058_u1 ( .a(FE_OFN237_n_9118), .b(g58058_sb), .o(g58058_da) );
na02s01 g58058_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__Q), .b(FE_OFN607_n_9904), .o(g58058_db) );
na02s01 g58058_u3 ( .a(g58058_da), .b(g58058_db), .o(n_9091) );
in01s01 g58059_u0 ( .a(FE_OFN1795_n_9904), .o(g58059_sb) );
na02f02 TIMEBOOST_cell_39109 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_10164), .o(TIMEBOOST_net_11793) );
na02s01 g58059_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__Q), .b(FE_OFN1795_n_9904), .o(g58059_db) );
na02m02 TIMEBOOST_cell_38826 ( .a(TIMEBOOST_net_11651), .b(g58472_sb), .o(n_8981) );
in01s01 g58060_u0 ( .a(FE_OFN606_n_9904), .o(g58060_sb) );
na02s01 TIMEBOOST_cell_36510 ( .a(TIMEBOOST_net_10493), .b(g65994_sb), .o(n_2147) );
na02s02 TIMEBOOST_cell_43356 ( .a(TIMEBOOST_net_13916), .b(FE_OFN709_n_8232), .o(TIMEBOOST_net_11032) );
na02s01 TIMEBOOST_cell_36511 ( .a(g58042_sb), .b(g58065_db), .o(TIMEBOOST_net_10494) );
na02s01 TIMEBOOST_cell_37472 ( .a(TIMEBOOST_net_10974), .b(FE_OFN717_n_8176), .o(TIMEBOOST_net_4098) );
na02f02 TIMEBOOST_cell_44313 ( .a(n_9788), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__Q), .o(TIMEBOOST_net_14395) );
na02s01 TIMEBOOST_cell_37474 ( .a(TIMEBOOST_net_10975), .b(FE_OFN717_n_8176), .o(TIMEBOOST_net_4164) );
in01s01 g58062_u0 ( .a(FE_OFN1795_n_9904), .o(g58062_sb) );
na02s01 TIMEBOOST_cell_9072 ( .a(pci_target_unit_fifos_pcir_data_in_163), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__Q), .o(TIMEBOOST_net_1103) );
na02f02 TIMEBOOST_cell_41666 ( .a(TIMEBOOST_net_13071), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_11735) );
na02s01 TIMEBOOST_cell_9073 ( .a(TIMEBOOST_net_1103), .b(FE_OFN945_n_2248), .o(TIMEBOOST_net_143) );
in01s01 g58063_u0 ( .a(FE_OFN606_n_9904), .o(g58063_sb) );
na04m04 TIMEBOOST_cell_35852 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_18__Q), .b(FE_OFN262_n_9851), .c(FE_OFN1439_n_9372), .d(g58464_sb), .o(n_9387) );
na02s01 g58063_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q), .b(FE_OFN606_n_9904), .o(g58063_db) );
na02s01 TIMEBOOST_cell_31921 ( .a(TIMEBOOST_net_9871), .b(g57904_db), .o(n_9222) );
na02s01 TIMEBOOST_cell_45581 ( .a(n_15567), .b(FE_OFN1648_n_9428), .o(TIMEBOOST_net_15029) );
na02s01 g58064_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__Q), .b(FE_OFN607_n_9904), .o(g58064_db) );
na02s01 TIMEBOOST_cell_17954 ( .a(n_4476), .b(FE_OFN1680_n_4655), .o(TIMEBOOST_net_4234) );
na02s01 TIMEBOOST_cell_16640 ( .a(pci_target_unit_fifos_pciw_addr_data_in_149), .b(g64159_sb), .o(TIMEBOOST_net_3577) );
na02s01 g58065_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__Q), .b(n_9904), .o(g58065_db) );
na02s01 TIMEBOOST_cell_16641 ( .a(TIMEBOOST_net_3577), .b(g64159_db), .o(n_4006) );
in01s01 g58066_u0 ( .a(FE_OFN606_n_9904), .o(g58066_sb) );
na02s01 g58066_u1 ( .a(FE_OFN252_n_9868), .b(g58066_sb), .o(g58066_da) );
na02s01 g58066_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__8__Q), .b(FE_OFN606_n_9904), .o(g58066_db) );
na02s01 g58066_u3 ( .a(g58066_da), .b(g58066_db), .o(n_9726) );
na02f02 TIMEBOOST_cell_42168 ( .a(TIMEBOOST_net_13322), .b(FE_OFN1396_n_8567), .o(TIMEBOOST_net_12266) );
na02s01 g58067_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__Q), .b(FE_OFN608_n_9904), .o(g58067_db) );
na02s02 TIMEBOOST_cell_17787 ( .a(TIMEBOOST_net_4150), .b(g62071_sb), .o(n_7826) );
in01s01 g58068_u0 ( .a(FE_OFN1793_n_9904), .o(g58068_sb) );
na02s02 TIMEBOOST_cell_37696 ( .a(TIMEBOOST_net_11086), .b(g61823_sb), .o(n_8142) );
na03f02 TIMEBOOST_cell_44447 ( .a(n_8558), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__Q), .c(FE_OFN1403_n_8567), .o(TIMEBOOST_net_14462) );
na03s02 TIMEBOOST_cell_37697 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__Q), .b(FE_OFN2084_n_8407), .c(n_1596), .o(TIMEBOOST_net_11087) );
in01s01 g58069_u0 ( .a(FE_OFN576_n_9902), .o(g58069_sb) );
na02s01 g58069_u1 ( .a(FE_OFN207_n_9865), .b(g58069_sb), .o(g58069_da) );
na02s01 g58069_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__Q), .b(FE_OFN576_n_9902), .o(g58069_db) );
na02s01 g58069_u3 ( .a(g58069_da), .b(g58069_db), .o(n_9723) );
in01s01 g58070_u0 ( .a(FE_OFN577_n_9902), .o(g58070_sb) );
na02m02 TIMEBOOST_cell_10314 ( .a(g54141_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_406), .o(TIMEBOOST_net_1724) );
na02s01 TIMEBOOST_cell_45650 ( .a(TIMEBOOST_net_15063), .b(g58207_db), .o(n_9579) );
na02s01 TIMEBOOST_cell_37476 ( .a(TIMEBOOST_net_10976), .b(g65829_sb), .o(TIMEBOOST_net_327) );
in01s01 g58071_u0 ( .a(FE_OFN575_n_9902), .o(g58071_sb) );
na02f02 TIMEBOOST_cell_37075 ( .a(TIMEBOOST_net_10239), .b(FE_OCP_RBN1998_n_13971), .o(TIMEBOOST_net_10776) );
na02f02 TIMEBOOST_cell_42462 ( .a(TIMEBOOST_net_13469), .b(g57064_sb), .o(n_10501) );
na02s01 TIMEBOOST_cell_37446 ( .a(TIMEBOOST_net_10961), .b(g58430_db), .o(n_8996) );
in01s01 g58072_u0 ( .a(FE_OFN574_n_9902), .o(g58072_sb) );
na02s01 g58072_u1 ( .a(FE_OFN209_n_9126), .b(g58072_sb), .o(g58072_da) );
na02s01 g58072_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__Q), .b(FE_OFN574_n_9902), .o(g58072_db) );
na02s01 g58072_u3 ( .a(g58072_da), .b(g58072_db), .o(n_9087) );
in01s01 g58073_u0 ( .a(FE_OFN577_n_9902), .o(g58073_sb) );
na02s01 g58073_u1 ( .a(FE_OFN211_n_9858), .b(g58073_sb), .o(g58073_da) );
na02s01 g58073_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__Q), .b(FE_OFN577_n_9902), .o(g58073_db) );
na02s01 g58073_u3 ( .a(g58073_da), .b(g58073_db), .o(n_9720) );
in01s01 g58074_u0 ( .a(FE_OFN576_n_9902), .o(g58074_sb) );
na02m02 TIMEBOOST_cell_38945 ( .a(wbu_sel_in_314), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_35__Q), .o(TIMEBOOST_net_11711) );
na02s01 g58074_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__Q), .b(FE_OFN576_n_9902), .o(g58074_db) );
na02f02 TIMEBOOST_cell_39110 ( .a(TIMEBOOST_net_11793), .b(FE_OFN1600_n_13995), .o(n_14472) );
in01s01 g58075_u0 ( .a(FE_OFN576_n_9902), .o(g58075_sb) );
na02s01 TIMEBOOST_cell_9195 ( .a(TIMEBOOST_net_1164), .b(g65712_db), .o(n_2198) );
na02s01 g58075_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__Q), .b(FE_OFN576_n_9902), .o(g58075_db) );
na02s02 TIMEBOOST_cell_37478 ( .a(TIMEBOOST_net_10977), .b(g65383_sb), .o(n_4245) );
in01s01 g58076_u0 ( .a(FE_OFN577_n_9902), .o(g58076_sb) );
na02s01 g58076_u1 ( .a(FE_OFN217_n_9889), .b(g58076_sb), .o(g58076_da) );
na02s01 g58076_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__Q), .b(FE_OFN577_n_9902), .o(g58076_db) );
na02s01 g58076_u3 ( .a(g58076_da), .b(g58076_db), .o(n_9718) );
in01s01 g58077_u0 ( .a(FE_OFN575_n_9902), .o(g58077_sb) );
na02s01 g58077_u1 ( .a(FE_OFN219_n_9853), .b(g58077_sb), .o(g58077_da) );
na02s01 g58077_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__Q), .b(FE_OFN575_n_9902), .o(g58077_db) );
na02s01 g58077_u3 ( .a(g58077_da), .b(g58077_db), .o(n_9717) );
in01s01 g58078_u0 ( .a(FE_OFN577_n_9902), .o(g58078_sb) );
na02s02 TIMEBOOST_cell_37448 ( .a(TIMEBOOST_net_10962), .b(FE_OFN1634_n_9531), .o(TIMEBOOST_net_4056) );
na02s01 TIMEBOOST_cell_45651 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__Q), .b(FE_OFN270_n_9836), .o(TIMEBOOST_net_15064) );
na02s02 TIMEBOOST_cell_10558 ( .a(pci_cbe_o_3_), .b(n_14389), .o(TIMEBOOST_net_1846) );
in01s01 g58079_u0 ( .a(FE_OFN577_n_9902), .o(g58079_sb) );
na02s02 TIMEBOOST_cell_37372 ( .a(TIMEBOOST_net_10924), .b(g58322_db), .o(n_9491) );
na02s02 TIMEBOOST_cell_45652 ( .a(TIMEBOOST_net_15064), .b(FE_OFN1690_n_9528), .o(TIMEBOOST_net_11161) );
na02s02 TIMEBOOST_cell_37374 ( .a(TIMEBOOST_net_10925), .b(g58431_db), .o(n_9416) );
in01s01 g58080_u0 ( .a(FE_OFN577_n_9902), .o(g58080_sb) );
na02s01 g58080_u1 ( .a(FE_OFN221_n_9846), .b(g58080_sb), .o(g58080_da) );
na02s01 g58080_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q), .b(FE_OFN577_n_9902), .o(g58080_db) );
na02s01 g58080_u3 ( .a(g58080_da), .b(g58080_db), .o(n_9714) );
in01s01 g58081_u0 ( .a(FE_OFN574_n_9902), .o(g58081_sb) );
na02s01 TIMEBOOST_cell_36388 ( .a(TIMEBOOST_net_10432), .b(g65700_db), .o(n_2202) );
na02s01 g58081_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__Q), .b(FE_OFN574_n_9902), .o(g58081_db) );
na02m02 TIMEBOOST_cell_38860 ( .a(TIMEBOOST_net_11668), .b(g58469_sb), .o(n_8983) );
in01s01 g58082_u0 ( .a(FE_OFN577_n_9902), .o(g58082_sb) );
na02s01 g58082_u1 ( .a(FE_OFN225_n_9122), .b(g58082_sb), .o(g58082_da) );
na02s01 g58082_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__Q), .b(FE_OFN577_n_9902), .o(g58082_db) );
na02s01 g58082_u3 ( .a(g58082_da), .b(g58082_db), .o(n_9085) );
in01s01 g58083_u0 ( .a(FE_OFN575_n_9902), .o(g58083_sb) );
na02s01 TIMEBOOST_cell_37698 ( .a(TIMEBOOST_net_11087), .b(g61826_sb), .o(n_8135) );
na02f02 TIMEBOOST_cell_41528 ( .a(TIMEBOOST_net_13002), .b(g57562_sb), .o(n_11190) );
na02s01 TIMEBOOST_cell_37376 ( .a(TIMEBOOST_net_10926), .b(g58429_db), .o(n_9418) );
in01s01 g58084_u0 ( .a(FE_OFN575_n_9902), .o(g58084_sb) );
na02s01 g58084_u1 ( .a(FE_OFN227_n_9841), .b(g58084_sb), .o(g58084_da) );
na02s01 g58084_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__Q), .b(FE_OFN575_n_9902), .o(g58084_db) );
na02s02 g58084_u3 ( .a(g58084_da), .b(g58084_db), .o(n_9711) );
na02s01 g58085_u1 ( .a(FE_OFN229_n_9120), .b(g58097_sb), .o(g58085_da) );
na02s01 g58085_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__Q), .b(FE_OFN574_n_9902), .o(g58085_db) );
na02s02 g58085_u3 ( .a(g58085_da), .b(g58085_db), .o(n_9084) );
in01s01 g58086_u0 ( .a(FE_OFN575_n_9902), .o(g58086_sb) );
na02s01 TIMEBOOST_cell_9662 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__Q), .b(g58432_sb), .o(TIMEBOOST_net_1398) );
na02s01 g58086_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__Q), .b(FE_OFN575_n_9902), .o(g58086_db) );
na02s02 TIMEBOOST_cell_9663 ( .a(TIMEBOOST_net_1398), .b(g58432_db), .o(n_8995) );
in01s01 g58087_u0 ( .a(FE_OFN577_n_9902), .o(g58087_sb) );
na02s01 g58087_u1 ( .a(FE_OFN233_n_9876), .b(g58087_sb), .o(g58087_da) );
na02s01 g58087_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__Q), .b(FE_OFN577_n_9902), .o(g58087_db) );
na02s01 g58087_u3 ( .a(g58087_da), .b(g58087_db), .o(n_9709) );
in01s01 g58088_u0 ( .a(FE_OFN576_n_9902), .o(g58088_sb) );
na02s01 TIMEBOOST_cell_37378 ( .a(TIMEBOOST_net_10927), .b(g64766_sb), .o(n_3782) );
na02s02 TIMEBOOST_cell_45653 ( .a(n_1750), .b(g60682_da), .o(TIMEBOOST_net_15065) );
na02f02 TIMEBOOST_cell_39112 ( .a(TIMEBOOST_net_11794), .b(FE_OFN1601_n_13995), .o(n_14514) );
in01s01 g58089_u0 ( .a(FE_OFN577_n_9902), .o(g58089_sb) );
na02s01 g58089_u1 ( .a(FE_OFN235_n_9834), .b(g58089_sb), .o(g58089_da) );
na02s01 g58089_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__Q), .b(FE_OFN577_n_9902), .o(g58089_db) );
na02s02 g58089_u3 ( .a(g58089_da), .b(g58089_db), .o(n_9707) );
in01s01 g58090_u0 ( .a(FE_OFN574_n_9902), .o(g58090_sb) );
na02s01 g58090_u1 ( .a(FE_OFN237_n_9118), .b(g58090_sb), .o(g58090_da) );
na02s01 g58090_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q), .b(FE_OFN574_n_9902), .o(g58090_db) );
na02s01 g58090_u3 ( .a(g58090_da), .b(g58090_db), .o(n_9083) );
in01s01 g58091_u0 ( .a(FE_OFN577_n_9902), .o(g58091_sb) );
na02s01 g58091_u1 ( .a(FE_OFN239_n_9832), .b(g58091_sb), .o(g58091_da) );
na02s01 g58091_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__Q), .b(FE_OFN577_n_9902), .o(g58091_db) );
na02s01 g58091_u3 ( .a(g58091_da), .b(g58091_db), .o(n_9706) );
in01s01 g58092_u0 ( .a(FE_OFN576_n_9902), .o(g58092_sb) );
na02s01 g58092_u1 ( .a(FE_OFN241_n_9830), .b(g58092_sb), .o(g58092_da) );
na02s01 g58092_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__Q), .b(FE_OFN576_n_9902), .o(g58092_db) );
na02s01 g58092_u3 ( .a(g58092_da), .b(g58092_db), .o(n_9705) );
in01s01 g58093_u0 ( .a(FE_OFN575_n_9902), .o(g58093_sb) );
na02s02 TIMEBOOST_cell_37380 ( .a(TIMEBOOST_net_10928), .b(g58120_sb), .o(n_9076) );
na02m02 TIMEBOOST_cell_32568 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q), .o(TIMEBOOST_net_10195) );
na02s02 TIMEBOOST_cell_37382 ( .a(TIMEBOOST_net_10929), .b(n_4479), .o(n_4262) );
in01s01 g58094_u0 ( .a(FE_OFN577_n_9902), .o(g58094_sb) );
na02s01 TIMEBOOST_cell_42700 ( .a(TIMEBOOST_net_13588), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_10046) );
na02s01 g58094_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__Q), .b(FE_OFN577_n_9902), .o(g58094_db) );
na02f02 TIMEBOOST_cell_40465 ( .a(n_17048), .b(n_4880), .o(TIMEBOOST_net_12471) );
in01s01 g58095_u0 ( .a(FE_OFN576_n_9902), .o(g58095_sb) );
na02s02 TIMEBOOST_cell_40468 ( .a(TIMEBOOST_net_12472), .b(n_8590), .o(TIMEBOOST_net_11485) );
na02s01 g58095_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__Q), .b(FE_OFN576_n_9902), .o(g58095_db) );
na02s01 TIMEBOOST_cell_31920 ( .a(FE_OFN203_n_9228), .b(g57904_sb), .o(TIMEBOOST_net_9871) );
in01s01 g58096_u0 ( .a(FE_OFN574_n_9902), .o(g58096_sb) );
na02f02 TIMEBOOST_cell_44164 ( .a(TIMEBOOST_net_14320), .b(FE_OFN1401_n_8567), .o(TIMEBOOST_net_13391) );
na02s01 g58096_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q), .b(FE_OFN574_n_9902), .o(g58096_db) );
na02m02 TIMEBOOST_cell_38862 ( .a(TIMEBOOST_net_11669), .b(g58457_sb), .o(n_9398) );
in01s01 g58097_u0 ( .a(FE_OFN574_n_9902), .o(g58097_sb) );
na02s01 g58097_u1 ( .a(FE_OFN250_n_9789), .b(g58097_sb), .o(g58097_da) );
na02s01 g58097_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__Q), .b(FE_OFN574_n_9902), .o(g58097_db) );
na02s02 g58097_u3 ( .a(g58097_da), .b(g58097_db), .o(n_9703) );
na02s02 TIMEBOOST_cell_37384 ( .a(TIMEBOOST_net_10930), .b(FE_OFN681_n_4460), .o(TIMEBOOST_net_9489) );
na02m02 TIMEBOOST_cell_32550 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__Q), .o(TIMEBOOST_net_10186) );
na03s02 TIMEBOOST_cell_38195 ( .a(TIMEBOOST_net_3994), .b(g64110_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__Q), .o(TIMEBOOST_net_11336) );
in01s01 g58099_u0 ( .a(FE_OFN534_n_9823), .o(g58099_sb) );
na02s01 g58099_u1 ( .a(FE_OFN252_n_9868), .b(g58099_sb), .o(g58099_da) );
na02s01 g58099_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__Q), .b(FE_OFN534_n_9823), .o(g58099_db) );
na02s01 g58099_u3 ( .a(g58099_da), .b(g58099_db), .o(n_9701) );
in01s01 g58100_u0 ( .a(FE_OFN535_n_9823), .o(g58100_sb) );
na02m02 TIMEBOOST_cell_44165 ( .a(n_9718), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__Q), .o(TIMEBOOST_net_14321) );
na02s01 g58100_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__Q), .b(FE_OFN535_n_9823), .o(g58100_db) );
na02s01 TIMEBOOST_cell_38728 ( .a(TIMEBOOST_net_11602), .b(g61870_db), .o(n_8094) );
in01s01 g58101_u0 ( .a(FE_OFN519_n_9697), .o(g58101_sb) );
na02s01 g58101_u1 ( .a(FE_OFN252_n_9868), .b(g58101_sb), .o(g58101_da) );
na02s01 g58101_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__Q), .b(FE_OFN519_n_9697), .o(g58101_db) );
na02s01 g58101_u3 ( .a(g58101_da), .b(g58101_db), .o(n_9698) );
in01s01 g58102_u0 ( .a(FE_OFN595_n_9694), .o(g58102_sb) );
na03s02 TIMEBOOST_cell_40469 ( .a(n_3956), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__Q), .c(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_12473) );
na02s01 g58102_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__Q), .b(FE_OFN595_n_9694), .o(g58102_db) );
na02s02 TIMEBOOST_cell_38068 ( .a(TIMEBOOST_net_11272), .b(FE_OFN877_g64577_p), .o(TIMEBOOST_net_4559) );
in01s01 g58103_u0 ( .a(FE_OFN588_n_9692), .o(g58103_sb) );
na02s02 TIMEBOOST_cell_40470 ( .a(TIMEBOOST_net_12473), .b(g62861_sb), .o(n_5244) );
na02s01 g58103_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__Q), .b(FE_OFN588_n_9692), .o(g58103_db) );
na03s02 TIMEBOOST_cell_40471 ( .a(n_366), .b(FE_OFN1127_g64577_p), .c(n_4733), .o(TIMEBOOST_net_12474) );
in01s01 g58104_u0 ( .a(FE_OFN587_n_9692), .o(g58104_sb) );
na02s01 g58104_u1 ( .a(FE_OFN243_n_9116), .b(g58104_sb), .o(g58104_da) );
na02s01 g58104_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__Q), .b(FE_OFN587_n_9692), .o(g58104_db) );
na02s01 g58104_u3 ( .a(g58104_da), .b(g58104_db), .o(n_9079) );
in01s01 g58105_u0 ( .a(FE_OFN1803_n_9690), .o(g58105_sb) );
na02s02 TIMEBOOST_cell_38451 ( .a(TIMEBOOST_net_9855), .b(FE_OFN1085_n_13221), .o(TIMEBOOST_net_11464) );
na02s01 TIMEBOOST_cell_18020 ( .a(pci_target_unit_fifos_pciw_addr_data_in_139), .b(g64100_sb), .o(TIMEBOOST_net_4267) );
na03s02 TIMEBOOST_cell_36889 ( .a(g58598_db), .b(pci_target_unit_fifos_pcir_flush_in), .c(g57780_da), .o(TIMEBOOST_net_10683) );
in01s01 g58106_u0 ( .a(FE_OFN602_n_9687), .o(g58106_sb) );
na02s01 TIMEBOOST_cell_9197 ( .a(TIMEBOOST_net_1165), .b(g65772_db), .o(n_2194) );
na02s01 g58106_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__Q), .b(FE_OFN602_n_9687), .o(g58106_db) );
na03s02 TIMEBOOST_cell_38057 ( .a(g64350_da), .b(g64350_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__Q), .o(TIMEBOOST_net_11267) );
in01s01 g58107_u0 ( .a(FE_OFN601_n_9687), .o(g58107_sb) );
na02s01 TIMEBOOST_cell_37386 ( .a(TIMEBOOST_net_10931), .b(FE_OFN686_n_4417), .o(TIMEBOOST_net_9486) );
na02s02 TIMEBOOST_cell_45399 ( .a(n_3725), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__Q), .o(TIMEBOOST_net_14938) );
na02s01 TIMEBOOST_cell_37388 ( .a(TIMEBOOST_net_10932), .b(FE_OFN685_n_4417), .o(TIMEBOOST_net_9498) );
in01s01 g58108_u0 ( .a(FE_OFN600_n_9687), .o(g58108_sb) );
na02s01 TIMEBOOST_cell_42766 ( .a(TIMEBOOST_net_13621), .b(FE_OFN233_n_9876), .o(TIMEBOOST_net_10044) );
na02m02 TIMEBOOST_cell_44375 ( .a(n_9128), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q), .o(TIMEBOOST_net_14426) );
na02s01 TIMEBOOST_cell_38640 ( .a(TIMEBOOST_net_11558), .b(g59112_sb), .o(n_8705) );
na02s01 g58109_u1 ( .a(FE_OFN209_n_9126), .b(FE_OFN599_n_9687), .o(g58109_da) );
na02s01 g58109_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__Q), .b(FE_OFN603_n_9687), .o(g58109_db) );
na02s01 g58109_u3 ( .a(g58109_da), .b(g58109_db), .o(n_9078) );
in01s01 g58110_u0 ( .a(FE_OFN601_n_9687), .o(g58110_sb) );
na02f02 TIMEBOOST_cell_38946 ( .a(TIMEBOOST_net_11711), .b(FE_OFN2155_n_16439), .o(TIMEBOOST_net_10737) );
na02s01 g58110_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__Q), .b(FE_OFN601_n_9687), .o(g58110_db) );
na02s01 TIMEBOOST_cell_39302 ( .a(TIMEBOOST_net_11889), .b(g65890_db), .o(n_1859) );
in01s01 g58111_u0 ( .a(FE_OFN602_n_9687), .o(g58111_sb) );
na02s01 g58111_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__Q), .b(FE_OFN602_n_9687), .o(g58111_db) );
na02s02 TIMEBOOST_cell_40410 ( .a(TIMEBOOST_net_12443), .b(FE_OFN262_n_9851), .o(n_9497) );
in01s01 g58112_u0 ( .a(FE_OFN602_n_9687), .o(g58112_sb) );
na02s01 TIMEBOOST_cell_39364 ( .a(TIMEBOOST_net_11920), .b(g61874_sb), .o(n_8084) );
na02s01 g58112_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__Q), .b(FE_OFN602_n_9687), .o(g58112_db) );
na02s02 TIMEBOOST_cell_40412 ( .a(TIMEBOOST_net_12444), .b(FE_OFN262_n_9851), .o(n_9447) );
in01s01 g58113_u0 ( .a(FE_OFN601_n_9687), .o(g58113_sb) );
na02s01 g58113_u1 ( .a(FE_OFN217_n_9889), .b(g58113_sb), .o(g58113_da) );
na02s01 g58113_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__Q), .b(FE_OFN601_n_9687), .o(g58113_db) );
na02s01 g58113_u3 ( .a(g58113_da), .b(g58113_db), .o(n_9682) );
in01s01 g58114_u0 ( .a(FE_OFN600_n_9687), .o(g58114_sb) );
na02s01 g58114_u1 ( .a(FE_OFN219_n_9853), .b(g58114_sb), .o(g58114_da) );
na02s01 g58114_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__Q), .b(FE_OFN600_n_9687), .o(g58114_db) );
na02s01 g58114_u3 ( .a(g58114_da), .b(g58114_db), .o(n_9680) );
in01s01 g58115_u0 ( .a(FE_OFN600_n_9687), .o(g58115_sb) );
na02f02 TIMEBOOST_cell_41052 ( .a(TIMEBOOST_net_12764), .b(g57398_sb), .o(n_10372) );
na02s01 g58115_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__Q), .b(FE_OFN600_n_9687), .o(g58115_db) );
na02s02 TIMEBOOST_cell_38196 ( .a(TIMEBOOST_net_11336), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_4617) );
in01s01 g58116_u0 ( .a(FE_OFN601_n_9687), .o(g58116_sb) );
na02s02 TIMEBOOST_cell_18937 ( .a(TIMEBOOST_net_4725), .b(g58446_sb), .o(n_9199) );
na02s02 TIMEBOOST_cell_45400 ( .a(TIMEBOOST_net_14938), .b(FE_OFN1248_n_4093), .o(TIMEBOOST_net_12608) );
na02s01 TIMEBOOST_cell_37220 ( .a(TIMEBOOST_net_10848), .b(FE_OFN2096_n_2520), .o(TIMEBOOST_net_10491) );
in01s01 g58117_u0 ( .a(FE_OFN602_n_9687), .o(g58117_sb) );
na02s02 TIMEBOOST_cell_37222 ( .a(TIMEBOOST_net_10849), .b(TIMEBOOST_net_9310), .o(TIMEBOOST_net_10090) );
na02s01 TIMEBOOST_cell_41951 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__Q), .b(n_4163), .o(TIMEBOOST_net_13214) );
na02s01 TIMEBOOST_cell_37224 ( .a(TIMEBOOST_net_10850), .b(FE_OFN2095_n_2520), .o(TIMEBOOST_net_9326) );
in01s01 g58118_u0 ( .a(FE_OFN601_n_9687), .o(g58118_sb) );
na02s02 TIMEBOOST_cell_40414 ( .a(TIMEBOOST_net_12445), .b(FE_OFN266_n_9884), .o(n_9495) );
na02s01 g58118_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__Q), .b(FE_OFN601_n_9687), .o(g58118_db) );
na02s01 TIMEBOOST_cell_9347 ( .a(TIMEBOOST_net_1240), .b(g60677_sb), .o(n_3589) );
in01s01 g58119_u0 ( .a(FE_OFN601_n_9687), .o(g58119_sb) );
na02s01 g58119_u1 ( .a(FE_OFN223_n_9844), .b(g58119_sb), .o(g58119_da) );
na02s01 g58119_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__Q), .b(FE_OFN601_n_9687), .o(g58119_db) );
na02s01 g58119_u3 ( .a(g58119_da), .b(g58119_db), .o(n_9673) );
in01s01 g58120_u0 ( .a(FE_OFN2254_n_9687), .o(g58120_sb) );
na02s01 TIMEBOOST_cell_17466 ( .a(n_4493), .b(FE_OFN642_n_4677), .o(TIMEBOOST_net_3990) );
na02s02 TIMEBOOST_cell_39716 ( .a(TIMEBOOST_net_12096), .b(g63146_sb), .o(n_5848) );
na02s01 TIMEBOOST_cell_39374 ( .a(TIMEBOOST_net_11925), .b(FE_OFN704_n_8069), .o(TIMEBOOST_net_4341) );
na02s01 g58121_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__Q), .b(FE_OFN600_n_9687), .o(g58121_db) );
na03s02 TIMEBOOST_cell_1112 ( .a(n_3215), .b(g63435_sb), .c(g63435_db), .o(n_4625) );
na02s02 TIMEBOOST_cell_40472 ( .a(TIMEBOOST_net_12474), .b(g63035_sb), .o(n_7126) );
na03s02 TIMEBOOST_cell_40473 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__Q), .b(FE_OFN1127_g64577_p), .c(g62749_sb), .o(TIMEBOOST_net_12475) );
in01s02 g58123_u0 ( .a(FE_OFN603_n_9687), .o(g58123_sb) );
na02s01 g58123_u1 ( .a(FE_OFN229_n_9120), .b(g58123_sb), .o(g58123_da) );
na02s01 g58123_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__Q), .b(FE_OFN603_n_9687), .o(g58123_db) );
na02s02 g58123_u3 ( .a(g58123_da), .b(g58123_db), .o(n_9075) );
in01s01 g58124_u0 ( .a(FE_OFN601_n_9687), .o(g58124_sb) );
na02s01 TIMEBOOST_cell_9349 ( .a(TIMEBOOST_net_1241), .b(g65286_sb), .o(TIMEBOOST_net_219) );
na02s01 g58124_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__Q), .b(FE_OFN601_n_9687), .o(g58124_db) );
na02s01 TIMEBOOST_cell_44822 ( .a(TIMEBOOST_net_14649), .b(g65694_db), .o(TIMEBOOST_net_266) );
in01s01 g58125_u0 ( .a(FE_OFN601_n_9687), .o(g58125_sb) );
na02s02 TIMEBOOST_cell_36671 ( .a(n_1606), .b(g61798_sb), .o(TIMEBOOST_net_10574) );
na02s01 g58125_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__Q), .b(FE_OFN601_n_9687), .o(g58125_db) );
na02s02 TIMEBOOST_cell_43411 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__Q), .b(n_3793), .o(TIMEBOOST_net_13944) );
in01s01 g58126_u0 ( .a(FE_OFN602_n_9687), .o(g58126_sb) );
na02f02 TIMEBOOST_cell_39376 ( .a(g54304_sb), .b(TIMEBOOST_net_11926), .o(TIMEBOOST_net_10576) );
na02s01 TIMEBOOST_cell_39378 ( .a(TIMEBOOST_net_11927), .b(g58211_da), .o(TIMEBOOST_net_10054) );
in01s01 g58127_u0 ( .a(FE_OFN2253_n_9687), .o(g58127_sb) );
na02s01 TIMEBOOST_cell_44925 ( .a(FE_OFN213_n_9124), .b(g58013_sb), .o(TIMEBOOST_net_14701) );
na02s02 g58127_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__Q), .b(FE_OFN2253_n_9687), .o(g58127_db) );
na02s02 TIMEBOOST_cell_39718 ( .a(TIMEBOOST_net_12097), .b(g62398_sb), .o(n_6804) );
in01s01 g58128_u0 ( .a(FE_OFN601_n_9687), .o(g58128_sb) );
na02s01 g58128_u1 ( .a(FE_OFN237_n_9118), .b(g58128_sb), .o(g58128_da) );
na02s01 g58128_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__Q), .b(FE_OFN601_n_9687), .o(g58128_db) );
na02s01 g58128_u3 ( .a(g58128_da), .b(g58128_db), .o(n_9074) );
in01s01 g58129_u0 ( .a(FE_OFN601_n_9687), .o(g58129_sb) );
na02s02 TIMEBOOST_cell_43412 ( .a(TIMEBOOST_net_13944), .b(n_6554), .o(TIMEBOOST_net_12201) );
na02s01 g58129_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__Q), .b(FE_OFN601_n_9687), .o(g58129_db) );
na02s01 TIMEBOOST_cell_39288 ( .a(TIMEBOOST_net_11882), .b(g65768_sb), .o(n_1664) );
in01s01 g58130_u0 ( .a(FE_OFN602_n_9687), .o(g58130_sb) );
na02s01 TIMEBOOST_cell_37700 ( .a(TIMEBOOST_net_11088), .b(g61704_sb), .o(n_8419) );
na02s01 g58130_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__Q), .b(FE_OFN602_n_9687), .o(g58130_db) );
na02s01 TIMEBOOST_cell_39290 ( .a(TIMEBOOST_net_11883), .b(g65771_db), .o(n_1602) );
na02s02 TIMEBOOST_cell_39380 ( .a(TIMEBOOST_net_11928), .b(n_2276), .o(TIMEBOOST_net_5313) );
na02s02 TIMEBOOST_cell_22293 ( .a(n_10180), .b(TIMEBOOST_net_6403), .o(n_11859) );
na02s02 TIMEBOOST_cell_39382 ( .a(TIMEBOOST_net_11929), .b(FE_OFN707_n_8119), .o(TIMEBOOST_net_4373) );
in01s01 g58132_u0 ( .a(FE_OFN601_n_9687), .o(g58132_sb) );
na02s01 TIMEBOOST_cell_40474 ( .a(TIMEBOOST_net_12475), .b(n_4527), .o(n_6132) );
na02s01 g58132_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__Q), .b(FE_OFN601_n_9687), .o(g58132_db) );
na02s02 TIMEBOOST_cell_31918 ( .a(FE_OFN201_n_9230), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__Q), .o(TIMEBOOST_net_9870) );
in01s01 g58133_u0 ( .a(FE_OFN602_n_9687), .o(g58133_sb) );
na02s01 g58133_u1 ( .a(FE_OFN245_n_9114), .b(g58133_sb), .o(g58133_da) );
na02s01 g58133_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__Q), .b(FE_OFN602_n_9687), .o(g58133_db) );
na02s01 g58133_u3 ( .a(g58133_da), .b(g58133_db), .o(n_9072) );
na02s01 TIMEBOOST_cell_37702 ( .a(TIMEBOOST_net_11089), .b(g61951_sb), .o(n_7923) );
na02s01 g58134_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q), .b(FE_OFN603_n_9687), .o(g58134_db) );
na02s02 TIMEBOOST_cell_39438 ( .a(TIMEBOOST_net_11957), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_4533) );
na02s01 g58135_u1 ( .a(FE_OFN250_n_9789), .b(g58123_sb), .o(g58135_da) );
na02s01 g58135_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__Q), .b(FE_OFN603_n_9687), .o(g58135_db) );
na02s02 g58135_u3 ( .a(g58135_da), .b(g58135_db), .o(n_9661) );
in01s01 g58136_u0 ( .a(FE_OFN602_n_9687), .o(g58136_sb) );
na02f02 TIMEBOOST_cell_39114 ( .a(TIMEBOOST_net_11795), .b(FE_OFN1602_n_13995), .o(n_14443) );
na02s01 g58136_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q), .b(FE_OFN602_n_9687), .o(g58136_db) );
na02s01 TIMEBOOST_cell_37704 ( .a(TIMEBOOST_net_11090), .b(g61914_sb), .o(n_7993) );
na02m02 TIMEBOOST_cell_41599 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_1__Q), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_13038) );
na02s01 TIMEBOOST_cell_43298 ( .a(TIMEBOOST_net_13887), .b(g62712_sb), .o(n_6146) );
na02s02 TIMEBOOST_cell_37706 ( .a(TIMEBOOST_net_11091), .b(g61790_sb), .o(n_8220) );
in01s01 g58138_u0 ( .a(FE_OFN519_n_9697), .o(g58138_sb) );
na02s01 g58138_u1 ( .a(FE_OFN207_n_9865), .b(g58138_sb), .o(g58138_da) );
na02s01 g58138_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__Q), .b(FE_OFN519_n_9697), .o(g58138_db) );
na02s01 g58138_u3 ( .a(g58138_da), .b(g58138_db), .o(n_9658) );
in01s01 g58139_u0 ( .a(FE_OFN517_n_9697), .o(g58139_sb) );
na02s01 TIMEBOOST_cell_37226 ( .a(TIMEBOOST_net_10851), .b(g65325_sb), .o(TIMEBOOST_net_3560) );
na02s01 TIMEBOOST_cell_15787 ( .a(TIMEBOOST_net_3150), .b(g67042_sb), .o(n_1275) );
na02s02 TIMEBOOST_cell_39384 ( .a(TIMEBOOST_net_11930), .b(FE_OFN713_n_8140), .o(TIMEBOOST_net_4374) );
in01s01 g58140_u0 ( .a(FE_OFN516_n_9697), .o(g58140_sb) );
na02s01 TIMEBOOST_cell_37228 ( .a(TIMEBOOST_net_10852), .b(FE_OFN634_n_4454), .o(TIMEBOOST_net_9337) );
na02s01 TIMEBOOST_cell_15788 ( .a(parchk_pci_ad_reg_in_1210), .b(g67042_db), .o(TIMEBOOST_net_3151) );
na02s01 TIMEBOOST_cell_37230 ( .a(TIMEBOOST_net_10853), .b(FE_OFN622_n_4409), .o(TIMEBOOST_net_9334) );
in01s01 g58141_u0 ( .a(FE_OFN515_n_9697), .o(g58141_sb) );
na02s01 g58141_u1 ( .a(FE_OFN209_n_9126), .b(g58141_sb), .o(g58141_da) );
na02s01 g58141_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__Q), .b(FE_OFN515_n_9697), .o(g58141_db) );
na02s01 g58141_u3 ( .a(g58141_da), .b(g58141_db), .o(n_9070) );
in01s01 g58142_u0 ( .a(FE_OFN517_n_9697), .o(g58142_sb) );
na02s01 g58142_u1 ( .a(FE_OFN211_n_9858), .b(g58142_sb), .o(g58142_da) );
na02s01 g58142_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__Q), .b(FE_OFN517_n_9697), .o(g58142_db) );
na02s01 g58142_u3 ( .a(g58142_da), .b(g58142_db), .o(n_9653) );
in01s01 g58143_u0 ( .a(FE_OFN518_n_9697), .o(g58143_sb) );
na02f02 TIMEBOOST_cell_43783 ( .a(n_9138), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__Q), .o(TIMEBOOST_net_14130) );
na02s01 g58143_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__Q), .b(FE_OFN518_n_9697), .o(g58143_db) );
na02s02 TIMEBOOST_cell_38730 ( .a(TIMEBOOST_net_11603), .b(g53925_sb), .o(n_13520) );
in01s01 g58144_u0 ( .a(FE_OFN518_n_9697), .o(g58144_sb) );
na02f02 TIMEBOOST_cell_43784 ( .a(TIMEBOOST_net_14130), .b(FE_OFN1377_n_8567), .o(TIMEBOOST_net_12867) );
na02s01 g58144_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__Q), .b(FE_OFN518_n_9697), .o(g58144_db) );
na02f02 TIMEBOOST_cell_39116 ( .a(TIMEBOOST_net_11796), .b(FE_OFN1599_n_13995), .o(g53159_p) );
in01s01 g58145_u0 ( .a(FE_OFN517_n_9697), .o(g58145_sb) );
na02s01 g58145_u1 ( .a(FE_OFN217_n_9889), .b(g58145_sb), .o(g58145_da) );
na02s01 g58145_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__Q), .b(FE_OFN517_n_9697), .o(g58145_db) );
na02s01 g58145_u3 ( .a(g58145_da), .b(g58145_db), .o(n_9649) );
in01s01 g58146_u0 ( .a(FE_OFN517_n_9697), .o(g58146_sb) );
na02s01 g58146_u1 ( .a(FE_OFN219_n_9853), .b(g58146_sb), .o(g58146_da) );
na02s01 g58146_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__Q), .b(FE_OFN517_n_9697), .o(g58146_db) );
na02s01 g58146_u3 ( .a(g58146_da), .b(g58146_db), .o(n_9648) );
in01s01 g58147_u0 ( .a(FE_OFN517_n_9697), .o(g58147_sb) );
na02s01 TIMEBOOST_cell_37232 ( .a(TIMEBOOST_net_10854), .b(g58070_sb), .o(TIMEBOOST_net_349) );
na02s01 TIMEBOOST_cell_15789 ( .a(TIMEBOOST_net_3151), .b(g67042_sb), .o(n_1276) );
na02s01 TIMEBOOST_cell_37234 ( .a(TIMEBOOST_net_10855), .b(g58060_sb), .o(TIMEBOOST_net_9592) );
in01s01 g58148_u0 ( .a(FE_OFN517_n_9697), .o(g58148_sb) );
na02s01 TIMEBOOST_cell_37236 ( .a(TIMEBOOST_net_10856), .b(g65792_db), .o(n_1594) );
na02s01 TIMEBOOST_cell_15790 ( .a(parchk_pci_ad_reg_in_1225), .b(g67085_db), .o(TIMEBOOST_net_3152) );
na02f02 TIMEBOOST_cell_41032 ( .a(TIMEBOOST_net_12754), .b(g57087_sb), .o(n_11655) );
in01s01 g58149_u0 ( .a(FE_OFN519_n_9697), .o(g58149_sb) );
na03s04 TIMEBOOST_cell_45401 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__Q), .b(n_3719), .c(FE_OFN1317_n_6624), .o(TIMEBOOST_net_14939) );
na02s01 TIMEBOOST_cell_15791 ( .a(TIMEBOOST_net_3152), .b(g67042_sb), .o(n_1431) );
na03m02 TIMEBOOST_cell_1126 ( .a(g59350_db), .b(g59350_sb), .c(n_7115), .o(n_7701) );
in01s01 g58150_u0 ( .a(FE_OFN518_n_9697), .o(g58150_sb) );
na02s01 g58150_u1 ( .a(FE_OFN221_n_9846), .b(g58150_sb), .o(g58150_da) );
na02s01 g58150_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__Q), .b(FE_OFN518_n_9697), .o(g58150_db) );
na02s01 g58150_u3 ( .a(g58150_da), .b(g58150_db), .o(n_9642) );
na02s01 g58151_u1 ( .a(FE_OFN223_n_9844), .b(g58161_sb), .o(g58151_da) );
na02s01 g58151_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__Q), .b(FE_OFN515_n_9697), .o(g58151_db) );
na02s01 g58151_u3 ( .a(g58151_da), .b(g58151_db), .o(n_9640) );
in01s01 g58152_u0 ( .a(FE_OFN517_n_9697), .o(g58152_sb) );
na02s01 g58152_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__Q), .b(FE_OFN517_n_9697), .o(g58152_db) );
na02s02 TIMEBOOST_cell_39720 ( .a(TIMEBOOST_net_12098), .b(g62637_sb), .o(n_6276) );
in01s01 g58153_u0 ( .a(FE_OFN516_n_9697), .o(g58153_sb) );
na02s03 TIMEBOOST_cell_30760 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_4_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_7_), .o(TIMEBOOST_net_9291) );
na02s01 TIMEBOOST_cell_15796 ( .a(parchk_pci_ad_reg_in_1223), .b(g67049_db), .o(TIMEBOOST_net_3155) );
na02f02 TIMEBOOST_cell_41616 ( .a(FE_OFN1441_n_9372), .b(TIMEBOOST_net_13046), .o(TIMEBOOST_net_11675) );
in01s01 g58154_u0 ( .a(FE_OFN516_n_9697), .o(g58154_sb) );
na02s01 g58154_u1 ( .a(FE_OFN227_n_9841), .b(g58154_sb), .o(g58154_da) );
na02s01 g58154_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__Q), .b(FE_OFN516_n_9697), .o(g58154_db) );
na02s02 g58154_u3 ( .a(g58154_da), .b(g58154_db), .o(n_9637) );
na02s01 g58155_u1 ( .a(FE_OFN229_n_9120), .b(g58141_sb), .o(g58155_da) );
na02s01 g58155_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__Q), .b(FE_OFN517_n_9697), .o(g58155_db) );
na02s02 g58155_u3 ( .a(g58155_da), .b(g58155_db), .o(n_9067) );
in01s01 g58156_u0 ( .a(FE_OFN516_n_9697), .o(g58156_sb) );
na02s01 TIMEBOOST_cell_44926 ( .a(TIMEBOOST_net_14701), .b(g58013_db), .o(n_9102) );
na02s01 g58156_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__Q), .b(FE_OFN516_n_9697), .o(g58156_db) );
na02s02 TIMEBOOST_cell_39722 ( .a(TIMEBOOST_net_12099), .b(g62470_sb), .o(n_6651) );
na02s01 g58157_u1 ( .a(FE_OFN233_n_9876), .b(g58154_sb), .o(g58157_da) );
na02s01 g58157_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__Q), .b(FE_OFN516_n_9697), .o(g58157_db) );
na02s01 g58157_u3 ( .a(g58157_da), .b(g58157_db), .o(n_9633) );
in01s01 g58158_u0 ( .a(FE_OFN518_n_9697), .o(g58158_sb) );
na02m02 TIMEBOOST_cell_45141 ( .a(TIMEBOOST_net_511), .b(g53940_sb), .o(TIMEBOOST_net_14809) );
na02m02 TIMEBOOST_cell_32560 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__Q), .o(TIMEBOOST_net_10191) );
na02m08 TIMEBOOST_cell_30772 ( .a(n_2557), .b(wbs_stb_i), .o(TIMEBOOST_net_9297) );
in01s01 g58159_u0 ( .a(FE_OFN517_n_9697), .o(g58159_sb) );
na02s01 g58159_u1 ( .a(FE_OFN235_n_9834), .b(g58159_sb), .o(g58159_da) );
na02s01 g58159_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__29__Q), .b(FE_OFN517_n_9697), .o(g58159_db) );
na02s02 g58159_u3 ( .a(g58159_da), .b(g58159_db), .o(n_9629) );
in01s01 g58160_u0 ( .a(FE_OFN515_n_9697), .o(g58160_sb) );
na02s01 g58160_u1 ( .a(FE_OFN237_n_9118), .b(g58160_sb), .o(g58160_da) );
na02s01 g58160_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__Q), .b(FE_OFN515_n_9697), .o(g58160_db) );
na02s01 g58160_u3 ( .a(g58160_da), .b(g58160_db), .o(n_9066) );
in01s01 g58161_u0 ( .a(FE_OFN515_n_9697), .o(g58161_sb) );
na02s02 TIMEBOOST_cell_37708 ( .a(TIMEBOOST_net_11092), .b(g61785_sb), .o(n_8234) );
na02f02 TIMEBOOST_cell_41190 ( .a(TIMEBOOST_net_12833), .b(g57338_sb), .o(n_11414) );
na02s01 TIMEBOOST_cell_37710 ( .a(TIMEBOOST_net_11093), .b(g61745_sb), .o(n_8327) );
in01s01 g58162_u0 ( .a(FE_OFN518_n_9697), .o(g58162_sb) );
na02s01 g58162_u1 ( .a(FE_OFN241_n_9830), .b(g58162_sb), .o(g58162_da) );
na02s01 g58162_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__Q), .b(FE_OFN518_n_9697), .o(g58162_db) );
na02s01 g58162_u3 ( .a(g58162_da), .b(g58162_db), .o(n_9626) );
in01s01 g58163_u0 ( .a(FE_OFN517_n_9697), .o(g58163_sb) );
na02s01 TIMEBOOST_cell_30780 ( .a(pci_inti_conf_int_in), .b(pci_inta_oe_o), .o(TIMEBOOST_net_9301) );
na03s01 TIMEBOOST_cell_34287 ( .a(n_3935), .b(g63020_sb), .c(g63020_db), .o(n_5207) );
na02s04 TIMEBOOST_cell_45402 ( .a(TIMEBOOST_net_14939), .b(g62519_sb), .o(n_6538) );
in01s01 g58164_u0 ( .a(FE_OFN515_n_9697), .o(g58164_sb) );
na02s01 g58164_u1 ( .a(FE_OFN243_n_9116), .b(g58164_sb), .o(g58164_da) );
na02s01 g58164_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__Q), .b(FE_OFN515_n_9697), .o(g58164_db) );
na02s01 g58164_u3 ( .a(g58164_da), .b(g58164_db), .o(n_9065) );
in01s01 g58165_u0 ( .a(FE_OFN518_n_9697), .o(g58165_sb) );
na03s02 TIMEBOOST_cell_40475 ( .a(n_3974), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__16__Q), .c(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_12476) );
na02s01 g58165_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__Q), .b(FE_OFN518_n_9697), .o(g58165_db) );
na02s02 TIMEBOOST_cell_40476 ( .a(TIMEBOOST_net_12476), .b(g62842_sb), .o(n_5288) );
na02s01 TIMEBOOST_cell_9676 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__Q), .b(g58313_sb), .o(TIMEBOOST_net_1405) );
na02s01 g58166_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__Q), .b(FE_OFN517_n_9697), .o(g58166_db) );
na02s01 TIMEBOOST_cell_17661 ( .a(TIMEBOOST_net_4087), .b(g65305_db), .o(n_4275) );
in01s01 g58167_u0 ( .a(FE_OFN517_n_9697), .o(g58167_sb) );
na02s01 g58167_u1 ( .a(FE_OFN250_n_9789), .b(g58167_sb), .o(g58167_da) );
na02s01 g58167_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__Q), .b(FE_OFN517_n_9697), .o(g58167_db) );
na02s02 g58167_u3 ( .a(g58167_da), .b(g58167_db), .o(n_9624) );
na02f02 TIMEBOOST_cell_39118 ( .a(TIMEBOOST_net_11797), .b(FE_OFN1600_n_13995), .o(n_14459) );
na02s01 g58168_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__Q), .b(FE_OFN516_n_9697), .o(g58168_db) );
na03f04 TIMEBOOST_cell_37111 ( .a(n_10991), .b(n_10216), .c(n_10221), .o(TIMEBOOST_net_10794) );
in01s01 g58169_u0 ( .a(FE_OFN587_n_9692), .o(g58169_sb) );
na02f02 TIMEBOOST_cell_39111 ( .a(FE_OFN1605_n_13997), .b(TIMEBOOST_net_10173), .o(TIMEBOOST_net_11794) );
na02s01 g58169_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__Q), .b(FE_OFN587_n_9692), .o(g58169_db) );
na02f02 TIMEBOOST_cell_38948 ( .a(TIMEBOOST_net_11712), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10729) );
in01s01 g58170_u0 ( .a(FE_OFN588_n_9692), .o(g58170_sb) );
na03s03 TIMEBOOST_cell_45403 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__Q), .b(n_4906), .c(FE_OFN1320_n_6436), .o(TIMEBOOST_net_14940) );
na03s02 TIMEBOOST_cell_40477 ( .a(n_384), .b(FE_OFN1127_g64577_p), .c(n_4722), .o(TIMEBOOST_net_12477) );
na02s01 TIMEBOOST_cell_41800 ( .a(TIMEBOOST_net_13138), .b(g62027_sb), .o(n_7842) );
in01s01 g58171_u0 ( .a(FE_OFN584_n_9692), .o(g58171_sb) );
na02s01 TIMEBOOST_cell_43046 ( .a(TIMEBOOST_net_13761), .b(g63194_sb), .o(n_4798) );
na02s01 TIMEBOOST_cell_15876 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_100), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3195) );
na03s02 TIMEBOOST_cell_41801 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__Q), .b(FE_OFN702_n_7845), .c(n_1853), .o(TIMEBOOST_net_13139) );
in01s01 g58172_u0 ( .a(FE_OFN585_n_9692), .o(g58172_sb) );
na02s02 TIMEBOOST_cell_40478 ( .a(TIMEBOOST_net_12477), .b(g63044_sb), .o(n_7123) );
na02s01 g58172_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__Q), .b(FE_OFN585_n_9692), .o(g58172_db) );
na02s01 TIMEBOOST_cell_31804 ( .a(configuration_wb_err_data_576), .b(parchk_pci_ad_out_in_1173), .o(TIMEBOOST_net_9813) );
in01s01 g58173_u0 ( .a(FE_OFN588_n_9692), .o(g58173_sb) );
na02s01 g58173_u1 ( .a(FE_OFN211_n_9858), .b(g58173_sb), .o(g58173_da) );
na02s01 g58173_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__Q), .b(FE_OFN588_n_9692), .o(g58173_db) );
na02s01 g58173_u3 ( .a(g58173_da), .b(g58173_db), .o(n_9617) );
in01s01 g58174_u0 ( .a(FE_OFN589_n_9692), .o(g58174_sb) );
na02s01 TIMEBOOST_cell_17628 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__Q), .b(g64322_sb), .o(TIMEBOOST_net_4071) );
na02s01 g58174_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__Q), .b(FE_OFN589_n_9692), .o(g58174_db) );
na02f02 TIMEBOOST_cell_38991 ( .a(TIMEBOOST_net_10101), .b(FE_OFN2158_n_16439), .o(TIMEBOOST_net_11734) );
in01s01 g58175_u0 ( .a(FE_OFN589_n_9692), .o(g58175_sb) );
na02f02 TIMEBOOST_cell_39117 ( .a(TIMEBOOST_net_10167), .b(FE_OFN1606_n_13997), .o(TIMEBOOST_net_11797) );
na02s01 g58175_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__Q), .b(FE_OFN589_n_9692), .o(g58175_db) );
na02m02 TIMEBOOST_cell_38732 ( .a(TIMEBOOST_net_11604), .b(g59763_sb), .o(n_7625) );
in01s01 g58176_u0 ( .a(FE_OFN587_n_9692), .o(g58176_sb) );
na02s01 TIMEBOOST_cell_40487 ( .a(wishbone_slave_unit_pcim_sm_data_in_647), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__Q), .o(TIMEBOOST_net_12482) );
na02s01 g58176_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__Q), .b(FE_OFN587_n_9692), .o(g58176_db) );
na02s01 TIMEBOOST_cell_31747 ( .a(TIMEBOOST_net_9784), .b(g61912_db), .o(n_7997) );
in01s01 g58177_u0 ( .a(FE_OFN588_n_9692), .o(g58177_sb) );
na02f02 TIMEBOOST_cell_41683 ( .a(FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__Q), .o(TIMEBOOST_net_13080) );
na02s02 TIMEBOOST_cell_40862 ( .a(TIMEBOOST_net_12669), .b(FE_OFN1330_n_13547), .o(TIMEBOOST_net_11624) );
na02s01 TIMEBOOST_cell_41802 ( .a(TIMEBOOST_net_13139), .b(g61861_sb), .o(n_8116) );
in01s01 g58178_u0 ( .a(FE_OFN587_n_9692), .o(g58178_sb) );
na02f02 TIMEBOOST_cell_42254 ( .a(TIMEBOOST_net_13365), .b(FE_OFN1424_n_8567), .o(TIMEBOOST_net_12324) );
na02s02 TIMEBOOST_cell_40863 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__Q), .b(n_13165), .o(TIMEBOOST_net_12670) );
na03s02 TIMEBOOST_cell_41803 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__Q), .b(FE_OFN702_n_7845), .c(n_1836), .o(TIMEBOOST_net_13140) );
in01s01 g58179_u0 ( .a(FE_OFN587_n_9692), .o(g58179_sb) );
na03s02 TIMEBOOST_cell_43047 ( .a(n_8590), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q), .c(g59082_sb), .o(TIMEBOOST_net_13762) );
na02s02 TIMEBOOST_cell_40864 ( .a(TIMEBOOST_net_12670), .b(FE_OFN1331_n_13547), .o(TIMEBOOST_net_11616) );
na02f02 TIMEBOOST_cell_44732 ( .a(TIMEBOOST_net_14604), .b(n_12056), .o(n_12765) );
in01s01 g58180_u0 ( .a(FE_OFN588_n_9692), .o(g58180_sb) );
na02s01 TIMEBOOST_cell_44927 ( .a(FE_OFN247_n_9112), .b(g58160_sb), .o(TIMEBOOST_net_14702) );
na02s01 g58180_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__Q), .b(FE_OFN588_n_9692), .o(g58180_db) );
na02s01 TIMEBOOST_cell_39724 ( .a(TIMEBOOST_net_12100), .b(g62389_sb), .o(n_6821) );
in01s01 g58181_u0 ( .a(FE_OFN585_n_9692), .o(g58181_sb) );
na02s01 g58181_u1 ( .a(FE_OFN223_n_9844), .b(g58181_sb), .o(g58181_da) );
na02s01 g58181_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__Q), .b(FE_OFN587_n_9692), .o(g58181_db) );
na02s01 g58181_u3 ( .a(g58181_da), .b(g58181_db), .o(n_9605) );
in01s01 g58182_u0 ( .a(FE_OFN588_n_9692), .o(g58182_sb) );
no02f02 TIMEBOOST_cell_36946 ( .a(TIMEBOOST_net_10711), .b(TIMEBOOST_net_6240), .o(FE_RN_589_0) );
na02s01 g58182_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__Q), .b(FE_OFN588_n_9692), .o(g58182_db) );
na02m02 TIMEBOOST_cell_40480 ( .a(TIMEBOOST_net_12478), .b(TIMEBOOST_net_558), .o(n_13434) );
in01s01 g58183_u0 ( .a(FE_OFN584_n_9692), .o(g58183_sb) );
na02m02 TIMEBOOST_cell_40482 ( .a(TIMEBOOST_net_12479), .b(TIMEBOOST_net_562), .o(n_13429) );
na02s01 g58183_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__Q), .b(FE_OFN584_n_9692), .o(g58183_db) );
na02m02 TIMEBOOST_cell_40479 ( .a(g54177_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_397), .o(TIMEBOOST_net_12478) );
in01s01 g58184_u0 ( .a(FE_OFN585_n_9692), .o(g58184_sb) );
na02s01 TIMEBOOST_cell_40484 ( .a(TIMEBOOST_net_12480), .b(g58330_db), .o(n_9215) );
na02s01 g58184_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__Q), .b(FE_OFN585_n_9692), .o(g58184_db) );
na02s01 TIMEBOOST_cell_16212 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(g65777_sb), .o(TIMEBOOST_net_3363) );
in01s01 g58185_u0 ( .a(FE_OFN584_n_9692), .o(g58185_sb) );
na02s01 TIMEBOOST_cell_39217 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__Q), .b(n_8407), .o(TIMEBOOST_net_11847) );
na02s01 g58185_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__Q), .b(FE_OFN584_n_9692), .o(g58185_db) );
na02s01 TIMEBOOST_cell_39248 ( .a(TIMEBOOST_net_11862), .b(g64153_db), .o(n_4012) );
in01s01 g58186_u0 ( .a(FE_OFN584_n_9692), .o(g58186_sb) );
na02s01 TIMEBOOST_cell_36512 ( .a(TIMEBOOST_net_10494), .b(FE_OFN250_n_9789), .o(n_9727) );
na02s01 g58186_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__Q), .b(FE_OFN584_n_9692), .o(g58186_db) );
na02s01 TIMEBOOST_cell_36513 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__Q), .b(FE_OFN623_n_4409), .o(TIMEBOOST_net_10495) );
in01s01 g58187_u0 ( .a(FE_OFN589_n_9692), .o(g58187_sb) );
na02s02 TIMEBOOST_cell_40865 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__Q), .b(n_13174), .o(TIMEBOOST_net_12671) );
na03m02 TIMEBOOST_cell_40883 ( .a(TIMEBOOST_net_464), .b(g52650_da), .c(g52402_sb), .o(TIMEBOOST_net_12680) );
in01s01 g58188_u0 ( .a(FE_OFN588_n_9692), .o(g58188_sb) );
na02s01 TIMEBOOST_cell_43468 ( .a(TIMEBOOST_net_13972), .b(FE_OFN1233_n_6391), .o(TIMEBOOST_net_12205) );
na02s01 g58188_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q), .b(FE_OFN588_n_9692), .o(g58188_db) );
na02s02 TIMEBOOST_cell_38198 ( .a(TIMEBOOST_net_11337), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_4623) );
in01s01 g58189_u0 ( .a(FE_OFN587_n_9692), .o(g58189_sb) );
na02s01 TIMEBOOST_cell_16213 ( .a(TIMEBOOST_net_3363), .b(g65777_db), .o(n_1601) );
na02s01 g58189_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__Q), .b(FE_OFN585_n_9692), .o(g58189_db) );
na02s01 TIMEBOOST_cell_45090 ( .a(TIMEBOOST_net_14783), .b(g57947_db), .o(n_9863) );
in01s01 g58190_u0 ( .a(FE_OFN585_n_9692), .o(g58190_sb) );
na02s01 TIMEBOOST_cell_36514 ( .a(TIMEBOOST_net_10495), .b(g64904_sb), .o(TIMEBOOST_net_9604) );
na02s01 TIMEBOOST_cell_36780 ( .a(TIMEBOOST_net_10628), .b(FE_OFN1126_g64577_p), .o(TIMEBOOST_net_4505) );
na02f01 TIMEBOOST_cell_36515 ( .a(TIMEBOOST_net_1211), .b(n_2795), .o(TIMEBOOST_net_10496) );
in01s01 g58191_u0 ( .a(FE_OFN589_n_9692), .o(g58191_sb) );
na02f02 TIMEBOOST_cell_43785 ( .a(TIMEBOOST_net_10044), .b(g57123_sb), .o(TIMEBOOST_net_14131) );
na02s01 g58191_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__Q), .b(FE_OFN589_n_9692), .o(g58191_db) );
na02s01 TIMEBOOST_cell_38734 ( .a(TIMEBOOST_net_11605), .b(g53898_sb), .o(n_13550) );
in01s01 g58192_u0 ( .a(FE_OFN587_n_9692), .o(g58192_sb) );
na02s01 TIMEBOOST_cell_43574 ( .a(TIMEBOOST_net_14025), .b(n_6431), .o(TIMEBOOST_net_12153) );
na02m02 TIMEBOOST_cell_40866 ( .a(TIMEBOOST_net_12671), .b(FE_OFN1331_n_13547), .o(TIMEBOOST_net_11610) );
na02s01 TIMEBOOST_cell_41730 ( .a(TIMEBOOST_net_13103), .b(g57896_db), .o(n_9139) );
in01s01 g58193_u0 ( .a(FE_OFN589_n_9692), .o(g58193_sb) );
na02s01 g58193_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__Q), .b(FE_OFN589_n_9692), .o(g58193_db) );
na02s01 TIMEBOOST_cell_16251 ( .a(TIMEBOOST_net_3382), .b(g64781_db), .o(n_3769) );
in01s01 g58194_u0 ( .a(FE_OFN585_n_9692), .o(g58194_sb) );
na02m06 TIMEBOOST_cell_17634 ( .a(pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_77), .b(n_532), .o(TIMEBOOST_net_4074) );
na02s01 g58194_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__Q), .b(FE_OFN585_n_9692), .o(g58194_db) );
na02f06 TIMEBOOST_cell_17635 ( .a(TIMEBOOST_net_4074), .b(FE_OFN2125_n_16497), .o(TIMEBOOST_net_573) );
in01s01 g58195_u0 ( .a(FE_OFN585_n_9692), .o(g58195_sb) );
na02s02 TIMEBOOST_cell_16252 ( .a(n_3755), .b(g64782_sb), .o(TIMEBOOST_net_3383) );
na02s01 g58195_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__Q), .b(FE_OFN585_n_9692), .o(g58195_db) );
na02s01 TIMEBOOST_cell_16253 ( .a(TIMEBOOST_net_3383), .b(g64782_db), .o(n_3768) );
in01s01 g58196_u0 ( .a(FE_OFN587_n_9692), .o(g58196_sb) );
na02s01 g58196_u1 ( .a(FE_OFN252_n_9868), .b(g58196_sb), .o(g58196_da) );
na02s01 g58196_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__Q), .b(FE_OFN589_n_9692), .o(g58196_db) );
na02s01 g58196_u3 ( .a(g58196_da), .b(g58196_db), .o(n_9590) );
in01s01 g58197_u0 ( .a(FE_OFN584_n_9692), .o(g58197_sb) );
na02s01 TIMEBOOST_cell_17636 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__Q), .b(g64236_sb), .o(TIMEBOOST_net_4075) );
na02s01 g58197_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__Q), .b(FE_OFN584_n_9692), .o(g58197_db) );
na02s01 TIMEBOOST_cell_37238 ( .a(TIMEBOOST_net_10857), .b(g65806_db), .o(n_1589) );
in01s01 g58198_u0 ( .a(FE_OFN595_n_9694), .o(g58198_sb) );
na02s01 g58198_u1 ( .a(FE_OFN207_n_9865), .b(g58198_sb), .o(g58198_da) );
na02s01 g58198_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__Q), .b(FE_OFN595_n_9694), .o(g58198_db) );
na02s01 g58198_u3 ( .a(g58198_da), .b(g58198_db), .o(n_9588) );
in01s01 g58199_u0 ( .a(FE_OFN596_n_9694), .o(g58199_sb) );
na02s01 TIMEBOOST_cell_43064 ( .a(TIMEBOOST_net_13770), .b(FE_OFN1219_n_6886), .o(TIMEBOOST_net_12023) );
na02s01 TIMEBOOST_cell_40486 ( .a(TIMEBOOST_net_12481), .b(FE_OFN1300_n_5763), .o(TIMEBOOST_net_11520) );
na02f01 TIMEBOOST_cell_36516 ( .a(TIMEBOOST_net_10496), .b(n_2778), .o(n_3281) );
in01s01 g58200_u0 ( .a(FE_OFN592_n_9694), .o(g58200_sb) );
na02f02 TIMEBOOST_cell_44748 ( .a(TIMEBOOST_net_14612), .b(n_12389), .o(n_12702) );
na02s01 TIMEBOOST_cell_40483 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__Q), .b(g58330_sb), .o(TIMEBOOST_net_12480) );
na02s01 TIMEBOOST_cell_43065 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__Q), .b(n_3558), .o(TIMEBOOST_net_13771) );
in01s01 g58201_u0 ( .a(FE_OFN593_n_9694), .o(g58201_sb) );
na02s01 g58201_u1 ( .a(FE_OFN209_n_9126), .b(g58201_sb), .o(g58201_da) );
na02s01 g58201_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__Q), .b(FE_OFN593_n_9694), .o(g58201_db) );
na02s01 g58201_u3 ( .a(g58201_da), .b(g58201_db), .o(n_9055) );
in01s01 g58202_u0 ( .a(FE_OFN596_n_9694), .o(g58202_sb) );
na02s01 g58202_u1 ( .a(FE_OFN211_n_9858), .b(g58202_sb), .o(g58202_da) );
na02s01 g58202_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__Q), .b(FE_OFN596_n_9694), .o(g58202_db) );
na02s01 g58202_u3 ( .a(g58202_da), .b(g58202_db), .o(n_9584) );
in01s01 g58203_u0 ( .a(FE_OFN597_n_9694), .o(g58203_sb) );
na02s01 TIMEBOOST_cell_17638 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__Q), .b(g64258_sb), .o(TIMEBOOST_net_4076) );
na02s01 g58203_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__Q), .b(FE_OFN597_n_9694), .o(g58203_db) );
in01s01 g58204_u0 ( .a(FE_OFN597_n_9694), .o(g58204_sb) );
na02f02 TIMEBOOST_cell_43786 ( .a(TIMEBOOST_net_14131), .b(FE_OFN1414_n_8567), .o(n_11623) );
na02s01 g58204_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__Q), .b(FE_OFN597_n_9694), .o(g58204_db) );
na02s02 TIMEBOOST_cell_38736 ( .a(TIMEBOOST_net_11606), .b(g53931_sb), .o(n_13514) );
in01s01 g58205_u0 ( .a(FE_OFN592_n_9694), .o(g58205_sb) );
na02s01 g58205_u1 ( .a(FE_OFN219_n_9853), .b(g58205_sb), .o(g58205_da) );
na02s01 g58205_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__Q), .b(FE_OFN592_n_9694), .o(g58205_db) );
na02s01 g58205_u3 ( .a(g58205_da), .b(g58205_db), .o(n_9582) );
in01s01 g58206_u0 ( .a(FE_OFN596_n_9694), .o(g58206_sb) );
na02f02 TIMEBOOST_cell_42282 ( .a(TIMEBOOST_net_13379), .b(g57343_sb), .o(n_11406) );
na02f02 TIMEBOOST_cell_42506 ( .a(TIMEBOOST_net_13491), .b(g57561_sb), .o(n_11191) );
na03f06 TIMEBOOST_cell_41673 ( .a(n_10575), .b(n_10572), .c(n_9988), .o(TIMEBOOST_net_13075) );
in01s01 g58207_u0 ( .a(FE_OFN595_n_9694), .o(g58207_sb) );
na03s02 TIMEBOOST_cell_43299 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__Q), .b(n_3516), .c(FE_OFN1219_n_6886), .o(TIMEBOOST_net_13888) );
na02s01 g58207_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__Q), .b(FE_OFN595_n_9694), .o(g58207_db) );
na02m02 TIMEBOOST_cell_45803 ( .a(n_9707), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__Q), .o(TIMEBOOST_net_15140) );
in01s01 g58208_u0 ( .a(FE_OFN595_n_9694), .o(g58208_sb) );
na03f06 TIMEBOOST_cell_33474 ( .a(FE_RN_535_0), .b(n_16474), .c(FE_RN_360_0), .o(n_16268) );
na02s01 g58208_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__Q), .b(FE_OFN595_n_9694), .o(g58208_db) );
na02s01 TIMEBOOST_cell_37712 ( .a(TIMEBOOST_net_11094), .b(g61819_sb), .o(n_8152) );
in01s01 g58209_u0 ( .a(FE_OFN597_n_9694), .o(g58209_sb) );
na02s01 g58209_u1 ( .a(FE_OFN221_n_9846), .b(g58209_sb), .o(g58209_da) );
na02s01 g58209_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__Q), .b(FE_OFN597_n_9694), .o(g58209_db) );
na02s01 g58209_u3 ( .a(g58209_da), .b(g58209_db), .o(n_9576) );
in01s01 g58210_u0 ( .a(FE_OFN595_n_9694), .o(g58210_sb) );
na02s01 TIMEBOOST_cell_40491 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__Q), .b(wishbone_slave_unit_pcim_sm_data_in_655), .o(TIMEBOOST_net_12484) );
na02s01 g58210_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN595_n_9694), .o(g58210_db) );
na02s01 TIMEBOOST_cell_40488 ( .a(TIMEBOOST_net_12482), .b(FE_OFN1301_n_5763), .o(TIMEBOOST_net_11521) );
in01s01 g58211_u0 ( .a(FE_OFN596_n_9694), .o(g58211_sb) );
na02s01 g58211_u1 ( .a(FE_OFN225_n_9122), .b(g58211_sb), .o(g58211_da) );
na02s01 g58211_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q), .b(FE_OFN596_n_9694), .o(g58211_db) );
na02f02 TIMEBOOST_cell_37140 ( .a(TIMEBOOST_net_10808), .b(n_12570), .o(n_12832) );
in01s01 g58212_u0 ( .a(FE_OFN592_n_9694), .o(g58212_sb) );
na02s01 TIMEBOOST_cell_37714 ( .a(TIMEBOOST_net_11095), .b(g61711_sb), .o(n_8404) );
na02s02 TIMEBOOST_cell_43233 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__Q), .b(n_4496), .o(TIMEBOOST_net_13855) );
na02s02 TIMEBOOST_cell_39472 ( .a(TIMEBOOST_net_11974), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_4688) );
in01s01 g58213_u0 ( .a(FE_OFN592_n_9694), .o(g58213_sb) );
na02s01 g58213_u1 ( .a(FE_OFN227_n_9841), .b(g58213_sb), .o(g58213_da) );
na02s01 g58213_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__Q), .b(FE_OFN592_n_9694), .o(g58213_db) );
na02s02 g58213_u3 ( .a(g58213_da), .b(g58213_db), .o(n_9572) );
in01s01 g58214_u0 ( .a(FE_OFN593_n_9694), .o(g58214_sb) );
na02s01 g58214_u1 ( .a(FE_OFN229_n_9120), .b(g58214_sb), .o(g58214_da) );
na02s01 g58214_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__Q), .b(FE_OFN593_n_9694), .o(g58214_db) );
na02s02 g58214_u3 ( .a(g58214_da), .b(g58214_db), .o(n_9052) );
in01s01 g58215_u0 ( .a(FE_OFN596_n_9694), .o(g58215_sb) );
na02m02 TIMEBOOST_cell_43787 ( .a(n_9550), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__Q), .o(TIMEBOOST_net_14132) );
na02s01 g58215_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__Q), .b(FE_OFN596_n_9694), .o(g58215_db) );
na02s02 TIMEBOOST_cell_38738 ( .a(TIMEBOOST_net_11607), .b(g53929_sb), .o(n_13516) );
in01s01 g58216_u0 ( .a(FE_OFN596_n_9694), .o(g58216_sb) );
na02s01 g58216_u1 ( .a(FE_OFN233_n_9876), .b(g58216_sb), .o(g58216_da) );
na02s01 g58216_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__Q), .b(FE_OFN596_n_9694), .o(g58216_db) );
na02s01 g58216_u3 ( .a(g58216_da), .b(g58216_db), .o(n_9570) );
in01s01 g58217_u0 ( .a(FE_OFN597_n_9694), .o(g58217_sb) );
na02s01 TIMEBOOST_cell_37716 ( .a(TIMEBOOST_net_11096), .b(g61998_sb), .o(n_7899) );
na02s01 TIMEBOOST_cell_40489 ( .a(wishbone_slave_unit_pcim_sm_data_in_661), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__Q), .o(TIMEBOOST_net_12483) );
na02f02 TIMEBOOST_cell_37117 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_10161), .o(TIMEBOOST_net_10797) );
in01s01 g58218_u0 ( .a(FE_OFN596_n_9694), .o(g58218_sb) );
na02s01 g58218_u1 ( .a(FE_OFN235_n_9834), .b(g58218_sb), .o(g58218_da) );
na02s01 g58218_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__Q), .b(FE_OFN596_n_9694), .o(g58218_db) );
na02s02 g58218_u3 ( .a(g58218_da), .b(g58218_db), .o(n_9568) );
in01s01 g58219_u0 ( .a(FE_OFN595_n_9694), .o(g58219_sb) );
na02s01 g58219_u1 ( .a(FE_OFN237_n_9118), .b(g58219_sb), .o(g58219_da) );
na02s01 g58219_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__Q), .b(FE_OFN595_n_9694), .o(g58219_db) );
na02s01 g58219_u3 ( .a(g58219_da), .b(g58219_db), .o(n_9051) );
in01s01 g58220_u0 ( .a(FE_OFN595_n_9694), .o(g58220_sb) );
na02s01 g58220_u1 ( .a(FE_OFN239_n_9832), .b(g58220_sb), .o(g58220_da) );
na02s01 g58220_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__Q), .b(FE_OFN595_n_9694), .o(g58220_db) );
na02s01 g58220_u3 ( .a(g58220_da), .b(g58220_db), .o(n_9567) );
in01s01 g58221_u0 ( .a(FE_OFN597_n_9694), .o(g58221_sb) );
na02s01 g58221_u1 ( .a(FE_OFN241_n_9830), .b(g58221_sb), .o(g58221_da) );
na02s01 g58221_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__Q), .b(FE_OFN597_n_9694), .o(g58221_db) );
na02s01 g58221_u3 ( .a(g58221_da), .b(g58221_db), .o(n_9565) );
in01s01 g58222_u0 ( .a(FE_OFN592_n_9694), .o(g58222_sb) );
na02s01 TIMEBOOST_cell_37718 ( .a(TIMEBOOST_net_11097), .b(g61719_sb), .o(n_8387) );
na02s01 TIMEBOOST_cell_40867 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__Q), .b(n_13325), .o(TIMEBOOST_net_12672) );
na02s01 TIMEBOOST_cell_37239 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(g65794_sb), .o(TIMEBOOST_net_10858) );
in01s01 g58223_u0 ( .a(FE_OFN595_n_9694), .o(g58223_sb) );
na02s01 g58223_u1 ( .a(FE_OFN243_n_9116), .b(g58223_sb), .o(g58223_da) );
na02s01 g58223_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__Q), .b(FE_OFN595_n_9694), .o(g58223_db) );
na02s01 g58223_u3 ( .a(g58223_da), .b(g58223_db), .o(n_9050) );
in01s01 g58224_u0 ( .a(FE_OFN597_n_9694), .o(g58224_sb) );
na02s01 TIMEBOOST_cell_16098 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__Q), .b(pci_target_unit_fifos_pciw_control_in_156), .o(TIMEBOOST_net_3306) );
na02s01 g58224_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__Q), .b(FE_OFN597_n_9694), .o(g58224_db) );
na02s01 TIMEBOOST_cell_16099 ( .a(TIMEBOOST_net_3306), .b(FE_OFN903_n_4736), .o(TIMEBOOST_net_1240) );
in01s01 g58225_u0 ( .a(FE_OFN593_n_9694), .o(g58225_sb) );
na02f02 TIMEBOOST_cell_44312 ( .a(TIMEBOOST_net_14394), .b(FE_OFN1421_n_8567), .o(TIMEBOOST_net_12685) );
na02s01 g58225_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q), .b(FE_OFN593_n_9694), .o(g58225_db) );
na02f02 TIMEBOOST_cell_37123 ( .a(n_13997), .b(TIMEBOOST_net_6244), .o(TIMEBOOST_net_10800) );
na02s01 g58226_u1 ( .a(FE_OFN250_n_9789), .b(g58214_sb), .o(g58226_da) );
na02s01 g58226_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__Q), .b(FE_OFN593_n_9694), .o(g58226_db) );
na02s02 g58226_u3 ( .a(g58226_da), .b(g58226_db), .o(n_9563) );
in01s01 g58227_u0 ( .a(FE_OFN595_n_9694), .o(g58227_sb) );
na02s02 TIMEBOOST_cell_39726 ( .a(TIMEBOOST_net_12101), .b(g62930_sb), .o(n_6021) );
na02s01 g58227_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q), .b(FE_OFN595_n_9694), .o(g58227_db) );
na02s02 TIMEBOOST_cell_37185 ( .a(g57797_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_1_), .o(TIMEBOOST_net_10831) );
in01s01 g58228_u0 ( .a(FE_OFN592_n_9694), .o(g58228_sb) );
na02s01 TIMEBOOST_cell_44928 ( .a(TIMEBOOST_net_14702), .b(g58166_db), .o(n_9063) );
na02s01 g58228_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__Q), .b(FE_OFN592_n_9694), .o(g58228_db) );
na02s01 TIMEBOOST_cell_39728 ( .a(TIMEBOOST_net_12102), .b(g62467_sb), .o(n_6659) );
in01s01 g58229_u0 ( .a(FE_OFN540_n_9690), .o(g58229_sb) );
na02s01 TIMEBOOST_cell_37720 ( .a(TIMEBOOST_net_11098), .b(g61728_sb), .o(n_8364) );
na02s02 TIMEBOOST_cell_40868 ( .a(TIMEBOOST_net_12672), .b(FE_OFN1330_n_13547), .o(TIMEBOOST_net_11615) );
na02s02 TIMEBOOST_cell_39474 ( .a(TIMEBOOST_net_11975), .b(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_4532) );
in01s01 g58230_u0 ( .a(FE_OFN539_n_9690), .o(g58230_sb) );
na02s01 TIMEBOOST_cell_40271 ( .a(n_3741), .b(g65047_db), .o(TIMEBOOST_net_12374) );
na02s01 g58230_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__Q), .b(FE_OFN539_n_9690), .o(g58230_db) );
na02s02 TIMEBOOST_cell_39730 ( .a(TIMEBOOST_net_12103), .b(g62521_sb), .o(n_6534) );
in01s01 g58231_u0 ( .a(FE_OFN1801_n_9690), .o(g58231_sb) );
na02s01 TIMEBOOST_cell_40331 ( .a(n_36), .b(FE_OFN620_n_4490), .o(TIMEBOOST_net_12404) );
na02s01 TIMEBOOST_cell_18022 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(g63538_sb), .o(TIMEBOOST_net_4268) );
na02s02 TIMEBOOST_cell_39732 ( .a(TIMEBOOST_net_12104), .b(g62499_sb), .o(n_6585) );
in01s01 g58232_u0 ( .a(FE_OFN540_n_9690), .o(g58232_sb) );
na02s01 g58232_u1 ( .a(FE_OFN211_n_9858), .b(g58232_sb), .o(g58232_da) );
na02s01 g58232_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__Q), .b(FE_OFN540_n_9690), .o(g58232_db) );
na02s01 g58232_u3 ( .a(g58232_da), .b(g58232_db), .o(n_9558) );
in01s01 g58233_u0 ( .a(FE_OFN543_n_9690), .o(g58233_sb) );
na02s01 TIMEBOOST_cell_17270 ( .a(n_3755), .b(FE_OFN651_n_4508), .o(TIMEBOOST_net_3892) );
na02s01 g58233_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__Q), .b(FE_OFN543_n_9690), .o(g58233_db) );
na02s01 TIMEBOOST_cell_17271 ( .a(TIMEBOOST_net_3892), .b(g65341_da), .o(n_3547) );
in01s01 g58234_u0 ( .a(FE_OFN543_n_9690), .o(g58234_sb) );
na02s01 g58234_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__Q), .b(FE_OFN543_n_9690), .o(g58234_db) );
na02s02 TIMEBOOST_cell_39734 ( .a(TIMEBOOST_net_12105), .b(g63190_sb), .o(n_5774) );
in01s01 g58235_u0 ( .a(FE_OFN1800_n_9690), .o(g58235_sb) );
na02s01 TIMEBOOST_cell_19885 ( .a(TIMEBOOST_net_5199), .b(g63163_sb), .o(n_5810) );
na02s01 TIMEBOOST_cell_18024 ( .a(pci_target_unit_fifos_pciw_addr_data_in_123), .b(g64094_sb), .o(TIMEBOOST_net_4269) );
na02f02 TIMEBOOST_cell_38950 ( .a(TIMEBOOST_net_11713), .b(FE_OFN2157_n_16439), .o(TIMEBOOST_net_10724) );
in01s01 g58236_u0 ( .a(FE_OFN540_n_9690), .o(g58236_sb) );
na02s01 TIMEBOOST_cell_31762 ( .a(configuration_wb_err_addr_543), .b(conf_wb_err_addr_in_952), .o(TIMEBOOST_net_9792) );
na02s01 g58236_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__Q), .b(FE_OFN540_n_9690), .o(g58236_db) );
na02s01 TIMEBOOST_cell_16256 ( .a(n_3783), .b(g64785_sb), .o(TIMEBOOST_net_3385) );
in01s01 g58237_u0 ( .a(FE_OFN542_n_9690), .o(g58237_sb) );
na02s02 TIMEBOOST_cell_37722 ( .a(TIMEBOOST_net_11099), .b(g61724_sb), .o(n_8373) );
na03s02 TIMEBOOST_cell_40629 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__Q), .b(n_3587), .c(FE_OFN1242_n_4092), .o(TIMEBOOST_net_12553) );
na02s01 TIMEBOOST_cell_37724 ( .a(TIMEBOOST_net_11100), .b(g61721_sb), .o(n_8382) );
in01s01 g58238_u0 ( .a(FE_OFN542_n_9690), .o(g58238_sb) );
na02m02 TIMEBOOST_cell_36673 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_794), .b(n_12595), .o(TIMEBOOST_net_10575) );
na02f02 TIMEBOOST_cell_40889 ( .a(n_8560), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__Q), .o(TIMEBOOST_net_12683) );
na02s03 TIMEBOOST_cell_45404 ( .a(TIMEBOOST_net_14940), .b(g62576_sb), .o(n_7377) );
in01s01 g58239_u0 ( .a(FE_OFN539_n_9690), .o(g58239_sb) );
na02f02 TIMEBOOST_cell_42284 ( .a(TIMEBOOST_net_13380), .b(g57425_sb), .o(n_10361) );
na02s02 TIMEBOOST_cell_40628 ( .a(TIMEBOOST_net_12552), .b(g62658_sb), .o(n_6228) );
na02s02 TIMEBOOST_cell_45405 ( .a(TIMEBOOST_net_5439), .b(FE_OFN1312_n_6624), .o(TIMEBOOST_net_14941) );
in01s01 g58240_u0 ( .a(FE_OFN1801_n_9690), .o(g58240_sb) );
na02s02 TIMEBOOST_cell_39736 ( .a(TIMEBOOST_net_12106), .b(g62505_sb), .o(n_6569) );
na02f02 TIMEBOOST_cell_44376 ( .a(TIMEBOOST_net_14426), .b(FE_OFN1412_n_8567), .o(TIMEBOOST_net_12721) );
na02s01 TIMEBOOST_cell_18559 ( .a(TIMEBOOST_net_4536), .b(g63188_sb), .o(n_4943) );
na02s01 g58241_u1 ( .a(FE_OFN221_n_9846), .b(g58237_sb), .o(g58241_da) );
na02s01 g58241_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__Q), .b(FE_OFN542_n_9690), .o(g58241_db) );
na02s01 g58241_u3 ( .a(g58241_da), .b(g58241_db), .o(n_9550) );
in01s01 g58242_u0 ( .a(FE_OFN1802_n_9690), .o(g58242_sb) );
na02m02 TIMEBOOST_cell_38951 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_1__Q), .o(TIMEBOOST_net_11714) );
na02s02 TIMEBOOST_cell_18026 ( .a(pci_target_unit_fifos_pciw_addr_data_in_142), .b(g64211_sb), .o(TIMEBOOST_net_4270) );
na02f02 TIMEBOOST_cell_39120 ( .a(TIMEBOOST_net_11798), .b(FE_OFN1602_n_13995), .o(n_14439) );
in01s01 g58243_u0 ( .a(FE_OFN542_n_9690), .o(g58243_sb) );
na02s01 g58243_u1 ( .a(FE_OFN225_n_9122), .b(g58243_sb), .o(g58243_da) );
na02s01 g58243_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__Q), .b(FE_OFN542_n_9690), .o(g58243_db) );
na02s01 g58243_u3 ( .a(g58243_da), .b(g58243_db), .o(n_9045) );
in01s01 g58244_u0 ( .a(FE_OFN540_n_9690), .o(g58244_sb) );
na02m02 TIMEBOOST_cell_40891 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__Q), .b(n_9022), .o(TIMEBOOST_net_12684) );
na02s01 TIMEBOOST_cell_15857 ( .a(TIMEBOOST_net_3185), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_386), .o(TIMEBOOST_net_83) );
na02m02 TIMEBOOST_cell_32538 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__Q), .o(TIMEBOOST_net_10180) );
na02s02 TIMEBOOST_cell_37540 ( .a(TIMEBOOST_net_11008), .b(FE_OFN2084_n_8407), .o(TIMEBOOST_net_4163) );
na02s01 g58245_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__Q), .b(FE_OFN540_n_9690), .o(g58245_db) );
na02s01 TIMEBOOST_cell_40341 ( .a(n_3774), .b(g64999_db), .o(TIMEBOOST_net_12409) );
na02s01 TIMEBOOST_cell_16258 ( .a(n_3749), .b(g64809_sb), .o(TIMEBOOST_net_3386) );
na02s01 g58246_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__Q), .b(FE_OFN539_n_9690), .o(g58246_db) );
na02s01 TIMEBOOST_cell_16259 ( .a(TIMEBOOST_net_3386), .b(g64809_db), .o(n_3750) );
na02f02 TIMEBOOST_cell_44448 ( .a(TIMEBOOST_net_14462), .b(g58590_sb), .o(n_8910) );
na02s01 g58247_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__Q), .b(FE_OFN540_n_9690), .o(g58247_db) );
na02s02 TIMEBOOST_cell_39738 ( .a(TIMEBOOST_net_12107), .b(g62443_sb), .o(n_6709) );
na02s01 g58248_u1 ( .a(FE_OFN233_n_9876), .b(g58238_sb), .o(g58248_da) );
na02s01 g58248_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__Q), .b(FE_OFN542_n_9690), .o(g58248_db) );
na02s01 g58248_u3 ( .a(g58248_da), .b(g58248_db), .o(n_9545) );
na02s01 TIMEBOOST_cell_30748 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .o(TIMEBOOST_net_9285) );
na02s01 TIMEBOOST_cell_40490 ( .a(TIMEBOOST_net_12483), .b(FE_OFN1301_n_5763), .o(TIMEBOOST_net_11522) );
na02s01 TIMEBOOST_cell_37240 ( .a(TIMEBOOST_net_10858), .b(g65794_db), .o(n_1663) );
na02s01 g58250_u1 ( .a(FE_OFN235_n_9834), .b(g58243_sb), .o(g58250_da) );
na02s01 g58250_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__Q), .b(FE_OFN542_n_9690), .o(g58250_db) );
na02s02 g58250_u3 ( .a(g58250_da), .b(g58250_db), .o(n_9543) );
in01s01 g58251_u0 ( .a(FE_OFN541_n_9690), .o(g58251_sb) );
na02s01 TIMEBOOST_cell_40439 ( .a(parchk_pci_ad_out_in_1184), .b(configuration_wb_err_data_587), .o(TIMEBOOST_net_12458) );
na02f02 TIMEBOOST_cell_38911 ( .a(n_3167), .b(wbu_addr_in_270), .o(TIMEBOOST_net_11694) );
na02s01 TIMEBOOST_cell_40492 ( .a(TIMEBOOST_net_12484), .b(FE_OFN1299_n_5763), .o(TIMEBOOST_net_11514) );
in01s01 g58252_u0 ( .a(FE_OFN543_n_9690), .o(g58252_sb) );
na02s01 g58252_u1 ( .a(FE_OFN241_n_9830), .b(g58252_sb), .o(g58252_da) );
na02s01 g58252_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__Q), .b(FE_OFN543_n_9690), .o(g58252_db) );
na02s01 g58252_u3 ( .a(g58252_da), .b(g58252_db), .o(n_9542) );
na02s02 TIMEBOOST_cell_19361 ( .a(TIMEBOOST_net_4937), .b(g60618_sb), .o(n_4836) );
na02s01 TIMEBOOST_cell_15877 ( .a(TIMEBOOST_net_3195), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_413), .o(TIMEBOOST_net_74) );
na02s02 TIMEBOOST_cell_39440 ( .a(TIMEBOOST_net_11958), .b(TIMEBOOST_net_4257), .o(TIMEBOOST_net_4607) );
in01s01 g58254_u0 ( .a(FE_OFN1803_n_9690), .o(g58254_sb) );
na03s02 TIMEBOOST_cell_38199 ( .a(TIMEBOOST_net_3684), .b(g64287_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__Q), .o(TIMEBOOST_net_11338) );
na02s01 TIMEBOOST_cell_18028 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(g64109_sb), .o(TIMEBOOST_net_4271) );
na02s02 TIMEBOOST_cell_39740 ( .a(TIMEBOOST_net_12108), .b(g62482_sb), .o(n_6623) );
in01s01 g58255_u0 ( .a(FE_OFN543_n_9690), .o(g58255_sb) );
na02s01 TIMEBOOST_cell_31760 ( .a(configuration_wb_err_data_599), .b(parchk_pci_ad_out_in_1196), .o(TIMEBOOST_net_9791) );
na02s01 g58255_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__Q), .b(FE_OFN543_n_9690), .o(g58255_db) );
na02s02 TIMEBOOST_cell_37542 ( .a(TIMEBOOST_net_11009), .b(FE_OFN704_n_8069), .o(TIMEBOOST_net_4130) );
in01s01 g58256_u0 ( .a(FE_OFN539_n_9690), .o(g58256_sb) );
na02s02 TIMEBOOST_cell_42130 ( .a(TIMEBOOST_net_13303), .b(g62917_sb), .o(n_6045) );
na02s01 g58256_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__Q), .b(FE_OFN539_n_9690), .o(g58256_db) );
na02s01 TIMEBOOST_cell_39292 ( .a(TIMEBOOST_net_11884), .b(g65735_db), .o(n_1608) );
in01s01 g58257_u0 ( .a(FE_OFN539_n_9690), .o(g58257_sb) );
na02s01 TIMEBOOST_cell_31758 ( .a(configuration_wb_err_data_573), .b(parchk_pci_ad_out_in_1170), .o(TIMEBOOST_net_9790) );
na02s01 g58257_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__Q), .b(FE_OFN539_n_9690), .o(g58257_db) );
na02s01 TIMEBOOST_cell_16260 ( .a(n_3780), .b(g65099_sb), .o(TIMEBOOST_net_3387) );
in01s01 g58258_u0 ( .a(FE_OFN1801_n_9690), .o(g58258_sb) );
na03s02 TIMEBOOST_cell_38399 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__Q), .b(FE_OFN1137_g64577_p), .c(n_3887), .o(TIMEBOOST_net_11438) );
na02s02 TIMEBOOST_cell_18030 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(g60675_sb), .o(TIMEBOOST_net_4272) );
na02s01 TIMEBOOST_cell_39742 ( .a(TIMEBOOST_net_12109), .b(g62597_sb), .o(n_6358) );
na02s01 TIMEBOOST_cell_9716 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__Q), .b(g63567_sb), .o(TIMEBOOST_net_1425) );
na02s01 g58259_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__Q), .b(FE_OFN540_n_9690), .o(g58259_db) );
na02s01 TIMEBOOST_cell_9717 ( .a(TIMEBOOST_net_1425), .b(g63567_db), .o(n_4595) );
in01s01 g58260_u0 ( .a(FE_OFN584_n_9692), .o(g58260_sb) );
na03s02 TIMEBOOST_cell_33406 ( .a(n_4447), .b(g64865_sb), .c(g64865_db), .o(n_4426) );
na02s01 TIMEBOOST_cell_15878 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_74), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3196) );
in01s02 g58261_u0 ( .a(FE_OFN1698_n_5751), .o(g58261_sb) );
in01s01 TIMEBOOST_cell_45899 ( .a(wbm_dat_i_0_), .o(TIMEBOOST_net_15206) );
na02s02 TIMEBOOST_cell_19128 ( .a(wbm_adr_o_29_), .b(FE_OFN1697_n_5751), .o(TIMEBOOST_net_4821) );
na02s02 TIMEBOOST_cell_19289 ( .a(TIMEBOOST_net_4901), .b(g60649_sb), .o(n_5676) );
in01s01 g58262_u0 ( .a(FE_OFN519_n_9697), .o(g58262_sb) );
na02s01 TIMEBOOST_cell_15879 ( .a(TIMEBOOST_net_3196), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_387), .o(TIMEBOOST_net_78) );
na02s01 g58262_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__Q), .b(FE_OFN519_n_9697), .o(g58262_db) );
na03s02 TIMEBOOST_cell_40631 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__Q), .b(n_1861), .c(FE_OFN1215_n_4151), .o(TIMEBOOST_net_12554) );
in01s01 g58263_u0 ( .a(FE_OFN1801_n_9690), .o(g58263_sb) );
na02f02 TIMEBOOST_cell_39121 ( .a(FE_OFN1605_n_13997), .b(TIMEBOOST_net_10178), .o(TIMEBOOST_net_11799) );
na02s02 TIMEBOOST_cell_18032 ( .a(pci_target_unit_fifos_pciw_addr_data_in_132), .b(g64080_sb), .o(TIMEBOOST_net_4273) );
na02s02 TIMEBOOST_cell_38200 ( .a(TIMEBOOST_net_11338), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_4611) );
in01s01 g58264_u0 ( .a(FE_OFN1632_n_9531), .o(g58264_sb) );
na02s01 TIMEBOOST_cell_16321 ( .a(TIMEBOOST_net_3417), .b(g66406_sb), .o(n_2498) );
na02s01 g58264_u2 ( .a(FE_OFN250_n_9789), .b(FE_OFN1632_n_9531), .o(g58264_db) );
na02f04 TIMEBOOST_cell_37028 ( .a(TIMEBOOST_net_10752), .b(g52524_sb), .o(n_13696) );
in01s01 g58265_u0 ( .a(FE_OFN1649_n_9428), .o(g58265_sb) );
na02s01 g58265_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__Q), .b(g58265_sb), .o(g58265_da) );
na02s01 g58265_u2 ( .a(FE_OFN239_n_9832), .b(FE_OFN1649_n_9428), .o(g58265_db) );
na02s01 g58265_u3 ( .a(g58265_da), .b(g58265_db), .o(n_9534) );
in01s01 g58266_u0 ( .a(FE_OFN579_n_9531), .o(g58266_sb) );
na02m02 TIMEBOOST_cell_31494 ( .a(n_1782), .b(TIMEBOOST_net_1652), .o(TIMEBOOST_net_9658) );
na02s01 g58266_u2 ( .a(FE_OFN231_n_9839), .b(FE_OFN579_n_9531), .o(g58266_db) );
na02s01 TIMEBOOST_cell_40494 ( .a(TIMEBOOST_net_12485), .b(FE_OFN1300_n_5763), .o(TIMEBOOST_net_11510) );
in01s01 g58267_u0 ( .a(FE_OFN1651_n_9428), .o(g58267_sb) );
na02f02 TIMEBOOST_cell_43932 ( .a(TIMEBOOST_net_14204), .b(FE_OFN1415_n_8567), .o(TIMEBOOST_net_12819) );
na02s01 g58267_u2 ( .a(FE_OFN205_n_9140), .b(FE_OFN1651_n_9428), .o(g58267_db) );
na02s02 TIMEBOOST_cell_40664 ( .a(TIMEBOOST_net_12570), .b(g62624_sb), .o(n_6308) );
in01s01 g58268_u0 ( .a(FE_OFN602_n_9687), .o(g58268_sb) );
na02s01 TIMEBOOST_cell_16646 ( .a(pci_target_unit_fifos_pciw_addr_data_in_146), .b(g64163_sb), .o(TIMEBOOST_net_3580) );
na02s01 g58268_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__Q), .b(FE_OFN602_n_9687), .o(g58268_db) );
na02s01 TIMEBOOST_cell_44929 ( .a(FE_OFN239_n_9832), .b(g57937_sb), .o(TIMEBOOST_net_14703) );
in01s01 g58269_u0 ( .a(FE_OFN602_n_9687), .o(g58269_sb) );
na02s01 g58269_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__Q), .b(FE_OFN602_n_9687), .o(g58269_db) );
na02s02 TIMEBOOST_cell_43550 ( .a(TIMEBOOST_net_14013), .b(FE_OFN1311_n_6624), .o(TIMEBOOST_net_12216) );
in01s01 g58270_u0 ( .a(FE_OFN602_n_9687), .o(g58270_sb) );
na02s03 TIMEBOOST_cell_45758 ( .a(TIMEBOOST_net_15117), .b(FE_OFN1326_n_13547), .o(TIMEBOOST_net_14950) );
na02s01 g58270_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q), .b(FE_OFN602_n_9687), .o(g58270_db) );
na02m02 TIMEBOOST_cell_44659 ( .a(n_9233), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__Q), .o(TIMEBOOST_net_14568) );
in01s01 g58271_u0 ( .a(FE_OFN569_n_9528), .o(g58271_sb) );
na02s01 TIMEBOOST_cell_44930 ( .a(TIMEBOOST_net_14703), .b(g57937_db), .o(n_9873) );
na02s01 g58271_u2 ( .a(FE_OFN207_n_9865), .b(FE_OFN569_n_9528), .o(g58271_db) );
na02s01 TIMEBOOST_cell_39744 ( .a(TIMEBOOST_net_12110), .b(g62549_sb), .o(n_6468) );
in01s01 g58272_u0 ( .a(FE_OFN1690_n_9528), .o(g58272_sb) );
na02f02 TIMEBOOST_cell_42464 ( .a(TIMEBOOST_net_13470), .b(g57413_sb), .o(n_10363) );
na02m04 TIMEBOOST_cell_10506 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__Q), .b(FE_OFN2059_n_13447), .o(TIMEBOOST_net_1820) );
na02m02 TIMEBOOST_cell_38935 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_0__Q), .o(TIMEBOOST_net_11706) );
in01s01 g58273_u0 ( .a(FE_OFN1687_n_9528), .o(g58273_sb) );
na02s02 TIMEBOOST_cell_45654 ( .a(TIMEBOOST_net_15065), .b(g62716_sb), .o(TIMEBOOST_net_10611) );
na02m02 TIMEBOOST_cell_43699 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__Q), .b(n_9737), .o(TIMEBOOST_net_14088) );
na03s02 TIMEBOOST_cell_38355 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__Q), .b(FE_OFN1124_g64577_p), .c(n_3997), .o(TIMEBOOST_net_11416) );
in01s01 g58274_u0 ( .a(FE_OFN1688_n_9528), .o(g58274_sb) );
na02s01 TIMEBOOST_cell_17498 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_127), .o(TIMEBOOST_net_4006) );
na02s01 g58274_u2 ( .a(FE_OFN209_n_9126), .b(FE_OFN1688_n_9528), .o(g58274_db) );
na02s02 TIMEBOOST_cell_17499 ( .a(TIMEBOOST_net_4006), .b(FE_OFN1076_n_4740), .o(TIMEBOOST_net_1689) );
in01s01 g58275_u0 ( .a(FE_OFN1687_n_9528), .o(g58275_sb) );
na02f02 TIMEBOOST_cell_43933 ( .a(n_9903), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__Q), .o(TIMEBOOST_net_14205) );
na02s01 g58275_u2 ( .a(FE_OFN211_n_9858), .b(FE_OFN1687_n_9528), .o(g58275_db) );
na02f02 TIMEBOOST_cell_43934 ( .a(TIMEBOOST_net_14205), .b(FE_OFN1421_n_8567), .o(TIMEBOOST_net_12813) );
in01s01 g58276_u0 ( .a(FE_OFN568_n_9528), .o(g58276_sb) );
na02s02 TIMEBOOST_cell_45204 ( .a(TIMEBOOST_net_14840), .b(FE_OFN1208_n_6356), .o(TIMEBOOST_net_12099) );
na02s01 g58276_u2 ( .a(FE_OFN213_n_9124), .b(FE_OFN568_n_9528), .o(g58276_db) );
na02s02 TIMEBOOST_cell_40666 ( .a(TIMEBOOST_net_12571), .b(g62352_sb), .o(n_6897) );
in01s01 g58277_u0 ( .a(FE_OFN568_n_9528), .o(g58277_sb) );
na02s02 TIMEBOOST_cell_17500 ( .a(pci_target_unit_fifos_pciw_addr_data_in_146), .b(g64134_sb), .o(TIMEBOOST_net_4007) );
na02s01 g58277_u2 ( .a(FE_OFN215_n_9856), .b(FE_OFN568_n_9528), .o(g58277_db) );
na02s02 TIMEBOOST_cell_44413 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_771), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_6__Q), .o(TIMEBOOST_net_14445) );
in01s01 g58278_u0 ( .a(FE_OFN1691_n_9528), .o(g58278_sb) );
na02s02 TIMEBOOST_cell_43388 ( .a(TIMEBOOST_net_13932), .b(n_6554), .o(TIMEBOOST_net_12155) );
na02s01 g58278_u2 ( .a(FE_OFN217_n_9889), .b(FE_OFN1691_n_9528), .o(g58278_db) );
na02s01 TIMEBOOST_cell_9401 ( .a(TIMEBOOST_net_1267), .b(g65715_sb), .o(n_1722) );
in01s01 g58279_u0 ( .a(FE_OFN1687_n_9528), .o(g58279_sb) );
na02s02 TIMEBOOST_cell_39746 ( .a(TIMEBOOST_net_12111), .b(g62970_sb), .o(n_5942) );
na02s01 g58279_u2 ( .a(FE_OFN219_n_9853), .b(FE_OFN1687_n_9528), .o(g58279_db) );
na02s02 TIMEBOOST_cell_17361 ( .a(TIMEBOOST_net_3937), .b(FE_OFN235_n_9834), .o(n_9438) );
in01s01 g58280_u0 ( .a(FE_OFN1690_n_9528), .o(g58280_sb) );
na02s02 TIMEBOOST_cell_42378 ( .a(TIMEBOOST_net_13427), .b(g54349_sb), .o(n_13093) );
na02m02 TIMEBOOST_cell_10510 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__Q), .b(n_504), .o(TIMEBOOST_net_1822) );
na02s01 TIMEBOOST_cell_44862 ( .a(TIMEBOOST_net_14669), .b(g58326_sb), .o(TIMEBOOST_net_11935) );
in01s01 g58281_u0 ( .a(FE_OFN1689_n_9528), .o(g58281_sb) );
na02f02 TIMEBOOST_cell_44749 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__Q), .b(FE_OFN1753_n_12086), .o(TIMEBOOST_net_14613) );
na02s01 TIMEBOOST_cell_43357 ( .a(n_2184), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__Q), .o(TIMEBOOST_net_13917) );
na02s02 TIMEBOOST_cell_38202 ( .a(TIMEBOOST_net_11339), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_4717) );
in01s01 g58282_u0 ( .a(FE_OFN569_n_9528), .o(g58282_sb) );
na02f02 TIMEBOOST_cell_38808 ( .a(TIMEBOOST_net_11642), .b(FE_OFN1428_n_8567), .o(n_11380) );
na02s02 TIMEBOOST_cell_10512 ( .a(n_526), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_1823) );
na02s02 TIMEBOOST_cell_37836 ( .a(TIMEBOOST_net_11156), .b(g58316_sb), .o(n_9496) );
in01s01 g58283_u0 ( .a(FE_OFN1690_n_9528), .o(g58283_sb) );
na02s01 TIMEBOOST_cell_17362 ( .a(FE_OFN215_n_9856), .b(FE_OFN1650_n_9428), .o(TIMEBOOST_net_3938) );
na02s01 g58283_u2 ( .a(FE_OFN221_n_9846), .b(FE_OFN1690_n_9528), .o(g58283_db) );
na02s01 TIMEBOOST_cell_17363 ( .a(TIMEBOOST_net_3938), .b(g58424_da), .o(n_9424) );
in01s01 g58284_u0 ( .a(FE_OFN1692_n_9528), .o(g58284_sb) );
na02s02 TIMEBOOST_cell_45205 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__26__Q), .b(n_4355), .o(TIMEBOOST_net_14841) );
na02s01 g58284_u2 ( .a(FE_OFN223_n_9844), .b(FE_OFN1692_n_9528), .o(g58284_db) );
na02s01 TIMEBOOST_cell_40496 ( .a(TIMEBOOST_net_12486), .b(FE_OFN1299_n_5763), .o(TIMEBOOST_net_11511) );
in01s01 g58285_u0 ( .a(FE_OFN1690_n_9528), .o(g58285_sb) );
na02s01 TIMEBOOST_cell_9408 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(g65737_sb), .o(TIMEBOOST_net_1271) );
na02s01 g58285_u2 ( .a(FE_OFN225_n_9122), .b(FE_OFN1690_n_9528), .o(g58285_db) );
na02s01 TIMEBOOST_cell_9409 ( .a(TIMEBOOST_net_1271), .b(g65737_db), .o(n_1933) );
in01s01 g58286_u0 ( .a(FE_OFN1687_n_9528), .o(g58286_sb) );
na03s02 TIMEBOOST_cell_38203 ( .a(TIMEBOOST_net_4038), .b(g64314_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__Q), .o(TIMEBOOST_net_11340) );
na02s02 TIMEBOOST_cell_10514 ( .a(n_213), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_1824) );
na02s02 TIMEBOOST_cell_37838 ( .a(TIMEBOOST_net_11157), .b(g58403_sb), .o(n_9434) );
in01s01 g58287_u0 ( .a(FE_OFN1687_n_9528), .o(g58287_sb) );
na02m02 TIMEBOOST_cell_43935 ( .a(n_9522), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__Q), .o(TIMEBOOST_net_14206) );
na02s01 g58287_u2 ( .a(FE_OFN227_n_9841), .b(FE_OFN1687_n_9528), .o(g58287_db) );
na02f02 TIMEBOOST_cell_43936 ( .a(TIMEBOOST_net_14206), .b(FE_OFN1383_n_8567), .o(TIMEBOOST_net_12968) );
in01s01 g58288_u0 ( .a(FE_OFN1688_n_9528), .o(g58288_sb) );
na02s01 TIMEBOOST_cell_9412 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(g65764_sb), .o(TIMEBOOST_net_1273) );
na02s01 g58288_u2 ( .a(FE_OFN229_n_9120), .b(FE_OFN1688_n_9528), .o(g58288_db) );
na02s01 TIMEBOOST_cell_9413 ( .a(TIMEBOOST_net_1273), .b(g65764_db), .o(n_1917) );
in01s01 g58289_u0 ( .a(FE_OFN1687_n_9528), .o(g58289_sb) );
na02s01 g58289_u2 ( .a(FE_OFN231_n_9839), .b(FE_OFN1687_n_9528), .o(g58289_db) );
na02s01 TIMEBOOST_cell_40498 ( .a(TIMEBOOST_net_12487), .b(FE_OFN1299_n_5763), .o(TIMEBOOST_net_11513) );
in01s01 g58290_u0 ( .a(FE_OFN1690_n_9528), .o(g58290_sb) );
na02s02 TIMEBOOST_cell_17502 ( .a(pci_target_unit_fifos_pciw_addr_data_in_144), .b(g64137_sb), .o(TIMEBOOST_net_4008) );
na02s01 g58290_u2 ( .a(FE_OFN233_n_9876), .b(FE_OFN1690_n_9528), .o(g58290_db) );
na02m02 TIMEBOOST_cell_44407 ( .a(n_9612), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__Q), .o(TIMEBOOST_net_14442) );
in01s01 g58291_u0 ( .a(FE_OFN1690_n_9528), .o(g58291_sb) );
na02s02 TIMEBOOST_cell_37450 ( .a(TIMEBOOST_net_10963), .b(FE_OFN1800_n_9690), .o(TIMEBOOST_net_4062) );
na02s01 TIMEBOOST_cell_10516 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_1__Q), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_1825) );
na02s02 TIMEBOOST_cell_37840 ( .a(TIMEBOOST_net_11158), .b(g58376_sb), .o(n_9453) );
in01s01 g58292_u0 ( .a(FE_OFN1690_n_9528), .o(g58292_sb) );
na02s01 TIMEBOOST_cell_17504 ( .a(pci_target_unit_fifos_pciw_addr_data_in_147), .b(g64173_sb), .o(TIMEBOOST_net_4009) );
na02s01 g58292_u2 ( .a(FE_OFN235_n_9834), .b(FE_OFN1690_n_9528), .o(g58292_db) );
na02s02 TIMEBOOST_cell_43642 ( .a(TIMEBOOST_net_14059), .b(FE_OFN1295_n_4098), .o(TIMEBOOST_net_12048) );
in01s01 g58293_u0 ( .a(FE_OFN1689_n_9528), .o(g58293_sb) );
na02s02 TIMEBOOST_cell_17506 ( .a(pci_target_unit_fifos_pciw_addr_data_in_149), .b(g64179_sb), .o(TIMEBOOST_net_4010) );
na02s01 g58293_u2 ( .a(FE_OFN237_n_9118), .b(FE_OFN1689_n_9528), .o(g58293_db) );
na02s01 TIMEBOOST_cell_44931 ( .a(FE_OFN233_n_9876), .b(g57933_sb), .o(TIMEBOOST_net_14704) );
in01s01 g58294_u0 ( .a(FE_OFN1691_n_9528), .o(g58294_sb) );
na02s01 TIMEBOOST_cell_17508 ( .a(n_3770), .b(FE_OFN643_n_4677), .o(TIMEBOOST_net_4011) );
na02s01 g58294_u2 ( .a(FE_OFN239_n_9832), .b(FE_OFN1691_n_9528), .o(g58294_db) );
na02s01 TIMEBOOST_cell_17509 ( .a(TIMEBOOST_net_4011), .b(g65287_da), .o(n_3581) );
in01s01 g58295_u0 ( .a(FE_OFN568_n_9528), .o(g58295_sb) );
na02s01 g58295_u2 ( .a(FE_OFN241_n_9830), .b(FE_OFN568_n_9528), .o(g58295_db) );
na02s01 TIMEBOOST_cell_40500 ( .a(TIMEBOOST_net_12488), .b(FE_OFN1300_n_5763), .o(TIMEBOOST_net_11512) );
in01s01 g58296_u0 ( .a(FE_OFN569_n_9528), .o(g58296_sb) );
na02s01 TIMEBOOST_cell_39249 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__Q), .b(FE_OFN653_n_4508), .o(TIMEBOOST_net_11863) );
na02m04 TIMEBOOST_cell_39035 ( .a(wbs_wbb3_2_wbb2_dat_o_i_115), .b(wbs_dat_o_16_), .o(TIMEBOOST_net_11756) );
na02s01 TIMEBOOST_cell_39250 ( .a(TIMEBOOST_net_11863), .b(g65422_sb), .o(TIMEBOOST_net_3639) );
in01s01 g58297_u0 ( .a(FE_OFN568_n_9528), .o(g58297_sb) );
na02s01 TIMEBOOST_cell_39251 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__Q), .b(FE_OFN1649_n_9428), .o(TIMEBOOST_net_11864) );
na02s01 g58297_u2 ( .a(FE_OFN203_n_9228), .b(FE_OFN568_n_9528), .o(g58297_db) );
na02s01 TIMEBOOST_cell_45747 ( .a(n_1955), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__Q), .o(TIMEBOOST_net_15112) );
in01s01 g58298_u0 ( .a(FE_OFN569_n_9528), .o(g58298_sb) );
na02f02 TIMEBOOST_cell_43788 ( .a(TIMEBOOST_net_14132), .b(FE_OFN1419_n_8567), .o(TIMEBOOST_net_12798) );
na02s01 g58298_u2 ( .a(FE_OFN205_n_9140), .b(FE_OFN569_n_9528), .o(g58298_db) );
na02m02 TIMEBOOST_cell_38828 ( .a(TIMEBOOST_net_11652), .b(g58463_sb), .o(n_9389) );
in01s01 g58299_u0 ( .a(FE_OFN1691_n_9528), .o(g58299_sb) );
na02s01 TIMEBOOST_cell_42720 ( .a(TIMEBOOST_net_13598), .b(g58053_sb), .o(TIMEBOOST_net_10956) );
na02s01 TIMEBOOST_cell_9202 ( .a(pci_target_unit_fifos_pcir_data_in_164), .b(g65789_sb), .o(TIMEBOOST_net_1168) );
na02s01 TIMEBOOST_cell_9203 ( .a(TIMEBOOST_net_1168), .b(g65789_db), .o(n_2189) );
in01s01 g58300_u0 ( .a(FE_OFN1689_n_9528), .o(g58300_sb) );
na02s02 TIMEBOOST_cell_42974 ( .a(TIMEBOOST_net_13725), .b(n_4608), .o(n_6967) );
na02s02 TIMEBOOST_cell_43358 ( .a(TIMEBOOST_net_13917), .b(FE_OFN2212_n_8407), .o(TIMEBOOST_net_11242) );
na02s02 TIMEBOOST_cell_38204 ( .a(TIMEBOOST_net_11340), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_4614) );
in01s01 g58301_u0 ( .a(FE_OFN1691_n_9528), .o(g58301_sb) );
na02f02 TIMEBOOST_cell_43804 ( .a(TIMEBOOST_net_14140), .b(FE_OFN1382_n_8567), .o(TIMEBOOST_net_12961) );
na02s01 g58301_u2 ( .a(FE_OFN243_n_9116), .b(FE_OFN1691_n_9528), .o(g58301_db) );
na02s01 TIMEBOOST_cell_40502 ( .a(TIMEBOOST_net_12489), .b(FE_OFN1301_n_5763), .o(TIMEBOOST_net_11502) );
in01s01 g58302_u0 ( .a(FE_OFN568_n_9528), .o(g58302_sb) );
na02f02 TIMEBOOST_cell_4105 ( .a(TIMEBOOST_net_632), .b(n_15695), .o(n_15698) );
na02s01 g58302_u2 ( .a(FE_OFN245_n_9114), .b(FE_OFN568_n_9528), .o(g58302_db) );
na02s01 TIMEBOOST_cell_43127 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__Q), .b(n_3726), .o(TIMEBOOST_net_13802) );
in01s01 g58303_u0 ( .a(FE_OFN1689_n_9528), .o(g58303_sb) );
na02s01 TIMEBOOST_cell_39215 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__Q), .b(n_8119), .o(TIMEBOOST_net_11846) );
na02s01 g58303_u2 ( .a(FE_OFN247_n_9112), .b(FE_OFN1689_n_9528), .o(g58303_db) );
na02s01 TIMEBOOST_cell_41806 ( .a(TIMEBOOST_net_13141), .b(g61862_sb), .o(n_8114) );
in01s01 g58304_u0 ( .a(FE_OFN1689_n_9528), .o(g58304_sb) );
na02s02 TIMEBOOST_cell_39748 ( .a(TIMEBOOST_net_12112), .b(g62356_sb), .o(n_6887) );
na02s01 g58304_u2 ( .a(FE_OFN250_n_9789), .b(FE_OFN1689_n_9528), .o(g58304_db) );
na02s01 TIMEBOOST_cell_17373 ( .a(TIMEBOOST_net_3943), .b(n_4450), .o(n_4395) );
in01s01 g58305_u0 ( .a(FE_OFN569_n_9528), .o(g58305_sb) );
na02m02 TIMEBOOST_cell_45142 ( .a(TIMEBOOST_net_14809), .b(g54174_da), .o(TIMEBOOST_net_10642) );
na02s01 g58305_u2 ( .a(FE_OFN252_n_9868), .b(FE_OFN569_n_9528), .o(g58305_db) );
na02s01 TIMEBOOST_cell_39750 ( .a(TIMEBOOST_net_12113), .b(g62392_sb), .o(n_6814) );
in01s01 g58306_u0 ( .a(FE_OFN1687_n_9528), .o(g58306_sb) );
na02s01 TIMEBOOST_cell_17376 ( .a(g65057_sb), .b(g65057_db), .o(TIMEBOOST_net_3945) );
na02f02 TIMEBOOST_cell_39123 ( .a(TIMEBOOST_net_10163), .b(FE_OFN1606_n_13997), .o(TIMEBOOST_net_11800) );
na02s01 TIMEBOOST_cell_17377 ( .a(TIMEBOOST_net_3945), .b(n_4450), .o(n_4319) );
in01s01 g58307_u0 ( .a(FE_OFN1657_n_9502), .o(g58307_sb) );
na02s01 g58307_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__Q), .b(g58307_sb), .o(g58307_da) );
na02s01 g58307_u2 ( .a(FE_OFN207_n_9865), .b(FE_OFN1657_n_9502), .o(g58307_db) );
na02s02 g58307_u3 ( .a(g58307_da), .b(g58307_db), .o(n_9504) );
in01s01 g58308_u0 ( .a(FE_OFN572_n_9502), .o(g58308_sb) );
na02m02 TIMEBOOST_cell_31493 ( .a(FE_OFN1147_n_13249), .b(TIMEBOOST_net_9657), .o(TIMEBOOST_net_4338) );
na03s02 TIMEBOOST_cell_45793 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__Q), .b(g63563_da), .c(g63563_db), .o(TIMEBOOST_net_15135) );
in01s01 g58309_u0 ( .a(FE_OFN1654_n_9502), .o(g58309_sb) );
na02m02 TIMEBOOST_cell_31492 ( .a(TIMEBOOST_net_1642), .b(wishbone_slave_unit_pcim_if_wbw_cbe_in), .o(TIMEBOOST_net_9657) );
na03s02 TIMEBOOST_cell_33402 ( .a(n_4479), .b(g64784_sb), .c(g64784_db), .o(n_4480) );
na02f02 TIMEBOOST_cell_38952 ( .a(TIMEBOOST_net_11714), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10730) );
in01s01 g58310_u0 ( .a(FE_OFN1655_n_9502), .o(g58310_sb) );
na02m02 TIMEBOOST_cell_43937 ( .a(n_9683), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__Q), .o(TIMEBOOST_net_14207) );
na02s01 g58310_u2 ( .a(FE_OFN209_n_9126), .b(FE_OFN1655_n_9502), .o(g58310_db) );
na02f04 TIMEBOOST_cell_37030 ( .a(TIMEBOOST_net_10753), .b(g52526_sb), .o(n_13794) );
in01s01 g58311_u0 ( .a(FE_OFN572_n_9502), .o(g58311_sb) );
na02s01 g58311_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__Q), .b(g58311_sb), .o(g58311_da) );
na02f02 TIMEBOOST_cell_43700 ( .a(TIMEBOOST_net_14088), .b(FE_OFN1349_n_8567), .o(TIMEBOOST_net_12994) );
na02s01 TIMEBOOST_cell_43359 ( .a(n_2177), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__Q), .o(TIMEBOOST_net_13918) );
in01s01 g58312_u0 ( .a(FE_OFN1656_n_9502), .o(g58312_sb) );
na02s01 g58312_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__Q), .b(g58312_sb), .o(g58312_da) );
na02s01 g58312_u2 ( .a(FE_OFN213_n_9124), .b(FE_OFN1656_n_9502), .o(g58312_db) );
na02s01 g58312_u3 ( .a(g58312_da), .b(g58312_db), .o(n_9025) );
in01s01 g58313_u0 ( .a(FE_OFN572_n_9502), .o(g58313_sb) );
na02s02 TIMEBOOST_cell_43146 ( .a(TIMEBOOST_net_13811), .b(FE_OFN1258_n_4143), .o(TIMEBOOST_net_12066) );
na02s01 TIMEBOOST_cell_17660 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__Q), .b(g65305_sb), .o(TIMEBOOST_net_4087) );
na02f04 TIMEBOOST_cell_37032 ( .a(TIMEBOOST_net_10754), .b(g52520_sb), .o(n_13738) );
in01s01 g58314_u0 ( .a(FE_OFN1654_n_9502), .o(g58314_sb) );
na02s02 TIMEBOOST_cell_45039 ( .a(n_2039), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__Q), .o(TIMEBOOST_net_14758) );
na02s01 g58314_u2 ( .a(FE_OFN219_n_9853), .b(FE_OFN1654_n_9502), .o(g58314_db) );
na02f02 TIMEBOOST_cell_36966 ( .a(TIMEBOOST_net_10721), .b(g58831_sb), .o(n_8606) );
in01s01 g58315_u0 ( .a(FE_OFN572_n_9502), .o(g58315_sb) );
na02m02 TIMEBOOST_cell_31486 ( .a(n_1823), .b(n_8498), .o(TIMEBOOST_net_9654) );
na02s02 TIMEBOOST_cell_19349 ( .a(TIMEBOOST_net_4931), .b(g60614_sb), .o(n_4840) );
na02s02 TIMEBOOST_cell_42050 ( .a(TIMEBOOST_net_13263), .b(g62615_sb), .o(n_6327) );
in01s01 g58316_u0 ( .a(FE_OFN572_n_9502), .o(g58316_sb) );
na02s01 TIMEBOOST_cell_31485 ( .a(TIMEBOOST_net_9653), .b(g65300_sb), .o(n_4190) );
na03f02 TIMEBOOST_cell_22252 ( .a(n_10032), .b(n_9262), .c(n_9261), .o(TIMEBOOST_net_6383) );
na03s01 TIMEBOOST_cell_33132 ( .a(g65780_da), .b(g61713_db), .c(TIMEBOOST_net_188), .o(n_8400) );
in01s01 g58317_u0 ( .a(FE_OFN1657_n_9502), .o(g58317_sb) );
na02s01 TIMEBOOST_cell_42865 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__Q), .b(FE_OFN540_n_9690), .o(TIMEBOOST_net_13671) );
na03s01 TIMEBOOST_cell_33131 ( .a(g65733_da), .b(g61705_db), .c(TIMEBOOST_net_187), .o(n_8417) );
na02s02 TIMEBOOST_cell_45406 ( .a(TIMEBOOST_net_14941), .b(g62955_sb), .o(n_5971) );
in01s01 g58318_u0 ( .a(FE_OFN1656_n_9502), .o(g58318_sb) );
na02s01 g58318_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__Q), .b(g58318_sb), .o(g58318_da) );
na02s01 g58318_u2 ( .a(FE_OFN221_n_9846), .b(FE_OFN1656_n_9502), .o(g58318_db) );
na02s01 g58318_u3 ( .a(g58318_da), .b(g58318_db), .o(n_9494) );
in01s01 g58319_u0 ( .a(FE_OFN572_n_9502), .o(g58319_sb) );
na02s01 TIMEBOOST_cell_31483 ( .a(TIMEBOOST_net_9652), .b(g65328_db), .o(n_3555) );
na02s01 g58319_u2 ( .a(FE_OFN223_n_9844), .b(FE_OFN572_n_9502), .o(g58319_db) );
na02s01 TIMEBOOST_cell_31482 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q), .b(g65328_sb), .o(TIMEBOOST_net_9652) );
in01s01 g58320_u0 ( .a(FE_OFN572_n_9502), .o(g58320_sb) );
na02s01 g58320_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__22__Q), .b(g58320_sb), .o(g58320_da) );
na02s01 g58320_u2 ( .a(FE_OFN225_n_9122), .b(FE_OFN572_n_9502), .o(g58320_db) );
na02s01 g58320_u3 ( .a(g58320_da), .b(g58320_db), .o(n_9024) );
in01s01 g58321_u0 ( .a(FE_OFN1654_n_9502), .o(g58321_sb) );
na02s02 TIMEBOOST_cell_41731 ( .a(FE_OFN219_n_9853), .b(g57922_sb), .o(TIMEBOOST_net_13104) );
in01s01 g58322_u0 ( .a(FE_OFN1654_n_9502), .o(g58322_sb) );
na02s02 TIMEBOOST_cell_39752 ( .a(TIMEBOOST_net_12114), .b(g62629_sb), .o(n_6297) );
na02s01 g58322_u2 ( .a(FE_OFN227_n_9841), .b(FE_OFN1654_n_9502), .o(g58322_db) );
na02s01 TIMEBOOST_cell_31481 ( .a(TIMEBOOST_net_9651), .b(g65307_db), .o(n_3572) );
in01s01 g58323_u0 ( .a(FE_OFN1655_n_9502), .o(g58323_sb) );
na02s01 TIMEBOOST_cell_31480 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__Q), .b(g65307_sb), .o(TIMEBOOST_net_9651) );
na02s01 g58323_u2 ( .a(FE_OFN229_n_9120), .b(FE_OFN1655_n_9502), .o(g58323_db) );
na02s01 TIMEBOOST_cell_31479 ( .a(TIMEBOOST_net_9650), .b(g65296_db), .o(n_3576) );
in01s01 g58324_u0 ( .a(FE_OFN572_n_9502), .o(g58324_sb) );
na02s01 g58324_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__Q), .b(g58324_sb), .o(g58324_da) );
na02s01 g58324_u2 ( .a(FE_OFN231_n_9839), .b(FE_OFN572_n_9502), .o(g58324_db) );
na02s02 g58324_u3 ( .a(g58324_da), .b(g58324_db), .o(n_9490) );
in01s01 g58325_u0 ( .a(FE_OFN572_n_9502), .o(g58325_sb) );
na02s01 g58325_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__Q), .b(g58325_sb), .o(g58325_da) );
na02s01 g58325_u2 ( .a(FE_OFN233_n_9876), .b(FE_OFN572_n_9502), .o(g58325_db) );
na02s01 g58325_u3 ( .a(g58325_da), .b(g58325_db), .o(n_9489) );
in01s01 g58326_u0 ( .a(FE_OFN1657_n_9502), .o(g58326_sb) );
na02s01 TIMEBOOST_cell_31478 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q), .b(g65296_sb), .o(TIMEBOOST_net_9650) );
na02s02 TIMEBOOST_cell_42994 ( .a(TIMEBOOST_net_13735), .b(g58293_db), .o(n_9031) );
na02s02 TIMEBOOST_cell_42995 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__Q), .b(g58362_sb), .o(TIMEBOOST_net_13736) );
in01s01 g58327_u0 ( .a(FE_OFN572_n_9502), .o(g58327_sb) );
na02s01 g58327_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__Q), .b(g58327_sb), .o(g58327_da) );
na02s01 g58327_u2 ( .a(FE_OFN235_n_9834), .b(FE_OFN572_n_9502), .o(g58327_db) );
na02s02 g58327_u3 ( .a(g58327_da), .b(g58327_db), .o(n_9487) );
in01s01 g58328_u0 ( .a(FE_OFN572_n_9502), .o(g58328_sb) );
na02s01 g58328_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__Q), .b(g58328_sb), .o(g58328_da) );
na02s01 g58328_u2 ( .a(FE_OFN239_n_9832), .b(FE_OFN572_n_9502), .o(g58328_db) );
na02s01 g58328_u3 ( .a(g58328_da), .b(g58328_db), .o(n_9486) );
in01s01 g58329_u0 ( .a(FE_OFN1656_n_9502), .o(g58329_sb) );
na02s01 g58329_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q), .b(g58329_sb), .o(g58329_da) );
na02s01 g58329_u2 ( .a(FE_OFN241_n_9830), .b(FE_OFN1656_n_9502), .o(g58329_db) );
na02s01 g58329_u3 ( .a(g58329_da), .b(g58329_db), .o(n_9485) );
in01s01 g58330_u0 ( .a(FE_OFN1657_n_9502), .o(g58330_sb) );
na02s02 TIMEBOOST_cell_31477 ( .a(TIMEBOOST_net_9649), .b(g65345_db), .o(n_3544) );
na02s01 g58330_u2 ( .a(FE_OFN201_n_9230), .b(FE_OFN1657_n_9502), .o(g58330_db) );
na02s01 TIMEBOOST_cell_31476 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__Q), .b(g65345_sb), .o(TIMEBOOST_net_9649) );
in01s01 g58331_u0 ( .a(FE_OFN1656_n_9502), .o(g58331_sb) );
in01s01 TIMEBOOST_cell_45879 ( .a(n_727), .o(TIMEBOOST_net_15186) );
na02s01 g58331_u2 ( .a(FE_OFN203_n_9228), .b(FE_OFN1656_n_9502), .o(g58331_db) );
na02f02 TIMEBOOST_cell_36968 ( .a(TIMEBOOST_net_10722), .b(g58822_sb), .o(n_8619) );
in01s01 g58332_u0 ( .a(FE_OFN1657_n_9502), .o(g58332_sb) );
na02f04 TIMEBOOST_cell_42817 ( .a(TIMEBOOST_net_1424), .b(n_2957), .o(TIMEBOOST_net_13647) );
na02s01 g58332_u2 ( .a(FE_OFN205_n_9140), .b(FE_OFN1657_n_9502), .o(g58332_db) );
na02f02 TIMEBOOST_cell_36936 ( .a(TIMEBOOST_net_10706), .b(g52607_sb), .o(n_10225) );
in01s01 g58333_u0 ( .a(FE_OFN1657_n_9502), .o(g58333_sb) );
na02m02 TIMEBOOST_cell_38949 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_11__Q), .o(TIMEBOOST_net_11713) );
na02s01 TIMEBOOST_cell_9204 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__Q), .b(pci_target_unit_fifos_pcir_data_in_185), .o(TIMEBOOST_net_1169) );
na02s01 TIMEBOOST_cell_9205 ( .a(TIMEBOOST_net_1169), .b(FE_OFN1786_n_1699), .o(TIMEBOOST_net_255) );
in01s01 g58334_u0 ( .a(FE_OFN1654_n_9502), .o(g58334_sb) );
na02s01 TIMEBOOST_cell_42791 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__Q), .b(g64332_sb), .o(TIMEBOOST_net_13634) );
na02s02 TIMEBOOST_cell_41732 ( .a(TIMEBOOST_net_13104), .b(g57922_db), .o(n_9888) );
na02m02 TIMEBOOST_cell_44239 ( .a(n_9765), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__Q), .o(TIMEBOOST_net_14358) );
in01s01 g58335_u0 ( .a(FE_OFN572_n_9502), .o(g58335_sb) );
na02s01 g58335_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__Q), .b(g58335_sb), .o(g58335_da) );
na02s01 g58335_u2 ( .a(FE_OFN243_n_9116), .b(FE_OFN572_n_9502), .o(g58335_db) );
na02s01 g58335_u3 ( .a(g58335_da), .b(g58335_db), .o(n_9021) );
in01s01 g58336_u0 ( .a(FE_OFN1656_n_9502), .o(g58336_sb) );
na03f02 TIMEBOOST_cell_8302 ( .a(n_9454), .b(FE_OFN1426_n_8567), .c(g57516_db), .o(n_11224) );
na02s01 g58336_u2 ( .a(FE_OFN245_n_9114), .b(FE_OFN1656_n_9502), .o(g58336_db) );
in01s01 g58337_u0 ( .a(FE_OFN1655_n_9502), .o(g58337_sb) );
na02s01 g58337_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__Q), .b(g58337_sb), .o(g58337_da) );
na02s01 g58337_u2 ( .a(FE_OFN247_n_9112), .b(FE_OFN1655_n_9502), .o(g58337_db) );
na02s02 g58337_u3 ( .a(g58337_da), .b(g58337_db), .o(n_9019) );
in01s01 g58338_u0 ( .a(FE_OFN1654_n_9502), .o(g58338_sb) );
na02s01 TIMEBOOST_cell_42792 ( .a(TIMEBOOST_net_13634), .b(g64332_db), .o(n_4728) );
na02s01 g58338_u2 ( .a(FE_OFN250_n_9789), .b(FE_OFN1654_n_9502), .o(g58338_db) );
na02s02 TIMEBOOST_cell_40724 ( .a(TIMEBOOST_net_12600), .b(g62503_sb), .o(n_6575) );
in01s01 g58339_u0 ( .a(FE_OFN1657_n_9502), .o(g58339_sb) );
na02s01 TIMEBOOST_cell_44932 ( .a(TIMEBOOST_net_14704), .b(g57933_db), .o(n_9877) );
na02s01 g58339_u2 ( .a(FE_OFN252_n_9868), .b(FE_OFN1657_n_9502), .o(g58339_db) );
na02s01 TIMEBOOST_cell_39754 ( .a(TIMEBOOST_net_12115), .b(g62391_sb), .o(n_6816) );
in01s01 g58340_u0 ( .a(FE_OFN1654_n_9502), .o(g58340_sb) );
na02s01 TIMEBOOST_cell_40504 ( .a(TIMEBOOST_net_12490), .b(FE_OFN1301_n_5763), .o(TIMEBOOST_net_11503) );
na02s01 g58340_u2 ( .a(FE_OFN254_n_9825), .b(FE_OFN1654_n_9502), .o(g58340_db) );
na02f02 TIMEBOOST_cell_43938 ( .a(TIMEBOOST_net_14207), .b(FE_OFN1384_n_8567), .o(TIMEBOOST_net_12801) );
in01s01 g58341_u0 ( .a(FE_OFN1670_n_9477), .o(g58341_sb) );
na02s02 TIMEBOOST_cell_10518 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_14__Q), .b(FE_OFN2072_n_15978), .o(TIMEBOOST_net_1826) );
na03s02 TIMEBOOST_cell_38201 ( .a(TIMEBOOST_net_4033), .b(g64297_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__Q), .o(TIMEBOOST_net_11339) );
na02s02 TIMEBOOST_cell_10519 ( .a(TIMEBOOST_net_1826), .b(FE_OFN1082_n_13221), .o(TIMEBOOST_net_558) );
in01s01 g58342_u0 ( .a(FE_OFN1666_n_9477), .o(g58342_sb) );
na02s01 TIMEBOOST_cell_45131 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__Q), .b(n_3204), .o(TIMEBOOST_net_14804) );
na02s02 TIMEBOOST_cell_45794 ( .a(TIMEBOOST_net_15135), .b(FE_OFN1094_g64577_p), .o(TIMEBOOST_net_6225) );
na02s02 TIMEBOOST_cell_42070 ( .a(TIMEBOOST_net_13273), .b(g62423_sb), .o(n_6749) );
in01s01 g58343_u0 ( .a(FE_OFN1666_n_9477), .o(g58343_sb) );
na02f02 TIMEBOOST_cell_39105 ( .a(TIMEBOOST_net_10168), .b(FE_OFN1606_n_13997), .o(TIMEBOOST_net_11791) );
na02s01 TIMEBOOST_cell_42090 ( .a(TIMEBOOST_net_13283), .b(TIMEBOOST_net_5279), .o(n_6548) );
na02s02 TIMEBOOST_cell_42996 ( .a(TIMEBOOST_net_13736), .b(g58362_db), .o(n_9014) );
in01s01 g58344_u0 ( .a(FE_OFN1668_n_9477), .o(g58344_sb) );
na02m02 TIMEBOOST_cell_38973 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_14__Q), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__Q), .o(TIMEBOOST_net_11725) );
na02s01 g58344_u2 ( .a(FE_OFN209_n_9126), .b(FE_OFN1668_n_9477), .o(g58344_db) );
na02s02 TIMEBOOST_cell_39416 ( .a(TIMEBOOST_net_11946), .b(g52626_da), .o(n_14680) );
in01s01 g58345_u0 ( .a(FE_OFN1666_n_9477), .o(g58345_sb) );
na02s02 TIMEBOOST_cell_17384 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__Q), .b(g64264_sb), .o(TIMEBOOST_net_3949) );
na02s01 g58345_u2 ( .a(FE_OFN211_n_9858), .b(FE_OFN1666_n_9477), .o(g58345_db) );
na02s02 TIMEBOOST_cell_17385 ( .a(TIMEBOOST_net_3949), .b(g64264_db), .o(n_3909) );
in01s01 g58346_u0 ( .a(FE_OFN548_n_9477), .o(g58346_sb) );
na02s02 TIMEBOOST_cell_39417 ( .a(TIMEBOOST_net_329), .b(g61864_sb), .o(TIMEBOOST_net_11947) );
na02s01 g58346_u2 ( .a(FE_OFN213_n_9124), .b(FE_OFN548_n_9477), .o(g58346_db) );
na02f02 TIMEBOOST_cell_38954 ( .a(TIMEBOOST_net_11715), .b(FE_OFN2155_n_16439), .o(TIMEBOOST_net_10731) );
in01s01 g58347_u0 ( .a(FE_OFN548_n_9477), .o(g58347_sb) );
na02s02 TIMEBOOST_cell_45210 ( .a(TIMEBOOST_net_14843), .b(FE_OFN1275_n_4096), .o(TIMEBOOST_net_12589) );
na02s01 g58347_u2 ( .a(FE_OFN215_n_9856), .b(FE_OFN548_n_9477), .o(g58347_db) );
na02s01 TIMEBOOST_cell_9455 ( .a(TIMEBOOST_net_1294), .b(g65761_sb), .o(n_1919) );
in01s01 g58348_u0 ( .a(FE_OFN1671_n_9477), .o(g58348_sb) );
na02s02 TIMEBOOST_cell_45143 ( .a(n_3893), .b(g63063_db), .o(TIMEBOOST_net_14810) );
na03s02 TIMEBOOST_cell_38105 ( .a(TIMEBOOST_net_4260), .b(g64082_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__Q), .o(TIMEBOOST_net_11291) );
na02s02 TIMEBOOST_cell_39756 ( .a(TIMEBOOST_net_12116), .b(g62678_sb), .o(n_6184) );
in01s01 g58349_u0 ( .a(FE_OFN1666_n_9477), .o(g58349_sb) );
na02s01 TIMEBOOST_cell_39424 ( .a(TIMEBOOST_net_11950), .b(g61992_sb), .o(n_7911) );
na02s01 g58349_u2 ( .a(FE_OFN219_n_9853), .b(FE_OFN1666_n_9477), .o(g58349_db) );
na02s01 TIMEBOOST_cell_9457 ( .a(TIMEBOOST_net_1295), .b(g66403_sb), .o(n_2537) );
in01s01 g58350_u0 ( .a(FE_OFN1666_n_9477), .o(g58350_sb) );
na02f02 TIMEBOOST_cell_38956 ( .a(TIMEBOOST_net_11716), .b(FE_OFN2156_n_16439), .o(TIMEBOOST_net_10732) );
na02s01 TIMEBOOST_cell_42596 ( .a(TIMEBOOST_net_13536), .b(g58417_db), .o(n_8999) );
na02f02 TIMEBOOST_cell_44240 ( .a(TIMEBOOST_net_14358), .b(FE_OFN1383_n_8567), .o(TIMEBOOST_net_13481) );
in01s01 g58351_u0 ( .a(FE_OFN1670_n_9477), .o(g58351_sb) );
na02s02 TIMEBOOST_cell_10522 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_22__Q), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_1828) );
na02f02 TIMEBOOST_cell_39122 ( .a(TIMEBOOST_net_11799), .b(FE_OFN1599_n_13995), .o(n_14444) );
na02s02 TIMEBOOST_cell_10523 ( .a(TIMEBOOST_net_1828), .b(FE_OFN1084_n_13221), .o(TIMEBOOST_net_562) );
in01s01 g58352_u0 ( .a(FE_OFN1666_n_9477), .o(g58352_sb) );
na02f02 TIMEBOOST_cell_38958 ( .a(TIMEBOOST_net_11717), .b(FE_OFN2157_n_16439), .o(TIMEBOOST_net_10733) );
na02s01 g58352_u2 ( .a(FE_OFN221_n_9846), .b(FE_OFN1666_n_9477), .o(g58352_db) );
na02s01 TIMEBOOST_cell_9461 ( .a(TIMEBOOST_net_1297), .b(g66406_sb), .o(n_2533) );
in01s01 g58353_u0 ( .a(FE_OFN1668_n_9477), .o(g58353_sb) );
na02f02 TIMEBOOST_cell_38960 ( .a(TIMEBOOST_net_11718), .b(FE_OFN2157_n_16439), .o(TIMEBOOST_net_10734) );
na02s01 g58353_u2 ( .a(FE_OFN223_n_9844), .b(FE_OFN1668_n_9477), .o(g58353_db) );
na02s01 TIMEBOOST_cell_9463 ( .a(TIMEBOOST_net_1298), .b(g66403_sb), .o(n_2531) );
in01s01 g58354_u0 ( .a(FE_OFN1666_n_9477), .o(g58354_sb) );
na02s01 TIMEBOOST_cell_17564 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__Q), .b(g64318_sb), .o(TIMEBOOST_net_4039) );
na02s01 g58354_u2 ( .a(FE_OFN225_n_9122), .b(FE_OFN1666_n_9477), .o(g58354_db) );
na02s01 TIMEBOOST_cell_39185 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__Q), .b(g65934_sb), .o(TIMEBOOST_net_11831) );
in01s01 g58355_u0 ( .a(FE_OFN1666_n_9477), .o(g58355_sb) );
na02f02 TIMEBOOST_cell_38962 ( .a(TIMEBOOST_net_11719), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10722) );
na02f04 TIMEBOOST_cell_44708 ( .a(TIMEBOOST_net_14592), .b(g52602_db), .o(n_10257) );
na03f04 TIMEBOOST_cell_44709 ( .a(n_15537), .b(n_15533), .c(n_15528), .o(TIMEBOOST_net_14593) );
in01s01 g58356_u0 ( .a(FE_OFN1666_n_9477), .o(g58356_sb) );
na02f02 TIMEBOOST_cell_38964 ( .a(TIMEBOOST_net_11720), .b(FE_OFN2155_n_16439), .o(TIMEBOOST_net_10725) );
na02s01 g58356_u2 ( .a(FE_OFN227_n_9841), .b(FE_OFN1666_n_9477), .o(g58356_db) );
na02s01 TIMEBOOST_cell_9469 ( .a(TIMEBOOST_net_1301), .b(g66415_sb), .o(n_2518) );
in01s01 g58357_u0 ( .a(FE_OFN1668_n_9477), .o(g58357_sb) );
na02s02 TIMEBOOST_cell_39324 ( .a(TIMEBOOST_net_11900), .b(g65369_da), .o(TIMEBOOST_net_5438) );
na02s01 g58357_u2 ( .a(FE_OFN229_n_9120), .b(FE_OFN1668_n_9477), .o(g58357_db) );
na02s01 TIMEBOOST_cell_9471 ( .a(TIMEBOOST_net_1302), .b(g66406_sb), .o(n_2517) );
in01s01 g58358_u0 ( .a(FE_OFN1666_n_9477), .o(g58358_sb) );
na02f02 TIMEBOOST_cell_38966 ( .a(TIMEBOOST_net_11721), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10735) );
na02s01 g58358_u2 ( .a(FE_OFN231_n_9839), .b(FE_OFN1666_n_9477), .o(g58358_db) );
na02s01 TIMEBOOST_cell_9473 ( .a(TIMEBOOST_net_1303), .b(g66406_sb), .o(n_2514) );
in01s01 g58359_u0 ( .a(FE_OFN1666_n_9477), .o(g58359_sb) );
na02s01 TIMEBOOST_cell_17566 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__28__Q), .b(g64319_sb), .o(TIMEBOOST_net_4040) );
na02s01 g58359_u2 ( .a(FE_OFN233_n_9876), .b(FE_OFN1666_n_9477), .o(g58359_db) );
na02f04 TIMEBOOST_cell_38799 ( .a(n_8563), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__Q), .o(TIMEBOOST_net_11638) );
in01s01 g58360_u0 ( .a(FE_OFN1666_n_9477), .o(g58360_sb) );
na02s01 TIMEBOOST_cell_17568 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__Q), .b(g64323_sb), .o(TIMEBOOST_net_4041) );
na02f02 TIMEBOOST_cell_43780 ( .a(TIMEBOOST_net_14128), .b(FE_OFN1412_n_8567), .o(TIMEBOOST_net_12714) );
na02s01 TIMEBOOST_cell_37242 ( .a(TIMEBOOST_net_10859), .b(FE_OFN666_n_4495), .o(TIMEBOOST_net_9380) );
in01s01 g58361_u0 ( .a(FE_OFN1666_n_9477), .o(g58361_sb) );
na02s01 TIMEBOOST_cell_17570 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__Q), .b(g65915_sb), .o(TIMEBOOST_net_4042) );
na02s01 g58361_u2 ( .a(FE_OFN235_n_9834), .b(FE_OFN1666_n_9477), .o(g58361_db) );
na02s01 TIMEBOOST_cell_43469 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q), .b(n_3555), .o(TIMEBOOST_net_13973) );
in01s01 g58362_u0 ( .a(FE_OFN1668_n_9477), .o(g58362_sb) );
na02f02 TIMEBOOST_cell_39124 ( .a(TIMEBOOST_net_11800), .b(FE_OFN1599_n_13995), .o(n_14474) );
na02s01 g58362_u2 ( .a(FE_OFN237_n_9118), .b(FE_OFN1668_n_9477), .o(g58362_db) );
na02s01 TIMEBOOST_cell_9481 ( .a(TIMEBOOST_net_1307), .b(g66415_sb), .o(n_2497) );
in01s01 g58363_u0 ( .a(FE_OFN1668_n_9477), .o(g58363_sb) );
na02f02 TIMEBOOST_cell_39126 ( .a(TIMEBOOST_net_11801), .b(FE_OFN1600_n_13995), .o(n_14448) );
na02s01 g58363_u2 ( .a(FE_OFN239_n_9832), .b(FE_OFN1668_n_9477), .o(g58363_db) );
na02s01 TIMEBOOST_cell_9483 ( .a(TIMEBOOST_net_1308), .b(g66406_sb), .o(n_2496) );
in01s01 g58364_u0 ( .a(FE_OFN548_n_9477), .o(g58364_sb) );
na02m02 TIMEBOOST_cell_9484 ( .a(n_2914), .b(n_1966), .o(TIMEBOOST_net_1309) );
na02s01 g58364_u2 ( .a(FE_OFN241_n_9830), .b(FE_OFN548_n_9477), .o(g58364_db) );
na02m02 TIMEBOOST_cell_9485 ( .a(TIMEBOOST_net_1309), .b(n_1965), .o(TIMEBOOST_net_191) );
in01s01 g58365_u0 ( .a(FE_OFN1671_n_9477), .o(g58365_sb) );
na02s01 TIMEBOOST_cell_43300 ( .a(TIMEBOOST_net_13888), .b(g62892_sb), .o(n_6093) );
na03s02 TIMEBOOST_cell_34253 ( .a(TIMEBOOST_net_9793), .b(FE_OFN1168_n_5592), .c(g62096_sb), .o(n_5608) );
na02m02 TIMEBOOST_cell_38943 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_25__Q), .o(TIMEBOOST_net_11710) );
in01s01 g58366_u0 ( .a(FE_OFN1670_n_9477), .o(g58366_sb) );
na02s01 TIMEBOOST_cell_42793 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__1__Q), .b(g63564_sb), .o(TIMEBOOST_net_13635) );
na03s02 TIMEBOOST_cell_38335 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__Q), .b(FE_OFN1129_g64577_p), .c(n_3910), .o(TIMEBOOST_net_11406) );
na02s01 TIMEBOOST_cell_38253 ( .a(n_271), .b(n_4726), .o(TIMEBOOST_net_11365) );
na02s01 g58367_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__Q), .b(FE_OFN1669_n_9477), .o(g58367_da) );
na02s01 TIMEBOOST_cell_17120 ( .a(pci_target_unit_del_sync_addr_in_226), .b(parchk_pci_ad_reg_in_1227), .o(TIMEBOOST_net_3817) );
na02s02 TIMEBOOST_cell_39545 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__Q), .b(g58290_sb), .o(TIMEBOOST_net_12011) );
in01s01 g58368_u0 ( .a(FE_OFN1668_n_9477), .o(g58368_sb) );
na02m02 TIMEBOOST_cell_38955 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_9__Q), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__Q), .o(TIMEBOOST_net_11716) );
na02s01 TIMEBOOST_cell_37244 ( .a(TIMEBOOST_net_10860), .b(FE_OFN665_n_4495), .o(TIMEBOOST_net_9378) );
na02s01 TIMEBOOST_cell_37246 ( .a(TIMEBOOST_net_10861), .b(FE_OFN665_n_4495), .o(TIMEBOOST_net_9377) );
in01s01 g58369_u0 ( .a(FE_OFN1667_n_9477), .o(g58369_sb) );
na02s01 TIMEBOOST_cell_17424 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__18__Q), .b(g64238_sb), .o(TIMEBOOST_net_3969) );
na02s01 g58369_u2 ( .a(FE_OFN243_n_9116), .b(FE_OFN1667_n_9477), .o(g58369_db) );
na02f02 TIMEBOOST_cell_37102 ( .a(TIMEBOOST_net_10789), .b(n_12572), .o(n_12834) );
in01s01 g58370_u0 ( .a(FE_OFN548_n_9477), .o(g58370_sb) );
na02s01 TIMEBOOST_cell_17426 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__Q), .b(g64240_sb), .o(TIMEBOOST_net_3970) );
na02s01 g58370_u2 ( .a(FE_OFN245_n_9114), .b(FE_OFN548_n_9477), .o(g58370_db) );
na02f02 TIMEBOOST_cell_37104 ( .a(FE_OFN1751_n_12086), .b(TIMEBOOST_net_10790), .o(TIMEBOOST_net_10278) );
in01s01 g58371_u0 ( .a(FE_OFN1668_n_9477), .o(g58371_sb) );
na02s01 TIMEBOOST_cell_9492 ( .a(pci_target_unit_fifos_pciw_addr_data_in_145), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__Q), .o(TIMEBOOST_net_1313) );
na02s01 g58371_u2 ( .a(FE_OFN247_n_9112), .b(FE_OFN1668_n_9477), .o(g58371_db) );
na02s01 TIMEBOOST_cell_9493 ( .a(TIMEBOOST_net_1313), .b(FE_OFN927_n_4730), .o(TIMEBOOST_net_248) );
in01s01 g58372_u0 ( .a(FE_OFN1668_n_9477), .o(g58372_sb) );
na02s01 TIMEBOOST_cell_9494 ( .a(pci_target_unit_fifos_pciw_addr_data_in_128), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__Q), .o(TIMEBOOST_net_1314) );
na02s01 g58372_u2 ( .a(FE_OFN250_n_9789), .b(FE_OFN1668_n_9477), .o(g58372_db) );
na02s01 TIMEBOOST_cell_9495 ( .a(TIMEBOOST_net_1314), .b(FE_OFN927_n_4730), .o(TIMEBOOST_net_249) );
in01s01 g58373_u0 ( .a(FE_OFN1670_n_9477), .o(g58373_sb) );
na02s01 TIMEBOOST_cell_10528 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_31__Q), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_1831) );
na03s02 TIMEBOOST_cell_38337 ( .a(n_4735), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q), .c(FE_OFN1119_g64577_p), .o(TIMEBOOST_net_11407) );
na02s01 TIMEBOOST_cell_10529 ( .a(TIMEBOOST_net_1831), .b(FE_OFN1082_n_13221), .o(TIMEBOOST_net_568) );
in01s01 g58374_u0 ( .a(FE_OFN1666_n_9477), .o(g58374_sb) );
na02s01 TIMEBOOST_cell_9496 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__Q), .b(g65373_sb), .o(TIMEBOOST_net_1315) );
na02s01 g58374_u2 ( .a(FE_OFN254_n_9825), .b(FE_OFN1666_n_9477), .o(g58374_db) );
na02s01 TIMEBOOST_cell_9497 ( .a(TIMEBOOST_net_1315), .b(g65373_db), .o(n_3530) );
in01s01 g58375_u0 ( .a(FE_OFN1635_n_9531), .o(g58375_sb) );
na02s02 TIMEBOOST_cell_42721 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__Q), .b(FE_OFN223_n_9844), .o(TIMEBOOST_net_13599) );
na02s01 TIMEBOOST_cell_9720 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__Q), .b(g65823_sb), .o(TIMEBOOST_net_1427) );
na02s01 TIMEBOOST_cell_9721 ( .a(TIMEBOOST_net_1427), .b(g65823_db), .o(n_1893) );
in01s01 g58376_u0 ( .a(FE_OFN580_n_9531), .o(g58376_sb) );
na02m02 TIMEBOOST_cell_43939 ( .a(n_9024), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__22__Q), .o(TIMEBOOST_net_14208) );
na02s02 TIMEBOOST_cell_37186 ( .a(TIMEBOOST_net_10831), .b(TIMEBOOST_net_3259), .o(TIMEBOOST_net_10091) );
na02s02 TIMEBOOST_cell_37188 ( .a(TIMEBOOST_net_10832), .b(TIMEBOOST_net_1134), .o(TIMEBOOST_net_10089) );
in01s01 g58377_u0 ( .a(FE_OFN579_n_9531), .o(g58377_sb) );
na02f02 TIMEBOOST_cell_43940 ( .a(TIMEBOOST_net_14208), .b(FE_OFN1385_n_8567), .o(TIMEBOOST_net_12802) );
na02m02 TIMEBOOST_cell_37190 ( .a(TIMEBOOST_net_10833), .b(n_2982), .o(TIMEBOOST_net_167) );
na02s01 TIMEBOOST_cell_37880 ( .a(TIMEBOOST_net_11178), .b(g57916_sb), .o(n_9893) );
in01s01 g58378_u0 ( .a(FE_OFN1632_n_9531), .o(g58378_sb) );
na02f02 TIMEBOOST_cell_40235 ( .a(FE_OFN1759_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__Q), .o(TIMEBOOST_net_12356) );
na02s01 g58378_u2 ( .a(FE_OFN209_n_9126), .b(FE_OFN1632_n_9531), .o(g58378_db) );
na02s02 TIMEBOOST_cell_39758 ( .a(TIMEBOOST_net_12117), .b(g62349_sb), .o(n_6902) );
in01s01 g58379_u0 ( .a(FE_OFN580_n_9531), .o(g58379_sb) );
na02s01 g58379_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__Q), .b(g58379_sb), .o(g58379_da) );
na02s01 g58379_u2 ( .a(FE_OFN211_n_9858), .b(FE_OFN580_n_9531), .o(g58379_db) );
na02s01 g58379_u3 ( .a(g58379_da), .b(g58379_db), .o(n_9451) );
in01s01 g58380_u0 ( .a(FE_OFN1634_n_9531), .o(g58380_sb) );
na02f02 TIMEBOOST_cell_38968 ( .a(TIMEBOOST_net_11722), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10716) );
na02s02 TIMEBOOST_cell_39760 ( .a(TIMEBOOST_net_12118), .b(g62413_sb), .o(n_6772) );
in01s01 g58381_u0 ( .a(FE_OFN1634_n_9531), .o(g58381_sb) );
na02s01 TIMEBOOST_cell_9982 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__Q), .b(g65282_sb), .o(TIMEBOOST_net_1558) );
na03s02 TIMEBOOST_cell_38177 ( .a(TIMEBOOST_net_4040), .b(g64319_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__28__Q), .o(TIMEBOOST_net_11327) );
na02f02 TIMEBOOST_cell_38907 ( .a(n_3346), .b(wbu_addr_in_266), .o(TIMEBOOST_net_11692) );
in01s01 g58382_u0 ( .a(FE_OFN1631_n_9531), .o(g58382_sb) );
na02s01 g58382_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__Q), .b(g58382_sb), .o(g58382_da) );
na02s01 g58382_u2 ( .a(FE_OFN217_n_9889), .b(FE_OFN1631_n_9531), .o(g58382_db) );
na02s01 g58382_u3 ( .a(g58382_da), .b(g58382_db), .o(n_9449) );
in01s01 g58383_u0 ( .a(FE_OFN579_n_9531), .o(g58383_sb) );
na02s01 TIMEBOOST_cell_37480 ( .a(TIMEBOOST_net_10978), .b(g65824_sb), .o(TIMEBOOST_net_1682) );
na02s01 g58383_u2 ( .a(FE_OFN219_n_9853), .b(FE_OFN579_n_9531), .o(g58383_db) );
na03s02 TIMEBOOST_cell_43301 ( .a(n_4288), .b(FE_OFN1202_n_4090), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__Q), .o(TIMEBOOST_net_13889) );
in01s01 g58384_u0 ( .a(FE_OFN580_n_9531), .o(g58384_sb) );
na02s01 TIMEBOOST_cell_43302 ( .a(TIMEBOOST_net_13889), .b(g62894_sb), .o(n_6089) );
na02s01 TIMEBOOST_cell_37192 ( .a(TIMEBOOST_net_10834), .b(g65711_db), .o(n_2199) );
na02s01 TIMEBOOST_cell_37194 ( .a(TIMEBOOST_net_10835), .b(g65775_db), .o(n_2192) );
in01s01 g58385_u0 ( .a(FE_OFN580_n_9531), .o(g58385_sb) );
na02s01 TIMEBOOST_cell_37196 ( .a(TIMEBOOST_net_10836), .b(g65678_db), .o(n_2211) );
na02m02 TIMEBOOST_cell_37198 ( .a(TIMEBOOST_net_10837), .b(TIMEBOOST_net_925), .o(TIMEBOOST_net_10710) );
in01s01 g58386_u0 ( .a(FE_OFN1635_n_9531), .o(g58386_sb) );
na02s02 TIMEBOOST_cell_44933 ( .a(FE_OFN231_n_9839), .b(g57932_sb), .o(TIMEBOOST_net_14705) );
na02s01 TIMEBOOST_cell_39458 ( .a(TIMEBOOST_net_11967), .b(g62805_sb), .o(n_5371) );
na02s02 TIMEBOOST_cell_39494 ( .a(TIMEBOOST_net_11985), .b(g63043_sb), .o(n_5166) );
in01s01 g58387_u0 ( .a(FE_OFN1635_n_9531), .o(g58387_sb) );
na02s01 TIMEBOOST_cell_45132 ( .a(TIMEBOOST_net_14804), .b(FE_OFN1125_g64577_p), .o(TIMEBOOST_net_11441) );
na02s01 g58387_u2 ( .a(FE_OFN221_n_9846), .b(FE_OFN1635_n_9531), .o(g58387_db) );
na02s01 TIMEBOOST_cell_39762 ( .a(TIMEBOOST_net_12119), .b(g62508_sb), .o(n_6563) );
in01s01 g58388_u0 ( .a(FE_OFN580_n_9531), .o(g58388_sb) );
na02s01 TIMEBOOST_cell_40506 ( .a(TIMEBOOST_net_12491), .b(FE_OFN1300_n_5763), .o(TIMEBOOST_net_11508) );
na02s01 g58388_u2 ( .a(FE_OFN223_n_9844), .b(FE_OFN580_n_9531), .o(g58388_db) );
na02s02 TIMEBOOST_cell_44934 ( .a(TIMEBOOST_net_14705), .b(g57932_db), .o(n_9878) );
in01s01 g58389_u0 ( .a(FE_OFN580_n_9531), .o(g58389_sb) );
na02s01 g58389_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__22__Q), .b(g58389_sb), .o(g58389_da) );
na02s01 g58389_u2 ( .a(FE_OFN225_n_9122), .b(FE_OFN580_n_9531), .o(g58389_db) );
na02s01 g58389_u3 ( .a(g58389_da), .b(g58389_db), .o(n_9007) );
in01s01 g58390_u0 ( .a(FE_OFN579_n_9531), .o(g58390_sb) );
na02s01 TIMEBOOST_cell_40508 ( .a(TIMEBOOST_net_12492), .b(FE_OFN1301_n_5763), .o(TIMEBOOST_net_11500) );
na02s01 TIMEBOOST_cell_37200 ( .a(TIMEBOOST_net_10838), .b(g65698_db), .o(n_2203) );
na02f04 TIMEBOOST_cell_11925 ( .a(TIMEBOOST_net_2529), .b(FE_RN_705_0), .o(FE_RN_707_0) );
in01s01 g58391_u0 ( .a(FE_OFN579_n_9531), .o(g58391_sb) );
na02s01 TIMEBOOST_cell_40509 ( .a(wishbone_slave_unit_pcim_sm_data_in_657), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__Q), .o(TIMEBOOST_net_12493) );
na02s01 g58391_u2 ( .a(FE_OFN227_n_9841), .b(FE_OFN579_n_9531), .o(g58391_db) );
na02s01 TIMEBOOST_cell_40510 ( .a(TIMEBOOST_net_12493), .b(FE_OFN1301_n_5763), .o(TIMEBOOST_net_11501) );
in01s01 g58392_u0 ( .a(FE_OFN1632_n_9531), .o(g58392_sb) );
na02s02 TIMEBOOST_cell_31468 ( .a(n_4493), .b(g64760_sb), .o(TIMEBOOST_net_9645) );
na02s01 g58392_u2 ( .a(FE_OFN229_n_9120), .b(FE_OFN1632_n_9531), .o(g58392_db) );
in01s01 g58393_u0 ( .a(FE_OFN580_n_9531), .o(g58393_sb) );
na02s01 g58393_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__Q), .b(g58393_sb), .o(g58393_da) );
na02s01 g58393_u2 ( .a(FE_OFN233_n_9876), .b(FE_OFN580_n_9531), .o(g58393_db) );
na02s01 g58393_u3 ( .a(g58393_da), .b(g58393_db), .o(n_9440) );
in01s01 g58394_u0 ( .a(FE_OFN1635_n_9531), .o(g58394_sb) );
na02m02 TIMEBOOST_cell_9988 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__Q), .b(n_13447), .o(TIMEBOOST_net_1561) );
na02s01 TIMEBOOST_cell_39335 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q), .b(g64230_sb), .o(TIMEBOOST_net_11906) );
na02f02 TIMEBOOST_cell_44518 ( .a(TIMEBOOST_net_14497), .b(FE_OFN2170_n_8567), .o(TIMEBOOST_net_13013) );
in01s01 g58395_u0 ( .a(FE_OFN580_n_9531), .o(g58395_sb) );
na02s01 TIMEBOOST_cell_44935 ( .a(FE_OFN215_n_9856), .b(g58144_sb), .o(TIMEBOOST_net_14706) );
na02s01 TIMEBOOST_cell_9722 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__Q), .b(g65819_sb), .o(TIMEBOOST_net_1428) );
na02s01 TIMEBOOST_cell_9723 ( .a(TIMEBOOST_net_1428), .b(g65819_db), .o(n_1897) );
in01s01 g58396_u0 ( .a(FE_OFN580_n_9531), .o(g58396_sb) );
na03f02 TIMEBOOST_cell_35989 ( .a(TIMEBOOST_net_10121), .b(n_13617), .c(g54490_sb), .o(n_13605) );
na02s01 g58396_u2 ( .a(FE_OFN237_n_9118), .b(FE_OFN1632_n_9531), .o(g58396_db) );
na02s02 TIMEBOOST_cell_39764 ( .a(TIMEBOOST_net_12120), .b(g62639_sb), .o(n_6271) );
in01s01 g58397_u0 ( .a(FE_OFN580_n_9531), .o(g58397_sb) );
na02s01 g58397_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__Q), .b(g58397_sb), .o(g58397_da) );
na02s01 g58397_u2 ( .a(FE_OFN239_n_9832), .b(FE_OFN580_n_9531), .o(g58397_db) );
na02s01 g58397_u3 ( .a(g58397_da), .b(g58397_db), .o(n_9437) );
in01s01 g58398_u0 ( .a(FE_OFN1634_n_9531), .o(g58398_sb) );
na02s01 TIMEBOOST_cell_42686 ( .a(TIMEBOOST_net_13581), .b(g64184_db), .o(n_3982) );
na02s01 g58398_u2 ( .a(FE_OFN241_n_9830), .b(FE_OFN1634_n_9531), .o(g58398_db) );
na02s02 TIMEBOOST_cell_45184 ( .a(TIMEBOOST_net_14830), .b(FE_OFN1275_n_4096), .o(TIMEBOOST_net_12642) );
in01s01 g58399_u0 ( .a(FE_OFN1631_n_9531), .o(g58399_sb) );
na02s01 g58399_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__Q), .b(g58399_sb), .o(g58399_da) );
na02s01 g58399_u2 ( .a(FE_OFN201_n_9230), .b(FE_OFN1631_n_9531), .o(g58399_db) );
na02s01 g58399_u3 ( .a(g58399_da), .b(g58399_db), .o(n_9209) );
in01s01 g58400_u0 ( .a(FE_OFN1634_n_9531), .o(g58400_sb) );
na02m02 TIMEBOOST_cell_9992 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__Q), .b(n_13447), .o(TIMEBOOST_net_1563) );
na02s02 TIMEBOOST_cell_38206 ( .a(TIMEBOOST_net_11341), .b(FE_OFN1135_g64577_p), .o(TIMEBOOST_net_4681) );
na02f02 TIMEBOOST_cell_44166 ( .a(TIMEBOOST_net_14321), .b(FE_OFN1376_n_8567), .o(TIMEBOOST_net_13392) );
in01s01 g58401_u0 ( .a(FE_OFN1631_n_9531), .o(g58401_sb) );
na02s01 TIMEBOOST_cell_44936 ( .a(TIMEBOOST_net_14706), .b(g58144_db), .o(n_9651) );
na02s02 TIMEBOOST_cell_40869 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__Q), .b(n_13180), .o(TIMEBOOST_net_12673) );
na02s01 TIMEBOOST_cell_40630 ( .a(TIMEBOOST_net_12553), .b(g63162_sb), .o(n_5812) );
in01s01 g58402_u0 ( .a(FE_OFN1631_n_9531), .o(g58402_sb) );
na02s01 TIMEBOOST_cell_42942 ( .a(TIMEBOOST_net_13709), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_11177) );
na02s02 TIMEBOOST_cell_40849 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__Q), .b(n_13169), .o(TIMEBOOST_net_12663) );
in01s01 g58403_u0 ( .a(FE_OFN579_n_9531), .o(g58403_sb) );
na02s02 TIMEBOOST_cell_39766 ( .a(TIMEBOOST_net_12121), .b(g62514_sb), .o(n_6550) );
na02s01 TIMEBOOST_cell_37726 ( .a(TIMEBOOST_net_11101), .b(g62070_sb), .o(n_7828) );
na02s02 TIMEBOOST_cell_16784 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_28__Q), .b(n_8884), .o(TIMEBOOST_net_3649) );
in01s01 g58404_u0 ( .a(FE_OFN580_n_9531), .o(g58404_sb) );
na02s01 g58404_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__Q), .b(g58404_sb), .o(g58404_da) );
na02s01 g58404_u2 ( .a(FE_OFN243_n_9116), .b(FE_OFN580_n_9531), .o(g58404_db) );
na02s01 g58404_u3 ( .a(g58404_da), .b(g58404_db), .o(n_9003) );
in01s01 g58405_u0 ( .a(FE_OFN1634_n_9531), .o(g58405_sb) );
na02m02 TIMEBOOST_cell_9994 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__Q), .b(n_13447), .o(TIMEBOOST_net_1564) );
na02s01 TIMEBOOST_cell_18034 ( .a(pci_target_unit_fifos_pciw_addr_data_in_128), .b(g64081_sb), .o(TIMEBOOST_net_4274) );
na02f02 TIMEBOOST_cell_9995 ( .a(TIMEBOOST_net_1564), .b(FE_OFN1150_n_13249), .o(TIMEBOOST_net_477) );
in01s01 g58406_u0 ( .a(FE_OFN1632_n_9531), .o(g58406_sb) );
na02s02 TIMEBOOST_cell_16350 ( .a(n_3752), .b(g64833_sb), .o(TIMEBOOST_net_3432) );
na02s01 g58406_u2 ( .a(FE_OFN247_n_9112), .b(FE_OFN1632_n_9531), .o(g58406_db) );
na02s02 TIMEBOOST_cell_16351 ( .a(TIMEBOOST_net_3432), .b(g64833_db), .o(n_3730) );
in01s01 g58407_u0 ( .a(FE_OFN1635_n_9531), .o(g58407_sb) );
na02m02 TIMEBOOST_cell_9996 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__Q), .b(n_13447), .o(TIMEBOOST_net_1565) );
na02s01 TIMEBOOST_cell_43075 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__Q), .b(n_3607), .o(TIMEBOOST_net_13776) );
na02s02 TIMEBOOST_cell_44421 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_796), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_31__Q), .o(TIMEBOOST_net_14449) );
in01s01 g58408_u0 ( .a(FE_OFN579_n_9531), .o(g58408_sb) );
na02m02 TIMEBOOST_cell_38977 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_22__Q), .o(TIMEBOOST_net_11727) );
na02s01 TIMEBOOST_cell_9724 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__Q), .b(g65811_sb), .o(TIMEBOOST_net_1429) );
na02s01 TIMEBOOST_cell_9725 ( .a(TIMEBOOST_net_1429), .b(g65811_db), .o(n_1903) );
in01s01 g58409_u0 ( .a(FE_OFN1656_n_9502), .o(g58409_sb) );
na02f02 TIMEBOOST_cell_39128 ( .a(TIMEBOOST_net_11802), .b(FE_OFN1600_n_13995), .o(n_16249) );
na02s01 g58409_u2 ( .a(FE_OFN215_n_9856), .b(FE_OFN1656_n_9502), .o(g58409_db) );
na02s01 TIMEBOOST_cell_17809 ( .a(TIMEBOOST_net_4161), .b(g61747_sb), .o(n_8323) );
in01s01 g58410_u0 ( .a(FE_OFN519_n_9697), .o(g58410_sb) );
na02s02 TIMEBOOST_cell_38425 ( .a(n_1293), .b(g63571_db), .o(TIMEBOOST_net_11451) );
na02s01 g58410_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__Q), .b(FE_OFN519_n_9697), .o(g58410_db) );
na02f02 TIMEBOOST_cell_38970 ( .a(TIMEBOOST_net_11723), .b(FE_OFN2156_n_16439), .o(TIMEBOOST_net_10717) );
in01s01 g58411_u0 ( .a(FE_OFN518_n_9697), .o(g58411_sb) );
na02s01 g58411_u1 ( .a(FE_OFN203_n_9228), .b(g58411_sb), .o(g58411_da) );
na02s01 g58411_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__Q), .b(FE_OFN518_n_9697), .o(g58411_db) );
na02s01 g58411_u3 ( .a(g58411_da), .b(g58411_db), .o(n_9206) );
in01s01 g58412_u0 ( .a(FE_OFN587_n_9692), .o(g58412_sb) );
na02m08 TIMEBOOST_cell_42544 ( .a(TIMEBOOST_net_13510), .b(g67082_sb), .o(TIMEBOOST_net_3206) );
na02s01 g58412_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__Q), .b(FE_OFN587_n_9692), .o(g58412_db) );
na03s02 TIMEBOOST_cell_38099 ( .a(TIMEBOOST_net_3967), .b(g60687_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__Q), .o(TIMEBOOST_net_11288) );
in01s01 g58413_u0 ( .a(FE_OFN589_n_9692), .o(g58413_sb) );
na02m02 TIMEBOOST_cell_42545 ( .a(n_13447), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__Q), .o(TIMEBOOST_net_13511) );
na02s01 g58413_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__Q), .b(FE_OFN589_n_9692), .o(g58413_db) );
na02s02 TIMEBOOST_cell_19341 ( .a(TIMEBOOST_net_4927), .b(g60637_sb), .o(n_5696) );
in01s01 g58414_u0 ( .a(FE_OFN587_n_9692), .o(g58414_sb) );
na02s01 TIMEBOOST_cell_16261 ( .a(TIMEBOOST_net_3387), .b(g65099_db), .o(n_3594) );
na02s01 g58414_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__Q), .b(FE_OFN587_n_9692), .o(g58414_db) );
na02s01 TIMEBOOST_cell_16262 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(g65668_sb), .o(TIMEBOOST_net_3388) );
in01s01 g58415_u0 ( .a(FE_OFN595_n_9694), .o(g58415_sb) );
in01s01 TIMEBOOST_cell_45892 ( .a(TIMEBOOST_net_15198), .o(TIMEBOOST_net_15199) );
na02s01 g58415_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__Q), .b(FE_OFN595_n_9694), .o(g58415_db) );
na02s01 TIMEBOOST_cell_38050 ( .a(TIMEBOOST_net_11263), .b(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_4591) );
in01s01 g58416_u0 ( .a(FE_OFN597_n_9694), .o(g58416_sb) );
na02s01 g58416_u1 ( .a(FE_OFN203_n_9228), .b(g58416_sb), .o(g58416_da) );
na02s01 g58416_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__Q), .b(FE_OFN597_n_9694), .o(g58416_db) );
na02s01 g58416_u3 ( .a(g58416_da), .b(g58416_db), .o(n_9202) );
in01s01 g58417_u0 ( .a(FE_OFN595_n_9694), .o(g58417_sb) );
na03s02 TIMEBOOST_cell_40633 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__Q), .b(n_4326), .c(FE_OFN1212_n_4151), .o(TIMEBOOST_net_12555) );
na02s01 g58417_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__34__Q), .b(FE_OFN595_n_9694), .o(g58417_db) );
na02s02 TIMEBOOST_cell_40870 ( .a(TIMEBOOST_net_12673), .b(FE_OFN1331_n_13547), .o(TIMEBOOST_net_11609) );
in01s01 g58418_u0 ( .a(FE_OFN1655_n_9502), .o(g58418_sb) );
na02s01 TIMEBOOST_cell_16352 ( .a(n_3780), .b(g64840_sb), .o(TIMEBOOST_net_3433) );
na02s01 g58418_u2 ( .a(FE_OFN237_n_9118), .b(FE_OFN1655_n_9502), .o(g58418_db) );
na02s01 TIMEBOOST_cell_16353 ( .a(TIMEBOOST_net_3433), .b(g64840_db), .o(n_3727) );
in01s01 g58419_u0 ( .a(FE_OFN1651_n_9428), .o(g58419_sb) );
na02s02 TIMEBOOST_cell_45722 ( .a(TIMEBOOST_net_15099), .b(FE_OFN1283_n_4097), .o(TIMEBOOST_net_12609) );
na02s01 g58419_u2 ( .a(FE_OFN207_n_9865), .b(FE_OFN1651_n_9428), .o(g58419_db) );
na02s02 TIMEBOOST_cell_16354 ( .a(n_3747), .b(g64899_sb), .o(TIMEBOOST_net_3434) );
in01s01 g58420_u0 ( .a(FE_OFN1650_n_9428), .o(g58420_sb) );
na02s01 TIMEBOOST_cell_16355 ( .a(TIMEBOOST_net_3434), .b(g64899_db), .o(n_3694) );
na02s01 TIMEBOOST_cell_20073 ( .a(TIMEBOOST_net_5293), .b(FE_OFN1125_g64577_p), .o(n_5474) );
na02s02 TIMEBOOST_cell_39768 ( .a(TIMEBOOST_net_12122), .b(g62418_sb), .o(n_6761) );
in01s01 g58421_u0 ( .a(FE_OFN523_n_9428), .o(g58421_sb) );
na02s02 TIMEBOOST_cell_16356 ( .a(n_3761), .b(g64900_sb), .o(TIMEBOOST_net_3435) );
na02s02 TIMEBOOST_cell_39770 ( .a(TIMEBOOST_net_12123), .b(g62713_sb), .o(n_6144) );
na02f02 TIMEBOOST_cell_36938 ( .a(TIMEBOOST_net_10707), .b(g52610_sb), .o(n_10199) );
in01s01 g58422_u0 ( .a(FE_OFN1648_n_9428), .o(g58422_sb) );
na02s01 TIMEBOOST_cell_16357 ( .a(TIMEBOOST_net_3435), .b(g64900_db), .o(n_3693) );
na02m02 TIMEBOOST_cell_45034 ( .a(TIMEBOOST_net_14755), .b(g59383_db), .o(n_4204) );
na02s01 TIMEBOOST_cell_16358 ( .a(n_3752), .b(g64906_sb), .o(TIMEBOOST_net_3436) );
in01s01 g58423_u0 ( .a(FE_OFN1650_n_9428), .o(g58423_sb) );
na02s01 g58423_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q), .b(g58423_sb), .o(g58423_da) );
na02s01 g58423_u2 ( .a(FE_OFN213_n_9124), .b(FE_OFN1650_n_9428), .o(g58423_db) );
na02s01 g58423_u3 ( .a(g58423_da), .b(g58423_db), .o(n_8997) );
in01s01 g58424_u0 ( .a(FE_OFN1650_n_9428), .o(g58424_sb) );
na02s01 g58424_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__15__Q), .b(g58424_sb), .o(g58424_da) );
na02s02 TIMEBOOST_cell_38647 ( .a(n_4024), .b(g62777_sb), .o(TIMEBOOST_net_11562) );
na02s01 TIMEBOOST_cell_39326 ( .a(TIMEBOOST_net_11901), .b(FE_OFN239_n_9832), .o(TIMEBOOST_net_11014) );
in01s01 g58425_u0 ( .a(FE_OFN523_n_9428), .o(g58425_sb) );
na02f02 TIMEBOOST_cell_36948 ( .a(TIMEBOOST_net_10712), .b(g58807_sb), .o(n_8634) );
na02s01 g58425_u2 ( .a(FE_OFN219_n_9853), .b(FE_OFN523_n_9428), .o(g58425_db) );
na02s01 TIMEBOOST_cell_31464 ( .a(FE_OFN205_n_9140), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__Q), .o(TIMEBOOST_net_9643) );
in01s01 g58426_u0 ( .a(FE_OFN1648_n_9428), .o(g58426_sb) );
na02s01 TIMEBOOST_cell_16359 ( .a(TIMEBOOST_net_3436), .b(g64906_db), .o(n_3690) );
na02f02 TIMEBOOST_cell_37082 ( .a(TIMEBOOST_net_10779), .b(FE_OFN1587_n_13736), .o(g53301_p) );
na02s02 TIMEBOOST_cell_38052 ( .a(TIMEBOOST_net_11264), .b(FE_OFN1135_g64577_p), .o(TIMEBOOST_net_4575) );
in01s01 g58427_u0 ( .a(FE_OFN1649_n_9428), .o(g58427_sb) );
na02s01 TIMEBOOST_cell_16360 ( .a(n_3749), .b(g64907_sb), .o(TIMEBOOST_net_3437) );
na02f02 TIMEBOOST_cell_36896 ( .a(TIMEBOOST_net_10686), .b(g58607_sb), .o(n_8900) );
na02f02 TIMEBOOST_cell_11947 ( .a(TIMEBOOST_net_2540), .b(n_8897), .o(n_9932) );
in01s01 g58428_u0 ( .a(FE_OFN1650_n_9428), .o(g58428_sb) );
na02s01 g58428_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__Q), .b(g58428_sb), .o(g58428_da) );
na02s01 g58428_u2 ( .a(FE_OFN221_n_9846), .b(FE_OFN1650_n_9428), .o(g58428_db) );
na02s01 g58428_u3 ( .a(g58428_da), .b(g58428_db), .o(n_9419) );
in01s01 g58429_u0 ( .a(FE_OFN1649_n_9428), .o(g58429_sb) );
na02s01 TIMEBOOST_cell_36519 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__Q), .b(FE_OFN555_n_9864), .o(TIMEBOOST_net_10498) );
na02s01 g58429_u2 ( .a(FE_OFN223_n_9844), .b(FE_OFN1649_n_9428), .o(g58429_db) );
na02s01 TIMEBOOST_cell_36518 ( .a(TIMEBOOST_net_10497), .b(FE_OFN223_n_9844), .o(n_9575) );
in01s01 g58430_u0 ( .a(FE_OFN1648_n_9428), .o(g58430_sb) );
na02s01 TIMEBOOST_cell_31461 ( .a(TIMEBOOST_net_9641), .b(g64973_sb), .o(n_4370) );
na02s01 g58430_u2 ( .a(FE_OFN225_n_9122), .b(FE_OFN1648_n_9428), .o(g58430_db) );
na02s01 TIMEBOOST_cell_36475 ( .a(TIMEBOOST_net_3332), .b(FE_OFN1003_n_2047), .o(TIMEBOOST_net_10476) );
in01s01 g58431_u0 ( .a(FE_OFN1648_n_9428), .o(g58431_sb) );
na02s02 TIMEBOOST_cell_31459 ( .a(TIMEBOOST_net_9640), .b(g64965_sb), .o(n_3655) );
na02s01 g58431_u2 ( .a(FE_OFN227_n_9841), .b(FE_OFN1648_n_9428), .o(g58431_db) );
na02s01 TIMEBOOST_cell_36473 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(g65763_db), .o(TIMEBOOST_net_10475) );
in01s01 g58432_u0 ( .a(FE_OFN1649_n_9428), .o(g58432_sb) );
na02s02 TIMEBOOST_cell_39772 ( .a(TIMEBOOST_net_12124), .b(g62711_sb), .o(n_6148) );
na02s01 g58432_u2 ( .a(FE_OFN229_n_9120), .b(FE_OFN1649_n_9428), .o(g58432_db) );
na02s02 TIMEBOOST_cell_40311 ( .a(g64804_sb), .b(g64804_db), .o(TIMEBOOST_net_12394) );
in01s01 g58433_u0 ( .a(FE_OFN1648_n_9428), .o(g58433_sb) );
na02s01 g58433_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__Q), .b(g58433_sb), .o(g58433_da) );
na02s01 g58433_u2 ( .a(FE_OFN231_n_9839), .b(FE_OFN1648_n_9428), .o(g58433_db) );
na02s02 g58433_u3 ( .a(g58433_da), .b(g58433_db), .o(n_9415) );
in01s01 g58434_u0 ( .a(FE_OFN1650_n_9428), .o(g58434_sb) );
na02s02 TIMEBOOST_cell_39774 ( .a(TIMEBOOST_net_12125), .b(g62584_sb), .o(n_6384) );
na02f02 TIMEBOOST_cell_37084 ( .a(TIMEBOOST_net_10780), .b(FE_OFN1587_n_13736), .o(g53255_p) );
na02f02 TIMEBOOST_cell_37086 ( .a(TIMEBOOST_net_10781), .b(FE_OFN1588_n_13736), .o(g53235_p) );
in01s01 g58435_u0 ( .a(FE_OFN1648_n_9428), .o(g58435_sb) );
na02s01 g58435_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__29__Q), .b(g58435_sb), .o(g58435_da) );
na02s01 g58435_u2 ( .a(FE_OFN235_n_9834), .b(FE_OFN1648_n_9428), .o(g58435_db) );
na02s02 g58435_u3 ( .a(g58435_da), .b(g58435_db), .o(n_9413) );
in01s01 g58436_u0 ( .a(FE_OFN1649_n_9428), .o(g58436_sb) );
na02s01 g58436_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__Q), .b(g58436_sb), .o(g58436_da) );
na02s01 g58436_u2 ( .a(FE_OFN237_n_9118), .b(FE_OFN1649_n_9428), .o(g58436_db) );
na02s01 g58436_u3 ( .a(g58436_da), .b(g58436_db), .o(n_8994) );
in01s01 g58437_u0 ( .a(FE_OFN1650_n_9428), .o(g58437_sb) );
na02s01 g58437_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__31__Q), .b(g58437_sb), .o(g58437_da) );
na02s01 g58437_u2 ( .a(FE_OFN241_n_9830), .b(FE_OFN1650_n_9428), .o(g58437_db) );
na02s02 TIMEBOOST_cell_37934 ( .a(TIMEBOOST_net_11205), .b(g58343_sb), .o(n_9476) );
in01s01 g58438_u0 ( .a(FE_OFN1651_n_9428), .o(g58438_sb) );
na02s01 TIMEBOOST_cell_44937 ( .a(FE_OFN213_n_9124), .b(g58074_sb), .o(TIMEBOOST_net_14707) );
na03s02 TIMEBOOST_cell_38185 ( .a(TIMEBOOST_net_4075), .b(g64236_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__Q), .o(TIMEBOOST_net_11331) );
na02s02 TIMEBOOST_cell_43482 ( .a(TIMEBOOST_net_13979), .b(FE_OFN1234_n_6391), .o(TIMEBOOST_net_12186) );
in01s01 g58439_u0 ( .a(FE_OFN1650_n_9428), .o(g58439_sb) );
na02s01 TIMEBOOST_cell_31278 ( .a(configuration_wb_err_cs_bit_564), .b(conf_wb_err_bc_in_846), .o(TIMEBOOST_net_9550) );
na02s01 g58439_u2 ( .a(FE_OFN203_n_9228), .b(FE_OFN1650_n_9428), .o(g58439_db) );
na02s02 TIMEBOOST_cell_43485 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__Q), .b(n_4299), .o(TIMEBOOST_net_13981) );
in01s01 g58440_u0 ( .a(FE_OFN1651_n_9428), .o(g58440_sb) );
na02m02 TIMEBOOST_cell_38740 ( .a(TIMEBOOST_net_11608), .b(g53908_sb), .o(n_13533) );
na02s01 TIMEBOOST_cell_9206 ( .a(pci_target_unit_fifos_pcir_data_in_163), .b(g65803_sb), .o(TIMEBOOST_net_1170) );
na02s01 TIMEBOOST_cell_9207 ( .a(TIMEBOOST_net_1170), .b(g65803_db), .o(n_2187) );
in01s01 g58441_u0 ( .a(FE_OFN523_n_9428), .o(g58441_sb) );
na02s02 TIMEBOOST_cell_39776 ( .a(TIMEBOOST_net_12126), .b(g62438_sb), .o(n_6720) );
na02s01 TIMEBOOST_cell_17976 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(g64205_sb), .o(TIMEBOOST_net_4245) );
na02f02 TIMEBOOST_cell_37088 ( .a(TIMEBOOST_net_10782), .b(FE_OFN1589_n_13736), .o(g53174_p) );
in01s01 g58442_u0 ( .a(FE_OFN1650_n_9428), .o(g58442_sb) );
na02s01 g58442_u2 ( .a(FE_OFN245_n_9114), .b(FE_OFN1650_n_9428), .o(g58442_db) );
na02s01 TIMEBOOST_cell_31276 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__Q), .o(TIMEBOOST_net_9549) );
in01s01 g58443_u0 ( .a(FE_OFN1649_n_9428), .o(g58443_sb) );
na02s01 g58443_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__Q), .b(g58443_sb), .o(g58443_da) );
na02s01 g58443_u2 ( .a(FE_OFN247_n_9112), .b(FE_OFN1649_n_9428), .o(g58443_db) );
na02s01 g58443_u3 ( .a(g58443_da), .b(g58443_db), .o(n_8992) );
in01s01 g58444_u0 ( .a(FE_OFN523_n_9428), .o(g58444_sb) );
na02s02 TIMEBOOST_cell_42915 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q), .b(FE_OFN1654_n_9502), .o(TIMEBOOST_net_13696) );
na02s01 g58444_u2 ( .a(FE_OFN250_n_9789), .b(FE_OFN523_n_9428), .o(g58444_db) );
na02s01 TIMEBOOST_cell_31274 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__Q), .o(TIMEBOOST_net_9548) );
in01s01 g58445_u0 ( .a(FE_OFN523_n_9428), .o(g58445_sb) );
na02s01 g58445_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__Q), .b(g58445_sb), .o(g58445_da) );
na02s01 g58445_u2 ( .a(FE_OFN254_n_9825), .b(FE_OFN523_n_9428), .o(g58445_db) );
na02s02 g58445_u3 ( .a(g58445_da), .b(g58445_db), .o(n_9408) );
in01s01 g58446_u0 ( .a(FE_OFN1801_n_9690), .o(g58446_sb) );
na02s01 TIMEBOOST_cell_39436 ( .a(TIMEBOOST_net_11956), .b(g61990_sb), .o(n_7915) );
na02m02 TIMEBOOST_cell_43002 ( .a(TIMEBOOST_net_13739), .b(TIMEBOOST_net_341), .o(TIMEBOOST_net_4780) );
na02s01 TIMEBOOST_cell_37248 ( .a(TIMEBOOST_net_10862), .b(FE_OFN665_n_4495), .o(TIMEBOOST_net_9376) );
in01s01 g58447_u0 ( .a(FE_OFN543_n_9690), .o(g58447_sb) );
na02s01 g58447_u1 ( .a(FE_OFN203_n_9228), .b(g58447_sb), .o(g58447_da) );
na02s01 g58447_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__Q), .b(FE_OFN543_n_9690), .o(g58447_db) );
na02s01 g58447_u3 ( .a(g58447_da), .b(g58447_db), .o(n_9198) );
in01s01 g58448_u0 ( .a(FE_OFN548_n_9477), .o(g58448_sb) );
na02s01 TIMEBOOST_cell_9498 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__Q), .o(TIMEBOOST_net_1316) );
na02s01 g58448_u2 ( .a(FE_OFN203_n_9228), .b(FE_OFN548_n_9477), .o(g58448_db) );
na02s01 TIMEBOOST_cell_9499 ( .a(TIMEBOOST_net_1316), .b(FE_OFN1017_n_2053), .o(TIMEBOOST_net_247) );
in01s01 g58449_u0 ( .a(FE_OFN1648_n_9428), .o(g58449_sb) );
na02s01 g58449_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q), .b(g58449_sb), .o(g58449_da) );
na02s01 g58449_u2 ( .a(FE_OFN233_n_9876), .b(FE_OFN1648_n_9428), .o(g58449_db) );
na02s01 g58449_u3 ( .a(g58449_da), .b(g58449_db), .o(n_9407) );
in01s01 g58450_u0 ( .a(FE_OFN1648_n_9428), .o(g58450_sb) );
na02s02 TIMEBOOST_cell_31273 ( .a(TIMEBOOST_net_9547), .b(FE_OFN948_n_2248), .o(TIMEBOOST_net_4022) );
na02f02 TIMEBOOST_cell_37062 ( .a(TIMEBOOST_net_10769), .b(n_12565), .o(n_12827) );
na02f02 TIMEBOOST_cell_37064 ( .a(TIMEBOOST_net_10770), .b(n_12566), .o(n_12828) );
in01s01 g58451_u0 ( .a(FE_OFN1649_n_9428), .o(g58451_sb) );
na03s02 TIMEBOOST_cell_8376 ( .a(TIMEBOOST_net_597), .b(n_8568), .c(n_8570), .o(n_8843) );
na02s01 g58451_u2 ( .a(FE_OFN209_n_9126), .b(FE_OFN1649_n_9428), .o(g58451_db) );
na02s01 TIMEBOOST_cell_31103 ( .a(TIMEBOOST_net_9462), .b(g64815_db), .o(n_3743) );
in01s01 g58452_u0 ( .a(FE_OFN1651_n_9428), .o(g58452_sb) );
na02s02 TIMEBOOST_cell_31263 ( .a(TIMEBOOST_net_9542), .b(FE_OFN948_n_2248), .o(TIMEBOOST_net_4017) );
na02s01 g58452_u2 ( .a(FE_OFN252_n_9868), .b(FE_OFN1651_n_9428), .o(g58452_db) );
na02s02 TIMEBOOST_cell_16564 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(g65672_sb), .o(TIMEBOOST_net_3539) );
in01s01 g58453_u0 ( .a(FE_OFN1651_n_9428), .o(g58453_sb) );
na02s01 TIMEBOOST_cell_31252 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__21__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_141), .o(TIMEBOOST_net_9537) );
na02s01 g58453_u2 ( .a(FE_OFN217_n_9889), .b(FE_OFN1651_n_9428), .o(g58453_db) );
na02s01 TIMEBOOST_cell_31251 ( .a(TIMEBOOST_net_9536), .b(g65048_db), .o(n_4324) );
in01s01 g58454_u0 ( .a(FE_OFN1649_n_9428), .o(g58454_sb) );
na02s01 TIMEBOOST_cell_31250 ( .a(n_4465), .b(g65048_sb), .o(TIMEBOOST_net_9536) );
na02s01 g58454_u2 ( .a(FE_OFN243_n_9116), .b(FE_OFN1649_n_9428), .o(g58454_db) );
na02s01 TIMEBOOST_cell_31249 ( .a(TIMEBOOST_net_9535), .b(g64757_db), .o(n_4499) );
in01m02 g58455_u0 ( .a(FE_OFN1437_n_9372), .o(g58455_sb) );
na02f02 TIMEBOOST_cell_41376 ( .a(TIMEBOOST_net_12926), .b(g57589_sb), .o(n_11162) );
na02m02 TIMEBOOST_cell_43941 ( .a(n_9085), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__Q), .o(TIMEBOOST_net_14209) );
na02s01 TIMEBOOST_cell_40632 ( .a(TIMEBOOST_net_12554), .b(g63153_sb), .o(n_5836) );
in01m02 g58456_u0 ( .a(FE_OFN1436_n_9372), .o(g58456_sb) );
na02m02 TIMEBOOST_cell_32756 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__Q), .o(TIMEBOOST_net_10289) );
na02s01 TIMEBOOST_cell_15882 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_79), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3198) );
na02s01 TIMEBOOST_cell_15883 ( .a(TIMEBOOST_net_3198), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_392), .o(TIMEBOOST_net_84) );
in01m02 g58457_u0 ( .a(FE_OFN1440_n_9372), .o(g58457_sb) );
na02f02 TIMEBOOST_cell_32755 ( .a(FE_OFN1741_n_11019), .b(TIMEBOOST_net_10288), .o(TIMEBOOST_net_6532) );
na02s01 TIMEBOOST_cell_15884 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_88), .b(FE_OFN2119_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3199) );
na02s02 TIMEBOOST_cell_44849 ( .a(n_3780), .b(g64768_sb), .o(TIMEBOOST_net_14663) );
in01m02 g58458_u0 ( .a(FE_OFN1440_n_9372), .o(g58458_sb) );
na02m02 TIMEBOOST_cell_32754 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__Q), .o(TIMEBOOST_net_10288) );
na02f04 TIMEBOOST_cell_41674 ( .a(TIMEBOOST_net_13075), .b(n_9992), .o(n_12135) );
na02s01 TIMEBOOST_cell_15846 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_95), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3180) );
in01m02 g58459_u0 ( .a(FE_OFN1439_n_9372), .o(g58459_sb) );
na02f02 TIMEBOOST_cell_32753 ( .a(FE_OFN1742_n_11019), .b(TIMEBOOST_net_10287), .o(TIMEBOOST_net_6531) );
na02f02 TIMEBOOST_cell_43942 ( .a(TIMEBOOST_net_14209), .b(FE_OFN1407_n_8567), .o(TIMEBOOST_net_12800) );
na02s01 TIMEBOOST_cell_15847 ( .a(TIMEBOOST_net_3180), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_408), .o(TIMEBOOST_net_85) );
in01m02 g58460_u0 ( .a(FE_OFN1436_n_9372), .o(g58460_sb) );
na02m02 TIMEBOOST_cell_32752 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q), .o(TIMEBOOST_net_10287) );
na02f02 TIMEBOOST_cell_41675 ( .a(n_14895), .b(n_13485), .o(TIMEBOOST_net_13076) );
na03s02 TIMEBOOST_cell_40635 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__5__Q), .b(n_3756), .c(FE_OFN1207_n_6356), .o(TIMEBOOST_net_12556) );
in01m02 g58461_u0 ( .a(FE_OFN1436_n_9372), .o(g58461_sb) );
na02f02 TIMEBOOST_cell_32751 ( .a(FE_OFN1742_n_11019), .b(TIMEBOOST_net_10286), .o(TIMEBOOST_net_6530) );
na02f02 TIMEBOOST_cell_43757 ( .a(n_9052), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__Q), .o(TIMEBOOST_net_14117) );
na02s02 TIMEBOOST_cell_40634 ( .a(TIMEBOOST_net_12555), .b(g62659_sb), .o(n_6226) );
in01m02 g58462_u0 ( .a(FE_OFN1436_n_9372), .o(g58462_sb) );
na02m02 TIMEBOOST_cell_32750 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__Q), .o(TIMEBOOST_net_10286) );
in01s01 TIMEBOOST_cell_32830 ( .a(TIMEBOOST_net_10331), .o(wbs_dat_i_10_) );
in01m02 g58463_u0 ( .a(FE_OFN1441_n_9372), .o(g58463_sb) );
na02f02 TIMEBOOST_cell_41378 ( .a(TIMEBOOST_net_12927), .b(g57462_sb), .o(n_11271) );
na02m02 TIMEBOOST_cell_42546 ( .a(TIMEBOOST_net_13511), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_396), .o(TIMEBOOST_net_9656) );
na02m02 TIMEBOOST_cell_42547 ( .a(n_13447), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__Q), .o(TIMEBOOST_net_13512) );
in01f02 g58464_u0 ( .a(FE_OFN1439_n_9372), .o(g58464_sb) );
na02m02 TIMEBOOST_cell_32748 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__Q), .o(TIMEBOOST_net_10285) );
na02f02 TIMEBOOST_cell_44750 ( .a(TIMEBOOST_net_14613), .b(n_12366), .o(n_12664) );
na02s02 TIMEBOOST_cell_32015 ( .a(TIMEBOOST_net_9918), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4900) );
in01m02 g58465_u0 ( .a(FE_OFN1441_n_9372), .o(g58465_sb) );
na02f02 TIMEBOOST_cell_32747 ( .a(FE_OFN1742_n_11019), .b(TIMEBOOST_net_10284), .o(TIMEBOOST_net_6528) );
na03s02 TIMEBOOST_cell_43303 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__Q), .b(n_3543), .c(FE_OFN1213_n_4151), .o(TIMEBOOST_net_13890) );
na02f02 TIMEBOOST_cell_41130 ( .a(TIMEBOOST_net_12803), .b(g57294_sb), .o(n_11458) );
in01m02 g58466_u0 ( .a(FE_OFN1437_n_9372), .o(g58466_sb) );
na02m02 TIMEBOOST_cell_32746 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__Q), .o(TIMEBOOST_net_10284) );
na02s01 TIMEBOOST_cell_44938 ( .a(TIMEBOOST_net_14707), .b(g58074_db), .o(n_9086) );
na02s01 TIMEBOOST_cell_15885 ( .a(TIMEBOOST_net_3199), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_401), .o(TIMEBOOST_net_82) );
in01m02 g58467_u0 ( .a(FE_OFN1436_n_9372), .o(g58467_sb) );
na02f02 TIMEBOOST_cell_32745 ( .a(FE_OCP_RBN1979_n_10273), .b(TIMEBOOST_net_10283), .o(TIMEBOOST_net_6498) );
na02s02 TIMEBOOST_cell_45211 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__Q), .b(n_4361), .o(TIMEBOOST_net_14844) );
na02s01 TIMEBOOST_cell_45185 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__Q), .b(n_4908), .o(TIMEBOOST_net_14831) );
in01m02 g58468_u0 ( .a(FE_OFN1441_n_9372), .o(g58468_sb) );
na02m02 TIMEBOOST_cell_32744 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__Q), .o(TIMEBOOST_net_10283) );
na02s02 TIMEBOOST_cell_3657 ( .a(TIMEBOOST_net_408), .b(FE_OFN268_n_9880), .o(n_9537) );
na02s02 TIMEBOOST_cell_45144 ( .a(TIMEBOOST_net_14810), .b(g63063_sb), .o(n_5124) );
in01m02 g58469_u0 ( .a(FE_OFN1439_n_9372), .o(g58469_sb) );
na03s03 TIMEBOOST_cell_45407 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__Q), .b(n_3537), .c(FE_OFN1320_n_6436), .o(TIMEBOOST_net_14942) );
na02s02 TIMEBOOST_cell_3659 ( .a(TIMEBOOST_net_409), .b(FE_OFN258_n_9862), .o(n_9503) );
na02s02 TIMEBOOST_cell_31457 ( .a(TIMEBOOST_net_9639), .b(g64867_db), .o(n_3713) );
in01m02 g58470_u0 ( .a(FE_OFN1439_n_9372), .o(g58470_sb) );
na02f02 TIMEBOOST_cell_41018 ( .a(TIMEBOOST_net_12747), .b(g57104_sb), .o(n_11641) );
na02s01 TIMEBOOST_cell_16040 ( .a(FE_OFN2094_n_2520), .b(g66426_db), .o(TIMEBOOST_net_3277) );
na02s02 TIMEBOOST_cell_31456 ( .a(n_3752), .b(g64867_sb), .o(TIMEBOOST_net_9639) );
in01m02 g58471_u0 ( .a(FE_OFN1440_n_9372), .o(g58471_sb) );
na02s03 TIMEBOOST_cell_45408 ( .a(TIMEBOOST_net_14942), .b(g62998_sb), .o(n_5886) );
na02s01 TIMEBOOST_cell_16038 ( .a(FE_OFN2094_n_2520), .b(g66417_db), .o(TIMEBOOST_net_3276) );
na02s01 TIMEBOOST_cell_36521 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__Q), .b(FE_OFN535_n_9823), .o(TIMEBOOST_net_10499) );
in01m02 g58472_u0 ( .a(FE_OFN1440_n_9372), .o(g58472_sb) );
na02f02 TIMEBOOST_cell_41020 ( .a(TIMEBOOST_net_12748), .b(g57509_sb), .o(n_11230) );
na02s01 TIMEBOOST_cell_42722 ( .a(TIMEBOOST_net_13599), .b(FE_OFN1802_n_9690), .o(TIMEBOOST_net_11023) );
na02s01 TIMEBOOST_cell_36520 ( .a(TIMEBOOST_net_10498), .b(g57964_sb), .o(TIMEBOOST_net_9755) );
in01m02 g58473_u0 ( .a(FE_OFN1441_n_9372), .o(g58473_sb) );
na02f02 TIMEBOOST_cell_32739 ( .a(n_12099), .b(TIMEBOOST_net_10280), .o(TIMEBOOST_net_6518) );
na02m02 TIMEBOOST_cell_43701 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__Q), .b(n_9741), .o(TIMEBOOST_net_14089) );
na02f02 TIMEBOOST_cell_36950 ( .a(TIMEBOOST_net_10713), .b(g58817_sb), .o(n_8624) );
in01m02 g58474_u0 ( .a(FE_OFN1439_n_9372), .o(g58474_sb) );
na02m02 TIMEBOOST_cell_32738 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__Q), .o(TIMEBOOST_net_10280) );
na02s01 TIMEBOOST_cell_44939 ( .a(FE_OFN241_n_9830), .b(g57938_sb), .o(TIMEBOOST_net_14708) );
na02s01 TIMEBOOST_cell_31452 ( .a(FE_OFN217_n_9889), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__Q), .o(TIMEBOOST_net_9637) );
in01m02 g58475_u0 ( .a(FE_OFN1436_n_9372), .o(g58475_sb) );
na02f02 TIMEBOOST_cell_41324 ( .a(TIMEBOOST_net_12900), .b(g57036_sb), .o(n_11696) );
na02m02 FE_RC_884_0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_965), .o(FE_RN_580_0) );
na02s02 TIMEBOOST_cell_31451 ( .a(TIMEBOOST_net_9636), .b(g64869_db), .o(n_4425) );
in01m02 g58476_u0 ( .a(FE_OFN1438_n_9372), .o(g58476_sb) );
na02m02 TIMEBOOST_cell_32736 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__Q), .o(TIMEBOOST_net_10279) );
na02s01 TIMEBOOST_cell_9316 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(g63548_sb), .o(TIMEBOOST_net_1225) );
na02s01 TIMEBOOST_cell_39778 ( .a(TIMEBOOST_net_12127), .b(g62668_sb), .o(n_6201) );
in01m02 g58477_u0 ( .a(FE_OFN1440_n_9372), .o(g58477_sb) );
na02f02 TIMEBOOST_cell_41326 ( .a(TIMEBOOST_net_12901), .b(g57504_sb), .o(n_11234) );
na02s02 TIMEBOOST_cell_43360 ( .a(TIMEBOOST_net_13918), .b(FE_OFN2212_n_8407), .o(TIMEBOOST_net_11243) );
na02f02 TIMEBOOST_cell_38972 ( .a(TIMEBOOST_net_11724), .b(FE_OFN2155_n_16439), .o(TIMEBOOST_net_10718) );
in01m02 g58478_u0 ( .a(FE_OFN1438_n_9372), .o(g58478_sb) );
na02s01 TIMEBOOST_cell_41919 ( .a(FE_OFN203_n_9228), .b(g57898_sb), .o(TIMEBOOST_net_13198) );
na02s01 TIMEBOOST_cell_9459 ( .a(TIMEBOOST_net_1296), .b(g66403_sb), .o(n_2534) );
in01m02 g58479_u0 ( .a(FE_OFN1436_n_9372), .o(g58479_sb) );
na02f02 TIMEBOOST_cell_41328 ( .a(TIMEBOOST_net_12902), .b(g57511_sb), .o(n_10321) );
na02s02 TIMEBOOST_cell_38208 ( .a(TIMEBOOST_net_11342), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_4662) );
na02s01 TIMEBOOST_cell_9467 ( .a(TIMEBOOST_net_1300), .b(g66403_sb), .o(n_2528) );
in01m02 g58480_u0 ( .a(FE_OFN1440_n_9372), .o(g58480_sb) );
na02m02 TIMEBOOST_cell_32732 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__Q), .o(TIMEBOOST_net_10277) );
na02s01 TIMEBOOST_cell_43361 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__Q), .b(n_3663), .o(TIMEBOOST_net_13919) );
in01m02 g58481_u0 ( .a(FE_OFN1438_n_9372), .o(g58481_sb) );
na02f02 TIMEBOOST_cell_32731 ( .a(FE_OFN2209_n_11027), .b(TIMEBOOST_net_10276), .o(TIMEBOOST_net_6474) );
na02s02 TIMEBOOST_cell_43362 ( .a(TIMEBOOST_net_13919), .b(n_6554), .o(TIMEBOOST_net_12183) );
na02s01 TIMEBOOST_cell_39328 ( .a(TIMEBOOST_net_11902), .b(g58332_db), .o(n_9022) );
in01m02 g58482_u0 ( .a(FE_OFN1439_n_9372), .o(g58482_sb) );
na02m02 TIMEBOOST_cell_32730 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__Q), .o(TIMEBOOST_net_10276) );
na02s02 TIMEBOOST_cell_43363 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__Q), .b(n_3527), .o(TIMEBOOST_net_13920) );
na02s02 TIMEBOOST_cell_16362 ( .a(n_3755), .b(g64915_sb), .o(TIMEBOOST_net_3438) );
in01m02 g58483_u0 ( .a(FE_OFN1440_n_9372), .o(g58483_sb) );
na02f02 TIMEBOOST_cell_41330 ( .a(TIMEBOOST_net_12903), .b(g57318_sb), .o(n_11433) );
na02m02 TIMEBOOST_cell_44377 ( .a(n_9104), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__Q), .o(TIMEBOOST_net_14427) );
na02s02 TIMEBOOST_cell_31450 ( .a(n_4444), .b(g64869_sb), .o(TIMEBOOST_net_9636) );
in01m02 g58484_u0 ( .a(FE_OFN1440_n_9372), .o(g58484_sb) );
na02m02 TIMEBOOST_cell_32728 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__Q), .o(TIMEBOOST_net_10275) );
na02f02 TIMEBOOST_cell_43758 ( .a(TIMEBOOST_net_14117), .b(FE_OFN1400_n_8567), .o(TIMEBOOST_net_12784) );
na02s01 TIMEBOOST_cell_16363 ( .a(TIMEBOOST_net_3438), .b(g64915_db), .o(n_3688) );
in01m02 g58485_u0 ( .a(FE_OFN1437_n_9372), .o(g58485_sb) );
na02f02 TIMEBOOST_cell_32727 ( .a(FE_OFN2210_n_11027), .b(TIMEBOOST_net_10274), .o(TIMEBOOST_net_6477) );
na02m02 TIMEBOOST_cell_36941 ( .a(g52485_da), .b(FE_OFN1025_n_11877), .o(TIMEBOOST_net_10709) );
in01m02 g58486_u0 ( .a(FE_OFN1440_n_9372), .o(g58486_sb) );
na02m02 TIMEBOOST_cell_32726 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__Q), .o(TIMEBOOST_net_10274) );
na02s01 g66424_u2 ( .a(parchk_pci_ad_reg_in_1228), .b(FE_OFN795_n_2520), .o(g66424_db) );
in01s01 g58487_u0 ( .a(FE_OFN1668_n_9477), .o(g58487_sb) );
na02f02 TIMEBOOST_cell_37066 ( .a(FE_OFN1588_n_13736), .b(TIMEBOOST_net_10771), .o(n_16229) );
na02s02 TIMEBOOST_cell_36898 ( .a(TIMEBOOST_net_10687), .b(g54364_sb), .o(TIMEBOOST_net_5591) );
in01s01 g58488_u0 ( .a(FE_OFN1651_n_9428), .o(g58488_sb) );
na02s01 TIMEBOOST_cell_31248 ( .a(n_4498), .b(g64757_sb), .o(TIMEBOOST_net_9535) );
na02f02 TIMEBOOST_cell_36900 ( .a(TIMEBOOST_net_10688), .b(FE_RN_571_0), .o(FE_RN_573_0) );
na02f02 TIMEBOOST_cell_36902 ( .a(TIMEBOOST_net_10689), .b(n_14399), .o(n_14628) );
in01f01 g58489_u0 ( .a(n_9144), .o(g58489_sb) );
na02f02 TIMEBOOST_cell_36940 ( .a(TIMEBOOST_net_10708), .b(g52612_sb), .o(n_10180) );
na02s01 TIMEBOOST_cell_44940 ( .a(TIMEBOOST_net_14708), .b(g57938_db), .o(n_9872) );
na02s01 TIMEBOOST_cell_31447 ( .a(TIMEBOOST_net_9634), .b(g65355_db), .o(n_4317) );
no02f01 g58490_u0 ( .a(n_397), .b(n_9144), .o(g58490_p) );
ao12f01 g58490_u1 ( .a(g58490_p), .b(n_397), .c(n_9144), .o(n_8917) );
no02s01 g58554_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN601_n_9687), .o(n_8971) );
no02s01 g58555_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN562_n_9895), .o(n_8970) );
no02s01 g58556_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN554_n_9864), .o(n_8968) );
no02s01 g58557_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN519_n_9697), .o(n_8967) );
no02s01 g58558_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN587_n_9692), .o(n_8966) );
no02s01 g58559_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN532_n_9823), .o(n_8965) );
no02s01 g58560_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN595_n_9694), .o(n_8964) );
no02s01 g58561_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN529_n_9899), .o(n_8963) );
no02s01 g58562_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN606_n_9904), .o(n_8962) );
no02s02 g58563_u0 ( .a(n_3024), .b(n_522), .o(n_3025) );
no02s02 g58564_u0 ( .a(n_2479), .b(FE_OFN778_n_4152), .o(n_3028) );
no02s01 g58565_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN1803_n_9690), .o(n_8961) );
no02s01 g58566_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN577_n_9902), .o(n_8960) );
na02s01 TIMEBOOST_cell_39780 ( .a(TIMEBOOST_net_12128), .b(g62890_sb), .o(n_6097) );
no02m02 g58568_u0 ( .a(n_4713), .b(FE_OFN1145_n_15261), .o(n_5754) );
na02f01 g58569_u0 ( .a(n_14967), .b(n_8493), .o(g58569_p) );
in01f01 g58569_u1 ( .a(g58569_p), .o(n_10787) );
no02m04 g58570_u0 ( .a(n_3073), .b(n_784), .o(n_3074) );
no02s02 g58571_u0 ( .a(n_2631), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8661) );
na02f02 g58572_u0 ( .a(n_1085), .b(n_9144), .o(n_9143) );
na02s01 TIMEBOOST_cell_31446 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__Q), .b(g65355_sb), .o(TIMEBOOST_net_9634) );
in01f01 g58574_u0 ( .a(FE_OFN1398_n_8567), .o(g58574_sb) );
na02f02 TIMEBOOST_cell_41132 ( .a(TIMEBOOST_net_12804), .b(g57306_sb), .o(n_11445) );
na03s02 TIMEBOOST_cell_4981 ( .a(g58115_sb), .b(g58121_db), .c(FE_OFN268_n_9880), .o(n_9671) );
na02s01 TIMEBOOST_cell_31445 ( .a(TIMEBOOST_net_9633), .b(g65294_db), .o(n_4281) );
na02s01 TIMEBOOST_cell_31444 ( .a(n_4280), .b(g65294_sb), .o(TIMEBOOST_net_9633) );
in01f02 g58576_u0 ( .a(FE_OFN1369_n_8567), .o(g58576_sb) );
na02s01 TIMEBOOST_cell_30812 ( .a(n_15390), .b(n_8678), .o(TIMEBOOST_net_9317) );
na02m02 TIMEBOOST_cell_43943 ( .a(n_9560), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__Q), .o(TIMEBOOST_net_14210) );
na02s01 TIMEBOOST_cell_31064 ( .a(n_4493), .b(g64996_sb), .o(TIMEBOOST_net_9443) );
na02f02 TIMEBOOST_cell_44519 ( .a(n_9708), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__Q), .o(TIMEBOOST_net_14498) );
na02m02 g58578_u0 ( .a(n_2351), .b(n_8572), .o(n_8574) );
na02s02 TIMEBOOST_cell_45409 ( .a(TIMEBOOST_net_5437), .b(FE_OFN1312_n_6624), .o(TIMEBOOST_net_14943) );
oa12s02 g58580_u0 ( .a(n_8680), .b(FE_OFN1437_n_9372), .c(wishbone_slave_unit_pcim_if_del_bc_in_383), .o(n_8796) );
na02f04 TIMEBOOST_cell_44710 ( .a(TIMEBOOST_net_14593), .b(n_15529), .o(n_15538) );
na02f02 TIMEBOOST_cell_12973 ( .a(TIMEBOOST_net_3053), .b(n_11916), .o(n_12633) );
in01m02 g58582_u1 ( .a(g58582_p), .o(n_8571) );
oa12f02 g58583_u0 ( .a(n_8749), .b(n_8750), .c(n_3022), .o(n_8752) );
oa12m02 g58584_u0 ( .a(n_8749), .b(n_8750), .c(n_67), .o(n_8751) );
ao12m02 g58585_u0 ( .a(n_4715), .b(conf_wb_err_addr_in_967), .c(FE_OFN1145_n_15261), .o(n_5753) );
in01f01 g58586_u0 ( .a(FE_OFN1394_n_8567), .o(g58586_sb) );
na02s01 TIMEBOOST_cell_42906 ( .a(TIMEBOOST_net_13691), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_11186) );
na02s01 TIMEBOOST_cell_45053 ( .a(n_2150), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__Q), .o(TIMEBOOST_net_14765) );
na02s01 TIMEBOOST_cell_36367 ( .a(FE_OFN945_n_2248), .b(g65849_sb), .o(TIMEBOOST_net_10422) );
in01f02 g58587_u0 ( .a(FE_OFN2185_n_8567), .o(g58587_sb) );
na02f02 TIMEBOOST_cell_32725 ( .a(FE_OFN2210_n_11027), .b(TIMEBOOST_net_10273), .o(TIMEBOOST_net_6483) );
na02f02 g55270_u0 ( .a(n_12362), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__Q), .o(n_12410) );
na02s02 TIMEBOOST_cell_43551 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__Q), .b(n_3520), .o(TIMEBOOST_net_14014) );
in01f02 g58588_u0 ( .a(FE_OFN2184_n_8567), .o(g58588_sb) );
na02m02 TIMEBOOST_cell_32724 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__Q), .o(TIMEBOOST_net_10273) );
na02s01 TIMEBOOST_cell_42912 ( .a(TIMEBOOST_net_13694), .b(g58049_db), .o(n_9740) );
na02f02 TIMEBOOST_cell_31441 ( .a(TIMEBOOST_net_9631), .b(FE_OFN1150_n_13249), .o(TIMEBOOST_net_4292) );
in01f01 g58589_u0 ( .a(FE_OFN1403_n_8567), .o(g58589_sb) );
na02m02 TIMEBOOST_cell_42548 ( .a(TIMEBOOST_net_13512), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_389), .o(TIMEBOOST_net_9655) );
na02s02 TIMEBOOST_cell_45040 ( .a(TIMEBOOST_net_14758), .b(FE_OFN719_n_8060), .o(TIMEBOOST_net_11255) );
na02f02 TIMEBOOST_cell_36904 ( .a(TIMEBOOST_net_10690), .b(n_3428), .o(n_4799) );
in01f01 g58590_u0 ( .a(FE_OFN1403_n_8567), .o(g58590_sb) );
na02m02 TIMEBOOST_cell_42169 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__Q), .b(n_9552), .o(TIMEBOOST_net_13323) );
na02s01 TIMEBOOST_cell_42687 ( .a(FE_OFN225_n_9122), .b(g57928_sb), .o(TIMEBOOST_net_13582) );
na02f04 TIMEBOOST_cell_36906 ( .a(TIMEBOOST_net_10691), .b(g58587_sb), .o(n_8916) );
in01f01 g58591_u0 ( .a(FE_OFN1403_n_8567), .o(g58591_sb) );
na02s02 TIMEBOOST_cell_42052 ( .a(TIMEBOOST_net_13264), .b(g62399_sb), .o(n_6801) );
na02m02 TIMEBOOST_cell_31436 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_405), .b(TIMEBOOST_net_1563), .o(TIMEBOOST_net_9629) );
na02s02 TIMEBOOST_cell_31435 ( .a(TIMEBOOST_net_9628), .b(g65297_db), .o(n_4279) );
in01f01 g58592_u0 ( .a(FE_OFN1394_n_8567), .o(g58592_sb) );
na02s01 TIMEBOOST_cell_36390 ( .a(TIMEBOOST_net_10433), .b(g65923_db), .o(n_1565) );
na02s01 TIMEBOOST_cell_45054 ( .a(TIMEBOOST_net_14765), .b(FE_OFN719_n_8060), .o(TIMEBOOST_net_11246) );
na03f02 TIMEBOOST_cell_22366 ( .a(n_10235), .b(n_9331), .c(n_9332), .o(TIMEBOOST_net_6440) );
in01f01 g58593_u0 ( .a(FE_OFN1403_n_8567), .o(g58593_sb) );
na03s02 TIMEBOOST_cell_33472 ( .a(FE_OFN229_n_9120), .b(g57994_sb), .c(g57994_db), .o(n_9108) );
na02s02 TIMEBOOST_cell_31434 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__Q), .b(g65297_sb), .o(TIMEBOOST_net_9628) );
na02s01 TIMEBOOST_cell_42936 ( .a(TIMEBOOST_net_13706), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_11195) );
in01f01 g58594_u0 ( .a(FE_OFN1394_n_8567), .o(g58594_sb) );
na02s01 TIMEBOOST_cell_43038 ( .a(TIMEBOOST_net_13757), .b(n_4637), .o(n_4639) );
na02s02 TIMEBOOST_cell_39782 ( .a(TIMEBOOST_net_12129), .b(g62950_sb), .o(n_5981) );
na02s01 TIMEBOOST_cell_41922 ( .a(TIMEBOOST_net_13199), .b(g58412_db), .o(n_9205) );
in01f02 g58595_u0 ( .a(FE_OFN2184_n_8567), .o(g58595_sb) );
na02f02 TIMEBOOST_cell_41332 ( .a(TIMEBOOST_net_12904), .b(g57383_sb), .o(n_11362) );
na02s01 TIMEBOOST_cell_41914 ( .a(TIMEBOOST_net_13195), .b(g58302_db), .o(n_9028) );
na02s01 TIMEBOOST_cell_41923 ( .a(FE_OFN203_n_9228), .b(g58413_sb), .o(TIMEBOOST_net_13200) );
in01f02 g58596_u0 ( .a(FE_OFN2185_n_8567), .o(g58596_sb) );
na02m02 TIMEBOOST_cell_32722 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__Q), .o(TIMEBOOST_net_10272) );
na02s02 TIMEBOOST_cell_43234 ( .a(TIMEBOOST_net_13855), .b(FE_OFN1253_n_4143), .o(TIMEBOOST_net_12118) );
na02f02 TIMEBOOST_cell_43702 ( .a(TIMEBOOST_net_14089), .b(FE_OFN1349_n_8567), .o(TIMEBOOST_net_13311) );
in01f01 g58597_u0 ( .a(FE_OFN1398_n_8567), .o(g58597_sb) );
na03s02 TIMEBOOST_cell_36841 ( .a(g64984_da), .b(g64984_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__Q), .o(TIMEBOOST_net_10659) );
na02s02 TIMEBOOST_cell_36840 ( .a(TIMEBOOST_net_10658), .b(FE_OFN1226_n_6391), .o(TIMEBOOST_net_5299) );
in01s01 g58598_u0 ( .a(n_8747), .o(g58598_sb) );
na02s02 g58598_u1 ( .a(n_1423), .b(g58598_sb), .o(g58598_da) );
na02s01 g58598_u2 ( .a(n_11), .b(n_8747), .o(g58598_db) );
na02f02 TIMEBOOST_cell_4115 ( .a(TIMEBOOST_net_637), .b(n_3403), .o(n_4807) );
no02f02 g58599_u0 ( .a(n_440), .b(n_14971), .o(g58599_p) );
ao12f02 g58599_u1 ( .a(g58599_p), .b(n_440), .c(n_14971), .o(n_8842) );
in01f01 g58600_u0 ( .a(n_14971), .o(g58600_sb) );
na02m02 TIMEBOOST_cell_44167 ( .a(n_9127), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__Q), .o(TIMEBOOST_net_14322) );
na02f01 g58600_u2 ( .a(n_1421), .b(n_14971), .o(g58600_db) );
na02s02 TIMEBOOST_cell_43618 ( .a(TIMEBOOST_net_14047), .b(FE_OFN1323_n_6436), .o(TIMEBOOST_net_12243) );
in01f01 g58601_u0 ( .a(n_14971), .o(g58601_sb) );
na02f02 TIMEBOOST_cell_43944 ( .a(TIMEBOOST_net_14210), .b(FE_OFN1422_n_8567), .o(TIMEBOOST_net_12965) );
na02m02 TIMEBOOST_cell_43945 ( .a(n_9437), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__Q), .o(TIMEBOOST_net_14211) );
na03f02 TIMEBOOST_cell_3888 ( .a(n_3390), .b(n_3052), .c(n_3259), .o(TIMEBOOST_net_524) );
na02f02 TIMEBOOST_cell_44314 ( .a(TIMEBOOST_net_14395), .b(FE_OFN1425_n_8567), .o(TIMEBOOST_net_12689) );
oa12f02 g58603_u0 ( .a(n_8954), .b(FE_OFN1398_n_8567), .c(n_8953), .o(n_9340) );
oa12m01 g58604_u0 ( .a(n_8682), .b(n_8747), .c(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(n_8794) );
in01s02 g58605_u0 ( .a(FE_OFN1144_n_15261), .o(g58605_sb) );
na02f02 TIMEBOOST_cell_44520 ( .a(TIMEBOOST_net_14498), .b(FE_OFN2177_n_8567), .o(TIMEBOOST_net_13020) );
na03s02 TIMEBOOST_cell_38151 ( .a(TIMEBOOST_net_3551), .b(g64361_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__Q), .o(TIMEBOOST_net_11314) );
na02s01 TIMEBOOST_cell_38210 ( .a(TIMEBOOST_net_11343), .b(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_4509) );
in01f02 g58606_u0 ( .a(FE_OFN2182_n_8567), .o(g58606_sb) );
na02f02 TIMEBOOST_cell_32721 ( .a(FE_OFN2210_n_11027), .b(TIMEBOOST_net_10271), .o(TIMEBOOST_net_6481) );
na02s02 TIMEBOOST_cell_22307 ( .a(TIMEBOOST_net_6410), .b(n_10263), .o(n_11870) );
na02s04 TIMEBOOST_cell_45813 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_26__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_791), .o(TIMEBOOST_net_15145) );
in01f01 g58607_u0 ( .a(FE_OFN1394_n_8567), .o(g58607_sb) );
na02s02 TIMEBOOST_cell_43144 ( .a(TIMEBOOST_net_13810), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_12069) );
na02s01 TIMEBOOST_cell_44792 ( .a(TIMEBOOST_net_14634), .b(g58163_sb), .o(TIMEBOOST_net_12446) );
na02f02 TIMEBOOST_cell_22367 ( .a(TIMEBOOST_net_6440), .b(n_11008), .o(n_12165) );
in01f01 g58608_u0 ( .a(FE_OFN1403_n_8567), .o(g58608_sb) );
na02s02 TIMEBOOST_cell_42054 ( .a(TIMEBOOST_net_13265), .b(g62928_sb), .o(n_6025) );
na02s01 TIMEBOOST_cell_36842 ( .a(TIMEBOOST_net_10659), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_5118) );
na02s02 TIMEBOOST_cell_43147 ( .a(n_4220), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__Q), .o(TIMEBOOST_net_13812) );
in01f02 g58609_u0 ( .a(FE_OFN2185_n_8567), .o(g58609_sb) );
na02m02 TIMEBOOST_cell_32720 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__Q), .o(TIMEBOOST_net_10271) );
na02f02 TIMEBOOST_cell_44726 ( .a(TIMEBOOST_net_14601), .b(n_14019), .o(n_14408) );
na02s01 TIMEBOOST_cell_44941 ( .a(FE_OFN207_n_9865), .b(g57914_sb), .o(TIMEBOOST_net_14709) );
in01f01 g58610_u0 ( .a(FE_OFN1394_n_8567), .o(g58610_sb) );
na02s01 TIMEBOOST_cell_36844 ( .a(TIMEBOOST_net_10660), .b(FE_OFN1166_n_5615), .o(n_4891) );
na03m02 TIMEBOOST_cell_34852 ( .a(n_13214), .b(TIMEBOOST_net_9985), .c(n_4192), .o(n_13509) );
na02s01 TIMEBOOST_cell_31272 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__Q), .o(TIMEBOOST_net_9547) );
in01s01 g58611_u0 ( .a(n_6986), .o(g58611_sb) );
na02s01 TIMEBOOST_cell_18665 ( .a(TIMEBOOST_net_4589), .b(g59379_sb), .o(n_7681) );
na02s02 TIMEBOOST_cell_38212 ( .a(TIMEBOOST_net_11344), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_4633) );
in01f02 g58612_u0 ( .a(n_16534), .o(n_8686) );
in01s01 g58613_u0 ( .a(n_16536), .o(n_8745) );
in01f02 g58616_u0 ( .a(FE_OFN1369_n_8567), .o(g58616_sb) );
na02s02 TIMEBOOST_cell_31271 ( .a(TIMEBOOST_net_9546), .b(FE_OFN948_n_2248), .o(TIMEBOOST_net_4021) );
na02f02 TIMEBOOST_cell_43946 ( .a(TIMEBOOST_net_14211), .b(FE_OFN1396_n_8567), .o(TIMEBOOST_net_12979) );
na02s01 TIMEBOOST_cell_31270 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__Q), .o(TIMEBOOST_net_9546) );
in01f02 g58617_u0 ( .a(FE_OFN1369_n_8567), .o(g58617_sb) );
na02f04 TIMEBOOST_cell_36908 ( .a(TIMEBOOST_net_10692), .b(g58596_sb), .o(n_9191) );
na02m02 TIMEBOOST_cell_43947 ( .a(n_9665), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__Q), .o(TIMEBOOST_net_14212) );
na02f02 TIMEBOOST_cell_22369 ( .a(TIMEBOOST_net_6441), .b(n_15611), .o(n_14104) );
in01s02 g58618_u0 ( .a(FE_OFN1369_n_8567), .o(g58618_sb) );
na02s02 TIMEBOOST_cell_31269 ( .a(TIMEBOOST_net_9545), .b(FE_OFN948_n_2248), .o(TIMEBOOST_net_4020) );
na02f02 TIMEBOOST_cell_43948 ( .a(TIMEBOOST_net_14212), .b(FE_OFN1392_n_8567), .o(TIMEBOOST_net_12878) );
na02s01 TIMEBOOST_cell_31268 ( .a(pci_target_unit_fifos_pcir_data_in_167), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__Q), .o(TIMEBOOST_net_9545) );
in01f02 g58619_u0 ( .a(FE_OFN1369_n_8567), .o(g58619_sb) );
na02s02 TIMEBOOST_cell_31267 ( .a(TIMEBOOST_net_9544), .b(FE_OFN948_n_2248), .o(TIMEBOOST_net_4019) );
na02s01 TIMEBOOST_cell_43304 ( .a(TIMEBOOST_net_13890), .b(g62974_sb), .o(n_5934) );
na02f02 TIMEBOOST_cell_44150 ( .a(TIMEBOOST_net_14313), .b(FE_OFN1381_n_8567), .o(TIMEBOOST_net_13388) );
in01f02 g58620_u0 ( .a(FE_OFN1398_n_8567), .o(g58620_sb) );
na03s01 TIMEBOOST_cell_5101 ( .a(g58056_sb), .b(g58056_db), .c(FE_OFN270_n_9836), .o(n_9733) );
na02s01 TIMEBOOST_cell_42676 ( .a(TIMEBOOST_net_13576), .b(g64914_db), .o(n_4397) );
na02s02 TIMEBOOST_cell_45655 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q), .b(n_4003), .o(TIMEBOOST_net_15066) );
in01f02 g58621_u0 ( .a(FE_OFN1398_n_8567), .o(g58621_sb) );
na02s01 TIMEBOOST_cell_44823 ( .a(TIMEBOOST_net_9322), .b(FE_OFN953_n_2055), .o(TIMEBOOST_net_14650) );
na02s01 TIMEBOOST_cell_30937 ( .a(TIMEBOOST_net_9379), .b(g64986_db), .o(n_3647) );
na02f02 TIMEBOOST_cell_44711 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__Q), .b(FE_OFN1746_n_12004), .o(TIMEBOOST_net_14594) );
in01m01 g58622_u0 ( .a(n_8747), .o(g58622_sb) );
na02s02 g58622_u1 ( .a(n_1079), .b(g58622_sb), .o(g58622_da) );
na02s01 g58622_u2 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_), .b(n_8747), .o(g58622_db) );
na02s01 TIMEBOOST_cell_17418 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__Q), .b(g64228_sb), .o(TIMEBOOST_net_3966) );
in01f02 g58624_u0 ( .a(n_15517), .o(n_8792) );
in01f04 g58628_u0 ( .a(n_15515), .o(n_8790) );
in01m01 g58630_u0 ( .a(n_8747), .o(g58630_sb) );
na03f06 TIMEBOOST_cell_37153 ( .a(n_12805), .b(n_12939), .c(n_12940), .o(TIMEBOOST_net_10815) );
na02m01 g58630_u2 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_), .b(n_8747), .o(g58630_db) );
na02s01 TIMEBOOST_cell_16808 ( .a(n_3770), .b(g64990_sb), .o(TIMEBOOST_net_3661) );
in01m01 g58631_u0 ( .a(n_8747), .o(g58631_sb) );
na02f02 TIMEBOOST_cell_4005 ( .a(TIMEBOOST_net_582), .b(n_13921), .o(n_14399) );
na02m01 g58631_u2 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_), .b(n_8747), .o(g58631_db) );
na02m02 TIMEBOOST_cell_41617 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_11__Q), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_13047) );
in01m01 g58632_u0 ( .a(n_8747), .o(g58632_sb) );
na02f02 TIMEBOOST_cell_4007 ( .a(TIMEBOOST_net_583), .b(n_13679), .o(n_13747) );
na02m01 g58632_u2 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_), .b(n_8747), .o(g58632_db) );
na02s01 TIMEBOOST_cell_17115 ( .a(TIMEBOOST_net_3814), .b(g52459_sb), .o(TIMEBOOST_net_3028) );
in01s01 g58633_u0 ( .a(n_8747), .o(g58633_sb) );
na02m02 TIMEBOOST_cell_19135 ( .a(TIMEBOOST_net_4824), .b(g63577_sb), .o(n_3426) );
na02s01 g58633_u2 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_0__Q), .b(n_8747), .o(g58633_db) );
na02s01 TIMEBOOST_cell_37728 ( .a(TIMEBOOST_net_11102), .b(g61759_sb), .o(n_8295) );
in01s01 g58634_u0 ( .a(n_8747), .o(g58634_sb) );
na03s02 TIMEBOOST_cell_43305 ( .a(n_4241), .b(FE_OFN1284_n_4097), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__Q), .o(TIMEBOOST_net_13891) );
na02s01 g58634_u2 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_2__Q), .b(n_8747), .o(g58634_db) );
na02s02 TIMEBOOST_cell_37868 ( .a(TIMEBOOST_net_11172), .b(g58088_sb), .o(n_9708) );
in01s01 g58635_u0 ( .a(n_8747), .o(g58635_sb) );
na02s01 TIMEBOOST_cell_44824 ( .a(TIMEBOOST_net_14650), .b(g65726_sb), .o(TIMEBOOST_net_269) );
na02s01 g58635_u2 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_1__Q), .b(n_8747), .o(g58635_db) );
na02s01 TIMEBOOST_cell_37884 ( .a(TIMEBOOST_net_11180), .b(g58237_sb), .o(n_9554) );
in01m01 g58636_u0 ( .a(FE_OFN1700_n_5751), .o(g58636_sb) );
na02m02 TIMEBOOST_cell_44651 ( .a(n_9748), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__10__Q), .o(TIMEBOOST_net_14564) );
na03f04 TIMEBOOST_cell_42549 ( .a(n_15598), .b(n_360), .c(FE_RN_633_0), .o(TIMEBOOST_net_13513) );
na02f02 TIMEBOOST_cell_40896 ( .a(TIMEBOOST_net_12686), .b(g57329_sb), .o(n_11420) );
ao12s02 g58637_u0 ( .a(n_8732), .b(n_3158), .c(n_1077), .o(n_8734) );
ao12s02 g58638_u0 ( .a(n_8732), .b(n_3156), .c(n_1260), .o(n_8733) );
ao12s02 g58639_u0 ( .a(n_8732), .b(n_2988), .c(n_1261), .o(n_8731) );
in01f01 g58640_u0 ( .a(n_14971), .o(g58640_sb) );
na02m02 TIMEBOOST_cell_43949 ( .a(n_9633), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__Q), .o(TIMEBOOST_net_14213) );
na02f02 TIMEBOOST_cell_43950 ( .a(TIMEBOOST_net_14213), .b(FE_OFN1414_n_8567), .o(TIMEBOOST_net_12877) );
in01f01 g58641_u0 ( .a(n_16076), .o(n_8897) );
in01f01 g58645_u0 ( .a(n_16550), .o(n_8896) );
in01f01 g58652_u0 ( .a(n_14971), .o(g58652_sb) );
na02f02 TIMEBOOST_cell_39130 ( .a(TIMEBOOST_net_11803), .b(FE_OFN1599_n_13995), .o(n_14437) );
na02s01 TIMEBOOST_cell_15823 ( .a(TIMEBOOST_net_3168), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_393), .o(TIMEBOOST_net_64) );
na02s02 TIMEBOOST_cell_39784 ( .a(TIMEBOOST_net_12130), .b(g62374_sb), .o(n_6855) );
in01f01 g58653_u0 ( .a(n_14971), .o(g58653_sb) );
na02s02 TIMEBOOST_cell_18669 ( .a(TIMEBOOST_net_4591), .b(g62727_sb), .o(n_5526) );
na02s02 TIMEBOOST_cell_45214 ( .a(TIMEBOOST_net_14845), .b(FE_OFN1285_n_4097), .o(TIMEBOOST_net_12127) );
na02s02 TIMEBOOST_cell_39786 ( .a(TIMEBOOST_net_12131), .b(g62388_sb), .o(n_6824) );
in01f01 g58654_u0 ( .a(n_14971), .o(g58654_sb) );
na02s01 TIMEBOOST_cell_18671 ( .a(TIMEBOOST_net_4592), .b(g62732_sb), .o(n_5515) );
na02s01 TIMEBOOST_cell_15881 ( .a(TIMEBOOST_net_3197), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_390), .o(TIMEBOOST_net_80) );
na02s02 TIMEBOOST_cell_39788 ( .a(TIMEBOOST_net_12132), .b(g62566_sb), .o(n_6425) );
in01f01 g58655_u0 ( .a(n_14971), .o(g58655_sb) );
na02s02 TIMEBOOST_cell_18673 ( .a(TIMEBOOST_net_4593), .b(g62747_sb), .o(n_5486) );
na02s01 TIMEBOOST_cell_15845 ( .a(TIMEBOOST_net_3179), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_391), .o(TIMEBOOST_net_81) );
na02f02 TIMEBOOST_cell_39131 ( .a(FE_OFN1605_n_13997), .b(TIMEBOOST_net_10170), .o(TIMEBOOST_net_11804) );
no02f03 g58656_u0 ( .a(n_676), .b(n_7094), .o(g58656_p) );
ao12f02 g58656_u1 ( .a(g58656_p), .b(n_676), .c(n_7094), .o(n_7724) );
no02m02 g58691_u0 ( .a(n_983), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8658) );
no02f08 g58692_u0 ( .a(n_8747), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_), .o(g58692_p) );
in01f06 g58692_u1 ( .a(g58692_p), .o(n_8657) );
no02s02 g58693_u0 ( .a(n_2965), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8656) );
na02s01 g58694_u0 ( .a(n_8566), .b(n_8728), .o(n_8730) );
no02s01 g58695_u0 ( .a(n_8566), .b(n_8728), .o(g58695_p) );
in01s02 g58695_u1 ( .a(g58695_p), .o(n_8727) );
no02s02 g58696_u0 ( .a(n_2422), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8655) );
na02f02 g58697_u0 ( .a(FE_OFN1398_n_8567), .b(n_8953), .o(n_8954) );
na02s02 TIMEBOOST_cell_43148 ( .a(TIMEBOOST_net_13812), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_12647) );
na02s02 TIMEBOOST_cell_36846 ( .a(TIMEBOOST_net_10661), .b(n_2407), .o(n_4861) );
na02f02 TIMEBOOST_cell_18237 ( .a(TIMEBOOST_net_4375), .b(FE_RN_437_0), .o(TIMEBOOST_net_652) );
na02f02 TIMEBOOST_cell_39132 ( .a(TIMEBOOST_net_11804), .b(FE_OFN1601_n_13995), .o(n_14441) );
na02f03 g58702_u0 ( .a(FE_OFN2185_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__Q), .o(n_8950) );
in01s03 g58706_u0 ( .a(FE_OFN256_n_8969), .o(n_8892) );
na02s02 g58708_u0 ( .a(n_8780), .b(n_8832), .o(n_8969) );
na02f02 g58709_u0 ( .a(FE_OFN2184_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__Q), .o(n_8949) );
na02f02 g58710_u0 ( .a(FE_OFN1402_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__Q), .o(n_8890) );
na02f02 g58711_u0 ( .a(FE_OFN1403_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__Q), .o(n_8889) );
na02f02 g58712_u0 ( .a(FE_OFN1403_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__Q), .o(n_8888) );
na02f02 g58713_u0 ( .a(FE_OFN1402_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__Q), .o(n_8947) );
na02f02 g58714_u0 ( .a(FE_OFN2184_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__Q), .o(n_8946) );
na02f02 g58715_u0 ( .a(FE_OFN1402_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__Q), .o(n_8945) );
na02f02 g58716_u0 ( .a(FE_OFN2184_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__Q), .o(n_8944) );
na03s02 TIMEBOOST_cell_38397 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__Q), .b(FE_OFN1133_g64577_p), .c(n_3918), .o(TIMEBOOST_net_11437) );
na02f02 g58718_u0 ( .a(FE_OFN1402_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__Q), .o(n_8943) );
na02f02 g58723_u0 ( .a(FE_OFN2184_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q), .o(n_8887) );
na02m01 g58724_u0 ( .a(n_8747), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(n_8682) );
na02f02 g58725_u0 ( .a(n_16332), .b(FE_OFN2093_n_2301), .o(n_8572) );
na02f08 g58727_u0 ( .a(n_8747), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q), .o(n_8653) );
no02m02 g58728_u0 ( .a(n_3496), .b(FE_OFN1144_n_15261), .o(n_4715) );
na02s02 TIMEBOOST_cell_42997 ( .a(FE_OFN227_n_9841), .b(g57930_sb), .o(TIMEBOOST_net_13737) );
no02s01 g58730_u0 ( .a(FE_OCP_DRV_N1950_n_8660), .b(wishbone_slave_unit_del_sync_comp_cycle_count_0_), .o(n_8652) );
no02s02 g58731_u0 ( .a(n_2996), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8651) );
no02s02 g58732_u0 ( .a(n_2731), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8650) );
no02s02 g58733_u0 ( .a(n_3184), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8649) );
no02s02 g58734_u0 ( .a(n_3209), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8648) );
no02s02 g58735_u0 ( .a(n_1422), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8647) );
no02s02 g58736_u0 ( .a(n_2023), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8646) );
no02s01 g58737_u0 ( .a(n_2326), .b(FE_OCP_DRV_N2262_n_8660), .o(n_8645) );
no02s02 g58738_u0 ( .a(n_1656), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8644) );
no02s02 g58739_u0 ( .a(n_2008), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8643) );
no02s02 g58740_u0 ( .a(n_2302), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8642) );
no02f03 g58741_u0 ( .a(FE_OFN1344_n_8567), .b(n_8489), .o(n_9144) );
no02f04 g58742_u0 ( .a(n_1110), .b(FE_OFN1398_n_8567), .o(g58742_p) );
in01f02 g58742_u1 ( .a(g58742_p), .o(n_9341) );
na02f02 g58744_u0 ( .a(n_16577), .b(n_16573), .o(g58744_p) );
in01f02 g58744_u1 ( .a(g58744_p), .o(n_8866) );
no02f04 g58745_u0 ( .a(n_8784), .b(n_16573), .o(n_8860) );
ao12s01 g58748_u0 ( .a(n_8782), .b(n_8831), .c(wishbone_slave_unit_wishbone_slave_d_incoming_reg_34__Q), .o(n_9140) );
na02s02 TIMEBOOST_cell_41970 ( .a(TIMEBOOST_net_13223), .b(g62667_sb), .o(n_6204) );
na02f02 TIMEBOOST_cell_42354 ( .a(TIMEBOOST_net_13415), .b(g57222_sb), .o(n_11533) );
ao12s02 g58751_u0 ( .a(n_8732), .b(n_1264), .c(n_3159), .o(n_8726) );
ao12s02 g58752_u0 ( .a(n_8732), .b(n_1259), .c(n_3076), .o(n_8725) );
ao12s02 g58753_u0 ( .a(n_8732), .b(n_1475), .c(n_2998), .o(n_8724) );
oa12s02 g58754_u0 ( .a(n_8597), .b(FE_OFN1437_n_9372), .c(wishbone_slave_unit_pcim_if_del_bc_in_382), .o(n_8723) );
na02s02 TIMEBOOST_cell_42998 ( .a(TIMEBOOST_net_13737), .b(g57930_db), .o(n_9879) );
ao12s01 g58756_u0 ( .a(n_8732), .b(n_2223), .c(n_2958), .o(n_8721) );
ao12m02 g58757_u0 ( .a(n_5750), .b(conf_wb_err_addr_in_970), .c(FE_OFN1145_n_15261), .o(n_7341) );
ao12m02 g58758_u0 ( .a(n_3501), .b(conf_wb_err_addr_in_963), .c(FE_OFN1145_n_15261), .o(n_4714) );
no02s01 g58759_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_8_), .b(n_2179), .o(g58759_p) );
ao12s01 g58759_u1 ( .a(g58759_p), .b(pci_target_unit_del_sync_comp_cycle_count_8_), .c(n_2179), .o(n_2479) );
no02m02 g58760_u0 ( .a(n_3359), .b(conf_wb_err_addr_in_971), .o(g58760_p) );
ao12m02 g58760_u1 ( .a(g58760_p), .b(conf_wb_err_addr_in_971), .c(n_3359), .o(n_4713) );
no02s01 g58761_u0 ( .a(n_882), .b(n_2175), .o(g58761_p) );
ao12s01 g58761_u1 ( .a(g58761_p), .b(n_882), .c(n_2175), .o(n_2631) );
ao12m02 g58762_u0 ( .a(n_3502), .b(conf_wb_err_addr_in_955), .c(FE_OFN1144_n_15261), .o(n_4712) );
no02f02 g58763_u0 ( .a(wbu_addr_in_279), .b(n_3489), .o(g58763_p) );
ao12f02 g58763_u1 ( .a(g58763_p), .b(wbu_addr_in_279), .c(n_3489), .o(n_4890) );
no02m02 g58764_u0 ( .a(n_3488), .b(wbm_adr_o_30_), .o(g58764_p) );
ao12m02 g58764_u1 ( .a(g58764_p), .b(wbm_adr_o_30_), .c(n_3488), .o(n_4889) );
na02s01 TIMEBOOST_cell_42086 ( .a(TIMEBOOST_net_13281), .b(n_6232), .o(TIMEBOOST_net_11566) );
na02f02 TIMEBOOST_cell_41658 ( .a(TIMEBOOST_net_13067), .b(g55852_sb), .o(TIMEBOOST_net_11702) );
in01s01 g58767_u0 ( .a(FE_OFN2054_n_8831), .o(g58767_sb) );
na03s02 TIMEBOOST_cell_33818 ( .a(FE_OFN231_n_9839), .b(g58232_sb), .c(g58247_db), .o(n_9546) );
na02s01 g58767_u2 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_0__Q), .b(FE_OFN2054_n_8831), .o(g58767_db) );
na02s01 TIMEBOOST_cell_41816 ( .a(TIMEBOOST_net_13146), .b(g58276_db), .o(n_9034) );
in01s02 g58768_u0 ( .a(n_8884), .o(g58768_sb) );
no02s01 TIMEBOOST_cell_15886 ( .a(n_1780), .b(n_692), .o(TIMEBOOST_net_3200) );
na02f02 TIMEBOOST_cell_41687 ( .a(n_12357), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__Q), .o(TIMEBOOST_net_13082) );
in01s01 g58769_u0 ( .a(n_8884), .o(g58769_sb) );
na02f02 TIMEBOOST_cell_43951 ( .a(n_9097), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__Q), .o(TIMEBOOST_net_14214) );
na02f02 TIMEBOOST_cell_41688 ( .a(TIMEBOOST_net_10310), .b(TIMEBOOST_net_13082), .o(n_12877) );
na02s01 TIMEBOOST_cell_42073 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__Q), .b(n_3507), .o(TIMEBOOST_net_13275) );
in01s01 g58770_u0 ( .a(n_8831), .o(g58770_sb) );
na02s02 TIMEBOOST_cell_38214 ( .a(TIMEBOOST_net_11345), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_4620) );
na02s01 g58770_u2 ( .a(n_8831), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_12__Q), .o(g58770_db) );
na02s02 TIMEBOOST_cell_42746 ( .a(TIMEBOOST_net_13611), .b(g58304_db), .o(n_9507) );
in01s01 g58771_u0 ( .a(FE_OFN2055_n_8831), .o(g58771_sb) );
na02s01 TIMEBOOST_cell_45084 ( .a(TIMEBOOST_net_14780), .b(FE_OFN270_n_9836), .o(TIMEBOOST_net_11196) );
na03s01 TIMEBOOST_cell_5926 ( .a(n_1918), .b(g61749_sb), .c(g61749_db), .o(n_8319) );
in01s01 g58772_u0 ( .a(FE_OFN2054_n_8831), .o(g58772_sb) );
na02s02 TIMEBOOST_cell_43039 ( .a(n_8526), .b(wishbone_slave_unit_fifos_outGreyCount_0_), .o(TIMEBOOST_net_13758) );
na02s01 TIMEBOOST_cell_40387 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__Q), .b(g64325_sb), .o(TIMEBOOST_net_12432) );
na02f02 TIMEBOOST_cell_42236 ( .a(TIMEBOOST_net_13356), .b(FE_OFN1422_n_8567), .o(TIMEBOOST_net_12313) );
in01s01 g58773_u0 ( .a(FE_OFN2054_n_8831), .o(g58773_sb) );
na02s02 TIMEBOOST_cell_22305 ( .a(n_10199), .b(TIMEBOOST_net_6409), .o(n_11861) );
na02s02 TIMEBOOST_cell_22289 ( .a(n_10279), .b(TIMEBOOST_net_6401), .o(n_11876) );
na02f02 TIMEBOOST_cell_44246 ( .a(TIMEBOOST_net_14361), .b(FE_OFN1408_n_8567), .o(TIMEBOOST_net_12985) );
in01s01 g58774_u0 ( .a(n_8831), .o(g58774_sb) );
na02s02 TIMEBOOST_cell_15815 ( .a(TIMEBOOST_net_3164), .b(n_261), .o(TIMEBOOST_net_125) );
na02s01 g58774_u2 ( .a(n_8831), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_16__Q), .o(g58774_db) );
na02f02 TIMEBOOST_cell_44378 ( .a(TIMEBOOST_net_14427), .b(FE_OFN1413_n_8567), .o(TIMEBOOST_net_12722) );
in01s01 g58775_u0 ( .a(n_8831), .o(g58775_sb) );
na02f02 TIMEBOOST_cell_42242 ( .a(TIMEBOOST_net_13359), .b(FE_OFN1408_n_8567), .o(TIMEBOOST_net_12316) );
na02s01 g58775_u2 ( .a(n_8831), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_17__Q), .o(g58775_db) );
na02s01 TIMEBOOST_cell_39496 ( .a(TIMEBOOST_net_11986), .b(g63438_sb), .o(n_4621) );
in01s02 g58776_u0 ( .a(n_8884), .o(g58776_sb) );
no02s01 TIMEBOOST_cell_15887 ( .a(TIMEBOOST_net_3200), .b(n_2354), .o(g65573_p) );
na03s02 TIMEBOOST_cell_5961 ( .a(n_4470), .b(g64947_sb), .c(g64947_db), .o(n_4380) );
na02f02 TIMEBOOST_cell_41689 ( .a(n_12357), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__Q), .o(TIMEBOOST_net_13083) );
in01s02 g58777_u0 ( .a(n_8884), .o(g58777_sb) );
na02s01 TIMEBOOST_cell_15888 ( .a(n_8876), .b(pci_target_unit_fifos_pcir_flush_in), .o(TIMEBOOST_net_3201) );
na02f02 TIMEBOOST_cell_42146 ( .a(TIMEBOOST_net_13311), .b(g57184_sb), .o(n_11570) );
na03s02 TIMEBOOST_cell_5964 ( .a(n_4482), .b(g64951_sb), .c(g64951_db), .o(n_4379) );
in01s01 g58778_u0 ( .a(n_8884), .o(g58778_sb) );
na02f02 TIMEBOOST_cell_43952 ( .a(TIMEBOOST_net_14214), .b(FE_OFN1416_n_8567), .o(TIMEBOOST_net_12876) );
na02s02 TIMEBOOST_cell_43040 ( .a(TIMEBOOST_net_13758), .b(n_8668), .o(n_8717) );
na02s02 TIMEBOOST_cell_42074 ( .a(TIMEBOOST_net_13275), .b(n_6431), .o(TIMEBOOST_net_11575) );
in01s01 g58779_u0 ( .a(FE_OFN2054_n_8831), .o(g58779_sb) );
na02s01 g58779_u2 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_20__Q), .b(FE_OFN2054_n_8831), .o(g58779_db) );
na02f02 TIMEBOOST_cell_22598 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__Q), .b(n_12183), .o(TIMEBOOST_net_6556) );
na02f02 TIMEBOOST_cell_42170 ( .a(TIMEBOOST_net_13323), .b(FE_OFN1390_n_8567), .o(TIMEBOOST_net_12268) );
na02s01 g58780_u2 ( .a(n_8831), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_21__Q), .o(g58780_db) );
na02f02 TIMEBOOST_cell_41684 ( .a(TIMEBOOST_net_13080), .b(TIMEBOOST_net_3121), .o(n_12499) );
na02m02 TIMEBOOST_cell_44257 ( .a(n_9409), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__Q), .o(TIMEBOOST_net_14367) );
na02s01 TIMEBOOST_cell_41758 ( .a(TIMEBOOST_net_13117), .b(g64946_db), .o(n_3669) );
na02m04 TIMEBOOST_cell_41759 ( .a(configuration_pci_err_data_509), .b(pciu_am1_in), .o(TIMEBOOST_net_13118) );
in01s02 g58782_u0 ( .a(n_8884), .o(g58782_sb) );
na02s02 TIMEBOOST_cell_43413 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__Q), .b(n_4431), .o(TIMEBOOST_net_13945) );
na02s01 TIMEBOOST_cell_45219 ( .a(n_38), .b(n_4390), .o(TIMEBOOST_net_14848) );
na02s02 TIMEBOOST_cell_43545 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__Q), .b(n_3569), .o(TIMEBOOST_net_14011) );
in01s01 g58783_u0 ( .a(n_8831), .o(g58783_sb) );
na02m02 TIMEBOOST_cell_42171 ( .a(n_9073), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__Q), .o(TIMEBOOST_net_13324) );
na02s01 TIMEBOOST_cell_44942 ( .a(TIMEBOOST_net_14709), .b(g57914_db), .o(n_9896) );
na02s01 TIMEBOOST_cell_45055 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__Q), .b(n_1748), .o(TIMEBOOST_net_14766) );
na02s02 TIMEBOOST_cell_42108 ( .a(TIMEBOOST_net_13292), .b(FE_OFN1314_n_6624), .o(TIMEBOOST_net_11599) );
in01s01 g58785_u0 ( .a(FE_OFN2055_n_8831), .o(g58785_sb) );
na02f02 TIMEBOOST_cell_41166 ( .a(TIMEBOOST_net_12821), .b(g57477_sb), .o(n_11260) );
na02m02 TIMEBOOST_cell_44661 ( .a(n_9229), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__Q), .o(TIMEBOOST_net_14569) );
na02s02 TIMEBOOST_cell_45410 ( .a(TIMEBOOST_net_14943), .b(g62912_sb), .o(n_6054) );
in01s01 g58786_u0 ( .a(FE_OFN2055_n_8831), .o(g58786_sb) );
na02s02 TIMEBOOST_cell_45411 ( .a(TIMEBOOST_net_5433), .b(FE_OFN1312_n_6624), .o(TIMEBOOST_net_14944) );
na02s01 g58786_u2 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_27__Q), .b(FE_OFN2055_n_8831), .o(g58786_db) );
na02s02 TIMEBOOST_cell_42082 ( .a(TIMEBOOST_net_13279), .b(n_6645), .o(TIMEBOOST_net_11567) );
in01s01 g58787_u0 ( .a(n_8884), .o(g58787_sb) );
na02m02 TIMEBOOST_cell_43953 ( .a(n_9706), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__Q), .o(TIMEBOOST_net_14215) );
na02f02 TIMEBOOST_cell_21551 ( .a(TIMEBOOST_net_6032), .b(n_3060), .o(n_4168) );
na02s02 TIMEBOOST_cell_43017 ( .a(n_3833), .b(g63051_sb), .o(TIMEBOOST_net_13747) );
in01s01 g58788_u0 ( .a(FE_OFN2054_n_8831), .o(g58788_sb) );
na02f02 TIMEBOOST_cell_22253 ( .a(TIMEBOOST_net_6383), .b(n_10035), .o(n_11845) );
na02f02 TIMEBOOST_cell_42380 ( .a(TIMEBOOST_net_13428), .b(g57200_sb), .o(n_10834) );
na02s01 TIMEBOOST_cell_15860 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_82), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3187) );
in01s01 g58789_u0 ( .a(n_8831), .o(g58789_sb) );
na02s01 TIMEBOOST_cell_18025 ( .a(TIMEBOOST_net_4269), .b(g64094_db), .o(n_4061) );
na02m02 TIMEBOOST_cell_42381 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__Q), .b(n_9012), .o(TIMEBOOST_net_13429) );
na03s02 TIMEBOOST_cell_38257 ( .a(TIMEBOOST_net_3978), .b(g64248_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__Q), .o(TIMEBOOST_net_11367) );
in01s01 g58790_u0 ( .a(FE_OFN2055_n_8831), .o(g58790_sb) );
na02f02 g55370_u0 ( .a(FE_OFN1751_n_12086), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__Q), .o(n_12062) );
na02s01 g58790_u2 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_30__Q), .b(FE_OFN2055_n_8831), .o(g58790_db) );
na02s02 TIMEBOOST_cell_42126 ( .a(TIMEBOOST_net_13301), .b(FE_OFN1323_n_6436), .o(TIMEBOOST_net_11596) );
in01s01 g58791_u0 ( .a(FE_OFN2054_n_8831), .o(g58791_sb) );
na02f02 TIMEBOOST_cell_44718 ( .a(TIMEBOOST_net_14597), .b(n_11995), .o(n_12712) );
na02s02 g58791_u2 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_31__Q), .b(FE_OFN2054_n_8831), .o(g58791_db) );
na03s02 TIMEBOOST_cell_226 ( .a(g65213_sb), .b(pci_target_unit_del_sync_addr_in_231), .c(g65213_db), .o(n_2674) );
in01s01 g58792_u0 ( .a(n_8884), .o(g58792_sb) );
na02f02 TIMEBOOST_cell_43954 ( .a(TIMEBOOST_net_14215), .b(FE_OFN1392_n_8567), .o(TIMEBOOST_net_12729) );
na02s01 TIMEBOOST_cell_44943 ( .a(FE_OFN207_n_9865), .b(g57946_sb), .o(TIMEBOOST_net_14710) );
na02s02 TIMEBOOST_cell_39404 ( .a(TIMEBOOST_net_11940), .b(FE_OFN266_n_9884), .o(n_9643) );
in01s01 g58793_u0 ( .a(n_8831), .o(g58793_sb) );
na02s02 TIMEBOOST_cell_42100 ( .a(TIMEBOOST_net_13288), .b(g62980_sb), .o(n_5922) );
na02s01 g58793_u2 ( .a(n_8831), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_4__Q), .o(g58793_db) );
na02f02 TIMEBOOST_cell_42172 ( .a(TIMEBOOST_net_13324), .b(FE_OFN1394_n_8567), .o(TIMEBOOST_net_12273) );
in01s01 g58794_u0 ( .a(n_8831), .o(g58794_sb) );
na02s02 TIMEBOOST_cell_43534 ( .a(TIMEBOOST_net_14005), .b(FE_OFN1310_n_6624), .o(TIMEBOOST_net_12252) );
na02s01 g58794_u2 ( .a(n_8831), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_5__Q), .o(g58794_db) );
na03s02 TIMEBOOST_cell_41811 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__14__Q), .b(g64273_da), .c(g64273_db), .o(TIMEBOOST_net_13144) );
in01s01 g58795_u0 ( .a(FE_OFN2055_n_8831), .o(g58795_sb) );
na02s01 g58795_u2 ( .a(n_8831), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_6__Q), .o(g58795_db) );
na02s02 TIMEBOOST_cell_43364 ( .a(TIMEBOOST_net_13920), .b(n_6232), .o(TIMEBOOST_net_12176) );
na02m02 TIMEBOOST_cell_42173 ( .a(n_9728), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q), .o(TIMEBOOST_net_13325) );
na02s01 g58796_u2 ( .a(n_8831), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_7__Q), .o(g58796_db) );
na02f02 TIMEBOOST_cell_42174 ( .a(TIMEBOOST_net_13325), .b(FE_OFN1399_n_8567), .o(TIMEBOOST_net_12274) );
in01s01 g58797_u0 ( .a(FE_OFN2054_n_8831), .o(g58797_sb) );
na02s01 TIMEBOOST_cell_40493 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__Q), .b(wishbone_slave_unit_pcim_sm_data_in_642), .o(TIMEBOOST_net_12485) );
na02s01 g58797_u2 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_8__Q), .b(FE_OFN2054_n_8831), .o(g58797_db) );
na02s01 TIMEBOOST_cell_40512 ( .a(TIMEBOOST_net_12494), .b(FE_OFN1299_n_5763), .o(TIMEBOOST_net_11506) );
in01s01 g58798_u0 ( .a(FE_OFN2055_n_8831), .o(g58798_sb) );
na02m02 TIMEBOOST_cell_16106 ( .a(n_8486), .b(n_12179), .o(TIMEBOOST_net_3310) );
na02f02 TIMEBOOST_cell_42382 ( .a(TIMEBOOST_net_13429), .b(FE_OFN2182_n_8567), .o(TIMEBOOST_net_12333) );
na02m02 TIMEBOOST_cell_16107 ( .a(n_14070), .b(TIMEBOOST_net_3310), .o(TIMEBOOST_net_705) );
in01m01 g58799_u0 ( .a(FE_OFN1700_n_5751), .o(g58799_sb) );
na02s02 TIMEBOOST_cell_44825 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__Q), .b(g64359_sb), .o(TIMEBOOST_net_14651) );
na02m02 TIMEBOOST_cell_43955 ( .a(n_8992), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__Q), .o(TIMEBOOST_net_14216) );
na02f02 TIMEBOOST_cell_43956 ( .a(TIMEBOOST_net_14216), .b(FE_OFN1412_n_8567), .o(TIMEBOOST_net_12875) );
in01s01 g58800_u0 ( .a(FE_OFN1697_n_5751), .o(g58800_sb) );
na02s01 TIMEBOOST_cell_44826 ( .a(TIMEBOOST_net_14651), .b(g64359_db), .o(n_3820) );
na02f02 TIMEBOOST_cell_43957 ( .a(n_9509), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__Q), .o(TIMEBOOST_net_14217) );
in01m02 g58801_u0 ( .a(FE_OFN2153_n_16439), .o(g58801_sb) );
na02s01 TIMEBOOST_cell_40636 ( .a(TIMEBOOST_net_12556), .b(g62715_sb), .o(n_6140) );
na03s02 TIMEBOOST_cell_5457 ( .a(n_4470), .b(g64793_sb), .c(g64793_db), .o(n_4471) );
na03s02 TIMEBOOST_cell_5458 ( .a(n_4493), .b(g64795_sb), .c(g64795_db), .o(n_4469) );
in01m02 g58802_u0 ( .a(FE_OFN2153_n_16439), .o(g58802_sb) );
na02s01 TIMEBOOST_cell_44944 ( .a(TIMEBOOST_net_14710), .b(g57946_db), .o(n_9866) );
na03s02 TIMEBOOST_cell_33819 ( .a(FE_OFN254_n_9825), .b(g58229_sb), .c(g58259_db), .o(n_9538) );
na03s02 TIMEBOOST_cell_5460 ( .a(n_4465), .b(g64802_sb), .c(g64802_db), .o(n_4466) );
in01m02 g58803_u0 ( .a(FE_OFN2157_n_16439), .o(g58803_sb) );
na02s02 TIMEBOOST_cell_40638 ( .a(TIMEBOOST_net_12557), .b(g63164_sb), .o(n_5808) );
na02m02 TIMEBOOST_cell_43522 ( .a(TIMEBOOST_net_13999), .b(TIMEBOOST_net_10049), .o(n_14814) );
na02s02 TIMEBOOST_cell_43523 ( .a(n_6986), .b(n_13447), .o(TIMEBOOST_net_14000) );
in01m02 g58804_u0 ( .a(FE_OFN2157_n_16439), .o(g58804_sb) );
na03s02 TIMEBOOST_cell_33820 ( .a(FE_OFN254_n_9825), .b(g57948_sb), .c(g57976_db), .o(n_9826) );
na02f02 TIMEBOOST_cell_45842 ( .a(TIMEBOOST_net_15159), .b(n_12567), .o(n_12829) );
in01f02 g58805_u0 ( .a(FE_OFN2153_n_16439), .o(g58805_sb) );
na02s01 TIMEBOOST_cell_40640 ( .a(TIMEBOOST_net_12558), .b(g62373_sb), .o(n_6857) );
na03s02 TIMEBOOST_cell_5465 ( .a(n_4479), .b(g64820_sb), .c(g64820_db), .o(n_4456) );
na02m02 TIMEBOOST_cell_41641 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_3__Q), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_13059) );
in01m02 g58806_u0 ( .a(FE_OFN2153_n_16439), .o(g58806_sb) );
na02s02 TIMEBOOST_cell_44945 ( .a(FE_OFN254_n_9825), .b(g57945_sb), .o(TIMEBOOST_net_14711) );
na03s02 TIMEBOOST_cell_33822 ( .a(FE_OFN231_n_9839), .b(g58086_sb), .c(g58086_db), .o(n_9710) );
na03s02 TIMEBOOST_cell_33823 ( .a(FE_OFN254_n_9825), .b(g58041_sb), .c(g58067_db), .o(n_9725) );
in01m02 g58807_u0 ( .a(FE_OFN2153_n_16439), .o(g58807_sb) );
na02s01 TIMEBOOST_cell_40642 ( .a(TIMEBOOST_net_12559), .b(g62887_sb), .o(n_6103) );
na03s02 TIMEBOOST_cell_33824 ( .a(FE_OFN213_n_9124), .b(g58203_sb), .c(g58203_db), .o(n_9054) );
na03s02 TIMEBOOST_cell_33825 ( .a(FE_OFN235_n_9834), .b(g58057_sb), .c(g58057_db), .o(n_9732) );
in01m02 g58808_u0 ( .a(FE_OFN2153_n_16439), .o(g58808_sb) );
na02f02 TIMEBOOST_cell_41676 ( .a(TIMEBOOST_net_13076), .b(n_14830), .o(n_14896) );
na03s01 TIMEBOOST_cell_5472 ( .a(n_4452), .b(g64845_sb), .c(g64845_db), .o(n_4437) );
in01f01 g58809_u0 ( .a(FE_OFN2158_n_16439), .o(g58809_sb) );
na02s01 TIMEBOOST_cell_40644 ( .a(TIMEBOOST_net_12560), .b(g62587_sb), .o(n_6376) );
na03s02 TIMEBOOST_cell_33827 ( .a(FE_OFN235_n_9834), .b(g57935_sb), .c(g57935_db), .o(n_9874) );
na02s02 TIMEBOOST_cell_30901 ( .a(TIMEBOOST_net_9361), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_3740) );
in01m02 g58810_u0 ( .a(FE_OFN2153_n_16439), .o(g58810_sb) );
na02s02 TIMEBOOST_cell_44946 ( .a(TIMEBOOST_net_14711), .b(g57945_db), .o(n_9867) );
na03s01 TIMEBOOST_cell_5475 ( .a(n_4479), .b(g64853_sb), .c(g64853_db), .o(n_4432) );
na02f02 TIMEBOOST_cell_42466 ( .a(TIMEBOOST_net_13471), .b(g57461_sb), .o(n_11273) );
in01f01 g58811_u0 ( .a(FE_OFN2158_n_16439), .o(g58811_sb) );
na02s02 TIMEBOOST_cell_40646 ( .a(TIMEBOOST_net_12561), .b(g62496_sb), .o(n_6592) );
na02s02 TIMEBOOST_cell_43093 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__Q), .b(g58294_sb), .o(TIMEBOOST_net_13785) );
na02s02 TIMEBOOST_cell_45656 ( .a(TIMEBOOST_net_15066), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_11426) );
in01m02 g58812_u0 ( .a(FE_OFN2153_n_16439), .o(g58812_sb) );
na03s02 TIMEBOOST_cell_5479 ( .a(n_4447), .b(g64885_sb), .c(g64885_db), .o(n_4415) );
na02s01 TIMEBOOST_cell_45145 ( .a(FE_OFN201_n_9230), .b(g57903_sb), .o(TIMEBOOST_net_14811) );
in01m02 g58813_u0 ( .a(FE_OFN2153_n_16439), .o(g58813_sb) );
na02s01 TIMEBOOST_cell_40648 ( .a(TIMEBOOST_net_12562), .b(g62714_sb), .o(n_6142) );
na02s01 TIMEBOOST_cell_30902 ( .a(pci_target_unit_pcit_if_strd_addr_in_691), .b(n_2512), .o(TIMEBOOST_net_9362) );
na03s02 TIMEBOOST_cell_5482 ( .a(n_4672), .b(g64892_sb), .c(g64892_db), .o(n_4412) );
in01m02 g58814_u0 ( .a(FE_OFN2157_n_16439), .o(g58814_sb) );
na02m02 TIMEBOOST_cell_43524 ( .a(TIMEBOOST_net_14000), .b(n_7618), .o(TIMEBOOST_net_11586) );
na02m02 TIMEBOOST_cell_42175 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__Q), .b(n_9740), .o(TIMEBOOST_net_13326) );
in01m02 g58815_u0 ( .a(FE_OFN2153_n_16439), .o(g58815_sb) );
na02s02 TIMEBOOST_cell_40650 ( .a(TIMEBOOST_net_12563), .b(g62544_sb), .o(n_7379) );
na02s01 TIMEBOOST_cell_44947 ( .a(g65333_da), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__Q), .o(TIMEBOOST_net_14712) );
na02s01 TIMEBOOST_cell_43525 ( .a(n_2004), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__Q), .o(TIMEBOOST_net_14001) );
in01f01 g58816_u0 ( .a(FE_OFN2158_n_16439), .o(g58816_sb) );
na02s01 TIMEBOOST_cell_44948 ( .a(TIMEBOOST_net_14712), .b(TIMEBOOST_net_3880), .o(TIMEBOOST_net_4815) );
na02f02 TIMEBOOST_cell_42176 ( .a(TIMEBOOST_net_13326), .b(FE_OFN1391_n_8567), .o(TIMEBOOST_net_12269) );
na02m02 TIMEBOOST_cell_42177 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__Q), .b(n_9678), .o(TIMEBOOST_net_13327) );
in01m02 g58817_u0 ( .a(FE_OFN2156_n_16439), .o(g58817_sb) );
na02s01 TIMEBOOST_cell_40652 ( .a(TIMEBOOST_net_12564), .b(g62586_sb), .o(n_6379) );
na03s02 TIMEBOOST_cell_5489 ( .a(n_4479), .b(g64911_sb), .c(g64911_db), .o(n_4401) );
na03s01 TIMEBOOST_cell_5490 ( .a(n_4672), .b(g64912_sb), .c(g64912_db), .o(n_4400) );
in01m02 g58818_u0 ( .a(FE_OFN2157_n_16439), .o(g58818_sb) );
na02s01 TIMEBOOST_cell_43108 ( .a(TIMEBOOST_net_13792), .b(FE_OFN1196_n_4090), .o(TIMEBOOST_net_12053) );
na02f02 TIMEBOOST_cell_44705 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__Q), .b(FE_OCP_RBN1962_FE_OFN1591_n_13741), .o(TIMEBOOST_net_14591) );
in01f01 g58819_u0 ( .a(FE_OFN2158_n_16439), .o(g58819_sb) );
na02s02 TIMEBOOST_cell_40654 ( .a(TIMEBOOST_net_12565), .b(g62620_sb), .o(n_6318) );
na03s02 TIMEBOOST_cell_5493 ( .a(n_4452), .b(g64922_sb), .c(g64922_db), .o(n_4393) );
na02s01 TIMEBOOST_cell_43526 ( .a(TIMEBOOST_net_14001), .b(FE_OFN719_n_8060), .o(TIMEBOOST_net_11257) );
in01f02 g58820_u0 ( .a(FE_OFN2153_n_16439), .o(g58820_sb) );
na02s02 TIMEBOOST_cell_44949 ( .a(FE_OFN215_n_9856), .b(g57952_sb), .o(TIMEBOOST_net_14713) );
na02s02 TIMEBOOST_cell_42986 ( .a(TIMEBOOST_net_13731), .b(TIMEBOOST_net_4247), .o(TIMEBOOST_net_4513) );
na02s02 TIMEBOOST_cell_43109 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__Q), .b(n_3680), .o(TIMEBOOST_net_13793) );
in01m02 g58821_u0 ( .a(FE_OFN2153_n_16439), .o(g58821_sb) );
na02s02 TIMEBOOST_cell_40656 ( .a(TIMEBOOST_net_12566), .b(g62492_sb), .o(n_6601) );
na03s02 TIMEBOOST_cell_5497 ( .a(n_4498), .b(g64933_sb), .c(g64933_db), .o(n_4386) );
na02s02 TIMEBOOST_cell_43110 ( .a(TIMEBOOST_net_13793), .b(FE_OFN1253_n_4143), .o(TIMEBOOST_net_12089) );
in01m02 g58822_u0 ( .a(FE_OFN2153_n_16439), .o(g58822_sb) );
na03s02 TIMEBOOST_cell_5499 ( .a(n_4645), .b(g64935_sb), .c(g64935_db), .o(n_4384) );
na02f02 TIMEBOOST_cell_44280 ( .a(TIMEBOOST_net_14378), .b(FE_OFN1411_n_8567), .o(TIMEBOOST_net_12817) );
in01m02 g58823_u0 ( .a(FE_OFN2156_n_16439), .o(g58823_sb) );
na02s01 TIMEBOOST_cell_40658 ( .a(TIMEBOOST_net_12567), .b(g62517_sb), .o(n_6543) );
na02s02 TIMEBOOST_cell_43568 ( .a(TIMEBOOST_net_14022), .b(FE_OFN1311_n_6624), .o(TIMEBOOST_net_12675) );
na02m02 TIMEBOOST_cell_44281 ( .a(n_9070), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__Q), .o(TIMEBOOST_net_14379) );
in01f01 g58824_u0 ( .a(FE_OFN2158_n_16439), .o(g58824_sb) );
na02s02 TIMEBOOST_cell_44827 ( .a(n_4444), .b(g64875_sb), .o(TIMEBOOST_net_14652) );
na02f02 TIMEBOOST_cell_44282 ( .a(TIMEBOOST_net_14379), .b(FE_OFN1381_n_8567), .o(TIMEBOOST_net_12815) );
na02s02 TIMEBOOST_cell_43569 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__Q), .b(n_4321), .o(TIMEBOOST_net_14023) );
in01m02 g58825_u0 ( .a(FE_OFN2153_n_16439), .o(g58825_sb) );
na02s02 TIMEBOOST_cell_37820 ( .a(TIMEBOOST_net_11148), .b(g58107_sb), .o(n_9686) );
na02m02 TIMEBOOST_cell_44283 ( .a(n_9027), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__Q), .o(TIMEBOOST_net_14380) );
na03s02 TIMEBOOST_cell_5506 ( .a(n_4465), .b(g64982_sb), .c(g64982_db), .o(n_4363) );
in01m02 g58826_u0 ( .a(FE_OFN2155_n_16439), .o(g58826_sb) );
na02s01 TIMEBOOST_cell_37823 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__Q), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_11150) );
na02f02 TIMEBOOST_cell_44284 ( .a(TIMEBOOST_net_14380), .b(FE_OFN1413_n_8567), .o(TIMEBOOST_net_13405) );
na02s02 TIMEBOOST_cell_43570 ( .a(TIMEBOOST_net_14023), .b(FE_OFN1313_n_6624), .o(TIMEBOOST_net_12242) );
in01m02 g58827_u0 ( .a(FE_OFN2155_n_16439), .o(g58827_sb) );
na02s02 TIMEBOOST_cell_37822 ( .a(TIMEBOOST_net_11149), .b(g58390_sb), .o(n_9442) );
na03s02 TIMEBOOST_cell_5509 ( .a(n_4442), .b(g64993_sb), .c(g64993_db), .o(n_4357) );
na02m02 TIMEBOOST_cell_44285 ( .a(n_9045), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__Q), .o(TIMEBOOST_net_14381) );
in01m02 g58828_u0 ( .a(FE_OFN2155_n_16439), .o(g58828_sb) );
na03s02 TIMEBOOST_cell_37619 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__Q), .b(FE_OFN2257_n_8060), .c(n_1957), .o(TIMEBOOST_net_11048) );
na02f02 TIMEBOOST_cell_42178 ( .a(TIMEBOOST_net_13327), .b(FE_OFN1387_n_8567), .o(TIMEBOOST_net_12276) );
na03s01 TIMEBOOST_cell_33847 ( .a(n_1948), .b(g61772_sb), .c(g61772_db), .o(n_8264) );
in01m02 g58829_u0 ( .a(FE_OFN2155_n_16439), .o(g58829_sb) );
na02m02 TIMEBOOST_cell_42179 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__Q), .b(n_9783), .o(TIMEBOOST_net_13328) );
na02f02 TIMEBOOST_cell_42180 ( .a(TIMEBOOST_net_13328), .b(FE_OFN1423_n_8567), .o(TIMEBOOST_net_12278) );
in01m02 g58830_u0 ( .a(FE_OFN2157_n_16439), .o(g58830_sb) );
na02s01 TIMEBOOST_cell_40686 ( .a(TIMEBOOST_net_12581), .b(g62895_sb), .o(n_6087) );
na02m02 TIMEBOOST_cell_42181 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__Q), .b(n_9478), .o(TIMEBOOST_net_13329) );
na02s02 TIMEBOOST_cell_43527 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__Q), .b(n_4389), .o(TIMEBOOST_net_14002) );
in01m02 g58831_u0 ( .a(FE_OFN2156_n_16439), .o(g58831_sb) );
na02m04 TIMEBOOST_cell_32224 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_17__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_782), .o(TIMEBOOST_net_10023) );
na02f02 TIMEBOOST_cell_42182 ( .a(TIMEBOOST_net_13329), .b(FE_OFN1419_n_8567), .o(TIMEBOOST_net_12275) );
na02m02 TIMEBOOST_cell_42183 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q), .b(n_9089), .o(TIMEBOOST_net_13330) );
in01m02 g58832_u0 ( .a(FE_OFN2155_n_16439), .o(g58832_sb) );
na02f02 TIMEBOOST_cell_32223 ( .a(TIMEBOOST_net_10022), .b(n_13922), .o(n_14619) );
na03s01 TIMEBOOST_cell_5519 ( .a(n_4645), .b(g65019_sb), .c(g65019_db), .o(n_4341) );
na03s01 TIMEBOOST_cell_5520 ( .a(n_4672), .b(g65028_sb), .c(g65028_db), .o(n_4337) );
in01m02 g58833_u0 ( .a(FE_OFN2156_n_16439), .o(g58833_sb) );
na02s02 TIMEBOOST_cell_43497 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__Q), .b(n_3544), .o(TIMEBOOST_net_13987) );
na03s02 TIMEBOOST_cell_5521 ( .a(n_4442), .b(g65029_sb), .c(g65029_db), .o(n_4336) );
na02s02 TIMEBOOST_cell_43528 ( .a(TIMEBOOST_net_14002), .b(FE_OFN1213_n_4151), .o(TIMEBOOST_net_12114) );
in01m02 g58834_u0 ( .a(FE_OFN2156_n_16439), .o(g58834_sb) );
na02s02 TIMEBOOST_cell_32033 ( .a(TIMEBOOST_net_9927), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_4909) );
na03s02 TIMEBOOST_cell_33853 ( .a(n_1930), .b(g61781_sb), .c(g61781_db), .o(n_8244) );
na03s02 TIMEBOOST_cell_5524 ( .a(n_4645), .b(g65034_sb), .c(g65034_db), .o(n_4333) );
in01f02 g58835_u0 ( .a(FE_OFN2153_n_16439), .o(g58835_sb) );
na02s01 TIMEBOOST_cell_32032 ( .a(configuration_pci_err_data_531), .b(wbm_dat_o_30_), .o(TIMEBOOST_net_9927) );
na03s02 TIMEBOOST_cell_33854 ( .a(n_1921), .b(g61768_sb), .c(g61768_db), .o(n_8274) );
na02s01 TIMEBOOST_cell_43032 ( .a(TIMEBOOST_net_13754), .b(g57894_db), .o(n_9231) );
in01m02 g58836_u0 ( .a(FE_OFN2157_n_16439), .o(g58836_sb) );
na02s02 TIMEBOOST_cell_32031 ( .a(TIMEBOOST_net_9926), .b(FE_OFN1185_n_3476), .o(TIMEBOOST_net_4908) );
na02f02 TIMEBOOST_cell_42184 ( .a(TIMEBOOST_net_13330), .b(FE_OFN1384_n_8567), .o(TIMEBOOST_net_12270) );
na02f02 TIMEBOOST_cell_42185 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__Q), .b(n_9716), .o(TIMEBOOST_net_13331) );
in01m02 g58837_u0 ( .a(FE_OFN1437_n_9372), .o(g58837_sb) );
na02f02 TIMEBOOST_cell_41334 ( .a(TIMEBOOST_net_12905), .b(g57525_sb), .o(n_11216) );
na02s02 TIMEBOOST_cell_43306 ( .a(TIMEBOOST_net_13891), .b(g62900_sb), .o(n_6077) );
na02s02 TIMEBOOST_cell_39790 ( .a(TIMEBOOST_net_12133), .b(g62414_sb), .o(n_6770) );
in01m02 g58838_u0 ( .a(FE_OFN1438_n_9372), .o(g58838_sb) );
na02m02 TIMEBOOST_cell_32718 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__Q), .o(TIMEBOOST_net_10270) );
na02s01 TIMEBOOST_cell_43235 ( .a(n_4423), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__Q), .o(TIMEBOOST_net_13856) );
na03f02 TIMEBOOST_cell_8343 ( .a(n_9201), .b(FE_OFN1426_n_8567), .c(g57585_db), .o(n_10800) );
in01m02 g58839_u0 ( .a(FE_OFN1438_n_9372), .o(g58839_sb) );
na02f02 TIMEBOOST_cell_32717 ( .a(FE_OFN1572_n_11027), .b(TIMEBOOST_net_10269), .o(TIMEBOOST_net_6479) );
na02s01 g66420_u2 ( .a(n_2509), .b(FE_OFN795_n_2520), .o(g66420_db) );
na02s02 TIMEBOOST_cell_44950 ( .a(TIMEBOOST_net_14713), .b(g57952_db), .o(n_9857) );
in01m02 g58840_u0 ( .a(FE_OFN1438_n_9372), .o(g58840_sb) );
na02m02 TIMEBOOST_cell_32716 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__Q), .o(TIMEBOOST_net_10269) );
na02s02 TIMEBOOST_cell_43365 ( .a(n_3672), .b(n_3673), .o(TIMEBOOST_net_13921) );
na02s01 TIMEBOOST_cell_42611 ( .a(FE_OFN245_n_9114), .b(g58034_sb), .o(TIMEBOOST_net_13544) );
in01m02 g58841_u0 ( .a(FE_OFN1438_n_9372), .o(g58841_sb) );
na02f02 TIMEBOOST_cell_21823 ( .a(TIMEBOOST_net_6168), .b(n_2829), .o(n_4169) );
na02s02 TIMEBOOST_cell_43366 ( .a(TIMEBOOST_net_13921), .b(n_6645), .o(TIMEBOOST_net_12177) );
na02s02 TIMEBOOST_cell_39792 ( .a(TIMEBOOST_net_12134), .b(g62380_sb), .o(n_6842) );
in01s02 g58842_u0 ( .a(FE_OFN21_n_9372), .o(g58842_sb) );
na02s01 TIMEBOOST_cell_18649 ( .a(TIMEBOOST_net_4581), .b(g63097_sb), .o(n_5060) );
na02f02 TIMEBOOST_cell_32715 ( .a(FE_OFN2209_n_11027), .b(TIMEBOOST_net_10268), .o(TIMEBOOST_net_6473) );
na02s02 TIMEBOOST_cell_38742 ( .a(TIMEBOOST_net_11609), .b(g53907_sb), .o(n_13534) );
in01m01 g58843_u0 ( .a(FE_OFN1700_n_5751), .o(g58843_sb) );
na03s02 TIMEBOOST_cell_37883 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__Q), .b(FE_OFN542_n_9690), .c(FE_OFN258_n_9862), .o(TIMEBOOST_net_11180) );
na02f02 TIMEBOOST_cell_43808 ( .a(TIMEBOOST_net_14142), .b(FE_OFN1411_n_8567), .o(TIMEBOOST_net_12959) );
na02s01 TIMEBOOST_cell_15849 ( .a(TIMEBOOST_net_3181), .b(n_1817), .o(TIMEBOOST_net_799) );
in01s02 g58855_u0 ( .a(pci_target_unit_wishbone_master_reset_rty_cnt), .o(n_8732) );
no02s02 g58859_u0 ( .a(FE_OFN1437_n_9372), .b(wishbone_slave_unit_pcim_if_del_bc_in), .o(n_8598) );
in01m01 g58860_u0 ( .a(n_8596), .o(n_8597) );
no02f01 g58861_u0 ( .a(n_8569), .b(wishbone_slave_unit_wishbone_slave_map), .o(n_8596) );
na02m01 g58862_u0 ( .a(n_8569), .b(wishbone_slave_unit_pcim_if_del_burst_in), .o(n_8570) );
in01s02 g58863_u0 ( .a(n_8782), .o(n_8832) );
no02m04 g58865_u0 ( .a(n_8831), .b(n_1323), .o(n_8782) );
no02s01 g58866_u0 ( .a(n_8665), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_35__Q), .o(n_8780) );
no02m02 g58871_u0 ( .a(FE_OFN1144_n_15261), .b(n_3206), .o(n_3502) );
no02m02 g58872_u0 ( .a(n_3210), .b(FE_OFN1144_n_15261), .o(n_3501) );
no02m02 g58873_u0 ( .a(n_4707), .b(FE_OFN1145_n_15261), .o(n_5750) );
na02s01 TIMEBOOST_cell_41733 ( .a(FE_OFN205_n_9140), .b(g57893_sb), .o(TIMEBOOST_net_13105) );
no02m01 g58875_u0 ( .a(n_8569), .b(n_665), .o(n_8568) );
na02f02 g58_u0 ( .a(n_15527), .b(n_15539), .o(n_15540) );
na03s02 TIMEBOOST_cell_37879 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__Q), .b(FE_OFN561_n_9895), .c(FE_OFN260_n_9860), .o(TIMEBOOST_net_11178) );
no02s02 g59072_u0 ( .a(n_3211), .b(FE_OFN778_n_4152), .o(n_3497) );
na02m02 TIMEBOOST_cell_42237 ( .a(n_9621), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__Q), .o(TIMEBOOST_net_13357) );
in01f02 g59074_u0 ( .a(n_16332), .o(n_8538) );
oa12m01 g59081_u0 ( .a(n_8668), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_1_), .c(n_8590), .o(n_8669) );
in01s01 g59082_u0 ( .a(n_8590), .o(g59082_sb) );
na02s02 TIMEBOOST_cell_43546 ( .a(TIMEBOOST_net_14011), .b(FE_OFN1317_n_6624), .o(TIMEBOOST_net_12255) );
na02m02 TIMEBOOST_cell_38971 ( .a(wbu_sel_in_312), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_33__Q), .o(TIMEBOOST_net_11724) );
na02f02 TIMEBOOST_cell_44724 ( .a(TIMEBOOST_net_14600), .b(n_12338), .o(n_16597) );
ao12s01 g59083_u0 ( .a(n_7720), .b(wishbone_slave_unit_del_sync_comp_done_reg_clr), .c(wishbone_slave_unit_del_sync_comp_done_reg_main), .o(n_8496) );
ao12s01 g59084_u0 ( .a(n_2877), .b(n_7704), .c(n_709), .o(n_8495) );
na02m02 TIMEBOOST_cell_43703 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__Q), .b(n_9443), .o(TIMEBOOST_net_14090) );
no02m02 g59086_u0 ( .a(n_3008), .b(conf_wb_err_addr_in_967), .o(g59086_p) );
ao12m02 g59086_u1 ( .a(g59086_p), .b(conf_wb_err_addr_in_967), .c(n_3008), .o(n_3496) );
oa12f02 g59087_u0 ( .a(n_3492), .b(n_3491), .c(wbu_addr_in_275), .o(n_4708) );
oa12f02 g59088_u0 ( .a(n_8492), .b(n_16876), .c(n_8564), .o(n_8565) );
in01m01 g59089_u0 ( .a(n_8590), .o(g59089_sb) );
na04f02 TIMEBOOST_cell_33547 ( .a(TIMEBOOST_net_3689), .b(n_3296), .c(n_3374), .d(n_3399), .o(n_5549) );
na02f04 TIMEBOOST_cell_42550 ( .a(TIMEBOOST_net_13513), .b(FE_RN_632_0), .o(FE_RN_636_0) );
na03s01 TIMEBOOST_cell_33546 ( .a(TIMEBOOST_net_246), .b(g61764_sb), .c(g61764_db), .o(n_8283) );
in01m02 g59090_u0 ( .a(FE_OCPN1847_n_14981), .o(g59090_sb) );
na02s02 TIMEBOOST_cell_3315 ( .a(TIMEBOOST_net_237), .b(n_4465), .o(n_4320) );
na02s01 TIMEBOOST_cell_37824 ( .a(TIMEBOOST_net_11150), .b(FE_OFN1666_n_9477), .o(TIMEBOOST_net_9710) );
na02s01 TIMEBOOST_cell_15889 ( .a(TIMEBOOST_net_3201), .b(g56933_sb), .o(TIMEBOOST_net_621) );
na02s01 TIMEBOOST_cell_3317 ( .a(TIMEBOOST_net_238), .b(n_4645), .o(n_4313) );
in01s01 TIMEBOOST_cell_45900 ( .a(TIMEBOOST_net_15206), .o(TIMEBOOST_net_15207) );
na02s01 TIMEBOOST_cell_15890 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__Q), .b(pci_target_unit_fifos_pcir_flush_in), .o(TIMEBOOST_net_3202) );
in01s01 g59092_u0 ( .a(n_4662), .o(g59092_sb) );
na02m02 TIMEBOOST_cell_39353 ( .a(TIMEBOOST_net_1561), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_398), .o(TIMEBOOST_net_11915) );
na02s01 TIMEBOOST_cell_38604 ( .a(TIMEBOOST_net_11540), .b(g62913_sb), .o(n_6053) );
na02f02 TIMEBOOST_cell_44650 ( .a(TIMEBOOST_net_14563), .b(FE_OFN2184_n_8567), .o(TIMEBOOST_net_13027) );
in01s01 g59093_u0 ( .a(FE_OFN1705_n_4868), .o(g59093_sb) );
na02s02 TIMEBOOST_cell_3705 ( .a(TIMEBOOST_net_432), .b(FE_OFN264_n_9849), .o(n_9420) );
na02f02 TIMEBOOST_cell_39134 ( .a(TIMEBOOST_net_11805), .b(FE_OFN1599_n_13995), .o(n_16225) );
na02s01 TIMEBOOST_cell_31266 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__Q), .o(TIMEBOOST_net_9544) );
oa12f01 g59094_u0 ( .a(n_8664), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_), .c(FE_OCPN1847_n_14981), .o(n_8765) );
no02s01 g59095_u0 ( .a(n_425), .b(n_8590), .o(g59095_p) );
ao12s01 g59095_u1 ( .a(g59095_p), .b(n_425), .c(n_8590), .o(n_8588) );
in01s01 g59096_u0 ( .a(FE_OFN1698_n_5751), .o(g59096_sb) );
in01s01 TIMEBOOST_cell_45901 ( .a(wbm_dat_i_10_), .o(TIMEBOOST_net_15208) );
na02s01 TIMEBOOST_cell_3441 ( .a(TIMEBOOST_net_300), .b(g58136_db), .o(n_9660) );
na03s02 TIMEBOOST_cell_34261 ( .a(TIMEBOOST_net_9814), .b(FE_OFN1171_n_5592), .c(g62128_sb), .o(n_5568) );
in01s01 g59097_u0 ( .a(n_14389), .o(g59097_sb) );
na02s02 TIMEBOOST_cell_42551 ( .a(n_1252), .b(n_1340), .o(TIMEBOOST_net_13514) );
na02s01 TIMEBOOST_cell_39794 ( .a(TIMEBOOST_net_12135), .b(g62546_sb), .o(n_6475) );
in01m02 g59098_u0 ( .a(FE_OCPN1847_n_14981), .o(g59098_sb) );
na02s02 TIMEBOOST_cell_3319 ( .a(TIMEBOOST_net_239), .b(n_4482), .o(n_4299) );
na02s02 TIMEBOOST_cell_44828 ( .a(TIMEBOOST_net_14652), .b(g64875_db), .o(n_4421) );
na02s01 TIMEBOOST_cell_31247 ( .a(TIMEBOOST_net_9534), .b(g65017_db), .o(n_4342) );
in01f02 g59099_u0 ( .a(n_16577), .o(n_8784) );
in01s01 g59102_u0 ( .a(n_16537), .o(n_8712) );
in01s01 g59105_u0 ( .a(n_16573), .o(n_8711) );
in01s01 g59109_u0 ( .a(FE_OCPN1847_n_14981), .o(g59109_sb) );
na02s02 TIMEBOOST_cell_16565 ( .a(TIMEBOOST_net_3539), .b(g65672_db), .o(n_2455) );
in01s01 TIMEBOOST_cell_45902 ( .a(TIMEBOOST_net_15208), .o(TIMEBOOST_net_15209) );
na02s02 TIMEBOOST_cell_31246 ( .a(n_4444), .b(g65017_sb), .o(TIMEBOOST_net_9534) );
in01m02 g59110_u0 ( .a(FE_OCPN1847_n_14981), .o(g59110_sb) );
na02s01 TIMEBOOST_cell_31245 ( .a(TIMEBOOST_net_9533), .b(g65014_db), .o(n_4344) );
na02s01 TIMEBOOST_cell_44829 ( .a(n_4476), .b(g64902_sb), .o(TIMEBOOST_net_14653) );
na02s01 TIMEBOOST_cell_3324 ( .a(n_4718), .b(n_2087), .o(TIMEBOOST_net_242) );
in01s01 g59111_u0 ( .a(FE_OCPN1847_n_14981), .o(g59111_sb) );
na02s01 TIMEBOOST_cell_3325 ( .a(TIMEBOOST_net_242), .b(n_3314), .o(n_3402) );
na03s02 TIMEBOOST_cell_37861 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__Q), .b(FE_OFN260_n_9860), .c(FE_OFN1687_n_9528), .o(TIMEBOOST_net_11169) );
na02f02 TIMEBOOST_cell_43704 ( .a(TIMEBOOST_net_14090), .b(FE_OFN1349_n_8567), .o(TIMEBOOST_net_13312) );
in01s01 g59112_u0 ( .a(FE_OCPN1847_n_14981), .o(g59112_sb) );
na02s04 TIMEBOOST_cell_3327 ( .a(n_2180), .b(TIMEBOOST_net_243), .o(n_3024) );
in01s01 TIMEBOOST_cell_45903 ( .a(wbm_dat_i_11_), .o(TIMEBOOST_net_15210) );
na03s02 TIMEBOOST_cell_43023 ( .a(n_4058), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__Q), .c(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_13750) );
in01s01 g59113_u0 ( .a(FE_OCPN1847_n_14981), .o(g59113_sb) );
na02m04 TIMEBOOST_cell_3329 ( .a(TIMEBOOST_net_244), .b(n_2176), .o(n_3073) );
na02s01 TIMEBOOST_cell_44830 ( .a(TIMEBOOST_net_14653), .b(g64902_db), .o(n_4408) );
na02f02 TIMEBOOST_cell_21809 ( .a(TIMEBOOST_net_6161), .b(g58588_sb), .o(n_8914) );
na02s01 TIMEBOOST_cell_3331 ( .a(TIMEBOOST_net_245), .b(g65876_sb), .o(n_1868) );
na02m02 TIMEBOOST_cell_20540 ( .a(g52441_sb), .b(g52441_db), .o(TIMEBOOST_net_5527) );
na03s02 TIMEBOOST_cell_37679 ( .a(n_1572), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__Q), .c(FE_OFN706_n_8119), .o(TIMEBOOST_net_11078) );
na02s01 TIMEBOOST_cell_17186 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__Q), .b(g65354_sb), .o(TIMEBOOST_net_3850) );
na02s01 TIMEBOOST_cell_32022 ( .a(configuration_pci_err_addr_480), .b(wbm_adr_o_10_), .o(TIMEBOOST_net_9922) );
na02s01 TIMEBOOST_cell_3335 ( .a(TIMEBOOST_net_247), .b(g65876_sb), .o(n_1899) );
in01s01 TIMEBOOST_cell_45904 ( .a(TIMEBOOST_net_15210), .o(TIMEBOOST_net_15211) );
na02s01 TIMEBOOST_cell_15891 ( .a(TIMEBOOST_net_3202), .b(g57780_sb), .o(TIMEBOOST_net_895) );
na02s01 TIMEBOOST_cell_3337 ( .a(TIMEBOOST_net_248), .b(g64286_sb), .o(n_3887) );
na02s01 TIMEBOOST_cell_44831 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__Q), .b(FE_OFN639_n_4669), .o(TIMEBOOST_net_14654) );
na02s01 TIMEBOOST_cell_15892 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__Q), .b(pci_target_unit_fifos_pcir_flush_in), .o(TIMEBOOST_net_3203) );
in01m02 g59118_u0 ( .a(FE_OCPN1847_n_14981), .o(g59118_sb) );
na02s01 TIMEBOOST_cell_3339 ( .a(TIMEBOOST_net_249), .b(g64286_sb), .o(n_3870) );
na02s01 TIMEBOOST_cell_44832 ( .a(TIMEBOOST_net_14654), .b(n_4442), .o(TIMEBOOST_net_10907) );
na02s02 TIMEBOOST_cell_3340 ( .a(n_2463), .b(n_2596), .o(TIMEBOOST_net_250) );
na02s02 TIMEBOOST_cell_3341 ( .a(TIMEBOOST_net_250), .b(n_2738), .o(n_2989) );
na03s02 TIMEBOOST_cell_37801 ( .a(n_1864), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__Q), .c(FE_OFN706_n_8119), .o(TIMEBOOST_net_11139) );
na02f02 TIMEBOOST_cell_44646 ( .a(TIMEBOOST_net_14561), .b(FE_OFN2190_n_8567), .o(TIMEBOOST_net_13493) );
na02m02 TIMEBOOST_cell_3343 ( .a(TIMEBOOST_net_251), .b(n_2738), .o(n_3174) );
na02s02 TIMEBOOST_cell_44951 ( .a(FE_OFN239_n_9832), .b(g57999_sb), .o(TIMEBOOST_net_14714) );
na02m02 TIMEBOOST_cell_32714 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__Q), .o(TIMEBOOST_net_10268) );
in01s01 g59121_u0 ( .a(FE_OFN1144_n_15261), .o(g59121_sb) );
na02s02 TIMEBOOST_cell_39330 ( .a(TIMEBOOST_net_11903), .b(FE_OFN699_n_7845), .o(TIMEBOOST_net_4106) );
na02s01 TIMEBOOST_cell_9940 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__8__Q), .b(g58407_sb), .o(TIMEBOOST_net_1537) );
na02s01 TIMEBOOST_cell_18837 ( .a(TIMEBOOST_net_4675), .b(g63125_sb), .o(n_5003) );
in01s02 g59122_u0 ( .a(n_8590), .o(g59122_sb) );
na02m02 TIMEBOOST_cell_37793 ( .a(FE_OFN1145_n_15261), .b(conf_wb_err_addr_in_959), .o(TIMEBOOST_net_11135) );
na02s01 TIMEBOOST_cell_36522 ( .a(TIMEBOOST_net_10499), .b(g57985_sb), .o(TIMEBOOST_net_4317) );
na02f02 TIMEBOOST_cell_36524 ( .a(TIMEBOOST_net_10500), .b(n_2389), .o(n_3125) );
in01s02 g59123_u0 ( .a(FE_OFN1697_n_5751), .o(g59123_sb) );
na03s02 TIMEBOOST_cell_43307 ( .a(n_3518), .b(FE_OFN1272_n_4096), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q), .o(TIMEBOOST_net_13892) );
na02s01 TIMEBOOST_cell_37789 ( .a(TIMEBOOST_net_9621), .b(FE_OFN1077_n_4740), .o(TIMEBOOST_net_11133) );
na02s01 TIMEBOOST_cell_37730 ( .a(TIMEBOOST_net_11103), .b(g62001_sb), .o(n_7893) );
no02f02 g59124_u0 ( .a(wbu_addr_in_267), .b(n_3203), .o(g59124_p) );
ao12f02 g59124_u1 ( .a(g59124_p), .b(wbu_addr_in_267), .c(n_3203), .o(n_4210) );
no02m02 g59125_u0 ( .a(n_3191), .b(wbm_adr_o_26_), .o(g59125_p) );
ao12m02 g59125_u1 ( .a(g59125_p), .b(wbm_adr_o_26_), .c(n_3191), .o(n_4209) );
in01s01 g59126_u0 ( .a(wbs_rty_o), .o(g59126_sb) );
na02f02 TIMEBOOST_cell_43958 ( .a(TIMEBOOST_net_14217), .b(FE_OFN1402_n_8567), .o(TIMEBOOST_net_12874) );
na02m01 g59126_u2 ( .a(n_15313), .b(wbs_rty_o), .o(g59126_db) );
na02s01 TIMEBOOST_cell_15792 ( .a(parchk_pci_ad_reg_in_1205), .b(g67083_db), .o(TIMEBOOST_net_3153) );
no02s02 g59127_u0 ( .a(conf_wb_err_addr_in_959), .b(n_3015), .o(g59127_p) );
ao12s02 g59127_u1 ( .a(g59127_p), .b(conf_wb_err_addr_in_959), .c(n_3015), .o(n_3493) );
no02f02 g59128_u0 ( .a(n_1407), .b(n_4704), .o(g59128_p) );
ao12f02 g59128_u1 ( .a(g59128_p), .b(n_1407), .c(n_4704), .o(n_7095) );
no02f03 g59129_u0 ( .a(parchk_pci_cbe_out_in), .b(n_4703), .o(g59129_p) );
in01s10 g59133_u0 ( .a(FE_OFN2054_n_8831), .o(n_8665) );
in01s10 g59141_u0 ( .a(n_8665), .o(n_8884) );
no02f01 g59161_u0 ( .a(n_8760), .b(FE_OCP_RBN2003_FE_OFN1026_n_16760), .o(n_14689) );
in01f08 g59169_u0 ( .a(n_8569), .o(n_9372) );
na02s02 TIMEBOOST_cell_43126 ( .a(TIMEBOOST_net_13801), .b(FE_OFN1253_n_4143), .o(TIMEBOOST_net_12104) );
na02s04 g59175_u0 ( .a(n_1095), .b(n_8590), .o(n_8668) );
na02m02 g59176_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_), .b(FE_OCPN1847_n_14981), .o(n_8664) );
na02f02 g59177_u0 ( .a(n_3491), .b(wbu_addr_in_275), .o(n_3492) );
no02s01 g59180_u0 ( .a(n_3185), .b(FE_OFN778_n_4152), .o(n_3490) );
no02s02 g59181_u0 ( .a(n_2327), .b(FE_OFN778_n_4152), .o(n_2774) );
na02m01 g59182_u0 ( .a(n_1064), .b(n_8493), .o(n_8494) );
na02f02 g59183_u0 ( .a(n_8493), .b(n_7114), .o(n_8492) );
na02f02 TIMEBOOST_cell_43705 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q), .b(n_9575), .o(TIMEBOOST_net_14091) );
na02m02 TIMEBOOST_cell_3983 ( .a(n_3189), .b(TIMEBOOST_net_571), .o(n_3190) );
na02s01 TIMEBOOST_cell_43367 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__Q), .b(n_4380), .o(TIMEBOOST_net_13922) );
no02f04 g59187_u0 ( .a(n_3193), .b(n_1286), .o(n_3489) );
na02f02 TIMEBOOST_cell_42286 ( .a(TIMEBOOST_net_13381), .b(g57424_sb), .o(n_11311) );
no02m04 g59189_u0 ( .a(n_3190), .b(n_876), .o(n_3488) );
na02s02 TIMEBOOST_cell_38216 ( .a(TIMEBOOST_net_11346), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_4661) );
na02m02 TIMEBOOST_cell_37103 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__Q), .o(TIMEBOOST_net_10790) );
na02s02 TIMEBOOST_cell_19281 ( .a(TIMEBOOST_net_4897), .b(g60636_sb), .o(n_5699) );
ao12s02 g59194_u0 ( .a(wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q), .b(n_7715), .c(n_169), .o(n_7720) );
no02s02 g59196_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_15_), .b(n_2491), .o(g59196_p) );
ao12s02 g59196_u1 ( .a(g59196_p), .b(pci_target_unit_del_sync_comp_cycle_count_15_), .c(n_2491), .o(n_3211) );
oa12s02 g59197_u0 ( .a(n_3201), .b(n_3200), .c(wbu_addr_in_271), .o(n_3487) );
no02f02 g59198_u0 ( .a(n_261), .b(n_3179), .o(g59198_p) );
ao12f02 g59198_u1 ( .a(g59198_p), .b(n_261), .c(n_3179), .o(n_4208) );
no02m02 g59199_u0 ( .a(n_2492), .b(conf_wb_err_addr_in_963), .o(g59199_p) );
ao12m02 g59199_u1 ( .a(g59199_p), .b(conf_wb_err_addr_in_963), .c(n_2492), .o(n_3210) );
ao12m02 g59200_u0 ( .a(n_4207), .b(conf_wb_err_addr_in_966), .c(FE_OFN1142_n_15261), .o(n_4886) );
no02m02 g59201_u0 ( .a(n_3353), .b(conf_wb_err_addr_in_970), .o(g59201_p) );
ao12m02 g59201_u1 ( .a(g59201_p), .b(conf_wb_err_addr_in_970), .c(n_3353), .o(n_4707) );
oa12m02 g59202_u0 ( .a(n_3198), .b(n_3197), .c(wbm_adr_o_18_), .o(n_3486) );
oa12s02 g59203_u0 ( .a(n_3196), .b(n_3195), .c(wbm_adr_o_22_), .o(n_3485) );
oa12m01 g59204_u0 ( .a(n_5739), .b(FE_OFN987_n_2696), .c(n_7717), .o(n_7719) );
oa12s06 g59205_u0 ( .a(n_5737), .b(FE_OFN985_n_2697), .c(n_7717), .o(n_7718) );
no02s02 g59206_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__Q), .b(n_2490), .o(g59206_p) );
ao12s02 g59206_u1 ( .a(g59206_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__Q), .c(n_2490), .o(n_3209) );
ao12m02 g59208_u0 ( .a(n_3199), .b(conf_wb_err_addr_in_947), .c(FE_OFN1143_n_15261), .o(n_3484) );
in01s02 g59209_u0 ( .a(n_8487), .o(n_8528) );
na03s02 TIMEBOOST_cell_6267 ( .a(FE_OFN231_n_9839), .b(g58025_sb), .c(g58025_db), .o(n_9765) );
in01s02 g59211_u0 ( .a(n_2179), .o(n_2180) );
na02m02 TIMEBOOST_cell_42383 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__Q), .b(n_9537), .o(TIMEBOOST_net_13430) );
oa12f02 g59213_u0 ( .a(n_1493), .b(FE_OFN562_n_9895), .c(n_8561), .o(n_8563) );
oa12f01 g59214_u0 ( .a(n_1806), .b(FE_OFN601_n_9687), .c(n_8561), .o(n_8562) );
oa12f02 g59215_u0 ( .a(n_1800), .b(FE_OFN554_n_9864), .c(n_8561), .o(n_8560) );
oa12f02 g59216_u0 ( .a(n_1821), .b(FE_OFN519_n_9697), .c(n_8561), .o(n_8559) );
oa12f02 g59217_u0 ( .a(n_1540), .b(FE_OFN587_n_9692), .c(n_8561), .o(n_8558) );
oa12f02 g59218_u0 ( .a(n_1542), .b(FE_OFN532_n_9823), .c(n_8561), .o(n_8557) );
oa12f01 g59219_u0 ( .a(n_1814), .b(FE_OFN595_n_9694), .c(n_8561), .o(n_8556) );
oa12f02 g59220_u0 ( .a(n_1820), .b(FE_OFN529_n_9899), .c(n_8561), .o(n_8555) );
oa12f01 g59221_u0 ( .a(n_1230), .b(FE_OFN1795_n_9904), .c(n_8561), .o(n_8554) );
oa12f02 g59222_u0 ( .a(n_1822), .b(FE_OFN1800_n_9690), .c(n_8561), .o(n_8553) );
oa12f02 g59223_u0 ( .a(n_1810), .b(FE_OFN577_n_9902), .c(n_8561), .o(n_8552) );
in01m02 g59224_u0 ( .a(n_2175), .o(n_2176) );
na02f02 TIMEBOOST_cell_42384 ( .a(TIMEBOOST_net_13430), .b(FE_OFN2191_n_8567), .o(TIMEBOOST_net_12332) );
in01s01 g59226_u0 ( .a(n_6986), .o(g59226_sb) );
na02s01 TIMEBOOST_cell_45056 ( .a(TIMEBOOST_net_14766), .b(FE_OFN720_n_8060), .o(TIMEBOOST_net_11240) );
na03m02 TIMEBOOST_cell_6629 ( .a(n_3347), .b(g59234_sb), .c(TIMEBOOST_net_584), .o(g53938_da) );
na02f02 TIMEBOOST_cell_36910 ( .a(TIMEBOOST_net_10693), .b(n_2823), .o(n_4683) );
no02m02 g59227_u0 ( .a(wbu_addr_in_263), .b(n_3202), .o(g59227_p) );
ao12m02 g59227_u1 ( .a(g59227_p), .b(wbu_addr_in_263), .c(n_3202), .o(n_3358) );
no02m02 g59228_u0 ( .a(n_3014), .b(conf_wb_err_addr_in_955), .o(g59228_p) );
ao12m02 g59228_u1 ( .a(g59228_p), .b(conf_wb_err_addr_in_955), .c(n_3014), .o(n_3206) );
no02s02 g59229_u0 ( .a(n_3189), .b(wbm_adr_o_14_), .o(g59229_p) );
ao12m02 g59229_u1 ( .a(g59229_p), .b(wbm_adr_o_14_), .c(n_3189), .o(n_3357) );
in01m01 g59230_u0 ( .a(FE_OFN1699_n_5751), .o(g59230_sb) );
na03s02 TIMEBOOST_cell_37731 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__Q), .b(FE_OFN701_n_7845), .c(n_1668), .o(TIMEBOOST_net_11104) );
no02f04 TIMEBOOST_cell_22412 ( .a(FE_RN_769_0), .b(FE_RN_768_0), .o(TIMEBOOST_net_6463) );
na02f04 TIMEBOOST_cell_22461 ( .a(TIMEBOOST_net_6487), .b(FE_OFN1753_n_12086), .o(n_12641) );
in01s01 g59231_u0 ( .a(FE_OFN1698_n_5751), .o(g59231_sb) );
na02s04 TIMEBOOST_cell_45817 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_22__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_787), .o(TIMEBOOST_net_15147) );
no02f04 TIMEBOOST_cell_22413 ( .a(FE_RN_767_0), .b(TIMEBOOST_net_6463), .o(n_14251) );
na02m02 TIMEBOOST_cell_44521 ( .a(n_9586), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__Q), .o(TIMEBOOST_net_14499) );
na02s02 TIMEBOOST_cell_30752 ( .a(g54160_sb), .b(wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_9287) );
na02s01 TIMEBOOST_cell_44877 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__Q), .b(g64280_sb), .o(TIMEBOOST_net_14677) );
na02s02 TIMEBOOST_cell_32021 ( .a(TIMEBOOST_net_9921), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4903) );
in01m02 g59232_u3 ( .a(g59232_p), .o(n_7716) );
oa12f02 g59233_u0 ( .a(n_8480), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__309), .c(FE_OFN1651_n_9428), .o(n_8551) );
in01s02 g59234_u0 ( .a(FE_OFN1145_n_15261), .o(g59234_sb) );
na02s02 TIMEBOOST_cell_45657 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__Q), .b(n_4042), .o(TIMEBOOST_net_15067) );
na02s01 TIMEBOOST_cell_17114 ( .a(wbs_adr_i_13_), .b(FE_OFN1022_n_11877), .o(TIMEBOOST_net_3814) );
na02f02 TIMEBOOST_cell_32713 ( .a(FE_OFN1572_n_11027), .b(TIMEBOOST_net_10267), .o(TIMEBOOST_net_6478) );
oa12f02 g59235_u0 ( .a(n_8485), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_11__465), .c(FE_OFN1691_n_9528), .o(n_8550) );
oa12m02 g59236_u0 ( .a(n_8484), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_13__543), .c(FE_OFN1655_n_9502), .o(n_8549) );
oa12f02 g59237_u0 ( .a(n_8482), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_14__582), .c(FE_OFN1667_n_9477), .o(n_8548) );
oa12f02 g59238_u0 ( .a(n_8481), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_15__621), .c(FE_OFN1631_n_9531), .o(n_8547) );
in01s01 g59239_u0 ( .a(FE_OFN999_n_15978), .o(g59239_sb) );
na02s01 g59239_u1 ( .a(conf_wb_err_bc_in_846), .b(g59239_sb), .o(g59239_da) );
na02m02 TIMEBOOST_cell_41647 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_14__Q), .b(FE_OFN213_n_9124), .o(TIMEBOOST_net_13062) );
na02s02 TIMEBOOST_cell_37906 ( .a(TIMEBOOST_net_11191), .b(g58212_sb), .o(n_9573) );
in01m01 g59240_u0 ( .a(FE_OFN1698_n_5751), .o(g59240_sb) );
na02s02 g59240_u1 ( .a(g59240_sb), .b(wbm_adr_o_6_), .o(g59240_da) );
na02s02 g59240_u2 ( .a(n_2486), .b(FE_OFN1698_n_5751), .o(g59240_db) );
na02m02 g59240_u3 ( .a(g59240_da), .b(g59240_db), .o(n_3356) );
na02s01 TIMEBOOST_cell_44844 ( .a(TIMEBOOST_net_14660), .b(g64862_db), .o(n_3716) );
in01f02 g59294_u0 ( .a(n_5747), .o(n_7092) );
no02f02 g59296_u0 ( .a(n_8759), .b(pci_target_unit_pcit_if_strd_bc_in_719), .o(g59296_p) );
in01f02 g59296_u1 ( .a(g59296_p), .o(n_8760) );
na02s01 g59297_u0 ( .a(n_8759), .b(wbm_adr_o_0_), .o(n_8880) );
na02s01 g59298_u0 ( .a(n_8759), .b(wbm_adr_o_1_), .o(n_8879) );
no02m02 g59299_u0 ( .a(n_3352), .b(FE_OFN1142_n_15261), .o(n_4207) );
na02f02 g59300_u0 ( .a(n_3202), .b(n_3194), .o(g59300_p) );
in01f02 g59300_u1 ( .a(g59300_p), .o(n_3203) );
in01f02 g59302_u0 ( .a(n_15188), .o(n_7712) );
na02s02 g59309_u0 ( .a(n_3200), .b(wbu_addr_in_271), .o(n_3201) );
in01f02 g59311_u0 ( .a(n_8582), .o(n_8527) );
na02f04 g59312_u0 ( .a(n_7027), .b(n_7624), .o(n_8582) );
na02f01 g59313_u0 ( .a(FE_OFN1691_n_9528), .b(n_8483), .o(n_8485) );
na02f01 g59314_u0 ( .a(FE_OFN1655_n_9502), .b(n_8483), .o(n_8484) );
na03m02 TIMEBOOST_cell_34426 ( .a(n_2698), .b(g59369_sb), .c(g59369_db), .o(n_7540) );
na02f01 g59316_u0 ( .a(FE_OFN1667_n_9477), .b(n_8483), .o(n_8482) );
na02f01 g59317_u0 ( .a(FE_OFN1631_n_9531), .b(n_8483), .o(n_8481) );
no02s01 g59318_u0 ( .a(n_2997), .b(FE_OFN778_n_4152), .o(n_3355) );
na02f01 g59319_u0 ( .a(FE_OFN1651_n_9428), .b(n_8483), .o(n_8480) );
no02m02 g59320_u0 ( .a(n_3014), .b(n_1119), .o(n_3015) );
no02m01 g59321_u0 ( .a(n_8759), .b(n_16738), .o(n_14688) );
no02m04 g59322_u0 ( .a(n_1410), .b(n_3014), .o(n_3013) );
no02f02 g59323_u0 ( .a(FE_OFN1143_n_15261), .b(n_2752), .o(n_3199) );
na02m02 g59324_u0 ( .a(wbm_adr_o_18_), .b(n_3197), .o(n_3198) );
na02m02 TIMEBOOST_cell_41657 ( .a(pci_target_unit_pci_target_sm_n_2), .b(n_9178), .o(TIMEBOOST_net_13067) );
na02s01 TIMEBOOST_cell_43308 ( .a(TIMEBOOST_net_13892), .b(g62923_sb), .o(n_6035) );
no02m06 g59327_u0 ( .a(n_7322), .b(n_3310), .o(n_8493) );
ao12f02 g59329_u0 ( .a(n_7552), .b(n_7309), .c(n_3036), .o(n_7824) );
in01s02 g59330_u0 ( .a(n_8590), .o(n_8526) );
na02f02 TIMEBOOST_cell_44308 ( .a(TIMEBOOST_net_14392), .b(FE_OFN1409_n_8567), .o(TIMEBOOST_net_12796) );
in01f04 g59331_u1 ( .a(g59331_p), .o(n_8590) );
ao12f02 g59332_u0 ( .a(n_7822), .b(n_7032), .c(n_3033), .o(n_7709) );
na02s02 g59333_u0 ( .a(n_3195), .b(wbm_adr_o_22_), .o(n_3196) );
ao12f02 g59334_u0 ( .a(n_7822), .b(n_7030), .c(n_3055), .o(n_7708) );
ao12f02 g59335_u0 ( .a(n_7822), .b(n_7029), .c(n_3072), .o(n_7707) );
ao12s02 g59336_u0 ( .a(n_2979), .b(n_7047), .c(pci_target_unit_wbm_sm_pci_tar_read_request), .o(n_7706) );
na03s02 TIMEBOOST_cell_38205 ( .a(g64272_da), .b(g64272_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__Q), .o(TIMEBOOST_net_11341) );
na02s02 TIMEBOOST_cell_37958 ( .a(TIMEBOOST_net_11217), .b(g58199_sb), .o(n_9586) );
in01f04 g59339_u0 ( .a(n_7704), .o(n_7705) );
na02s01 TIMEBOOST_cell_30742 ( .a(pci_ad_i_12_), .b(parchk_pci_ad_reg_in_1216), .o(TIMEBOOST_net_9282) );
ao12f02 g59341_u0 ( .a(n_7822), .b(n_7308), .c(n_2768), .o(n_7823) );
na02s01 TIMEBOOST_cell_43236 ( .a(TIMEBOOST_net_13856), .b(FE_OFN1284_n_4097), .o(TIMEBOOST_net_12599) );
in01f02 g59344_u1 ( .a(g59344_p), .o(n_7551) );
na03f06 TIMEBOOST_cell_45843 ( .a(n_11121), .b(n_11120), .c(n_11119), .o(TIMEBOOST_net_15160) );
in01f02 g59345_u1 ( .a(g59345_p), .o(n_7550) );
na02m02 TIMEBOOST_cell_43959 ( .a(n_9468), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__Q), .o(TIMEBOOST_net_14218) );
in01f02 g59346_u1 ( .a(g59346_p), .o(n_7548) );
na02s01 TIMEBOOST_cell_30904 ( .a(pci_target_unit_pcit_if_strd_addr_in_692), .b(n_2541), .o(TIMEBOOST_net_9363) );
in01f02 g59347_u1 ( .a(g59347_p), .o(n_7547) );
ao12f02 g59348_u0 ( .a(n_12595), .b(n_7220), .c(n_3051), .o(n_7702) );
in01s01 g59350_u0 ( .a(FE_OFN1189_n_5742), .o(g59350_sb) );
na02m02 TIMEBOOST_cell_15924 ( .a(n_1441), .b(n_529), .o(TIMEBOOST_net_3219) );
na02m01 g59350_u2 ( .a(wishbone_slave_unit_wishbone_slave_del_completion_allow), .b(FE_OFN1189_n_5742), .o(g59350_db) );
na02s01 TIMEBOOST_cell_22286 ( .a(g52467_da), .b(FE_OFN1022_n_11877), .o(TIMEBOOST_net_6400) );
na02m02 g59351_u0 ( .a(n_7315), .b(n_1105), .o(n_8529) );
na02m02 TIMEBOOST_cell_32514 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q), .o(TIMEBOOST_net_10168) );
na02s01 TIMEBOOST_cell_42584 ( .a(TIMEBOOST_net_13530), .b(g65878_sb), .o(TIMEBOOST_net_252) );
ao12s01 g59354_u0 ( .a(n_7324), .b(pci_target_unit_del_sync_comp_done_reg_clr), .c(n_2146), .o(n_7699) );
ao12s02 g59355_u0 ( .a(n_7684), .b(n_1069), .c(n_7529), .o(n_7698) );
no02m04 g59356_u0 ( .a(n_3197), .b(n_1356), .o(n_3191) );
na02s01 TIMEBOOST_cell_36526 ( .a(TIMEBOOST_net_10501), .b(FE_OFN243_n_9116), .o(TIMEBOOST_net_3792) );
oa12m02 g59358_u0 ( .a(n_7079), .b(n_7078), .c(wishbone_slave_unit_pci_initiator_if_read_count_3_), .o(n_7544) );
no02f02 g59359_u0 ( .a(n_7325), .b(n_4188), .o(n_7697) );
ao12f02 g59361_u0 ( .a(n_1536), .b(n_7538), .c(n_3386), .o(n_7543) );
ao12f01 g59362_u0 ( .a(n_7316), .b(n_2999), .c(n_15407), .o(n_7695) );
oa12m01 g59363_u0 ( .a(n_7816), .b(n_6943), .c(FE_OCPN1875_n_14526), .o(n_8525) );
no02s02 g59364_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_14_), .b(n_2478), .o(g59364_p) );
ao12s02 g59364_u1 ( .a(g59364_p), .b(pci_target_unit_del_sync_comp_cycle_count_14_), .c(n_2478), .o(n_3185) );
ao12m02 g59365_u0 ( .a(n_3354), .b(conf_wb_err_addr_in_962), .c(FE_OFN1142_n_15261), .o(n_4206) );
oa12m02 g59366_u0 ( .a(n_5735), .b(FE_OFN1188_n_5742), .c(FE_OFN983_n_2700), .o(n_7542) );
no02s02 g59367_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q), .b(n_2474), .o(g59367_p) );
ao12s02 g59367_u1 ( .a(g59367_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q), .c(n_2474), .o(n_3184) );
in01m01 g59368_u0 ( .a(FE_OFN1188_n_5742), .o(g59368_sb) );
na02f02 TIMEBOOST_cell_37142 ( .a(TIMEBOOST_net_10809), .b(FE_RN_847_0), .o(n_14591) );
na02m01 g59368_u2 ( .a(FE_OFN1188_n_5742), .b(wishbone_slave_unit_wishbone_slave_img_hit_0_), .o(g59368_db) );
na02f02 TIMEBOOST_cell_37144 ( .a(n_14549), .b(TIMEBOOST_net_10810), .o(n_14594) );
in01m01 g59369_u0 ( .a(FE_OFN1188_n_5742), .o(g59369_sb) );
na02f02 TIMEBOOST_cell_37146 ( .a(n_14550), .b(TIMEBOOST_net_10811), .o(n_14595) );
na02m01 g59369_u2 ( .a(FE_OFN1188_n_5742), .b(wishbone_slave_unit_wishbone_slave_img_hit_1_), .o(g59369_db) );
na02s01 TIMEBOOST_cell_39294 ( .a(TIMEBOOST_net_11885), .b(g65736_db), .o(n_1607) );
in01s01 g59370_u0 ( .a(FE_OFN1126_g64577_p), .o(g59370_sb) );
na02m02 TIMEBOOST_cell_32712 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__Q), .o(TIMEBOOST_net_10267) );
na02f02 TIMEBOOST_cell_38790 ( .a(TIMEBOOST_net_11633), .b(g57395_db), .o(n_11347) );
na02f04 TIMEBOOST_cell_32711 ( .a(FE_OFN1568_n_11027), .b(TIMEBOOST_net_10266), .o(TIMEBOOST_net_6487) );
in01s01 g59371_u0 ( .a(FE_OFN1126_g64577_p), .o(g59371_sb) );
na02m04 TIMEBOOST_cell_32710 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__Q), .o(TIMEBOOST_net_10266) );
na02f02 TIMEBOOST_cell_38792 ( .a(TIMEBOOST_net_11634), .b(FE_OFN1389_n_8567), .o(n_11468) );
na02f02 TIMEBOOST_cell_32709 ( .a(FE_OFN1572_n_11027), .b(TIMEBOOST_net_10265), .o(TIMEBOOST_net_6486) );
in01s01 g59372_u0 ( .a(FE_OFN1128_g64577_p), .o(g59372_sb) );
na02m02 TIMEBOOST_cell_32708 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__Q), .o(TIMEBOOST_net_10265) );
na02f02 TIMEBOOST_cell_44693 ( .a(n_580), .b(n_14971), .o(TIMEBOOST_net_14585) );
na02f02 TIMEBOOST_cell_41336 ( .a(TIMEBOOST_net_12906), .b(g57319_sb), .o(n_11432) );
in01s01 g59373_u0 ( .a(FE_OFN1126_g64577_p), .o(g59373_sb) );
na02m02 TIMEBOOST_cell_32706 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__Q), .o(TIMEBOOST_net_10264) );
na02f02 TIMEBOOST_cell_38974 ( .a(TIMEBOOST_net_11725), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10719) );
na02s02 TIMEBOOST_cell_43585 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__Q), .b(n_4415), .o(TIMEBOOST_net_14031) );
no02f02 g59374_u0 ( .a(n_3170), .b(wbm_adr_o_29_), .o(g59374_p) );
ao12f02 g59374_u1 ( .a(g59374_p), .b(wbm_adr_o_29_), .c(n_3170), .o(n_4205) );
na02s02 TIMEBOOST_cell_39796 ( .a(TIMEBOOST_net_12136), .b(g63187_sb), .o(n_5778) );
ao22m02 g59376_u0 ( .a(n_9175), .b(n_7684), .c(n_7039), .d(n_2763), .o(n_7685) );
no02s02 g59377_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_7_), .b(n_1716), .o(g59377_p) );
ao12s02 g59377_u1 ( .a(g59377_p), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_7_), .c(n_1716), .o(n_2559) );
in01s01 g59378_u0 ( .a(FE_OFN1126_g64577_p), .o(g59378_sb) );
na02s02 TIMEBOOST_cell_45412 ( .a(TIMEBOOST_net_14944), .b(g62547_sb), .o(n_6473) );
na02s02 TIMEBOOST_cell_43580 ( .a(TIMEBOOST_net_14028), .b(FE_OFN1317_n_6624), .o(TIMEBOOST_net_12232) );
na02f02 TIMEBOOST_cell_41340 ( .a(TIMEBOOST_net_12908), .b(g57435_sb), .o(n_10357) );
in01s01 g59379_u0 ( .a(FE_OFN1132_g64577_p), .o(g59379_sb) );
na03s04 TIMEBOOST_cell_45413 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__Q), .b(n_3733), .c(FE_OFN1319_n_6436), .o(TIMEBOOST_net_14945) );
in01s01 TIMEBOOST_cell_45917 ( .a(wbm_dat_i_18_), .o(TIMEBOOST_net_15224) );
na02f02 TIMEBOOST_cell_41342 ( .a(TIMEBOOST_net_12909), .b(g57459_sb), .o(n_11274) );
in01s01 g59380_u0 ( .a(FE_OFN1132_g64577_p), .o(g59380_sb) );
na02s04 TIMEBOOST_cell_45414 ( .a(TIMEBOOST_net_14945), .b(g62453_sb), .o(n_6691) );
na02f04 TIMEBOOST_cell_41760 ( .a(TIMEBOOST_net_13118), .b(FE_OFN1063_n_15808), .o(TIMEBOOST_net_11136) );
na02f02 TIMEBOOST_cell_41344 ( .a(TIMEBOOST_net_12910), .b(g57570_sb), .o(n_11181) );
in01s01 g59381_u0 ( .a(FE_OFN1126_g64577_p), .o(g59381_sb) );
na02s02 TIMEBOOST_cell_45415 ( .a(n_1602), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__Q), .o(TIMEBOOST_net_14946) );
na02s02 g59381_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__Q), .b(FE_OFN1126_g64577_p), .o(g59381_db) );
na02f02 TIMEBOOST_cell_41346 ( .a(TIMEBOOST_net_12911), .b(g57261_sb), .o(n_10419) );
in01m01 g59382_u0 ( .a(FE_OFN1699_n_5751), .o(g59382_sb) );
na02s01 TIMEBOOST_cell_42701 ( .a(FE_OFN209_n_9126), .b(g57980_sb), .o(TIMEBOOST_net_13589) );
na02f02 TIMEBOOST_cell_37151 ( .a(n_16260), .b(n_16255), .o(TIMEBOOST_net_10814) );
na02f02 TIMEBOOST_cell_37148 ( .a(TIMEBOOST_net_10812), .b(n_14544), .o(n_14589) );
in01m01 g59383_u0 ( .a(FE_OFN1145_n_15261), .o(g59383_sb) );
na02s01 TIMEBOOST_cell_18839 ( .a(TIMEBOOST_net_4676), .b(g62828_sb), .o(n_5320) );
na02s02 g59383_u2 ( .a(conf_wb_err_addr_in_954), .b(FE_OFN1145_n_15261), .o(g59383_db) );
na02s01 TIMEBOOST_cell_18841 ( .a(TIMEBOOST_net_4677), .b(g63130_sb), .o(n_4991) );
in01s01 g59384_u0 ( .a(n_4936), .o(g59384_sb) );
na02s01 TIMEBOOST_cell_36804 ( .a(TIMEBOOST_net_10640), .b(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_4711) );
in01s01 TIMEBOOST_cell_45914 ( .a(TIMEBOOST_net_15220), .o(TIMEBOOST_net_15221) );
na02s02 TIMEBOOST_cell_36782 ( .a(TIMEBOOST_net_10629), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_4653) );
no02s01 g59385_u0 ( .a(wbu_addr_in_259), .b(n_2762), .o(g59385_p) );
ao12m01 g59385_u1 ( .a(g59385_p), .b(wbu_addr_in_259), .c(n_2762), .o(n_3006) );
no02m01 g59386_u0 ( .a(n_2761), .b(wbm_adr_o_10_), .o(g59386_p) );
ao12s02 g59386_u1 ( .a(g59386_p), .b(wbm_adr_o_10_), .c(n_2761), .o(n_3005) );
in01m01 g59387_u0 ( .a(FE_OFN1699_n_5751), .o(g59387_sb) );
na02f02 TIMEBOOST_cell_39137 ( .a(n_10763), .b(FE_RN_480_0), .o(TIMEBOOST_net_11807) );
na03s02 TIMEBOOST_cell_37689 ( .a(n_1869), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__Q), .c(FE_OFN714_n_8140), .o(TIMEBOOST_net_11083) );
na02s01 TIMEBOOST_cell_37732 ( .a(TIMEBOOST_net_11104), .b(g61830_sb), .o(n_8125) );
no02f02 g59388_u0 ( .a(n_1406), .b(n_4702), .o(g59388_p) );
ao12f02 g59388_u1 ( .a(g59388_p), .b(n_1406), .c(n_4702), .o(n_4704) );
no02s01 g59389_u0 ( .a(n_2769), .b(conf_wb_err_addr_in_951), .o(g59389_p) );
ao12s01 g59389_u1 ( .a(g59389_p), .b(conf_wb_err_addr_in_951), .c(n_2769), .o(n_2770) );
no02m02 g59588_u0 ( .a(FE_OFN1189_n_5742), .b(n_2933), .o(n_5745) );
oa12s02 g59589_u0 ( .a(n_4859), .b(n_1660), .c(n_5229), .o(n_7333) );
in01f04 g59591_u0 ( .a(n_16437), .o(n_17032) );
in01f04 g59593_u0 ( .a(n_8483), .o(n_8561) );
in01f01 g59594_u0 ( .a(n_8489), .o(n_8483) );
na02f06 g59595_u0 ( .a(n_16435), .b(n_6943), .o(n_8489) );
na02s01 g59596_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1183), .o(n_7673) );
na02s01 g59597_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1184), .o(n_7672) );
na02s01 g59598_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1185), .o(n_7671) );
na02s01 g59599_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1186), .o(n_7669) );
na02s01 g59600_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_5_), .o(n_7535) );
na02m01 g59601_u0 ( .a(FE_OFN1710_n_4868), .b(parchk_pci_ad_out_in_1168), .o(n_7667) );
na02s01 g59602_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_4_), .o(n_7534) );
na02s01 g59603_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1187), .o(n_7666) );
na02s01 g59604_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_2_), .o(n_7532) );
na02s01 g59605_u0 ( .a(FE_OFN1709_n_4868), .b(pci_ad_o_29_), .o(n_7665) );
na02s01 g59606_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1188), .o(n_7664) );
na02s01 g59607_u0 ( .a(FE_OFN1706_n_4868), .b(parchk_pci_ad_out_in_1189), .o(n_7663) );
na02s01 g59608_u0 ( .a(FE_OFN1706_n_4868), .b(parchk_pci_ad_out_in_1190), .o(n_7661) );
na02s01 g59610_u0 ( .a(FE_OFN1710_n_4868), .b(parchk_pci_ad_out_in_1192), .o(n_7658) );
na02s01 g59611_u0 ( .a(FE_OFN1710_n_4868), .b(parchk_pci_ad_out_in_1193), .o(n_7657) );
na02s01 g59612_u0 ( .a(FE_OFN1709_n_4868), .b(parchk_pci_ad_out_in_1194), .o(n_7656) );
na02s01 g59613_u0 ( .a(FE_OFN1709_n_4868), .b(parchk_pci_ad_out_in_1195), .o(n_7655) );
na02s01 g59614_u0 ( .a(FE_OFN1709_n_4868), .b(parchk_pci_ad_out_in_1196), .o(n_7654) );
na02s01 g59615_u0 ( .a(FE_OFN1710_n_4868), .b(parchk_pci_ad_out_in_1169), .o(n_7653) );
na02s01 g59616_u0 ( .a(FE_OFN1709_n_4868), .b(parchk_pci_ad_out_in_1197), .o(n_7652) );
na02s01 g59617_u0 ( .a(FE_OFN1710_n_4868), .b(parchk_pci_ad_out_in_1170), .o(n_7651) );
na02s01 g59618_u0 ( .a(FE_OFN1705_n_4868), .b(parchk_pci_ad_out_in_1171), .o(n_7650) );
na02s01 g59619_u0 ( .a(FE_OFN1705_n_4868), .b(parchk_pci_ad_out_in_1172), .o(n_7649) );
na02f01 g59620_u0 ( .a(FE_OFN1705_n_4868), .b(parchk_pci_ad_out_in_1173), .o(n_7648) );
na02s02 g59621_u0 ( .a(FE_OFN1705_n_4868), .b(parchk_pci_ad_out_in_1174), .o(n_7647) );
na02f06 g59622_u0 ( .a(n_2762), .b(n_2755), .o(g59622_p) );
in01f06 g59622_u1 ( .a(g59622_p), .o(n_3202) );
na02m02 g59623_u0 ( .a(n_7530), .b(n_7529), .o(g59623_p) );
in01m02 g59623_u1 ( .a(g59623_p), .o(n_7531) );
na02s02 g59624_u0 ( .a(FE_OFN1708_n_4868), .b(parchk_pci_ad_out_in_1175), .o(n_7528) );
na02f02 TIMEBOOST_cell_39136 ( .a(TIMEBOOST_net_11806), .b(FE_OFN1601_n_13995), .o(g53275_p) );
na02s02 g59626_u0 ( .a(FE_OFN1708_n_4868), .b(parchk_pci_ad_out_in_1176), .o(n_7646) );
na02m04 g59627_u0 ( .a(n_2761), .b(n_2756), .o(g59627_p) );
in01m04 g59627_u1 ( .a(g59627_p), .o(n_3189) );
na02s01 g59628_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_26_), .o(n_7527) );
na02s01 g59629_u0 ( .a(FE_OFN1706_n_4868), .b(pci_ad_o_23_), .o(n_7525) );
na02s01 g59630_u0 ( .a(FE_OFN1706_n_4868), .b(pci_ad_o_20_), .o(n_7524) );
na02s01 g59632_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_0_), .o(n_7523) );
na02s01 g59633_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_13_), .o(n_7522) );
na02s01 g59634_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_14_), .o(n_7521) );
na02s01 g59635_u0 ( .a(FE_OFN1706_n_4868), .b(pci_ad_o_15_), .o(n_7519) );
na02s01 g59636_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_17_), .o(n_7518) );
na02s01 g59637_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_18_), .o(n_7645) );
na02s01 g59638_u0 ( .a(FE_OFN1706_n_4868), .b(pci_ad_o_19_), .o(n_7643) );
na02s01 g59639_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_1_), .o(n_7517) );
na02s01 g59640_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_21_), .o(n_7516) );
na02s01 g59641_u0 ( .a(FE_OFN1706_n_4868), .b(pci_ad_o_22_), .o(n_7515) );
na02s01 g59642_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_24_), .o(n_7514) );
na02s01 g59643_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_25_), .o(n_7642) );
na02s01 g59644_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_27_), .o(n_7640) );
na02s01 g59645_u0 ( .a(FE_OFN1709_n_4868), .b(pci_ad_o_28_), .o(n_7639) );
na02s01 g59646_u0 ( .a(FE_OFN1709_n_4868), .b(pci_ad_o_30_), .o(n_7513) );
na02s01 g59647_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_3_), .o(n_7512) );
na02s01 g59648_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_6_), .o(n_7511) );
na02s01 g59649_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_7_), .o(n_7638) );
na02s01 g59650_u0 ( .a(FE_OFN1708_n_4868), .b(pci_ad_o_8_), .o(n_7510) );
na02s01 g59651_u0 ( .a(FE_OFN1708_n_4868), .b(pci_ad_o_9_), .o(n_7637) );
na02m08 g59652_u0 ( .a(n_2769), .b(n_1270), .o(n_3014) );
no02m02 g59653_u0 ( .a(n_2986), .b(FE_OFN1142_n_15261), .o(n_3354) );
na02s01 TIMEBOOST_cell_40668 ( .a(TIMEBOOST_net_12572), .b(g63156_sb), .o(n_5827) );
no02s01 g59655_u0 ( .a(n_2304), .b(FE_OFN778_n_4152), .o(n_2757) );
na02s01 g59656_u0 ( .a(FE_OFN1708_n_4868), .b(pci_ad_o_10_), .o(n_7636) );
na02s01 g59657_u0 ( .a(FE_OFN1708_n_4868), .b(pci_ad_o_11_), .o(n_7509) );
na02s01 g59658_u0 ( .a(FE_OFN1189_n_5742), .b(n_7329), .o(n_7330) );
no02f01 g59659_u0 ( .a(n_16435), .b(n_2134), .o(g59659_p) );
in01m02 g59659_u1 ( .a(g59659_p), .o(n_7508) );
na03s02 TIMEBOOST_cell_38051 ( .a(g64329_da), .b(g64329_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__Q), .o(TIMEBOOST_net_11264) );
no02s02 g59664_u0 ( .a(FE_OFN1189_n_5742), .b(n_1826), .o(n_5743) );
na02s01 g59665_u0 ( .a(FE_OFN1189_n_5742), .b(wishbone_slave_unit_wishbone_slave_img_hit_2_), .o(g59665_p) );
in01s01 g59665_u1 ( .a(g59665_p), .o(n_5741) );
na02s01 g59666_u0 ( .a(FE_OFN1189_n_5742), .b(wishbone_slave_unit_wishbone_slave_img_hit_3_), .o(g59666_p) );
in01s01 g59666_u1 ( .a(g59666_p), .o(n_5740) );
na02s02 g59667_u0 ( .a(n_5725), .b(pciu_cache_lsize_not_zero_in), .o(n_7717) );
na02s01 g59668_u0 ( .a(FE_OFN1188_n_5742), .b(wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q), .o(n_5739) );
na02s01 g59669_u0 ( .a(FE_OFN1188_n_5742), .b(wishbone_slave_unit_wishbone_slave_pref_en_reg_Q), .o(n_5737) );
na02s01 g59670_u0 ( .a(FE_OFN1189_n_5742), .b(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(g59670_p) );
in01s01 g59670_u1 ( .a(g59670_p), .o(n_5736) );
na02s01 g59671_u0 ( .a(FE_OFN1710_n_4868), .b(parchk_pci_ad_out_in), .o(n_7635) );
na02m01 g59672_u0 ( .a(FE_OFN1188_n_5742), .b(wishbone_slave_unit_wishbone_slave_map), .o(n_5735) );
na02m01 g59673_u0 ( .a(FE_OFN1189_n_5742), .b(wishbone_slave_unit_wishbone_slave_img_wallow), .o(n_7326) );
na02s01 g59674_u0 ( .a(FE_OFN1189_n_5742), .b(wishbone_slave_unit_wishbone_slave_img_hit_4_), .o(g59674_p) );
in01s01 g59674_u1 ( .a(g59674_p), .o(n_5733) );
na02s01 TIMEBOOST_cell_42028 ( .a(TIMEBOOST_net_13252), .b(g62551_sb), .o(n_6463) );
na02s02 g59676_u0 ( .a(FE_OFN1708_n_4868), .b(parchk_pci_ad_out_in_1177), .o(n_7634) );
na02s02 g59677_u0 ( .a(FE_OFN1708_n_4868), .b(parchk_pci_ad_out_in_1178), .o(n_7633) );
ao12f02 g59678_u0 ( .a(n_7552), .b(n_4691), .c(n_2906), .o(n_7091) );
na02s02 g59679_u0 ( .a(FE_OFN1708_n_4868), .b(parchk_pci_ad_out_in_1179), .o(n_7632) );
na02s02 g59681_u0 ( .a(FE_OFN1708_n_4868), .b(parchk_pci_ad_out_in_1180), .o(n_7631) );
na02s01 g59682_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1181), .o(n_7630) );
na02s01 g59683_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_16_), .o(n_7629) );
na02s01 g59684_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1182), .o(n_7628) );
na02s01 g59685_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_12_), .o(n_7505) );
na03s02 TIMEBOOST_cell_6341 ( .a(n_4450), .b(FE_OFN643_n_4677), .c(g65275_da), .o(n_4289) );
na03s02 TIMEBOOST_cell_33806 ( .a(FE_OFN231_n_9839), .b(g57995_sb), .c(g57995_db), .o(n_9800) );
na02s02 TIMEBOOST_cell_45416 ( .a(TIMEBOOST_net_14946), .b(FE_OFN1812_n_7845), .o(TIMEBOOST_net_11385) );
na02f02 TIMEBOOST_cell_13018 ( .a(FE_OCP_RBN1978_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__Q), .o(TIMEBOOST_net_3076) );
na02s02 TIMEBOOST_cell_30907 ( .a(TIMEBOOST_net_9364), .b(FE_OFN784_n_2678), .o(TIMEBOOST_net_3752) );
na02f02 TIMEBOOST_cell_42468 ( .a(TIMEBOOST_net_13472), .b(g57234_sb), .o(n_10833) );
no02m02 g59694_u0 ( .a(FE_OFN1189_n_5742), .b(n_2709), .o(n_5732) );
ao12f02 g59695_u0 ( .a(n_12595), .b(n_4819), .c(n_3066), .o(n_7084) );
ao12f02 g59696_u0 ( .a(n_7552), .b(n_4820), .c(n_3064), .o(n_7083) );
ao12f02 g59697_u0 ( .a(n_7552), .b(n_4823), .c(n_3061), .o(n_7082) );
ao12f02 g59698_u0 ( .a(n_7552), .b(n_4824), .c(n_3045), .o(n_7081) );
ao12f02 g59699_u0 ( .a(n_7552), .b(n_4825), .c(n_3059), .o(n_7080) );
in01f10 g59702_u0 ( .a(n_8759), .o(n_14839) );
in01m10 g59716_u0 ( .a(n_8759), .o(n_8757) );
in01f08 g59717_u0 ( .a(n_14837), .o(n_8759) );
in01f04 g59718_u0 ( .a(n_16475), .o(n_14837) );
na02s02 TIMEBOOST_cell_37882 ( .a(TIMEBOOST_net_11179), .b(g58234_sb), .o(n_9544) );
in01f02 g59721_u1 ( .a(g59721_p), .o(n_7821) );
ao12s01 g59723_u0 ( .a(wbu_pci_drcomp_pending_in), .b(pci_target_unit_del_sync_comp_in), .c(pci_target_unit_wbm_sm_pci_tar_read_request), .o(n_7324) );
na02s01 TIMEBOOST_cell_45128 ( .a(TIMEBOOST_net_14802), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_11415) );
na02f02 TIMEBOOST_cell_42498 ( .a(TIMEBOOST_net_13487), .b(g57547_sb), .o(n_10306) );
ao12m01 g59726_u0 ( .a(n_3157), .b(n_2289), .c(wbm_rty_i), .o(n_2998) );
ao12f02 g59727_u0 ( .a(n_7822), .b(n_4899), .c(n_3043), .o(n_7320) );
na02f02 TIMEBOOST_cell_44719 ( .a(TIMEBOOST_net_10238), .b(FE_OCP_RBN1999_n_13971), .o(TIMEBOOST_net_14598) );
na02s01 TIMEBOOST_cell_42702 ( .a(TIMEBOOST_net_13589), .b(g57980_db), .o(n_9111) );
in01f01 g59730_u0 ( .a(n_7715), .o(n_7317) );
oa12f02 g59731_u0 ( .a(n_3402), .b(n_4717), .c(n_2888), .o(n_7715) );
na02m02 TIMEBOOST_cell_41663 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_13__Q), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__Q), .o(TIMEBOOST_net_13070) );
na02f02 TIMEBOOST_cell_41134 ( .a(TIMEBOOST_net_12805), .b(g57314_sb), .o(n_11437) );
oa12f01 g59734_u0 ( .a(n_2616), .b(FE_OCPN1836_n_16798), .c(n_1435), .o(n_7316) );
oa12s01 g59735_u0 ( .a(n_7313), .b(n_7818), .c(n_8540), .o(n_7627) );
na02s02 TIMEBOOST_cell_45658 ( .a(TIMEBOOST_net_15067), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_11427) );
na02f02 TIMEBOOST_cell_42148 ( .a(TIMEBOOST_net_13312), .b(g57529_sb), .o(n_11212) );
oa12m01 g59738_u0 ( .a(n_7311), .b(n_1758), .c(n_3123), .o(n_7626) );
oa12s02 g59739_u0 ( .a(n_7074), .b(FE_OFN732_n_7498), .c(n_2075), .o(n_7500) );
oa12s02 g59740_u0 ( .a(n_7073), .b(FE_OFN732_n_7498), .c(n_2067), .o(n_7499) );
oa12s02 g59741_u0 ( .a(n_7071), .b(FE_OFN732_n_7498), .c(n_2077), .o(n_7497) );
oa12s02 g59742_u0 ( .a(n_7475), .b(n_7818), .c(n_8517), .o(n_7820) );
oa12s02 g59743_u0 ( .a(n_7069), .b(FE_OFN732_n_7498), .c(n_2082), .o(n_7496) );
oa12s02 g59744_u0 ( .a(n_7070), .b(FE_OFN732_n_7498), .c(n_2069), .o(n_7495) );
oa12m01 g59745_u0 ( .a(n_7068), .b(n_7498), .c(n_2076), .o(n_7494) );
oa12s01 g59746_u0 ( .a(n_7474), .b(n_7818), .c(n_2464), .o(n_7819) );
oa12s02 g59747_u0 ( .a(n_7067), .b(n_7498), .c(n_2068), .o(n_7493) );
oa12s01 g59748_u0 ( .a(n_7472), .b(n_7818), .c(n_2319), .o(n_7817) );
oa12s01 g59749_u0 ( .a(n_7066), .b(n_7498), .c(n_2083), .o(n_7492) );
oa12s01 g59750_u0 ( .a(n_7064), .b(n_7498), .c(n_2286), .o(n_7491) );
oa12s01 g59751_u0 ( .a(n_7063), .b(n_7498), .c(n_2080), .o(n_7490) );
oa12m01 g59752_u0 ( .a(n_7062), .b(n_7498), .c(n_2079), .o(n_7489) );
oa12s01 g59753_u0 ( .a(n_7061), .b(n_7498), .c(n_2072), .o(n_7488) );
oa12s01 g59754_u0 ( .a(n_7060), .b(n_7498), .c(n_2070), .o(n_7487) );
oa12s01 g59755_u0 ( .a(n_7059), .b(n_7498), .c(n_8540), .o(n_7486) );
oa12s02 g59756_u0 ( .a(n_7057), .b(FE_OFN732_n_7498), .c(n_1737), .o(n_7485) );
oa12m01 g59757_u0 ( .a(n_7058), .b(n_7498), .c(n_3280), .o(n_7484) );
oa12s02 g59758_u0 ( .a(n_7613), .b(n_8476), .c(n_8517), .o(n_8478) );
oa12m01 g59759_u0 ( .a(n_7610), .b(n_8476), .c(n_2319), .o(n_8477) );
oa12m01 g59760_u0 ( .a(n_7612), .b(n_8476), .c(n_2464), .o(n_8474) );
no02m02 g59761_u0 ( .a(n_2983), .b(conf_wb_err_addr_in_966), .o(g59761_p) );
ao12m02 g59761_u1 ( .a(g59761_p), .b(conf_wb_err_addr_in_966), .c(n_2983), .o(n_3352) );
oa12m02 g59762_u0 ( .a(n_2992), .b(n_2991), .c(wbu_addr_in_274), .o(n_3351) );
in01m02 g59763_u0 ( .a(FE_OFN1330_n_13547), .o(g59763_sb) );
na02f02 TIMEBOOST_cell_43960 ( .a(TIMEBOOST_net_14218), .b(FE_OFN1392_n_8567), .o(TIMEBOOST_net_12873) );
na02s01 TIMEBOOST_cell_37960 ( .a(TIMEBOOST_net_11218), .b(g58148_sb), .o(n_9645) );
na02s02 TIMEBOOST_cell_19283 ( .a(TIMEBOOST_net_4898), .b(g60642_sb), .o(n_5687) );
oa12s01 g59764_u0 ( .a(n_7815), .b(n_8521), .c(n_2464), .o(n_8523) );
ao12f02 g59765_u0 ( .a(n_4696), .b(wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q), .c(FE_OFN1144_n_15261), .o(n_5731) );
oa12m01 g59766_u0 ( .a(n_7814), .b(n_8521), .c(n_2319), .o(n_8522) );
ao12f02 g59767_u0 ( .a(n_3475), .b(conf_wb_err_addr_in_969), .c(FE_OFN1144_n_15261), .o(n_4700) );
ao12s02 g59768_u0 ( .a(n_3172), .b(conf_wb_err_addr_in_950), .c(FE_OFN1142_n_15261), .o(n_3479) );
oa12s02 g59769_u0 ( .a(n_2990), .b(n_2989), .c(wbm_adr_o_17_), .o(n_3350) );
na02s01 TIMEBOOST_cell_15893 ( .a(TIMEBOOST_net_3203), .b(g57780_sb), .o(TIMEBOOST_net_896) );
na02s01 TIMEBOOST_cell_36392 ( .a(TIMEBOOST_net_10434), .b(g65802_db), .o(n_2188) );
na02s01 TIMEBOOST_cell_36394 ( .a(TIMEBOOST_net_10435), .b(g65891_db), .o(n_1573) );
oa12s02 g59771_u0 ( .a(n_3455), .b(n_2034), .c(n_4662), .o(n_4202) );
oa12f01 g59772_u0 ( .a(FE_OCPN1875_n_14526), .b(n_7096), .c(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(n_7816) );
oa12s02 g59773_u0 ( .a(n_3175), .b(n_3174), .c(wbm_adr_o_25_), .o(n_3478) );
oa12s02 g59774_u0 ( .a(n_7055), .b(FE_OFN732_n_7498), .c(n_1743), .o(n_7483) );
oa12s02 g59775_u0 ( .a(n_7054), .b(FE_OFN732_n_7498), .c(n_2041), .o(n_7482) );
oa12s02 g59776_u0 ( .a(n_7053), .b(FE_OFN732_n_7498), .c(n_2040), .o(n_7481) );
oa12s02 g59777_u0 ( .a(n_7052), .b(FE_OFN732_n_7498), .c(n_1746), .o(n_7480) );
oa12s02 g59778_u0 ( .a(n_7051), .b(FE_OFN732_n_7498), .c(n_2052), .o(n_7479) );
oa12s02 g59779_u0 ( .a(n_7050), .b(FE_OFN732_n_7498), .c(n_1740), .o(n_7478) );
oa12s02 g59780_u0 ( .a(n_7049), .b(FE_OFN732_n_7498), .c(n_2074), .o(n_7477) );
oa12s02 g59781_u0 ( .a(n_7048), .b(FE_OFN732_n_7498), .c(n_2084), .o(n_7476) );
na02f02 TIMEBOOST_cell_43961 ( .a(n_8993), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__Q), .o(TIMEBOOST_net_14219) );
no02s02 g59783_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_11_), .b(n_2421), .o(g59783_p) );
ao12s02 g59783_u1 ( .a(g59783_p), .b(pci_target_unit_del_sync_comp_cycle_count_11_), .c(n_2421), .o(n_2997) );
ao12s02 g59784_u0 ( .a(n_3173), .b(conf_wb_err_addr_in_946), .c(FE_OFN1143_n_15261), .o(n_3477) );
no02s02 g59785_u0 ( .a(n_193), .b(n_2425), .o(g59785_p) );
ao12s02 g59785_u1 ( .a(g59785_p), .b(n_193), .c(n_2425), .o(n_2996) );
ao22m02 g59786_u0 ( .a(n_5642), .b(n_13447), .c(FE_OFN1619_n_1787), .d(conf_wb_err_bc_in_846), .o(n_7315) );
na02f02 TIMEBOOST_cell_41104 ( .a(TIMEBOOST_net_12790), .b(g57556_sb), .o(n_10804) );
in01s02 g59788_u0 ( .a(n_4883), .o(n_5730) );
ao22s02 g59789_u0 ( .a(n_925), .b(n_72), .c(n_4694), .d(configuration_icr_bit_2967), .o(n_4883) );
no02s01 g59790_u0 ( .a(n_2035), .b(conf_wb_err_addr_in_947), .o(g59790_p) );
ao12s01 g59790_u1 ( .a(g59790_p), .b(conf_wb_err_addr_in_947), .c(n_2035), .o(n_2752) );
no02s01 g59791_u0 ( .a(wbu_addr_in_255), .b(n_2487), .o(g59791_p) );
ao12s01 g59791_u1 ( .a(g59791_p), .b(wbu_addr_in_255), .c(n_2487), .o(n_2488) );
ao22m02 g59792_u0 ( .a(n_2405), .b(n_7078), .c(n_2014), .d(n_5228), .o(n_7079) );
no02s01 g59793_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_4_), .b(n_1693), .o(g59793_p) );
ao12s01 g59793_u1 ( .a(g59793_p), .b(pci_target_unit_del_sync_comp_cycle_count_4_), .c(n_1693), .o(n_2327) );
no02s01 g59794_u0 ( .a(n_2485), .b(wbm_adr_o_6_), .o(g59794_p) );
ao12s01 g59794_u1 ( .a(g59794_p), .b(wbm_adr_o_6_), .c(n_2485), .o(n_2486) );
no02s01 g59795_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_4_), .b(n_1695), .o(g59795_p) );
ao12s01 g59795_u1 ( .a(g59795_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_4_), .c(n_1695), .o(n_2326) );
in01s01 g59796_u0 ( .a(n_13547), .o(g59796_sb) );
na02s02 TIMEBOOST_cell_42552 ( .a(TIMEBOOST_net_13514), .b(n_1354), .o(TIMEBOOST_net_10385) );
na02s01 g59796_u2 ( .a(n_5641), .b(n_13547), .o(g59796_db) );
na02s01 TIMEBOOST_cell_44952 ( .a(TIMEBOOST_net_14714), .b(g57999_db), .o(n_9794) );
in01s01 g59797_u0 ( .a(FE_OFN1698_n_5751), .o(g59797_sb) );
na02m02 TIMEBOOST_cell_44733 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__Q), .b(FE_OFN1734_n_16317), .o(TIMEBOOST_net_14605) );
na03s01 TIMEBOOST_cell_33545 ( .a(n_1913), .b(g61740_sb), .c(g61740_db), .o(n_8337) );
na03s02 TIMEBOOST_cell_33544 ( .a(n_2006), .b(g61738_sb), .c(g61738_db), .o(n_8341) );
in01s02 g59798_u0 ( .a(FE_OFN1700_n_5751), .o(g59798_sb) );
na02s04 TIMEBOOST_cell_45818 ( .a(TIMEBOOST_net_15147), .b(FE_OFN2135_n_13124), .o(TIMEBOOST_net_14989) );
na02f02 TIMEBOOST_cell_43962 ( .a(TIMEBOOST_net_14219), .b(FE_OFN1384_n_8567), .o(TIMEBOOST_net_13014) );
na02s02 TIMEBOOST_cell_43237 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__Q), .b(n_3769), .o(TIMEBOOST_net_13857) );
in01m02 g59799_u0 ( .a(FE_OFN1083_n_13221), .o(g59799_sb) );
na02m02 g59799_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__Q), .b(g59799_sb), .o(g59799_da) );
na02s02 TIMEBOOST_cell_42553 ( .a(n_1170), .b(n_2136), .o(TIMEBOOST_net_13515) );
na02s02 TIMEBOOST_cell_43389 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__Q), .b(n_3572), .o(TIMEBOOST_net_13933) );
in01m01 g59800_u0 ( .a(FE_OFN1697_n_5751), .o(g59800_sb) );
na02s01 TIMEBOOST_cell_42703 ( .a(FE_OFN250_n_9789), .b(g58005_sb), .o(TIMEBOOST_net_13590) );
na02s02 TIMEBOOST_cell_10369 ( .a(TIMEBOOST_net_1751), .b(g62019_sb), .o(n_7857) );
na02s02 TIMEBOOST_cell_38218 ( .a(TIMEBOOST_net_11347), .b(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_4624) );
in01m01 g59801_u0 ( .a(FE_OFN1697_n_5751), .o(g59801_sb) );
na02m02 TIMEBOOST_cell_44734 ( .a(TIMEBOOST_net_14605), .b(n_12267), .o(n_12696) );
na02f02 TIMEBOOST_cell_42470 ( .a(TIMEBOOST_net_13473), .b(g57094_sb), .o(n_10845) );
na02s02 TIMEBOOST_cell_39442 ( .a(TIMEBOOST_net_11959), .b(TIMEBOOST_net_4271), .o(TIMEBOOST_net_4596) );
no02s02 g59802_u0 ( .a(conf_wb_err_addr_in_958), .b(n_2751), .o(g59802_p) );
ao12s02 g59802_u1 ( .a(g59802_p), .b(conf_wb_err_addr_in_958), .c(n_2751), .o(n_3347) );
no02m02 g59803_u0 ( .a(wbu_addr_in_266), .b(n_2968), .o(g59803_p) );
ao12m02 g59803_u1 ( .a(g59803_p), .b(wbu_addr_in_266), .c(n_2968), .o(n_3346) );
in01m01 g59804_u0 ( .a(n_7618), .o(g59804_sb) );
na02s06 g59804_u1 ( .a(n_16867), .b(g59804_sb), .o(g59804_da) );
na02s02 TIMEBOOST_cell_42554 ( .a(TIMEBOOST_net_13515), .b(n_1160), .o(TIMEBOOST_net_87) );
na02s02 TIMEBOOST_cell_19355 ( .a(TIMEBOOST_net_4934), .b(g60633_sb), .o(n_5703) );
in01m02 g59805_u0 ( .a(n_7618), .o(g59805_sb) );
na02m06 g59805_u1 ( .a(n_16860), .b(g59805_sb), .o(g59805_da) );
na03f04 TIMEBOOST_cell_42555 ( .a(n_3404), .b(n_290), .c(FE_RN_623_0), .o(TIMEBOOST_net_13516) );
na02s02 TIMEBOOST_cell_19357 ( .a(TIMEBOOST_net_4935), .b(g60641_sb), .o(n_5688) );
in01m01 g59806_u0 ( .a(n_7618), .o(g59806_sb) );
na02s04 TIMEBOOST_cell_45814 ( .a(TIMEBOOST_net_15145), .b(FE_OFN2136_n_13124), .o(TIMEBOOST_net_14987) );
na02f04 TIMEBOOST_cell_42556 ( .a(TIMEBOOST_net_13516), .b(FE_RN_622_0), .o(FE_RN_626_0) );
na02s02 TIMEBOOST_cell_19359 ( .a(TIMEBOOST_net_4936), .b(g60612_sb), .o(n_4842) );
in01m01 g59807_u0 ( .a(n_7618), .o(g59807_sb) );
na02s06 g59807_u1 ( .a(n_696), .b(g59807_sb), .o(g59807_da) );
na02m02 TIMEBOOST_cell_32512 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__21__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__21__Q), .o(TIMEBOOST_net_10167) );
na02s02 TIMEBOOST_cell_37908 ( .a(TIMEBOOST_net_11192), .b(g58222_sb), .o(n_9564) );
in01m01 g59808_u0 ( .a(n_7618), .o(g59808_sb) );
na02s02 TIMEBOOST_cell_43414 ( .a(TIMEBOOST_net_13945), .b(n_6554), .o(TIMEBOOST_net_12199) );
na02s02 TIMEBOOST_cell_42557 ( .a(n_2872), .b(n_1968), .o(TIMEBOOST_net_13517) );
na02f02 TIMEBOOST_cell_42186 ( .a(TIMEBOOST_net_13331), .b(FE_OFN1389_n_8567), .o(TIMEBOOST_net_12277) );
in01m01 g59809_u0 ( .a(n_7618), .o(g59809_sb) );
na02s03 TIMEBOOST_cell_44772 ( .a(TIMEBOOST_net_14624), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_13__Q), .o(TIMEBOOST_net_10829) );
na03s02 TIMEBOOST_cell_39443 ( .a(TIMEBOOST_net_4264), .b(g64088_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__Q), .o(TIMEBOOST_net_11960) );
na02s01 TIMEBOOST_cell_45582 ( .a(TIMEBOOST_net_15029), .b(g58426_sb), .o(TIMEBOOST_net_13160) );
in01f02 g59_u0 ( .a(n_15538), .o(n_15539) );
na02s02 TIMEBOOST_cell_45417 ( .a(n_1608), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__Q), .o(TIMEBOOST_net_14947) );
in01s01 TIMEBOOST_cell_45923 ( .a(wbm_dat_i_20_), .o(TIMEBOOST_net_15230) );
na02s02 TIMEBOOST_cell_43609 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__8__Q), .b(n_4363), .o(TIMEBOOST_net_14043) );
na02f02 TIMEBOOST_cell_44662 ( .a(TIMEBOOST_net_14569), .b(FE_OFN1417_n_8567), .o(TIMEBOOST_net_12794) );
na02s02 g60264_u0 ( .a(n_7072), .b(pciu_bar1_in_389), .o(n_7074) );
na02s02 g60265_u0 ( .a(n_7072), .b(pciu_bar1_in_390), .o(n_7073) );
na02s02 g60266_u0 ( .a(n_7072), .b(pciu_bar1_in_391), .o(n_7071) );
na02s02 g60267_u0 ( .a(n_7072), .b(pciu_bar1_in_392), .o(n_7070) );
na02s02 g60268_u0 ( .a(n_7072), .b(pciu_bar1_in_393), .o(n_7069) );
na02s02 g60269_u0 ( .a(n_7072), .b(pciu_bar1_in_394), .o(n_7068) );
na02m02 g60270_u0 ( .a(n_7473), .b(configuration_icr_bit2_0), .o(n_7475) );
na02s02 g60271_u0 ( .a(n_7065), .b(pciu_bar1_in_395), .o(n_7067) );
na02s02 g60272_u0 ( .a(n_7065), .b(pciu_bar1_in_396), .o(n_7066) );
na02s02 g60273_u0 ( .a(n_7473), .b(configuration_icr_bit_2961), .o(n_7474) );
na02s02 g60274_u0 ( .a(n_7065), .b(pciu_bar1_in_397), .o(n_7064) );
na02s02 g60275_u0 ( .a(n_7473), .b(configuration_icr_bit_2967), .o(n_7472) );
na02m02 g60276_u0 ( .a(n_7065), .b(pciu_bar1_in_398), .o(n_7063) );
na02m02 g60277_u0 ( .a(n_7065), .b(pciu_bar1_in_399), .o(n_7062) );
oa12s01 g60278_u0 ( .a(pci_resi_conf_soft_res_in), .b(n_7818), .c(n_8511), .o(n_7313) );
na02s02 g60279_u0 ( .a(n_7065), .b(pciu_bar1_in_400), .o(n_7061) );
na02s02 g60280_u0 ( .a(n_7065), .b(pciu_bar1_in_401), .o(n_7060) );
na02s02 g60281_u0 ( .a(n_7065), .b(pciu_bar1_in_402), .o(n_7059) );
na02s02 g60282_u0 ( .a(n_7056), .b(pciu_bar1_in), .o(n_7058) );
na02s02 g60283_u0 ( .a(n_7056), .b(pciu_bar1_in_380), .o(n_7057) );
na02s02 g60284_u0 ( .a(n_7611), .b(wbu_mrl_en_in_141), .o(n_7613) );
na02s02 g60285_u0 ( .a(n_7611), .b(wbu_pref_en_in_136), .o(n_7612) );
na02s02 g60286_u0 ( .a(n_7611), .b(n_14907), .o(n_7610) );
na02s02 g60287_u0 ( .a(n_7813), .b(pciu_pref_en_in_320), .o(n_7815) );
na02s02 g60288_u0 ( .a(n_7813), .b(n_14910), .o(n_7814) );
na02s02 g60289_u0 ( .a(n_7056), .b(pciu_bar1_in_381), .o(n_7055) );
na02s02 g60290_u0 ( .a(n_7056), .b(pciu_bar1_in_382), .o(n_7054) );
na02m02 g60291_u0 ( .a(n_7056), .b(pciu_bar1_in_383), .o(n_7053) );
na02s02 g60292_u0 ( .a(n_7056), .b(pciu_bar1_in_384), .o(n_7052) );
na02s02 g60293_u0 ( .a(n_7056), .b(pciu_bar1_in_385), .o(n_7051) );
na02s02 g60294_u0 ( .a(n_7056), .b(pciu_bar1_in_386), .o(n_7050) );
na02m02 g60295_u0 ( .a(n_7072), .b(pciu_bar1_in_387), .o(n_7049) );
na02s02 g60296_u0 ( .a(n_7072), .b(pciu_bar1_in_388), .o(n_7048) );
na02s02 g60297_u0 ( .a(n_3174), .b(wbm_adr_o_25_), .o(n_3175) );
no02s02 g60298_u0 ( .a(pci_target_unit_del_sync_comp_in), .b(n_4177), .o(g60298_p) );
in01s02 g60298_u1 ( .a(g60298_p), .o(n_7047) );
na02s02 TIMEBOOST_cell_45745 ( .a(n_3645), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__Q), .o(TIMEBOOST_net_15111) );
na03s02 TIMEBOOST_cell_42029 ( .a(n_50), .b(n_4398), .c(FE_OFN1241_n_4092), .o(TIMEBOOST_net_13253) );
no02m02 g60303_u0 ( .a(n_2476), .b(n_2750), .o(n_2993) );
na02f04 g60304_u0 ( .a(n_2306), .b(n_2487), .o(g60304_p) );
in01f04 g60304_u1 ( .a(g60304_p), .o(n_2762) );
ao12f02 g60305_u0 ( .a(n_7552), .b(n_4803), .c(n_2853), .o(n_7046) );
ao12f02 g60306_u0 ( .a(n_12595), .b(n_4802), .c(n_2848), .o(n_7045) );
na02f01 g60307_u0 ( .a(FE_OCPN1836_n_16798), .b(n_7044), .o(g60307_p) );
in01f02 g60307_u1 ( .a(g60307_p), .o(n_7529) );
na02m02 g60308_u0 ( .a(n_2991), .b(wbu_addr_in_274), .o(n_2992) );
in01s02 g60309_u0 ( .a(n_7310), .o(n_7311) );
na02f01 g60310_u0 ( .a(FE_OCPN1836_n_16798), .b(n_9175), .o(g60310_p) );
in01m02 g60310_u1 ( .a(g60310_p), .o(n_7310) );
na02s01 TIMEBOOST_cell_30746 ( .a(FE_OFN2114_wishbone_slave_unit_pci_initiator_if_data_source), .b(wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_9284) );
na02f02 g60312_u0 ( .a(n_2343), .b(n_16452), .o(n_7043) );
in01m01 g60314_u0 ( .a(n_7040), .o(n_7039) );
na02f02 g60315_u0 ( .a(n_16798), .b(n_15407), .o(n_7040) );
no02m08 g60318_u0 ( .a(n_2035), .b(n_1972), .o(n_2769) );
na02m04 g60319_u0 ( .a(n_2305), .b(n_2485), .o(g60319_p) );
in01m04 g60319_u1 ( .a(g60319_p), .o(n_2761) );
no02f02 g60320_u0 ( .a(n_3344), .b(FE_OFN1144_n_15261), .o(n_3475) );
na02s02 g60321_u0 ( .a(n_1715), .b(n_1714), .o(g60321_p) );
in01s02 g60321_u1 ( .a(g60321_p), .o(n_1716) );
no02m02 g60322_u0 ( .a(n_4162), .b(FE_OFN1144_n_15261), .o(n_4696) );
no02s02 g60323_u0 ( .a(n_2272), .b(FE_OFN1143_n_15261), .o(n_3173) );
no02s02 g60324_u0 ( .a(n_2981), .b(FE_OFN1142_n_15261), .o(n_3172) );
na02s02 g60325_u0 ( .a(n_2989), .b(wbm_adr_o_17_), .o(n_2990) );
no02s01 g60326_u0 ( .a(n_2024), .b(FE_OFN778_n_4152), .o(n_2748) );
na04s02 TIMEBOOST_cell_34191 ( .a(g64330_da), .b(g64330_db), .c(g63126_sb), .d(g63126_db), .o(n_5001) );
in01f01 g60328_u0 ( .a(n_15446), .o(n_7038) );
na02m02 g60330_u0 ( .a(FE_OCPN1836_n_16798), .b(pci_target_unit_pci_target_sm_cnf_progress), .o(g60330_p) );
in01m02 g60330_u1 ( .a(g60330_p), .o(n_7684) );
no02f02 g60331_u0 ( .a(n_5728), .b(n_7031), .o(n_7309) );
no02s02 g60333_u0 ( .a(n_2964), .b(FE_OFN778_n_4152), .o(n_3171) );
in01s02 g60335_u0 ( .a(FE_OFN1188_n_5742), .o(n_5725) );
na03s02 TIMEBOOST_cell_45659 ( .a(configuration_wb_err_data_590), .b(parchk_pci_ad_out_in_1187), .c(g62091_sb), .o(TIMEBOOST_net_15068) );
na02f02 TIMEBOOST_cell_41642 ( .a(FE_OFN1440_n_9372), .b(TIMEBOOST_net_13059), .o(TIMEBOOST_net_11656) );
in01f02 g60339_u1 ( .a(g60339_p), .o(n_7307) );
ao12f02 g60340_u0 ( .a(n_5643), .b(n_16000), .c(n_2856), .o(n_7033) );
na02s01 TIMEBOOST_cell_37734 ( .a(TIMEBOOST_net_11105), .b(g61926_sb), .o(n_7971) );
na02s01 TIMEBOOST_cell_37736 ( .a(TIMEBOOST_net_11106), .b(g61813_sb), .o(n_8166) );
oa12s01 g60343_u0 ( .a(n_4591), .b(n_3437), .c(n_4869), .o(n_4870) );
na02f02 TIMEBOOST_cell_41558 ( .a(TIMEBOOST_net_13017), .b(g57199_sb), .o(n_10835) );
no02s02 g60345_u0 ( .a(n_1191), .b(n_4694), .o(g60345_p) );
in01s02 g60345_u1 ( .a(g60345_p), .o(n_4695) );
oa12s01 g60346_u0 ( .a(n_4080), .b(n_3289), .c(n_15856), .o(n_4693) );
no02f04 g60347_u0 ( .a(n_2874), .b(n_1353), .o(n_3170) );
no02f02 g60348_u0 ( .a(n_4856), .b(n_7031), .o(n_7032) );
no02f02 g60349_u0 ( .a(n_4857), .b(n_7031), .o(n_7030) );
no02f02 g60350_u0 ( .a(n_4858), .b(n_7031), .o(n_7029) );
ao12m01 g60353_u0 ( .a(n_3157), .b(n_2451), .c(wbm_rty_i), .o(n_2988) );
oa12s01 g60354_u0 ( .a(FE_OFN1083_n_13221), .b(n_4719), .c(FE_OCPN1839_n_1238), .o(n_7028) );
oa12m01 g60355_u0 ( .a(n_8451), .b(n_8450), .c(n_8540), .o(n_8520) );
oa12s02 g60356_u0 ( .a(n_8447), .b(n_8446), .c(n_8517), .o(n_8519) );
oa12s02 g60357_u0 ( .a(n_7789), .b(n_8468), .c(n_8517), .o(n_8470) );
oa12s02 g60358_u0 ( .a(n_8515), .b(n_8514), .c(n_8540), .o(n_8542) );
oa12m01 g60359_u0 ( .a(n_8513), .b(n_8512), .c(n_8540), .o(n_8541) );
oa12s02 g60360_u0 ( .a(n_7790), .b(n_8468), .c(n_8540), .o(n_8469) );
oa12s02 g60361_u0 ( .a(n_7788), .b(n_8465), .c(n_8517), .o(n_8467) );
oa12m01 g60362_u0 ( .a(n_7787), .b(n_8465), .c(n_8540), .o(n_8466) );
oa12s01 g60363_u0 ( .a(n_7786), .b(n_7785), .c(n_3280), .o(n_8464) );
oa12s02 g60364_u0 ( .a(n_8445), .b(n_8444), .c(n_8517), .o(n_8518) );
oa12f01 g60365_u0 ( .a(n_2135), .b(n_4816), .c(n_4853), .o(n_7027) );
ao12f08 g60398_u0 ( .a(n_2951), .b(n_3408), .c(FE_OFN191_n_1193), .o(n_4868) );
oa12m01 g60399_u0 ( .a(n_8449), .b(n_8540), .c(FE_OFN2086_n_8448), .o(n_8516) );
oa12s02 g60400_u0 ( .a(n_4211), .b(FE_OFN1183_n_3476), .c(wbm_sel_o_0_), .o(n_4867) );
oa12s02 g60401_u0 ( .a(n_4212), .b(FE_OFN1183_n_3476), .c(wbm_sel_o_1_), .o(n_4866) );
oa12s02 g60402_u0 ( .a(n_4213), .b(FE_OFN1181_n_3476), .c(wbm_sel_o_2_), .o(n_4864) );
oa12s02 g60403_u0 ( .a(n_4216), .b(FE_OFN1181_n_3476), .c(wbm_sel_o_3_), .o(n_4863) );
ao12f02 g60404_u0 ( .a(n_3376), .b(conf_wb_err_addr_in_965), .c(FE_OFN1143_n_15261), .o(n_4201) );
ao12m02 g60405_u0 ( .a(n_4504), .b(conf_wb_err_addr_in_968), .c(FE_OFN1145_n_15261), .o(n_4862) );
oa12s02 g60406_u0 ( .a(n_5758), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q), .c(n_15741), .o(n_7300) );
in01s01 g60407_u0 ( .a(n_7078), .o(g60407_sb) );
na02f02 TIMEBOOST_cell_32511 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_10166), .o(TIMEBOOST_net_6337) );
na02s01 TIMEBOOST_cell_9140 ( .a(pci_target_unit_fifos_pciw_cbe_in_152), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__Q), .o(TIMEBOOST_net_1137) );
na02f02 TIMEBOOST_cell_42999 ( .a(n_2615), .b(n_3293), .o(TIMEBOOST_net_13738) );
na02s02 TIMEBOOST_cell_43539 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__Q), .b(n_4221), .o(TIMEBOOST_net_14008) );
na02s01 TIMEBOOST_cell_9142 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q), .o(TIMEBOOST_net_1138) );
na02m02 TIMEBOOST_cell_30796 ( .a(wbu_addr_in), .b(g58767_sb), .o(TIMEBOOST_net_9309) );
in01s01 g60409_u0 ( .a(n_7078), .o(g60409_sb) );
na02s01 TIMEBOOST_cell_36541 ( .a(TIMEBOOST_net_9321), .b(FE_OFN951_n_2055), .o(TIMEBOOST_net_10509) );
na02s01 TIMEBOOST_cell_18000 ( .a(pci_target_unit_fifos_pciw_addr_data_in_143), .b(g64103_sb), .o(TIMEBOOST_net_4257) );
na02s01 TIMEBOOST_cell_18639 ( .a(TIMEBOOST_net_4576), .b(g63066_sb), .o(n_5118) );
oa12m01 g60410_u0 ( .a(n_4811), .b(n_4197), .c(FE_OFN1171_n_5592), .o(n_5718) );
oa12s01 g60411_u0 ( .a(n_7339), .b(n_3251), .c(n_7608), .o(n_7609) );
ao12f02 g60412_u0 ( .a(n_4198), .b(FE_OFN1612_n_2122), .c(wishbone_slave_unit_pcim_sm_data_in), .o(n_4692) );
ao12f02 g60413_u0 ( .a(n_3375), .b(conf_wb_err_addr_in_957), .c(FE_OFN1144_n_15261), .o(n_4200) );
no02m02 g60414_u0 ( .a(wbm_adr_o_21_), .b(n_2456), .o(g60414_p) );
ao12m02 g60414_u1 ( .a(g60414_p), .b(wbm_adr_o_21_), .c(n_2456), .o(n_2987) );
no02m02 g60415_u0 ( .a(n_2459), .b(conf_wb_err_addr_in_962), .o(g60415_p) );
ao12m02 g60415_u1 ( .a(g60415_p), .b(conf_wb_err_addr_in_962), .c(n_2459), .o(n_2986) );
in01s01 g60416_u0 ( .a(n_7019), .o(n_7298) );
ao22s01 g60417_u0 ( .a(n_7007), .b(n_14922), .c(FE_OFN1159_n_15325), .d(n_7241), .o(n_7019) );
in01s02 g60418_u0 ( .a(n_7018), .o(n_7297) );
ao22s02 g60419_u0 ( .a(n_7015), .b(n_14932), .c(FE_OFN1158_n_15325), .d(n_7295), .o(n_7018) );
in01s01 g60420_u0 ( .a(n_7812), .o(n_8463) );
ao22s01 g60421_u0 ( .a(n_7810), .b(configuration_interrupt_line), .c(n_7809), .d(n_7806), .o(n_7812) );
in01s01 g60422_u0 ( .a(n_7811), .o(n_8462) );
ao22s01 g60423_u0 ( .a(n_7810), .b(configuration_interrupt_line_37), .c(n_7809), .d(n_7802), .o(n_7811) );
in01s01 g60424_u0 ( .a(n_7808), .o(n_8461) );
ao22s01 g60425_u0 ( .a(n_7810), .b(configuration_interrupt_line_38), .c(n_7809), .d(n_7800), .o(n_7808) );
in01s02 g60426_u0 ( .a(n_7807), .o(n_8460) );
ao22m02 g60427_u0 ( .a(n_7804), .b(wbu_mrl_en_in_142), .c(n_7803), .d(n_7806), .o(n_7807) );
in01s02 g60428_u0 ( .a(n_7805), .o(n_8459) );
ao22m02 g60429_u0 ( .a(n_7804), .b(wbu_pref_en_in_137), .c(n_7803), .d(n_7802), .o(n_7805) );
in01s02 g60430_u0 ( .a(n_7801), .o(n_8458) );
ao22m02 g60431_u0 ( .a(n_7804), .b(n_14906), .c(n_7803), .d(n_7800), .o(n_7801) );
in01s01 g60432_u0 ( .a(n_7799), .o(n_8457) );
ao22s01 g60433_u0 ( .a(n_7810), .b(configuration_interrupt_line_42), .c(n_7792), .d(n_7809), .o(n_7799) );
in01m02 g60434_u0 ( .a(n_7296), .o(n_7470) );
ao22m02 g60435_u0 ( .a(n_7293), .b(pciu_am1_in_538), .c(n_16916), .d(n_7295), .o(n_7296) );
in01s01 g60436_u0 ( .a(n_7469), .o(n_7607) );
ao22s01 g60437_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in), .c(n_7466), .d(n_7289), .o(n_7469) );
in01s01 g60438_u0 ( .a(n_7468), .o(n_7606) );
ao22s01 g60439_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_243), .c(n_7466), .d(n_7231), .o(n_7468) );
in01s01 g60440_u0 ( .a(n_7465), .o(n_7605) );
ao22s01 g60441_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_244), .c(n_7466), .d(n_7282), .o(n_7465) );
in01m02 g60442_u0 ( .a(n_7294), .o(n_7464) );
ao22m02 g60443_u0 ( .a(n_7293), .b(pciu_am1_in_539), .c(n_16916), .d(n_7291), .o(n_7294) );
in01s01 g60444_u0 ( .a(n_7463), .o(n_7604) );
ao22s01 g60445_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_245), .c(n_7466), .d(n_7279), .o(n_7463) );
in01m02 g60446_u0 ( .a(n_7462), .o(n_7603) );
ao22m02 g60447_u0 ( .a(n_7420), .b(pciu_bar0_in_364), .c(n_15931), .d(n_7272), .o(n_7462) );
in01s01 g60448_u0 ( .a(n_7461), .o(n_7602) );
ao22s01 g60449_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_246), .c(n_7466), .d(n_7426), .o(n_7461) );
in01m02 g60450_u0 ( .a(n_7290), .o(n_7460) );
ao22m02 g60451_u0 ( .a(n_7283), .b(pciu_am1_in), .c(n_16916), .d(n_7289), .o(n_7290) );
in01s01 g60452_u0 ( .a(n_7459), .o(n_7601) );
ao22s01 g60453_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_247), .c(n_7466), .d(n_7424), .o(n_7459) );
in01m02 g60454_u0 ( .a(n_7288), .o(n_7458) );
ao22m02 g60455_u0 ( .a(n_7273), .b(pciu_am1_in_531), .c(n_16916), .d(n_7287), .o(n_7288) );
in01s01 g60456_u0 ( .a(n_7457), .o(n_7600) );
ao22s01 g60457_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_248), .c(n_7466), .d(n_7422), .o(n_7457) );
in01m02 g60458_u0 ( .a(n_7286), .o(n_7456) );
ao22m02 g60459_u0 ( .a(n_7293), .b(pciu_am1_in_535), .c(n_16916), .d(n_7285), .o(n_7286) );
in01s01 g60460_u0 ( .a(n_7455), .o(n_7599) );
ao22s01 g60461_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_249), .c(n_7466), .d(n_7440), .o(n_7455) );
in01s01 g60462_u0 ( .a(n_7454), .o(n_7598) );
ao22s01 g60463_u0 ( .a(n_7437), .b(configuration_cache_line_size_reg), .c(n_7466), .d(n_7806), .o(n_7454) );
in01m02 g60464_u0 ( .a(n_7284), .o(n_7453) );
ao22m02 g60465_u0 ( .a(n_7283), .b(pciu_am1_in_519), .c(n_16916), .d(n_7282), .o(n_7284) );
in01s02 g60466_u0 ( .a(n_7016), .o(n_7281) );
ao22s02 g60467_u0 ( .a(n_7015), .b(n_14930), .c(FE_OFN1158_n_15325), .d(n_7239), .o(n_7016) );
in01m02 g60468_u0 ( .a(n_7280), .o(n_7452) );
ao22m02 g60469_u0 ( .a(n_7283), .b(pciu_am1_in_520), .c(n_16916), .d(n_7279), .o(n_7280) );
in01m02 g60470_u0 ( .a(n_7278), .o(n_7451) );
ao22m02 g60471_u0 ( .a(n_7283), .b(pciu_am1_in_521), .c(n_16916), .d(n_7426), .o(n_7278) );
in01m02 g60472_u0 ( .a(n_7277), .o(n_7450) );
ao22m02 g60473_u0 ( .a(n_7283), .b(pciu_am1_in_522), .c(n_16916), .d(n_7424), .o(n_7277) );
in01m02 g60474_u0 ( .a(n_7276), .o(n_7449) );
ao22m02 g60475_u0 ( .a(n_7283), .b(pciu_am1_in_523), .c(n_16916), .d(n_7422), .o(n_7276) );
in01m02 g60476_u0 ( .a(n_7275), .o(n_7448) );
ao22m02 g60477_u0 ( .a(n_7283), .b(pciu_am1_in_524), .c(n_16916), .d(n_7440), .o(n_7275) );
in01m02 g60478_u0 ( .a(n_7274), .o(n_7447) );
ao22m02 g60479_u0 ( .a(n_7273), .b(pciu_am1_in_525), .c(n_16916), .d(n_7272), .o(n_7274) );
in01s02 g60480_u0 ( .a(n_7014), .o(n_7271) );
ao22s02 g60481_u0 ( .a(n_7012), .b(n_14913), .c(FE_OFN1159_n_15325), .d(n_7282), .o(n_7014) );
in01m02 g60482_u0 ( .a(n_7270), .o(n_7446) );
ao22m02 g60483_u0 ( .a(n_7273), .b(pciu_am1_in_526), .c(n_16916), .d(n_7269), .o(n_7270) );
in01m02 g60484_u0 ( .a(n_7268), .o(n_7445) );
ao22m02 g60485_u0 ( .a(n_7273), .b(pciu_am1_in_527), .c(n_16916), .d(n_7267), .o(n_7268) );
in01m02 g60486_u0 ( .a(n_7266), .o(n_7444) );
ao22m02 g60487_u0 ( .a(n_7273), .b(pciu_am1_in_529), .c(n_16916), .d(n_7265), .o(n_7266) );
in01s02 g60488_u0 ( .a(n_7013), .o(n_7264) );
ao22s02 g60489_u0 ( .a(n_7012), .b(n_14914), .c(FE_OFN1159_n_15325), .d(n_7279), .o(n_7013) );
in01s02 g60490_u0 ( .a(n_7011), .o(n_7263) );
ao22s02 g60491_u0 ( .a(n_7012), .b(n_14915), .c(FE_OFN1159_n_15325), .d(n_7426), .o(n_7011) );
in01s01 g60492_u0 ( .a(n_7010), .o(n_7262) );
ao22s02 g60493_u0 ( .a(n_7012), .b(n_14916), .c(FE_OFN1159_n_15325), .d(n_7424), .o(n_7010) );
in01s01 g60494_u0 ( .a(n_7009), .o(n_7261) );
ao22s02 g60495_u0 ( .a(n_7012), .b(n_14917), .c(FE_OFN1159_n_15325), .d(n_7422), .o(n_7009) );
in01m02 g60496_u0 ( .a(n_7260), .o(n_7443) );
ao22m02 g60497_u0 ( .a(n_7273), .b(pciu_am1_in_530), .c(n_16916), .d(n_7259), .o(n_7260) );
in01m02 g60498_u0 ( .a(n_7442), .o(n_7597) );
ao22m02 g60499_u0 ( .a(n_7427), .b(pciu_bar0_in_363), .c(n_15931), .d(n_7440), .o(n_7442) );
in01s02 g60500_u0 ( .a(n_7008), .o(n_7258) );
ao22s02 g60501_u0 ( .a(n_7007), .b(n_14919), .c(FE_OFN1159_n_15325), .d(n_7272), .o(n_7008) );
in01s02 g60502_u0 ( .a(n_7006), .o(n_7257) );
ao22s02 g60503_u0 ( .a(n_7007), .b(n_14920), .c(FE_OFN1159_n_15325), .d(n_7269), .o(n_7006) );
in01s02 g60504_u0 ( .a(n_7005), .o(n_7256) );
ao22s02 g60505_u0 ( .a(n_7007), .b(n_14921), .c(FE_OFN1159_n_15325), .d(n_7267), .o(n_7005) );
in01m02 g60506_u0 ( .a(n_7255), .o(n_7439) );
ao22m02 g60507_u0 ( .a(n_7273), .b(pciu_am1_in_532), .c(n_16916), .d(n_7254), .o(n_7255) );
in01s02 g60508_u0 ( .a(n_7004), .o(n_7253) );
ao22s02 g60509_u0 ( .a(n_7007), .b(n_14923), .c(FE_OFN1159_n_15325), .d(n_7265), .o(n_7004) );
in01s02 g60510_u0 ( .a(n_7003), .o(n_7252) );
ao22s02 g60511_u0 ( .a(n_7007), .b(n_14924), .c(FE_OFN1159_n_15325), .d(n_7259), .o(n_7003) );
in01s02 g60512_u0 ( .a(n_7002), .o(n_7251) );
ao22s02 g60513_u0 ( .a(n_7007), .b(n_14925), .c(FE_OFN1158_n_15325), .d(n_7287), .o(n_7002) );
in01s01 g60514_u0 ( .a(n_7438), .o(n_7596) );
ao22s02 g60515_u0 ( .a(n_7437), .b(configuration_cache_line_size_reg_2996), .c(n_7466), .d(n_7802), .o(n_7438) );
in01m02 g60516_u0 ( .a(n_7250), .o(n_7436) );
ao22m02 g60517_u0 ( .a(n_7293), .b(pciu_am1_in_533), .c(n_16916), .d(n_7249), .o(n_7250) );
in01s02 g60518_u0 ( .a(n_7001), .o(n_7248) );
ao22s02 g60519_u0 ( .a(n_7007), .b(n_14926), .c(FE_OFN1158_n_15325), .d(n_7254), .o(n_7001) );
in01s02 g60520_u0 ( .a(n_7000), .o(n_7247) );
ao22s02 g60521_u0 ( .a(n_7015), .b(n_14927), .c(FE_OFN1158_n_15325), .d(n_7249), .o(n_7000) );
in01s01 g60522_u0 ( .a(n_6999), .o(n_7246) );
ao22s01 g60523_u0 ( .a(n_7015), .b(n_14928), .c(FE_OFN1158_n_15325), .d(n_7244), .o(n_6999) );
in01m02 g60524_u0 ( .a(n_7245), .o(n_7435) );
ao22m02 g60525_u0 ( .a(n_7293), .b(pciu_am1_in_534), .c(n_16916), .d(n_7244), .o(n_7245) );
in01s02 g60526_u0 ( .a(n_6998), .o(n_7243) );
ao22s02 g60527_u0 ( .a(n_7015), .b(n_14929), .c(FE_OFN1158_n_15325), .d(n_7285), .o(n_6998) );
in01s01 g60528_u0 ( .a(n_7434), .o(n_7595) );
ao22s01 g60529_u0 ( .a(n_7437), .b(wbu_cache_line_size_in_206), .c(n_7466), .d(n_7800), .o(n_7434) );
in01m02 g60530_u0 ( .a(n_7242), .o(n_7433) );
ao22m02 g60531_u0 ( .a(n_7273), .b(pciu_am1_in_528), .c(n_16916), .d(n_7241), .o(n_7242) );
in01m02 g60532_u0 ( .a(n_7240), .o(n_7432) );
ao22m02 g60533_u0 ( .a(n_7293), .b(pciu_am1_in_536), .c(n_16916), .d(n_7239), .o(n_7240) );
in01s02 g60534_u0 ( .a(n_6997), .o(n_7238) );
ao22s02 g60535_u0 ( .a(n_7015), .b(n_14934), .c(FE_OFN1158_n_15325), .d(n_6996), .o(n_6997) );
in01s02 g60536_u0 ( .a(n_6995), .o(n_7237) );
ao22s02 g60537_u0 ( .a(n_7012), .b(n_14911), .c(FE_OFN1159_n_15325), .d(n_7289), .o(n_6995) );
in01m02 g60538_u0 ( .a(n_6994), .o(n_7236) );
ao22m02 g60539_u0 ( .a(n_7012), .b(n_14912), .c(FE_OFN1159_n_15325), .d(n_7231), .o(n_6994) );
in01m02 g60540_u0 ( .a(n_7235), .o(n_7431) );
ao22m02 g60541_u0 ( .a(n_7293), .b(pciu_am1_in_537), .c(n_16916), .d(n_7234), .o(n_7235) );
na02f02 TIMEBOOST_cell_39155 ( .a(FE_OFN1559_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__31__Q), .o(TIMEBOOST_net_11816) );
in01m02 g60543_u0 ( .a(n_7233), .o(n_7430) );
ao22m02 g60544_u0 ( .a(n_7293), .b(pciu_am1_in_540), .c(n_16916), .d(n_6996), .o(n_7233) );
in01m02 g60545_u0 ( .a(n_7232), .o(n_7429) );
ao22m02 g60546_u0 ( .a(n_7283), .b(pciu_am1_in_518), .c(n_16916), .d(n_7231), .o(n_7232) );
in01m02 g60547_u0 ( .a(n_7428), .o(n_7594) );
ao22m02 g60548_u0 ( .a(n_7427), .b(pciu_bar0_in), .c(n_15931), .d(n_7426), .o(n_7428) );
in01m02 g60549_u0 ( .a(n_7425), .o(n_7593) );
ao22m02 g60550_u0 ( .a(n_7427), .b(pciu_bar0_in_361), .c(n_15931), .d(n_7424), .o(n_7425) );
in01m02 g60551_u0 ( .a(n_7423), .o(n_7592) );
ao22m02 g60552_u0 ( .a(n_7427), .b(pciu_bar0_in_362), .c(n_15931), .d(n_7422), .o(n_7423) );
in01m02 g60553_u0 ( .a(n_7421), .o(n_7591) );
ao22m02 g60554_u0 ( .a(n_7420), .b(pciu_bar0_in_366), .c(n_15931), .d(n_7267), .o(n_7421) );
in01s01 g60555_u0 ( .a(n_7419), .o(n_7590) );
ao22s02 g60556_u0 ( .a(n_7437), .b(wbu_cache_line_size_in_210), .c(n_7792), .d(n_7466), .o(n_7419) );
no02s01 g60557_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_7_), .b(n_2295), .o(g60557_p) );
ao12s01 g60557_u1 ( .a(g60557_p), .b(pci_target_unit_del_sync_comp_cycle_count_7_), .c(n_2295), .o(n_2304) );
in01m02 g60558_u0 ( .a(n_7418), .o(n_7589) );
ao22m02 g60559_u0 ( .a(n_7420), .b(pciu_bar0_in_365), .c(n_15931), .d(n_7269), .o(n_7418) );
in01m02 g60560_u0 ( .a(n_7417), .o(n_7588) );
ao22m02 g60561_u0 ( .a(n_7420), .b(pciu_bar0_in_367), .c(n_15931), .d(n_7241), .o(n_7417) );
in01m02 g60562_u0 ( .a(n_7416), .o(n_7587) );
ao22m02 g60563_u0 ( .a(n_7420), .b(pciu_bar0_in_368), .c(n_15931), .d(n_7265), .o(n_7416) );
in01m02 g60564_u0 ( .a(n_7415), .o(n_7586) );
ao22m02 g60565_u0 ( .a(n_7420), .b(pciu_bar0_in_369), .c(n_15931), .d(n_7259), .o(n_7415) );
in01m02 g60566_u0 ( .a(n_7414), .o(n_7585) );
ao22m02 g60567_u0 ( .a(n_7420), .b(pciu_bar0_in_370), .c(n_15931), .d(n_7287), .o(n_7414) );
in01m02 g60568_u0 ( .a(n_7413), .o(n_7584) );
ao22s02 g60569_u0 ( .a(n_7420), .b(pciu_bar0_in_371), .c(n_15931), .d(n_7254), .o(n_7413) );
in01m02 g60570_u0 ( .a(n_7412), .o(n_7583) );
ao22m02 g60571_u0 ( .a(n_7410), .b(pciu_bar0_in_372), .c(n_15931), .d(n_7249), .o(n_7412) );
in01m02 g60572_u0 ( .a(n_7411), .o(n_7582) );
ao22m02 g60573_u0 ( .a(n_7410), .b(pciu_bar0_in_373), .c(n_15931), .d(n_7244), .o(n_7411) );
in01m02 g60574_u0 ( .a(n_7798), .o(n_8456) );
ao22s02 g60575_u0 ( .a(n_7796), .b(configuration_sync_command_bit0), .c(n_7795), .d(n_7806), .o(n_7798) );
in01m02 g60576_u0 ( .a(n_7409), .o(n_7581) );
ao22m02 g60577_u0 ( .a(n_7410), .b(pciu_bar0_in_374), .c(n_15931), .d(n_7285), .o(n_7409) );
in01m02 g60578_u0 ( .a(n_7408), .o(n_7580) );
ao22m02 g60579_u0 ( .a(n_7410), .b(pciu_bar0_in_375), .c(n_15931), .d(n_7239), .o(n_7408) );
in01m02 g60580_u0 ( .a(n_7407), .o(n_7579) );
ao22m02 g60581_u0 ( .a(n_7410), .b(pciu_bar0_in_376), .c(n_15931), .d(n_7234), .o(n_7407) );
in01m02 g60582_u0 ( .a(n_7406), .o(n_7578) );
ao22m02 g60583_u0 ( .a(n_7410), .b(pciu_bar0_in_377), .c(n_15931), .d(n_7295), .o(n_7406) );
in01m02 g60584_u0 ( .a(n_7405), .o(n_7577) );
ao22m02 g60585_u0 ( .a(n_7410), .b(pciu_bar0_in_378), .c(n_15931), .d(n_7291), .o(n_7405) );
na02s02 TIMEBOOST_cell_42056 ( .a(TIMEBOOST_net_13266), .b(g62581_sb), .o(n_6390) );
in01s01 g60587_u0 ( .a(n_7797), .o(n_8455) );
ao22s02 g60588_u0 ( .a(n_7796), .b(configuration_sync_command_bit1), .c(n_7795), .d(n_7802), .o(n_7797) );
in01m02 g60589_u0 ( .a(n_7404), .o(n_7576) );
ao22m02 g60590_u0 ( .a(n_7410), .b(pciu_bar0_in_379), .c(n_15931), .d(n_6996), .o(n_7404) );
no02s01 g60591_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_7_), .b(n_2275), .o(g60591_p) );
ao12s01 g60591_u1 ( .a(g60591_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_7_), .c(n_2275), .o(n_2302) );
in01s01 g60592_u0 ( .a(n_7794), .o(n_8454) );
ao22s01 g60593_u0 ( .a(n_7796), .b(configuration_command_bit), .c(n_7795), .d(n_7800), .o(n_7794) );
in01s01 g60595_u0 ( .a(n_7793), .o(n_8453) );
ao22s01 g60596_u0 ( .a(n_7796), .b(configuration_sync_command_bit6), .c(n_7795), .d(n_7792), .o(n_7793) );
in01s02 g60597_u0 ( .a(n_6993), .o(n_7229) );
ao22s02 g60598_u0 ( .a(n_7015), .b(n_14931), .c(FE_OFN1158_n_15325), .d(n_7234), .o(n_6993) );
in01s02 g60599_u0 ( .a(n_6992), .o(n_7228) );
ao22s02 g60600_u0 ( .a(n_7012), .b(n_14918), .c(FE_OFN1159_n_15325), .d(n_7440), .o(n_6992) );
in01s02 g60601_u0 ( .a(n_6991), .o(n_7227) );
ao22s02 g60602_u0 ( .a(n_7015), .b(n_14933), .c(FE_OFN1158_n_15325), .d(n_7291), .o(n_6991) );
in01s01 g60603_u0 ( .a(n_6986), .o(g60603_sb) );
na02f02 TIMEBOOST_cell_42238 ( .a(TIMEBOOST_net_13357), .b(FE_OFN1404_n_8567), .o(TIMEBOOST_net_12314) );
na02s01 TIMEBOOST_cell_36528 ( .a(TIMEBOOST_net_10502), .b(g65705_db), .o(n_1948) );
na02s01 TIMEBOOST_cell_42879 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__Q), .b(FE_OFN551_n_9864), .o(TIMEBOOST_net_13678) );
in01s01 g60604_u0 ( .a(FE_OFN1183_n_3476), .o(g60604_sb) );
na02s01 TIMEBOOST_cell_2909 ( .a(TIMEBOOST_net_34), .b(n_1187), .o(n_1425) );
na02f02 TIMEBOOST_cell_40399 ( .a(FE_RN_47_0), .b(n_2409), .o(TIMEBOOST_net_12438) );
na02s01 TIMEBOOST_cell_2910 ( .a(n_261), .b(wbu_addr_in_277), .o(TIMEBOOST_net_35) );
in01s01 g60605_u0 ( .a(FE_OFN1179_n_3476), .o(g60605_sb) );
na02s02 TIMEBOOST_cell_2911 ( .a(TIMEBOOST_net_35), .b(n_1285), .o(n_1286) );
na02s02 TIMEBOOST_cell_39798 ( .a(TIMEBOOST_net_12137), .b(g62479_sb), .o(n_7383) );
na02s01 TIMEBOOST_cell_2912 ( .a(pci_target_unit_del_sync_comp_cycle_count_7_), .b(pci_target_unit_del_sync_comp_cycle_count_8_), .o(TIMEBOOST_net_36) );
in01s01 g60606_u0 ( .a(FE_OFN1185_n_3476), .o(g60606_sb) );
na02s01 TIMEBOOST_cell_2913 ( .a(TIMEBOOST_net_36), .b(n_1690), .o(n_878) );
na02s02 TIMEBOOST_cell_39800 ( .a(TIMEBOOST_net_12138), .b(g62565_sb), .o(n_6427) );
na02f04 TIMEBOOST_cell_2914 ( .a(FE_RN_518_0), .b(FE_RN_521_0), .o(TIMEBOOST_net_37) );
in01s01 g60607_u0 ( .a(FE_OFN1185_n_3476), .o(g60607_sb) );
na02f04 TIMEBOOST_cell_2915 ( .a(TIMEBOOST_net_37), .b(FE_RN_516_0), .o(n_3334) );
na02s02 TIMEBOOST_cell_39802 ( .a(TIMEBOOST_net_12139), .b(g62706_sb), .o(n_6154) );
na02f01 TIMEBOOST_cell_2916 ( .a(n_15680), .b(n_16871), .o(TIMEBOOST_net_38) );
in01s01 g60608_u0 ( .a(FE_OFN1185_n_3476), .o(g60608_sb) );
na02f02 TIMEBOOST_cell_2917 ( .a(TIMEBOOST_net_38), .b(n_16860), .o(n_1805) );
na02s01 TIMEBOOST_cell_44953 ( .a(FE_OFN215_n_9856), .b(g58014_sb), .o(TIMEBOOST_net_14715) );
in01s01 g60609_u0 ( .a(FE_OFN1179_n_3476), .o(g60609_sb) );
na02s01 TIMEBOOST_cell_39804 ( .a(TIMEBOOST_net_12140), .b(n_1650), .o(n_8178) );
na02s01 TIMEBOOST_cell_40700 ( .a(TIMEBOOST_net_12588), .b(g62603_sb), .o(n_6345) );
na02s01 TIMEBOOST_cell_2920 ( .a(n_513), .b(n_1285), .o(TIMEBOOST_net_40) );
in01s01 g60610_u0 ( .a(FE_OFN1185_n_3476), .o(g60610_sb) );
na02m02 TIMEBOOST_cell_2921 ( .a(TIMEBOOST_net_40), .b(n_2237), .o(n_1372) );
na02s01 TIMEBOOST_cell_39460 ( .a(TIMEBOOST_net_11968), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_4583) );
na02s01 TIMEBOOST_cell_2922 ( .a(n_1689), .b(wishbone_slave_unit_del_sync_comp_cycle_count_7_), .o(TIMEBOOST_net_41) );
in01s01 g60611_u0 ( .a(FE_OFN1185_n_3476), .o(g60611_sb) );
na02s01 TIMEBOOST_cell_2923 ( .a(TIMEBOOST_net_41), .b(n_882), .o(n_883) );
na02s02 TIMEBOOST_cell_43498 ( .a(TIMEBOOST_net_13987), .b(FE_OFN1236_n_6391), .o(TIMEBOOST_net_12200) );
na02s02 TIMEBOOST_cell_45660 ( .a(TIMEBOOST_net_15068), .b(FE_OFN1164_n_5615), .o(n_5616) );
in01s01 g60612_u0 ( .a(FE_OFN1185_n_3476), .o(g60612_sb) );
na02s02 TIMEBOOST_cell_38220 ( .a(TIMEBOOST_net_11348), .b(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_4565) );
na02s02 TIMEBOOST_cell_40383 ( .a(n_4473), .b(g64831_db), .o(TIMEBOOST_net_12430) );
na03s02 TIMEBOOST_cell_38403 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__Q), .b(FE_OFN1116_g64577_p), .c(n_4020), .o(TIMEBOOST_net_11440) );
in01s01 g60613_u0 ( .a(FE_OFN1185_n_3476), .o(g60613_sb) );
na02s02 TIMEBOOST_cell_2927 ( .a(TIMEBOOST_net_43), .b(n_1437), .o(n_2018) );
na02s02 TIMEBOOST_cell_40385 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__Q), .b(g64257_sb), .o(TIMEBOOST_net_12431) );
na02s01 TIMEBOOST_cell_2928 ( .a(pci_target_unit_wishbone_master_rty_counter_5_), .b(pci_target_unit_wishbone_master_rty_counter_4_), .o(TIMEBOOST_net_44) );
in01s01 g60614_u0 ( .a(FE_OFN1179_n_3476), .o(g60614_sb) );
na02m02 TIMEBOOST_cell_2929 ( .a(TIMEBOOST_net_44), .b(n_907), .o(n_2001) );
na02m02 TIMEBOOST_cell_38953 ( .a(wbu_sel_in), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_32__Q), .o(TIMEBOOST_net_11715) );
na02s02 TIMEBOOST_cell_45418 ( .a(TIMEBOOST_net_14947), .b(FE_OFN1812_n_7845), .o(TIMEBOOST_net_11386) );
in01s01 g60615_u0 ( .a(FE_OFN1183_n_3476), .o(g60615_sb) );
na02f02 TIMEBOOST_cell_41348 ( .a(TIMEBOOST_net_12912), .b(g57352_sb), .o(n_11396) );
na02f02 TIMEBOOST_cell_2932 ( .a(n_2215), .b(n_1998), .o(TIMEBOOST_net_46) );
in01s01 g60616_u0 ( .a(FE_OFN1185_n_3476), .o(g60616_sb) );
na02f04 TIMEBOOST_cell_2933 ( .a(TIMEBOOST_net_46), .b(n_2214), .o(n_2701) );
na02s01 TIMEBOOST_cell_2934 ( .a(n_1416), .b(n_561), .o(TIMEBOOST_net_47) );
in01s01 g60617_u0 ( .a(FE_OFN1184_n_3476), .o(g60617_sb) );
na02s01 TIMEBOOST_cell_2935 ( .a(TIMEBOOST_net_47), .b(n_1175), .o(n_1417) );
na03s02 TIMEBOOST_cell_34288 ( .a(n_3940), .b(g63016_sb), .c(g63016_db), .o(n_5216) );
na02f08 TIMEBOOST_cell_2936 ( .a(n_15330), .b(n_2092), .o(TIMEBOOST_net_48) );
in01s01 g60618_u0 ( .a(FE_OFN1179_n_3476), .o(g60618_sb) );
na02f08 TIMEBOOST_cell_2937 ( .a(TIMEBOOST_net_48), .b(n_16936), .o(n_3395) );
na03s01 TIMEBOOST_cell_34289 ( .a(n_3830), .b(g63013_sb), .c(g63013_db), .o(n_5223) );
na02f02 TIMEBOOST_cell_44168 ( .a(TIMEBOOST_net_14322), .b(FE_OFN1370_n_8567), .o(TIMEBOOST_net_13393) );
in01s01 g60619_u0 ( .a(FE_OFN1179_n_3476), .o(g60619_sb) );
no02f10 TIMEBOOST_cell_2939 ( .a(TIMEBOOST_net_49), .b(n_15999), .o(n_16000) );
na02s02 TIMEBOOST_cell_45041 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__Q), .b(n_1873), .o(TIMEBOOST_net_14759) );
na02m02 TIMEBOOST_cell_41589 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_0__Q), .b(FE_OFN207_n_9865), .o(TIMEBOOST_net_13033) );
in01s01 g60620_u0 ( .a(FE_OFN1180_n_3476), .o(g60620_sb) );
na02f02 TIMEBOOST_cell_44292 ( .a(TIMEBOOST_net_14384), .b(FE_OFN1425_n_8567), .o(TIMEBOOST_net_12690) );
na02s02 TIMEBOOST_cell_19136 ( .a(wbm_adr_o_25_), .b(FE_OFN1697_n_5751), .o(TIMEBOOST_net_4825) );
na02m01 TIMEBOOST_cell_2942 ( .a(wbs_ack_o), .b(n_16818), .o(TIMEBOOST_net_51) );
in01s01 g60621_u0 ( .a(FE_OFN1181_n_3476), .o(g60621_sb) );
na02s02 TIMEBOOST_cell_2943 ( .a(TIMEBOOST_net_51), .b(n_1349), .o(n_1963) );
na04s02 TIMEBOOST_cell_34291 ( .a(wbs_dat_i_25_), .b(g63592_sb), .c(g63592_db), .d(TIMEBOOST_net_4400), .o(n_7203) );
na03s02 TIMEBOOST_cell_6426 ( .a(g52628_db), .b(g52628_sb), .c(pci_target_unit_pcit_if_strd_addr_in_699), .o(n_14678) );
in01s01 g60622_u0 ( .a(FE_OFN1180_n_3476), .o(g60622_sb) );
na02m02 TIMEBOOST_cell_43963 ( .a(n_9133), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__Q), .o(TIMEBOOST_net_14220) );
na03s02 TIMEBOOST_cell_39441 ( .a(g64109_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__Q), .c(FE_OFN877_g64577_p), .o(TIMEBOOST_net_11959) );
na02s01 TIMEBOOST_cell_43024 ( .a(TIMEBOOST_net_13750), .b(g62739_sb), .o(n_5501) );
in01s01 g60623_u0 ( .a(FE_OFN1180_n_3476), .o(g60623_sb) );
na02f04 TIMEBOOST_cell_2947 ( .a(TIMEBOOST_net_53), .b(n_1074), .o(n_2440) );
na02s01 TIMEBOOST_cell_44850 ( .a(TIMEBOOST_net_14663), .b(g64768_db), .o(n_3781) );
na02s02 TIMEBOOST_cell_43540 ( .a(TIMEBOOST_net_14008), .b(FE_OFN1313_n_6624), .o(TIMEBOOST_net_12247) );
in01s01 g60624_u0 ( .a(FE_OFN1181_n_3476), .o(g60624_sb) );
na02s01 TIMEBOOST_cell_39806 ( .a(TIMEBOOST_net_12141), .b(n_1592), .o(n_8186) );
na02s02 TIMEBOOST_cell_44851 ( .a(n_4672), .b(g64762_sb), .o(TIMEBOOST_net_14664) );
na02s02 TIMEBOOST_cell_40811 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__Q), .b(n_3602), .o(TIMEBOOST_net_12644) );
in01s01 g60625_u0 ( .a(FE_OFN1181_n_3476), .o(g60625_sb) );
na02s01 TIMEBOOST_cell_32020 ( .a(configuration_pci_err_data_522), .b(wbm_dat_o_21_), .o(TIMEBOOST_net_9921) );
na03s02 TIMEBOOST_cell_39445 ( .a(TIMEBOOST_net_4274), .b(g64081_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__Q), .o(TIMEBOOST_net_11961) );
na02f02 TIMEBOOST_cell_44300 ( .a(TIMEBOOST_net_14388), .b(FE_OFN1420_n_8567), .o(TIMEBOOST_net_12739) );
in01s01 g60626_u0 ( .a(FE_OFN1182_n_3476), .o(g60626_sb) );
na02s02 TIMEBOOST_cell_22287 ( .a(TIMEBOOST_net_6400), .b(n_10237), .o(n_11866) );
na02f02 TIMEBOOST_cell_44320 ( .a(TIMEBOOST_net_14398), .b(FE_OFN1383_n_8567), .o(TIMEBOOST_net_12319) );
na02f02 TIMEBOOST_cell_41028 ( .a(TIMEBOOST_net_12752), .b(g57580_sb), .o(n_11171) );
in01s01 g60627_u0 ( .a(FE_OFN1181_n_3476), .o(g60627_sb) );
na02s02 TIMEBOOST_cell_41720 ( .a(TIMEBOOST_net_13098), .b(g64783_db), .o(n_3767) );
na03s02 TIMEBOOST_cell_39447 ( .a(TIMEBOOST_net_3682), .b(g64279_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__Q), .o(TIMEBOOST_net_11962) );
na02s01 TIMEBOOST_cell_41761 ( .a(g64971_db), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q), .o(TIMEBOOST_net_13119) );
in01s01 g60628_u0 ( .a(FE_OFN1181_n_3476), .o(g60628_sb) );
na02s02 TIMEBOOST_cell_45419 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__Q), .b(n_3605), .o(TIMEBOOST_net_14948) );
na02s02 TIMEBOOST_cell_19146 ( .a(wbm_adr_o_24_), .b(FE_OFN1697_n_5751), .o(TIMEBOOST_net_4830) );
na02s01 TIMEBOOST_cell_42610 ( .a(TIMEBOOST_net_13543), .b(FE_OFN223_n_9844), .o(n_9713) );
in01s01 g60629_u0 ( .a(FE_OFN1182_n_3476), .o(g60629_sb) );
na02f02 TIMEBOOST_cell_41350 ( .a(TIMEBOOST_net_12913), .b(g57336_sb), .o(n_10393) );
na02s02 TIMEBOOST_cell_45420 ( .a(TIMEBOOST_net_14948), .b(FE_OFN1261_n_4143), .o(TIMEBOOST_net_12678) );
in01s01 g60630_u0 ( .a(FE_OFN1180_n_3476), .o(g60630_sb) );
na02s01 TIMEBOOST_cell_2957 ( .a(TIMEBOOST_net_58), .b(g54209_sb), .o(n_13181) );
na02m02 TIMEBOOST_cell_44307 ( .a(n_9555), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__Q), .o(TIMEBOOST_net_14392) );
na04s02 TIMEBOOST_cell_6761 ( .a(configuration_wb_err_data_598), .b(FE_OFN1163_n_5615), .c(parchk_pci_ad_out_in_1195), .d(g62099_sb), .o(n_5604) );
in01s01 g60631_u0 ( .a(FE_OFN1180_n_3476), .o(g60631_sb) );
na02f02 TIMEBOOST_cell_3041 ( .a(TIMEBOOST_net_100), .b(n_2701), .o(n_2702) );
na02m02 TIMEBOOST_cell_19152 ( .a(FE_OFN1698_n_5751), .b(wbm_adr_o_30_), .o(TIMEBOOST_net_4833) );
na03s04 TIMEBOOST_cell_3042 ( .a(pciu_pciif_stop_reg_in), .b(wishbone_slave_unit_pci_initiator_sm_transfer), .c(wishbone_slave_unit_pci_initiator_sm_timeout), .o(TIMEBOOST_net_101) );
in01s01 g60632_u0 ( .a(FE_OFN1186_n_3476), .o(g60632_sb) );
na02m02 TIMEBOOST_cell_3043 ( .a(TIMEBOOST_net_101), .b(n_2132), .o(n_2378) );
na02s02 TIMEBOOST_cell_19154 ( .a(wbm_adr_o_22_), .b(FE_OFN1697_n_5751), .o(TIMEBOOST_net_4834) );
na02s02 TIMEBOOST_cell_36848 ( .a(TIMEBOOST_net_10662), .b(n_2418), .o(n_4860) );
in01s01 g60633_u0 ( .a(FE_OFN1179_n_3476), .o(g60633_sb) );
na02s01 TIMEBOOST_cell_2959 ( .a(TIMEBOOST_net_59), .b(g54205_sb), .o(n_13180) );
na02s02 TIMEBOOST_cell_19156 ( .a(parchk_pci_cbe_out_in), .b(FE_OFN1705_n_4868), .o(TIMEBOOST_net_4835) );
na02f02 TIMEBOOST_cell_44338 ( .a(TIMEBOOST_net_14407), .b(FE_OFN1401_n_8567), .o(TIMEBOOST_net_12858) );
in01s01 g60634_u0 ( .a(FE_OFN1179_n_3476), .o(g60634_sb) );
na02s01 TIMEBOOST_cell_2961 ( .a(TIMEBOOST_net_60), .b(g54205_sb), .o(n_13179) );
na02s02 TIMEBOOST_cell_19158 ( .a(parchk_pci_cbe_out_in_1204), .b(FE_OFN1705_n_4868), .o(TIMEBOOST_net_4836) );
na02m02 TIMEBOOST_cell_44339 ( .a(n_9557), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__Q), .o(TIMEBOOST_net_14408) );
in01s01 g60635_u0 ( .a(FE_OFN1179_n_3476), .o(g60635_sb) );
na02s01 TIMEBOOST_cell_2963 ( .a(TIMEBOOST_net_61), .b(g54171_sb), .o(n_13178) );
na02s02 TIMEBOOST_cell_19160 ( .a(parchk_pci_cbe_out_in_1203), .b(FE_OFN1705_n_4868), .o(TIMEBOOST_net_4837) );
na02s02 TIMEBOOST_cell_43634 ( .a(TIMEBOOST_net_14055), .b(FE_OFN2104_g64577_p), .o(TIMEBOOST_net_11408) );
in01s01 g60636_u0 ( .a(FE_OFN1183_n_3476), .o(g60636_sb) );
na02s01 TIMEBOOST_cell_2965 ( .a(TIMEBOOST_net_62), .b(g54171_sb), .o(n_13177) );
na02s02 TIMEBOOST_cell_19162 ( .a(parchk_pci_cbe_out_in_1202), .b(FE_OFN1705_n_4868), .o(TIMEBOOST_net_4838) );
na02f02 TIMEBOOST_cell_44340 ( .a(TIMEBOOST_net_14408), .b(FE_OFN1384_n_8567), .o(TIMEBOOST_net_12791) );
in01s01 g60637_u0 ( .a(FE_OFN1183_n_3476), .o(g60637_sb) );
na02s01 TIMEBOOST_cell_2967 ( .a(TIMEBOOST_net_63), .b(g54209_sb), .o(n_13175) );
na03s01 TIMEBOOST_cell_39465 ( .a(TIMEBOOST_net_3966), .b(g64228_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__Q), .o(TIMEBOOST_net_11971) );
na04s02 TIMEBOOST_cell_6751 ( .a(configuration_wb_err_cs_bit_567), .b(FE_OFN1163_n_5615), .c(parchk_pci_cbe_out_in), .d(g62075_sb), .o(n_5636) );
in01s01 g60638_u0 ( .a(FE_OFN1183_n_3476), .o(g60638_sb) );
na02s01 TIMEBOOST_cell_2969 ( .a(TIMEBOOST_net_64), .b(g54205_sb), .o(n_13185) );
na03s02 TIMEBOOST_cell_39463 ( .a(TIMEBOOST_net_3970), .b(g64240_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__Q), .o(TIMEBOOST_net_11970) );
na04s02 TIMEBOOST_cell_6753 ( .a(configuration_wb_err_data), .b(FE_OFN1163_n_5615), .c(parchk_pci_ad_out_in), .d(g62079_sb), .o(n_5631) );
in01m01 g60639_u0 ( .a(FE_OFN1183_n_3476), .o(g60639_sb) );
na02s01 TIMEBOOST_cell_2971 ( .a(TIMEBOOST_net_65), .b(g54171_sb), .o(n_13184) );
na03s02 TIMEBOOST_cell_37739 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__Q), .b(FE_OFN712_n_8140), .c(n_1599), .o(TIMEBOOST_net_11108) );
na02s01 TIMEBOOST_cell_43107 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__Q), .b(n_4412), .o(TIMEBOOST_net_13792) );
in01m01 g60640_u0 ( .a(FE_OFN1182_n_3476), .o(g60640_sb) );
na02s01 TIMEBOOST_cell_2973 ( .a(TIMEBOOST_net_66), .b(g54216_sb), .o(n_13106) );
na02f02 TIMEBOOST_cell_39139 ( .a(FE_OFN1762_n_10780), .b(TIMEBOOST_net_10250), .o(TIMEBOOST_net_11808) );
na02s02 TIMEBOOST_cell_42966 ( .a(TIMEBOOST_net_13721), .b(g54201_db), .o(n_13418) );
in01s01 g60641_u0 ( .a(FE_OFN1179_n_3476), .o(g60641_sb) );
na02s01 TIMEBOOST_cell_2975 ( .a(TIMEBOOST_net_67), .b(g54209_sb), .o(n_13174) );
na03s02 TIMEBOOST_cell_38191 ( .a(g64288_da), .b(g64288_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__Q), .o(TIMEBOOST_net_11334) );
na02f02 TIMEBOOST_cell_42958 ( .a(TIMEBOOST_net_13717), .b(TIMEBOOST_net_492), .o(n_13360) );
in01s01 g60642_u0 ( .a(FE_OFN1185_n_3476), .o(g60642_sb) );
na02s01 TIMEBOOST_cell_2977 ( .a(TIMEBOOST_net_68), .b(g54216_sb), .o(n_13173) );
na03s02 TIMEBOOST_cell_38231 ( .a(TIMEBOOST_net_3708), .b(g64282_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__Q), .o(TIMEBOOST_net_11354) );
na02f02 TIMEBOOST_cell_42472 ( .a(TIMEBOOST_net_13474), .b(g57566_sb), .o(n_10296) );
in01s01 g60643_u0 ( .a(FE_OFN1185_n_3476), .o(g60643_sb) );
na02s01 TIMEBOOST_cell_2979 ( .a(TIMEBOOST_net_69), .b(g54219_sb), .o(n_13172) );
na02s01 TIMEBOOST_cell_43478 ( .a(TIMEBOOST_net_13977), .b(FE_OFN1236_n_6391), .o(TIMEBOOST_net_12182) );
na02f02 TIMEBOOST_cell_40898 ( .a(TIMEBOOST_net_12687), .b(g57519_sb), .o(n_10317) );
in01s01 g60644_u0 ( .a(FE_OFN1185_n_3476), .o(g60644_sb) );
na02s01 TIMEBOOST_cell_2981 ( .a(TIMEBOOST_net_70), .b(g54167_sb), .o(n_13171) );
na02m02 TIMEBOOST_cell_44169 ( .a(n_9796), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__Q), .o(TIMEBOOST_net_14323) );
na02m02 TIMEBOOST_cell_44221 ( .a(n_8998), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__Q), .o(TIMEBOOST_net_14349) );
in01s01 g60645_u0 ( .a(FE_OFN1185_n_3476), .o(g60645_sb) );
na02s01 TIMEBOOST_cell_2983 ( .a(TIMEBOOST_net_71), .b(g54205_sb), .o(n_13170) );
na02s02 TIMEBOOST_cell_43479 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__Q), .b(n_4270), .o(TIMEBOOST_net_13978) );
na02s02 TIMEBOOST_cell_43094 ( .a(TIMEBOOST_net_13785), .b(g58294_db), .o(n_9511) );
in01s01 g60646_u0 ( .a(FE_OFN1179_n_3476), .o(g60646_sb) );
na02s01 TIMEBOOST_cell_2985 ( .a(TIMEBOOST_net_72), .b(g54209_sb), .o(n_13169) );
na02f02 TIMEBOOST_cell_39141 ( .a(FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__Q), .o(TIMEBOOST_net_11809) );
na02s01 TIMEBOOST_cell_45421 ( .a(TIMEBOOST_net_4810), .b(FE_OFN1200_n_4090), .o(TIMEBOOST_net_14949) );
in01s01 g60647_u0 ( .a(FE_OFN1185_n_3476), .o(g60647_sb) );
na02s01 TIMEBOOST_cell_2987 ( .a(TIMEBOOST_net_73), .b(g54219_sb), .o(n_13168) );
na02s01 TIMEBOOST_cell_37203 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(g65674_sb), .o(TIMEBOOST_net_10840) );
na02s01 TIMEBOOST_cell_31146 ( .a(n_3741), .b(g65066_sb), .o(TIMEBOOST_net_9484) );
in01s01 g60648_u0 ( .a(FE_OFN1184_n_3476), .o(g60648_sb) );
na02s01 TIMEBOOST_cell_2989 ( .a(TIMEBOOST_net_74), .b(g54207_sb), .o(n_13105) );
na02s02 TIMEBOOST_cell_20673 ( .a(TIMEBOOST_net_5593), .b(n_4871), .o(n_4873) );
na02s01 TIMEBOOST_cell_31145 ( .a(TIMEBOOST_net_9483), .b(g65007_db), .o(n_3638) );
in01s01 g60649_u0 ( .a(FE_OFN1185_n_3476), .o(g60649_sb) );
na02s01 TIMEBOOST_cell_2991 ( .a(TIMEBOOST_net_75), .b(g54205_sb), .o(n_13167) );
na02s02 TIMEBOOST_cell_20671 ( .a(TIMEBOOST_net_5592), .b(n_4871), .o(n_4872) );
na03s02 TIMEBOOST_cell_45661 ( .a(configuration_wb_err_data_601), .b(parchk_pci_ad_out_in_1198), .c(g62103_sb), .o(TIMEBOOST_net_15069) );
in01s01 g60650_u0 ( .a(FE_OFN1185_n_3476), .o(g60650_sb) );
na02s01 TIMEBOOST_cell_2993 ( .a(TIMEBOOST_net_76), .b(g54167_sb), .o(n_13182) );
na02s01 TIMEBOOST_cell_43077 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__Q), .b(n_4284), .o(TIMEBOOST_net_13777) );
na02f02 TIMEBOOST_cell_42474 ( .a(TIMEBOOST_net_13475), .b(g57542_sb), .o(n_10812) );
in01s01 g60651_u0 ( .a(FE_OFN1183_n_3476), .o(g60651_sb) );
na02s01 TIMEBOOST_cell_2995 ( .a(TIMEBOOST_net_77), .b(g54207_sb), .o(n_13183) );
na03s02 TIMEBOOST_cell_38081 ( .a(TIMEBOOST_net_3470), .b(g64333_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__Q), .o(TIMEBOOST_net_11279) );
na02s01 TIMEBOOST_cell_31144 ( .a(n_3774), .b(g65007_sb), .o(TIMEBOOST_net_9483) );
in01s01 g60652_u0 ( .a(FE_OFN1185_n_3476), .o(g60652_sb) );
na02s01 TIMEBOOST_cell_2997 ( .a(TIMEBOOST_net_78), .b(g54219_sb), .o(n_13166) );
na03s02 TIMEBOOST_cell_38083 ( .a(TIMEBOOST_net_3995), .b(g64133_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__Q), .o(TIMEBOOST_net_11280) );
na02f02 TIMEBOOST_cell_37806 ( .a(TIMEBOOST_net_11141), .b(FE_OFN2126_n_16497), .o(n_12981) );
in01m01 g60653_u0 ( .a(FE_OFN1184_n_3476), .o(g60653_sb) );
na02s01 TIMEBOOST_cell_2999 ( .a(TIMEBOOST_net_79), .b(g54205_sb), .o(n_13165) );
na03s02 TIMEBOOST_cell_38085 ( .a(TIMEBOOST_net_4256), .b(g65251_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__Q), .o(TIMEBOOST_net_11281) );
na02m02 TIMEBOOST_cell_44301 ( .a(n_9142), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__Q), .o(TIMEBOOST_net_14389) );
in01s01 g60654_u0 ( .a(FE_OFN1180_n_3476), .o(g60654_sb) );
na02s01 TIMEBOOST_cell_3001 ( .a(TIMEBOOST_net_80), .b(g54219_sb), .o(n_13163) );
na03s02 TIMEBOOST_cell_38087 ( .a(TIMEBOOST_net_4272), .b(g60675_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__Q), .o(TIMEBOOST_net_11282) );
na02s02 TIMEBOOST_cell_43076 ( .a(TIMEBOOST_net_13776), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_12033) );
in01s01 g60655_u0 ( .a(FE_OFN1185_n_3476), .o(g60655_sb) );
na02s01 TIMEBOOST_cell_3003 ( .a(TIMEBOOST_net_81), .b(g54205_sb), .o(n_13162) );
na03s02 TIMEBOOST_cell_38089 ( .a(TIMEBOOST_net_4254), .b(g64140_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__Q), .o(TIMEBOOST_net_11283) );
na03m02 TIMEBOOST_cell_32955 ( .a(g58795_db), .b(wbu_addr_in_255), .c(g58795_sb), .o(n_9112) );
in01s01 g60656_u0 ( .a(FE_OFN1181_n_3476), .o(g60656_sb) );
na02s01 TIMEBOOST_cell_3005 ( .a(TIMEBOOST_net_82), .b(g54167_sb), .o(n_13228) );
na02s02 TIMEBOOST_cell_44418 ( .a(TIMEBOOST_net_14447), .b(FE_OFN1305_n_13124), .o(TIMEBOOST_net_13423) );
na02s02 TIMEBOOST_cell_45662 ( .a(TIMEBOOST_net_15069), .b(FE_OFN1164_n_5615), .o(n_5598) );
in01s01 g60657_u0 ( .a(FE_OFN1180_n_3476), .o(g60657_sb) );
na02s01 TIMEBOOST_cell_3007 ( .a(TIMEBOOST_net_83), .b(g54171_sb), .o(n_13223) );
na02s02 TIMEBOOST_cell_42558 ( .a(TIMEBOOST_net_13517), .b(n_1969), .o(TIMEBOOST_net_251) );
na02s01 TIMEBOOST_cell_44847 ( .a(n_3739), .b(g64874_sb), .o(TIMEBOOST_net_14662) );
in01s01 g60658_u0 ( .a(FE_OFN1179_n_3476), .o(g60658_sb) );
na02s01 TIMEBOOST_cell_3009 ( .a(TIMEBOOST_net_84), .b(g54219_sb), .o(n_13161) );
na02s02 TIMEBOOST_cell_37741 ( .a(FE_OFN207_n_9865), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q), .o(TIMEBOOST_net_11109) );
na02s01 TIMEBOOST_cell_41721 ( .a(n_3792), .b(g64829_sb), .o(TIMEBOOST_net_13099) );
in01s01 g60659_u0 ( .a(FE_OFN1181_n_3476), .o(g60659_sb) );
na02s01 TIMEBOOST_cell_3011 ( .a(TIMEBOOST_net_85), .b(g54219_sb), .o(n_13104) );
na02m02 TIMEBOOST_cell_19196 ( .a(n_4806), .b(pciu_bar0_in_371), .o(TIMEBOOST_net_4855) );
na03s02 TIMEBOOST_cell_3012 ( .a(n_1209), .b(n_1167), .c(n_1080), .o(TIMEBOOST_net_86) );
in01s01 g60660_u0 ( .a(FE_OFN1182_n_3476), .o(g60660_sb) );
na02s02 TIMEBOOST_cell_3013 ( .a(TIMEBOOST_net_86), .b(n_1207), .o(n_2232) );
na03s02 TIMEBOOST_cell_38073 ( .a(g64192_da), .b(g64192_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__Q), .o(TIMEBOOST_net_11275) );
na02f02 TIMEBOOST_cell_44644 ( .a(TIMEBOOST_net_14560), .b(FE_OFN2180_n_8567), .o(TIMEBOOST_net_13497) );
in01s01 g60661_u0 ( .a(FE_OFN1182_n_3476), .o(g60661_sb) );
na02s02 TIMEBOOST_cell_3015 ( .a(TIMEBOOST_net_87), .b(n_1168), .o(n_3080) );
na03s02 TIMEBOOST_cell_38067 ( .a(g64177_da), .b(g64177_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__Q), .o(TIMEBOOST_net_11272) );
na02s01 TIMEBOOST_cell_45422 ( .a(TIMEBOOST_net_14949), .b(g62651_sb), .o(n_6243) );
in01s01 g60662_u0 ( .a(FE_OFN1182_n_3476), .o(g60662_sb) );
na02f02 TIMEBOOST_cell_41352 ( .a(TIMEBOOST_net_12914), .b(g57452_sb), .o(n_11282) );
na02m02 TIMEBOOST_cell_39351 ( .a(TIMEBOOST_net_1565), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_393), .o(TIMEBOOST_net_11914) );
na02s02 TIMEBOOST_cell_36707 ( .a(TIMEBOOST_net_333), .b(g61904_sb), .o(TIMEBOOST_net_10592) );
in01s01 g60663_u0 ( .a(FE_OFN1180_n_3476), .o(g60663_sb) );
na02f02 TIMEBOOST_cell_43964 ( .a(TIMEBOOST_net_14220), .b(FE_OFN1407_n_8567), .o(TIMEBOOST_net_12807) );
na03s02 TIMEBOOST_cell_38065 ( .a(g64284_da), .b(g64284_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__Q), .o(TIMEBOOST_net_11271) );
na03s02 TIMEBOOST_cell_3020 ( .a(n_1343), .b(n_1344), .c(n_1253), .o(TIMEBOOST_net_90) );
in01s01 g60664_u0 ( .a(FE_OFN1183_n_3476), .o(g60664_sb) );
na02s02 TIMEBOOST_cell_3021 ( .a(TIMEBOOST_net_90), .b(n_1341), .o(n_2401) );
na03s02 TIMEBOOST_cell_39453 ( .a(TIMEBOOST_net_4037), .b(g64312_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__Q), .o(TIMEBOOST_net_11965) );
in01s01 g60665_u0 ( .a(FE_OFN1180_n_3476), .o(g60665_sb) );
na02f02 TIMEBOOST_cell_40932 ( .a(TIMEBOOST_net_12704), .b(g57247_sb), .o(n_10424) );
in01s01 TIMEBOOST_cell_45893 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_), .o(TIMEBOOST_net_15200) );
na02s01 TIMEBOOST_cell_36706 ( .a(TIMEBOOST_net_10591), .b(g61889_db), .o(n_8052) );
in01s01 g60666_u0 ( .a(FE_OFN1181_n_3476), .o(g60666_sb) );
na02f02 TIMEBOOST_cell_40900 ( .a(TIMEBOOST_net_12688), .b(g57122_sb), .o(n_11624) );
na02f02 TIMEBOOST_cell_39097 ( .a(FE_OCP_RBN1995_n_13971), .b(TIMEBOOST_net_10231), .o(TIMEBOOST_net_11787) );
na03s02 TIMEBOOST_cell_38165 ( .a(TIMEBOOST_net_3545), .b(g64336_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__28__Q), .o(TIMEBOOST_net_11321) );
in01s02 g60667_u0 ( .a(FE_OFN1180_n_3476), .o(g60667_sb) );
na02s01 TIMEBOOST_cell_3027 ( .a(TIMEBOOST_net_93), .b(n_9175), .o(n_2276) );
na02s01 TIMEBOOST_cell_45046 ( .a(TIMEBOOST_net_14761), .b(FE_OFN719_n_8060), .o(TIMEBOOST_net_11252) );
na02f03 TIMEBOOST_cell_3028 ( .a(n_16496), .b(n_978), .o(TIMEBOOST_net_94) );
in01s01 g60668_u0 ( .a(FE_OFN1180_n_3476), .o(g60668_sb) );
na02f06 TIMEBOOST_cell_3029 ( .a(TIMEBOOST_net_94), .b(n_2887), .o(n_15929) );
na02s01 TIMEBOOST_cell_45047 ( .a(n_2033), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__Q), .o(TIMEBOOST_net_14762) );
na02m04 TIMEBOOST_cell_3030 ( .a(n_1165), .b(n_994), .o(TIMEBOOST_net_95) );
in01s01 g60669_u0 ( .a(FE_OFN1179_n_3476), .o(g60669_sb) );
na02m04 TIMEBOOST_cell_3031 ( .a(TIMEBOOST_net_95), .b(n_1669), .o(n_2011) );
na03s02 TIMEBOOST_cell_39455 ( .a(TIMEBOOST_net_3963), .b(g64250_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q), .o(TIMEBOOST_net_11966) );
na02s02 TIMEBOOST_cell_36784 ( .a(TIMEBOOST_net_10630), .b(FE_OFN1134_g64577_p), .o(TIMEBOOST_net_4672) );
in01s01 g60670_u0 ( .a(FE_OFN1183_n_3476), .o(g60670_sb) );
na02s01 TIMEBOOST_cell_3033 ( .a(TIMEBOOST_net_96), .b(n_1632), .o(n_1990) );
na02s01 TIMEBOOST_cell_44793 ( .a(n_3739), .b(g64819_sb), .o(TIMEBOOST_net_14635) );
na02s02 TIMEBOOST_cell_42132 ( .a(TIMEBOOST_net_13304), .b(g62918_sb), .o(n_6043) );
in01s01 g60671_u0 ( .a(n_6986), .o(g60671_sb) );
na02s01 TIMEBOOST_cell_44954 ( .a(TIMEBOOST_net_14715), .b(g58014_db), .o(n_9779) );
na02s02 TIMEBOOST_cell_36530 ( .a(TIMEBOOST_net_10503), .b(FE_OFN1797_n_2299), .o(TIMEBOOST_net_9541) );
na02s01 TIMEBOOST_cell_36532 ( .a(TIMEBOOST_net_10504), .b(g64351_sb), .o(n_3827) );
in01s01 g60672_u0 ( .a(n_6986), .o(g60672_sb) );
na02s01 TIMEBOOST_cell_45133 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__Q), .b(n_3815), .o(TIMEBOOST_net_14805) );
na02s01 TIMEBOOST_cell_36396 ( .a(TIMEBOOST_net_10436), .b(g65699_db), .o(n_2058) );
na03f06 TIMEBOOST_cell_1806 ( .a(n_16268), .b(n_16511), .c(n_15217), .o(FE_RN_302_0) );
in01s01 g60673_u0 ( .a(FE_OFN1183_n_3476), .o(g60673_sb) );
na02s02 TIMEBOOST_cell_41884 ( .a(TIMEBOOST_net_13180), .b(FE_OFN1189_n_5742), .o(TIMEBOOST_net_11390) );
in01s01 TIMEBOOST_cell_45894 ( .a(TIMEBOOST_net_15200), .o(TIMEBOOST_net_15201) );
na02f02 TIMEBOOST_cell_41318 ( .a(TIMEBOOST_net_12897), .b(g57120_sb), .o(n_11625) );
in01s01 g60674_u0 ( .a(n_6986), .o(g60674_sb) );
na02s01 TIMEBOOST_cell_44955 ( .a(FE_OFN247_n_9112), .b(g58096_sb), .o(TIMEBOOST_net_14716) );
na02f02 TIMEBOOST_cell_36912 ( .a(TIMEBOOST_net_10694), .b(g52604_sb), .o(n_10247) );
na02f02 TIMEBOOST_cell_36914 ( .a(TIMEBOOST_net_10695), .b(g52594_sb), .o(n_10279) );
in01s01 g60675_u0 ( .a(FE_OFN923_n_4740), .o(g60675_sb) );
na02s01 TIMEBOOST_cell_39808 ( .a(TIMEBOOST_net_12142), .b(n_1611), .o(n_8193) );
na02s01 g60675_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__Q), .b(FE_OFN923_n_4740), .o(g60675_db) );
na02s02 TIMEBOOST_cell_18461 ( .a(TIMEBOOST_net_4487), .b(g62865_sb), .o(n_5235) );
in01s01 g60676_u0 ( .a(FE_OFN1046_n_16657), .o(g60676_sb) );
na02s01 g60676_u1 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(g60676_sb), .o(g60676_da) );
na02s01 g60676_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__Q), .b(FE_OFN1046_n_16657), .o(g60676_db) );
na02s02 TIMEBOOST_cell_38587 ( .a(TIMEBOOST_net_9957), .b(FE_OFN1185_n_3476), .o(TIMEBOOST_net_11532) );
in01s01 g60677_u0 ( .a(FE_OFN903_n_4736), .o(g60677_sb) );
na02s01 g60677_u1 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(g60677_sb), .o(g60677_da) );
na02s01 g60677_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__Q), .b(FE_OFN903_n_4736), .o(g60677_db) );
in01s01 g60678_u0 ( .a(FE_OFN1012_n_4734), .o(g60678_sb) );
na02s01 g60678_u1 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(g60678_sb), .o(g60678_da) );
na02s01 g60678_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__Q), .b(FE_OFN1012_n_4734), .o(g60678_db) );
no02f04 TIMEBOOST_cell_22291 ( .a(TIMEBOOST_net_6402), .b(n_13577), .o(g53017_p) );
in01m02 g60679_u0 ( .a(FE_OFN1700_n_5751), .o(g60679_sb) );
na02m02 g60679_u1 ( .a(wbm_adr_o_27_), .b(g60679_sb), .o(g60679_da) );
no02f04 TIMEBOOST_cell_19043 ( .a(TIMEBOOST_net_4778), .b(FE_RN_374_0), .o(TIMEBOOST_net_910) );
na02s01 TIMEBOOST_cell_3563 ( .a(TIMEBOOST_net_361), .b(FE_OFN260_n_9860), .o(n_9685) );
oa12s01 g60680_u0 ( .a(n_7369), .b(n_3316), .c(n_7608), .o(n_7791) );
in01s01 g60681_u0 ( .a(FE_OFN1697_n_5751), .o(g60681_sb) );
na03s02 TIMEBOOST_cell_39451 ( .a(TIMEBOOST_net_3688), .b(g64268_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__Q), .o(TIMEBOOST_net_11964) );
na02f02 TIMEBOOST_cell_42187 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__Q), .b(n_9643), .o(TIMEBOOST_net_13332) );
na02m02 TIMEBOOST_cell_22370 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__Q), .o(TIMEBOOST_net_6442) );
in01s01 g60682_u0 ( .a(n_6986), .o(g60682_sb) );
na02s01 g60682_u1 ( .a(wbu_latency_tim_val_in_246), .b(g60682_sb), .o(g60682_da) );
na02s01 TIMEBOOST_cell_15894 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__Q), .b(pci_target_unit_fifos_pcir_flush_in), .o(TIMEBOOST_net_3204) );
na02f04 TIMEBOOST_cell_37150 ( .a(TIMEBOOST_net_10813), .b(n_12378), .o(n_12813) );
ao12f02 g60684_u0 ( .a(n_4855), .b(FE_OFN1006_n_16288), .c(configuration_pci_err_addr_479), .o(n_7220) );
ao12f02 g60685_u0 ( .a(n_4799), .b(configuration_wb_err_data), .c(FE_OFN1071_n_15729), .o(n_6983) );
in01s01 g60686_u0 ( .a(FE_OFN1036_n_4732), .o(g60686_sb) );
na02s01 g60686_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__Q), .b(g60686_sb), .o(g60686_da) );
na02s01 g60686_u2 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(FE_OFN1036_n_4732), .o(g60686_db) );
na03s02 TIMEBOOST_cell_38179 ( .a(TIMEBOOST_net_4039), .b(g64318_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__Q), .o(TIMEBOOST_net_11328) );
in01s01 g60687_u0 ( .a(FE_OFN1059_n_4727), .o(g60687_sb) );
na02s02 TIMEBOOST_cell_38383 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_), .b(g63559_db), .o(TIMEBOOST_net_11430) );
na02s01 g60687_u2 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(FE_OFN1059_n_4727), .o(g60687_db) );
na02s02 TIMEBOOST_cell_38222 ( .a(TIMEBOOST_net_11349), .b(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_4556) );
in01s01 g60688_u0 ( .a(n_4730), .o(g60688_sb) );
na02s02 TIMEBOOST_cell_43561 ( .a(n_156), .b(n_4405), .o(TIMEBOOST_net_14019) );
na03s02 TIMEBOOST_cell_34247 ( .a(TIMEBOOST_net_9799), .b(FE_OFN1174_n_5592), .c(g62073_sb), .o(n_5638) );
na02f02 TIMEBOOST_cell_41690 ( .a(TIMEBOOST_net_10311), .b(TIMEBOOST_net_13083), .o(n_12874) );
in01s01 g60689_u0 ( .a(n_4725), .o(g60689_sb) );
na02s02 TIMEBOOST_cell_38224 ( .a(TIMEBOOST_net_11350), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_4500) );
na02s03 TIMEBOOST_cell_45424 ( .a(TIMEBOOST_net_14950), .b(g53903_sb), .o(n_13538) );
na02s02 TIMEBOOST_cell_38226 ( .a(TIMEBOOST_net_11351), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_4563) );
in01s01 g60690_u0 ( .a(n_6986), .o(g60690_sb) );
na02f02 TIMEBOOST_cell_37052 ( .a(FE_OFN1593_n_13741), .b(TIMEBOOST_net_10764), .o(g53258_p) );
na02f02 TIMEBOOST_cell_36970 ( .a(TIMEBOOST_net_10723), .b(g58825_sb), .o(n_8616) );
in01m01 g60691_u0 ( .a(FE_OFN1699_n_5751), .o(g60691_sb) );
na02s02 TIMEBOOST_cell_45753 ( .a(n_4421), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__Q), .o(TIMEBOOST_net_15115) );
na02s01 TIMEBOOST_cell_37155 ( .a(pci_target_unit_wbm_sm_pci_tar_read_request), .b(pci_target_unit_del_sync_comp_rty_exp_clr), .o(TIMEBOOST_net_10816) );
na02f02 TIMEBOOST_cell_37152 ( .a(n_16258), .b(TIMEBOOST_net_10814), .o(n_16261) );
in01s01 g60692_u0 ( .a(n_7608), .o(g60692_sb) );
na02f02 TIMEBOOST_cell_37068 ( .a(TIMEBOOST_net_10772), .b(FE_OFN1589_n_13736), .o(n_16252) );
na02s01 g60692_u2 ( .a(n_3449), .b(n_7608), .o(g60692_db) );
na02f02 TIMEBOOST_cell_36916 ( .a(TIMEBOOST_net_10696), .b(g52617_sb), .o(n_10139) );
no02s01 g60693_u0 ( .a(wbu_addr_in_262), .b(n_2970), .o(g60693_p) );
ao12s02 g60693_u1 ( .a(g60693_p), .b(wbu_addr_in_262), .c(n_2970), .o(n_3169) );
no02s02 g60694_u0 ( .a(wbm_adr_o_13_), .b(n_2873), .o(g60694_p) );
ao12s02 g60694_u1 ( .a(g60694_p), .b(wbm_adr_o_13_), .c(n_2873), .o(n_3168) );
no02m02 g60695_u0 ( .a(wbu_addr_in_270), .b(n_2462), .o(g60695_p) );
ao12m02 g60695_u1 ( .a(g60695_p), .b(wbu_addr_in_270), .c(n_2462), .o(n_3167) );
no02m01 g60696_u0 ( .a(conf_wb_err_addr_in_954), .b(n_2460), .o(g60696_p) );
ao12m01 g60696_u1 ( .a(g60696_p), .b(conf_wb_err_addr_in_954), .c(n_2460), .o(n_3345) );
na02s01 TIMEBOOST_cell_21937 ( .a(TIMEBOOST_net_6225), .b(g61955_sb), .o(n_6963) );
na02s02 TIMEBOOST_cell_40871 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__Q), .b(n_13181), .o(TIMEBOOST_net_12674) );
na02s01 TIMEBOOST_cell_36320 ( .a(TIMEBOOST_net_10398), .b(g65955_db), .o(n_2166) );
na02s01 TIMEBOOST_cell_16791 ( .a(TIMEBOOST_net_3652), .b(g65374_sb), .o(n_3529) );
na02f02 TIMEBOOST_cell_44297 ( .a(TIMEBOOST_net_10045), .b(g57158_sb), .o(TIMEBOOST_net_14387) );
no02f02 g61546_u0 ( .a(n_4167), .b(n_3227), .o(n_4691) );
na03s03 TIMEBOOST_cell_45777 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__0__Q), .b(n_4364), .c(FE_OFN1316_n_6624), .o(TIMEBOOST_net_15127) );
na02f02 TIMEBOOST_cell_42288 ( .a(TIMEBOOST_net_13382), .b(g57397_sb), .o(n_11344) );
na03s02 TIMEBOOST_cell_33344 ( .a(g65011_sb), .b(g65011_db), .c(n_4450), .o(n_4347) );
na02s02 TIMEBOOST_cell_42981 ( .a(TIMEBOOST_net_4298), .b(FE_OFN2212_n_8407), .o(TIMEBOOST_net_13729) );
oa12m02 g61555_u0 ( .a(n_14909), .b(n_8450), .c(n_8511), .o(n_8451) );
oa12m01 g61556_u0 ( .a(n_14908), .b(FE_OFN2086_n_8448), .c(n_8511), .o(n_8449) );
oa12m01 g61557_u0 ( .a(configuration_pci_err_cs_bit0), .b(n_8446), .c(n_3030), .o(n_8447) );
oa12s02 g61558_u0 ( .a(wbu_bar1_in), .b(n_8468), .c(n_8511), .o(n_7790) );
no02m02 g61559_u0 ( .a(n_2735), .b(n_2750), .o(n_2751) );
oa12s02 g61560_u0 ( .a(wbu_am1_in), .b(n_8514), .c(n_8511), .o(n_8515) );
oa12m01 g61561_u0 ( .a(wbu_map_in_131), .b(n_8468), .c(n_3030), .o(n_7789) );
oa12m01 g61562_u0 ( .a(wbu_map_in_132), .b(n_8465), .c(n_3030), .o(n_7788) );
oa12s02 g61563_u0 ( .a(wbu_bar2_in), .b(n_8465), .c(n_8511), .o(n_7787) );
no02f02 g61564_u0 ( .a(n_4165), .b(n_16168), .o(n_4744) );
oa12s02 g61565_u0 ( .a(wbu_am2_in), .b(n_8512), .c(n_8511), .o(n_8513) );
oa12s02 g61566_u0 ( .a(configuration_sync_command_bit8), .b(n_7785), .c(n_2651), .o(n_7786) );
oa12m02 g61567_u0 ( .a(configuration_wb_err_cs_bit0), .b(n_8444), .c(n_3030), .o(n_8445) );
na02m02 TIMEBOOST_cell_42243 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__Q), .b(n_9696), .o(TIMEBOOST_net_13360) );
na02m02 g61569_u0 ( .a(n_2967), .b(n_2970), .o(g61569_p) );
in01m02 g61569_u1 ( .a(g61569_p), .o(n_2968) );
na02m04 g61570_u0 ( .a(n_1971), .b(n_2970), .o(g61570_p) );
in01f02 g61570_u1 ( .a(g61570_p), .o(n_2971) );
na02s01 g61571_u0 ( .a(n_4666), .b(n_7608), .o(n_7369) );
no02m02 g61572_u0 ( .a(n_7818), .b(n_3030), .o(g61572_p) );
in01s02 g61572_u1 ( .a(g61572_p), .o(n_7473) );
no02f02 g61573_u0 ( .a(n_4172), .b(n_7031), .o(n_4819) );
no02f02 g61574_u0 ( .a(n_4171), .b(n_7031), .o(n_4820) );
no02m02 g61575_u0 ( .a(n_7498), .b(n_8511), .o(g61575_p) );
in01m04 g61575_u1 ( .a(g61575_p), .o(n_7065) );
no02f02 g61576_u0 ( .a(n_5549), .b(n_4146), .o(n_7213) );
no02f02 g61577_u0 ( .a(n_4170), .b(n_7031), .o(n_4823) );
no02f02 g61578_u0 ( .a(n_4169), .b(n_7031), .o(n_4824) );
no02s04 g61579_u0 ( .a(FE_OFN1180_n_3476), .b(n_200), .o(n_4694) );
no02f02 g61580_u0 ( .a(n_4168), .b(n_7031), .o(n_4825) );
no02m02 g61581_u0 ( .a(n_8476), .b(n_3030), .o(g61581_p) );
in01m02 g61581_u1 ( .a(g61581_p), .o(n_7611) );
na02f02 g61582_u0 ( .a(n_4155), .b(n_2768), .o(g61582_p) );
in01f02 g61582_u1 ( .a(g61582_p), .o(n_4826) );
in01f02 g61583_u0 ( .a(n_15377), .o(n_7567) );
in01f02 g61586_u0 ( .a(n_7216), .o(n_13814) );
in01f04 g61587_u0 ( .a(n_6989), .o(n_7216) );
in01f02 g61589_u0 ( .a(n_15467), .o(n_6989) );
no02f02 g61593_u0 ( .a(n_4786), .b(n_4812), .o(n_5717) );
na02s01 g61594_u0 ( .a(n_7738), .b(n_1759), .o(n_8472) );
ao12f02 g61595_u0 ( .a(n_7552), .b(n_4780), .c(n_3393), .o(n_7075) );
na03s02 TIMEBOOST_cell_39457 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q), .b(FE_OFN1134_g64577_p), .c(n_4013), .o(TIMEBOOST_net_11967) );
no02m01 g61597_u0 ( .a(FE_OFN1183_n_3476), .b(n_3342), .o(g61597_p) );
in01m02 g61597_u1 ( .a(g61597_p), .o(n_4871) );
na02f02 g54970_u0 ( .a(n_12468), .b(n_12410), .o(n_16601) );
na02s02 g61599_u0 ( .a(FE_OFN1183_n_3476), .b(configuration_pci_err_cs_bit_467), .o(n_4211) );
na02s02 g61600_u0 ( .a(FE_OFN1183_n_3476), .b(configuration_pci_err_cs_bit_468), .o(n_4212) );
na02s02 g61601_u0 ( .a(FE_OFN1181_n_3476), .b(configuration_pci_err_cs_bit_469), .o(n_4213) );
na02s02 g61602_u0 ( .a(FE_OFN1181_n_3476), .b(configuration_pci_err_cs_bit_470), .o(n_4216) );
na03s02 TIMEBOOST_cell_37735 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__Q), .b(FE_OFN710_n_8232), .c(n_1665), .o(TIMEBOOST_net_11106) );
na02f02 TIMEBOOST_cell_44224 ( .a(TIMEBOOST_net_14350), .b(FE_OFN1423_n_8567), .o(TIMEBOOST_net_12783) );
no02m02 g61606_u0 ( .a(n_8521), .b(n_3030), .o(g61606_p) );
in01m02 g61606_u1 ( .a(g61606_p), .o(n_7813) );
no02m02 g61608_u0 ( .a(n_3153), .b(FE_OFN1144_n_15261), .o(n_3375) );
no02f02 g61609_u0 ( .a(n_3154), .b(FE_OFN1143_n_15261), .o(n_3376) );
no02m02 g61610_u0 ( .a(n_3467), .b(FE_OFN1145_n_15261), .o(n_4504) );
na02m02 g61611_u0 ( .a(n_2460), .b(n_2475), .o(n_2476) );
na02s02 TIMEBOOST_cell_43562 ( .a(TIMEBOOST_net_14019), .b(FE_OFN1236_n_6391), .o(TIMEBOOST_net_12163) );
na02f02 TIMEBOOST_cell_38864 ( .a(TIMEBOOST_net_11670), .b(g58467_sb), .o(n_9381) );
ao12s01 g61614_u0 ( .a(n_7608), .b(n_2807), .c(n_3166), .o(n_7401) );
na02s01 TIMEBOOST_cell_42621 ( .a(n_3780), .b(g64798_sb), .o(TIMEBOOST_net_13549) );
in01s01 g61616_u0 ( .a(n_5228), .o(n_5229) );
na02s02 g61617_u0 ( .a(n_7078), .b(n_692), .o(g61617_p) );
in01s02 g61617_u1 ( .a(g61617_p), .o(n_5228) );
na03s02 TIMEBOOST_cell_43547 ( .a(n_4506), .b(FE_OFN1273_n_4096), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__Q), .o(TIMEBOOST_net_14012) );
na04f04 TIMEBOOST_cell_36219 ( .a(n_14566), .b(n_14475), .c(n_14957), .d(n_14956), .o(n_14611) );
na02f02 TIMEBOOST_cell_42188 ( .a(TIMEBOOST_net_13332), .b(FE_OFN1411_n_8567), .o(TIMEBOOST_net_12283) );
in01m01 g61618_u3 ( .a(g61618_p), .o(n_7115) );
na02f02 TIMEBOOST_cell_42290 ( .a(TIMEBOOST_net_13383), .b(g57292_sb), .o(n_11460) );
na02s01 g61620_u0 ( .a(n_7608), .b(n_16512), .o(n_7339) );
no02f02 g61621_u0 ( .a(n_4197), .b(n_1258), .o(n_4198) );
na02m02 g61622_u0 ( .a(n_15689), .b(n_7622), .o(g61622_p) );
in01m02 g61622_u1 ( .a(g61622_p), .o(n_4822) );
no02s06 g61636_u0 ( .a(n_7498), .b(n_2651), .o(g61636_p) );
in01m04 g61636_u1 ( .a(g61636_p), .o(n_7056) );
no02m02 g61637_u0 ( .a(n_7498), .b(n_2648), .o(g61637_p) );
in01m04 g61637_u1 ( .a(g61637_p), .o(n_7072) );
in01f01 g61641_u0 ( .a(n_16452), .o(n_7096) );
na02s02 TIMEBOOST_cell_43387 ( .a(n_4273), .b(n_4274), .o(TIMEBOOST_net_13932) );
na02m02 TIMEBOOST_cell_32510 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__Q), .o(TIMEBOOST_net_10166) );
no02s01 g61647_u0 ( .a(n_2284), .b(n_1551), .o(n_2285) );
oa12s02 g61649_u0 ( .a(n_7743), .b(FE_OFN1169_n_5592), .c(n_24), .o(n_8510) );
na02m02 TIMEBOOST_cell_41643 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_16__Q), .b(FE_OFN217_n_9889), .o(TIMEBOOST_net_13060) );
na02s01 g61651_u0 ( .a(n_7734), .b(conf_target_abort_recv_in), .o(n_8509) );
ao12f02 g61652_u0 ( .a(n_4808), .b(n_14928), .c(FE_OCPN1900_n_16810), .o(n_6978) );
na02s02 TIMEBOOST_cell_43238 ( .a(TIMEBOOST_net_13857), .b(FE_OFN1279_n_4097), .o(TIMEBOOST_net_12039) );
no02f01 g61654_u0 ( .a(n_6944), .b(n_7398), .o(g61654_p) );
in01f01 g61654_u1 ( .a(g61654_p), .o(n_7399) );
na02s03 TIMEBOOST_cell_45426 ( .a(TIMEBOOST_net_14951), .b(g53924_sb), .o(n_13468) );
oa12s02 g61656_u0 ( .a(n_7742), .b(n_369), .c(FE_OFN1169_n_5592), .o(n_8508) );
na02s01 g61657_u0 ( .a(n_2352), .b(n_3498), .o(n_3499) );
na02m02 TIMEBOOST_cell_44293 ( .a(n_9529), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__Q), .o(TIMEBOOST_net_14385) );
in01s01 g61660_u0 ( .a(n_2420), .o(n_2421) );
no02s02 g61661_u0 ( .a(n_1389), .b(n_2295), .o(n_2420) );
na02s01 g61662_u0 ( .a(n_2369), .b(n_3363), .o(n_3364) );
na02m02 g61663_u0 ( .a(n_2359), .b(n_4894), .o(n_4895) );
na02s01 g61664_u0 ( .a(n_7737), .b(n_2494), .o(n_8506) );
na02f02 TIMEBOOST_cell_42292 ( .a(TIMEBOOST_net_13384), .b(g57465_sb), .o(n_11266) );
in01s02 g61666_u0 ( .a(n_3392), .o(n_3832) );
ao12s02 g61667_u0 ( .a(n_3391), .b(n_3160), .c(n_4078), .o(n_3392) );
na02s01 TIMEBOOST_cell_41712 ( .a(TIMEBOOST_net_13094), .b(g58772_sb), .o(TIMEBOOST_net_9311) );
na02f02 TIMEBOOST_cell_41590 ( .a(TIMEBOOST_net_13033), .b(FE_OFN1436_n_9372), .o(TIMEBOOST_net_11654) );
ao12s01 g61670_u0 ( .a(n_3157), .b(n_1662), .c(wbm_rty_i), .o(n_3076) );
ao12f01 g61671_u0 ( .a(n_4896), .b(n_1200), .c(pci_target_unit_wishbone_master_c_state_2_), .o(n_4897) );
ao12f02 g61672_u0 ( .a(n_4683), .b(FE_OFN1006_n_16288), .c(configuration_pci_err_addr_480), .o(n_4899) );
in01s01 g61673_u0 ( .a(n_2424), .o(n_2425) );
no02s02 g61674_u0 ( .a(n_1392), .b(n_2275), .o(n_2424) );
na02s01 g61675_u0 ( .a(n_2371), .b(n_4894), .o(n_5640) );
in01s01 g61676_u0 ( .a(FE_OFN1166_n_5615), .o(g61676_sb) );
na03s02 TIMEBOOST_cell_41985 ( .a(n_3732), .b(FE_OFN1193_n_6935), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__Q), .o(TIMEBOOST_net_13231) );
na02s02 TIMEBOOST_cell_43619 ( .a(n_4396), .b(n_4397), .o(TIMEBOOST_net_14048) );
na02s01 TIMEBOOST_cell_41986 ( .a(TIMEBOOST_net_13231), .b(g62456_sb), .o(n_6684) );
oa12f01 g61677_u0 ( .a(n_4718), .b(n_4680), .c(n_3480), .o(n_4717) );
oa12s01 g61678_u0 ( .a(n_7565), .b(n_8440), .c(n_4784), .o(n_8442) );
oa12s01 g61679_u0 ( .a(n_7564), .b(n_8440), .c(n_4785), .o(n_8441) );
oa12s01 g61680_u0 ( .a(n_7562), .b(n_8440), .c(n_4782), .o(n_8439) );
oa12s01 g61681_u0 ( .a(n_7561), .b(n_8440), .c(n_4781), .o(n_8438) );
oa12s01 g61684_u0 ( .a(n_7559), .b(n_8440), .c(n_4629), .o(n_8437) );
oa12s01 g61685_u0 ( .a(n_7560), .b(n_8440), .c(n_4631), .o(n_8436) );
oa12s01 g61686_u0 ( .a(n_7558), .b(n_8440), .c(n_4633), .o(n_8434) );
ao12f02 g61687_u0 ( .a(n_3339), .b(conf_wb_err_addr_in_960), .c(FE_OFN1142_n_15261), .o(n_4161) );
ao12m02 g61688_u0 ( .a(n_3468), .b(conf_wb_err_addr_in_964), .c(FE_OFN1145_n_15261), .o(n_4668) );
no02m02 g61689_u0 ( .a(n_3141), .b(wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q), .o(g61689_p) );
ao12m02 g61689_u1 ( .a(g61689_p), .b(wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q), .c(n_3141), .o(n_4162) );
oa12s02 g61690_u0 ( .a(n_7731), .b(n_1755), .c(FE_OFN2079_n_8069), .o(n_8502) );
ao12m02 g61691_u0 ( .a(n_3338), .b(conf_wb_err_addr_in_961), .c(FE_OFN1144_n_15261), .o(n_3474) );
oa12s01 g61692_u0 ( .a(n_7557), .b(n_8440), .c(n_4628), .o(n_8433) );
no02f02 g61693_u0 ( .a(n_2939), .b(n_1461), .o(g61693_p) );
ao12f02 g61693_u1 ( .a(g61693_p), .b(n_1461), .c(n_2939), .o(n_3466) );
oa12s02 g61694_u0 ( .a(n_4813), .b(FE_OFN1169_n_5592), .c(n_2494), .o(n_6218) );
ao12s01 g61695_u0 ( .a(n_7571), .b(configuration_sync_isr_2_delayed_bckp_bit), .c(configuration_sync_isr_2_sync_bckp_bit), .o(n_8432) );
ao12s01 g61696_u0 ( .a(n_7574), .b(configuration_sync_pci_err_cs_8_delayed_bckp_bit), .c(configuration_sync_pci_err_cs_8_sync_bckp_bit), .o(n_8431) );
in01s01 g61697_u0 ( .a(FE_OFN1095_g64577_p), .o(g61697_sb) );
na02s01 TIMEBOOST_cell_36385 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(g65719_sb), .o(TIMEBOOST_net_10431) );
na02s01 g61697_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__Q), .b(FE_OFN1095_g64577_p), .o(g61697_db) );
na02s01 TIMEBOOST_cell_36398 ( .a(TIMEBOOST_net_10437), .b(g65745_db), .o(n_2195) );
in01s01 g61698_u0 ( .a(FE_OFN1097_g64577_p), .o(g61698_sb) );
na02s02 TIMEBOOST_cell_36806 ( .a(TIMEBOOST_net_10641), .b(n_8757), .o(TIMEBOOST_net_532) );
na02s01 g61698_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__Q), .b(FE_OFN1097_g64577_p), .o(g61698_db) );
na02s01 TIMEBOOST_cell_36400 ( .a(TIMEBOOST_net_10438), .b(g65941_db), .o(n_1653) );
in01s01 g61699_u0 ( .a(FE_OFN720_n_8060), .o(g61699_sb) );
na02m01 TIMEBOOST_cell_37738 ( .a(TIMEBOOST_net_11107), .b(n_16748), .o(TIMEBOOST_net_464) );
na02s01 TIMEBOOST_cell_39810 ( .a(TIMEBOOST_net_12143), .b(n_1612), .o(n_8150) );
na02f02 TIMEBOOST_cell_39138 ( .a(TIMEBOOST_net_11807), .b(n_12587), .o(n_12849) );
in01s01 g61700_u0 ( .a(FE_OFN2081_n_8176), .o(g61700_sb) );
na02s02 TIMEBOOST_cell_19957 ( .a(TIMEBOOST_net_5235), .b(g62537_sb), .o(n_6495) );
na02f02 TIMEBOOST_cell_44653 ( .a(n_9002), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__Q), .o(TIMEBOOST_net_14565) );
na02f02 TIMEBOOST_cell_41554 ( .a(TIMEBOOST_net_13015), .b(g57558_sb), .o(n_10803) );
in01s01 g61701_u0 ( .a(FE_OFN720_n_8060), .o(g61701_sb) );
na02f02 TIMEBOOST_cell_39140 ( .a(TIMEBOOST_net_11808), .b(FE_OFN1583_n_12306), .o(n_12754) );
na02s02 TIMEBOOST_cell_38228 ( .a(TIMEBOOST_net_11352), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_4485) );
na02s02 TIMEBOOST_cell_38230 ( .a(TIMEBOOST_net_11353), .b(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_4665) );
in01s01 g61702_u0 ( .a(n_8176), .o(g61702_sb) );
na02s01 TIMEBOOST_cell_45057 ( .a(FE_OFN268_n_9880), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__Q), .o(TIMEBOOST_net_14767) );
na02s01 TIMEBOOST_cell_44878 ( .a(TIMEBOOST_net_14677), .b(g64280_db), .o(n_3893) );
na02s02 TIMEBOOST_cell_39812 ( .a(TIMEBOOST_net_12144), .b(g62656_sb), .o(n_6231) );
in01s01 g61703_u0 ( .a(n_8407), .o(g61703_sb) );
na02s01 TIMEBOOST_cell_16694 ( .a(n_3792), .b(g64917_sb), .o(TIMEBOOST_net_3604) );
na02f02 TIMEBOOST_cell_40421 ( .a(TIMEBOOST_net_1740), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_394), .o(TIMEBOOST_net_12449) );
na02s02 TIMEBOOST_cell_16832 ( .a(n_3774), .b(g64796_sb), .o(TIMEBOOST_net_3673) );
in01s01 g61704_u0 ( .a(FE_OFN716_n_8176), .o(g61704_sb) );
na03s02 TIMEBOOST_cell_38227 ( .a(TIMEBOOST_net_4010), .b(g64179_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__Q), .o(TIMEBOOST_net_11352) );
na02s01 TIMEBOOST_cell_36402 ( .a(TIMEBOOST_net_10439), .b(g65688_db), .o(n_2208) );
na02f02 TIMEBOOST_cell_41182 ( .a(TIMEBOOST_net_12829), .b(g57282_sb), .o(n_11473) );
in01s01 g61705_u0 ( .a(n_7102), .o(g61705_sb) );
na02s01 TIMEBOOST_cell_43043 ( .a(TIMEBOOST_net_9868), .b(FE_OFN1634_n_9531), .o(TIMEBOOST_net_13760) );
na02s01 g61705_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__Q), .b(n_7102), .o(g61705_db) );
na02s01 TIMEBOOST_cell_31420 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q), .o(TIMEBOOST_net_9621) );
in01s01 g61706_u0 ( .a(FE_OFN714_n_8140), .o(g61706_sb) );
na02f02 TIMEBOOST_cell_44663 ( .a(n_9204), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__Q), .o(TIMEBOOST_net_14570) );
no02f04 TIMEBOOST_cell_22414 ( .a(FE_RN_811_0), .b(FE_RN_812_0), .o(TIMEBOOST_net_6464) );
na02f02 TIMEBOOST_cell_38976 ( .a(TIMEBOOST_net_11726), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10720) );
in01s01 g61707_u0 ( .a(n_8272), .o(g61707_sb) );
na02s01 TIMEBOOST_cell_36322 ( .a(TIMEBOOST_net_10399), .b(g65964_db), .o(n_2159) );
na02s01 g61707_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__Q), .b(n_8272), .o(g61707_db) );
na02f02 g55413_u0 ( .a(FE_OFN1583_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__Q), .o(n_12312) );
in01s01 g61708_u0 ( .a(n_8069), .o(g61708_sb) );
na02s01 TIMEBOOST_cell_37976 ( .a(TIMEBOOST_net_11226), .b(n_4598), .o(n_6961) );
na03s02 TIMEBOOST_cell_40433 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__Q), .b(FE_OFN1120_g64577_p), .c(g63045_sb), .o(TIMEBOOST_net_12455) );
na02s02 TIMEBOOST_cell_39814 ( .a(TIMEBOOST_net_12145), .b(g62534_sb), .o(n_6504) );
in01s01 g61709_u0 ( .a(n_8407), .o(g61709_sb) );
na02s02 TIMEBOOST_cell_42109 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__Q), .b(g58448_sb), .o(TIMEBOOST_net_13293) );
no02f08 TIMEBOOST_cell_44762 ( .a(TIMEBOOST_net_14619), .b(FE_RN_820_0), .o(FE_RN_822_0) );
na02s01 TIMEBOOST_cell_16789 ( .a(TIMEBOOST_net_3651), .b(g65295_sb), .o(n_3577) );
in01s01 g61710_u0 ( .a(n_8140), .o(g61710_sb) );
na02f02 TIMEBOOST_cell_44254 ( .a(TIMEBOOST_net_14365), .b(FE_OFN1385_n_8567), .o(TIMEBOOST_net_12916) );
na02s02 TIMEBOOST_cell_40407 ( .a(n_2153), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__Q), .o(TIMEBOOST_net_12442) );
na02s02 TIMEBOOST_cell_39816 ( .a(TIMEBOOST_net_12146), .b(g62469_sb), .o(n_6654) );
in01s01 g61711_u0 ( .a(FE_OFN702_n_7845), .o(g61711_sb) );
na02s02 TIMEBOOST_cell_42360 ( .a(TIMEBOOST_net_13418), .b(g54366_sb), .o(n_13076) );
na02s01 TIMEBOOST_cell_44848 ( .a(TIMEBOOST_net_14662), .b(g64874_db), .o(n_3710) );
na02s01 TIMEBOOST_cell_18593 ( .a(TIMEBOOST_net_4553), .b(g63432_sb), .o(n_4627) );
in01s01 g61712_u0 ( .a(FE_OFN707_n_8119), .o(g61712_sb) );
na02s02 TIMEBOOST_cell_43582 ( .a(TIMEBOOST_net_14029), .b(FE_OFN1322_n_6436), .o(TIMEBOOST_net_12219) );
na02s02 TIMEBOOST_cell_43470 ( .a(TIMEBOOST_net_13973), .b(FE_OFN2063_n_6391), .o(TIMEBOOST_net_12149) );
na03s03 TIMEBOOST_cell_45427 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__Q), .b(n_13171), .c(FE_OFN1332_n_13547), .o(TIMEBOOST_net_14952) );
na02s01 TIMEBOOST_cell_40257 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__Q), .b(n_8069), .o(TIMEBOOST_net_12367) );
na02s01 g61713_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__Q), .b(n_7102), .o(g61713_db) );
in01s01 g61714_u0 ( .a(FE_OFN1812_n_7845), .o(g61714_sb) );
na02m01 TIMEBOOST_cell_37737 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_55), .b(n_14837), .o(TIMEBOOST_net_11107) );
na02s01 TIMEBOOST_cell_36534 ( .a(TIMEBOOST_net_10505), .b(g65754_db), .o(n_1921) );
na02s01 g64972_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__Q), .b(FE_OFN1807_n_4501), .o(g64972_db) );
in01s01 g61715_u0 ( .a(n_8232), .o(g61715_sb) );
na02s02 TIMEBOOST_cell_45186 ( .a(TIMEBOOST_net_14831), .b(FE_OFN365_n_4093), .o(TIMEBOOST_net_12088) );
na02s03 TIMEBOOST_cell_45761 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__Q), .b(n_13223), .o(TIMEBOOST_net_15119) );
na02s02 TIMEBOOST_cell_39818 ( .a(TIMEBOOST_net_12147), .b(g62432_sb), .o(n_6733) );
in01s01 g61716_u0 ( .a(FE_OFN720_n_8060), .o(g61716_sb) );
na02f02 TIMEBOOST_cell_39142 ( .a(TIMEBOOST_net_11809), .b(TIMEBOOST_net_3086), .o(n_12720) );
na03s01 TIMEBOOST_cell_38123 ( .a(g64147_da), .b(g64147_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__28__Q), .o(TIMEBOOST_net_11300) );
na02m02 TIMEBOOST_cell_38866 ( .a(TIMEBOOST_net_11671), .b(g58466_sb), .o(n_9383) );
in01s02 g61717_u0 ( .a(n_8232), .o(g61717_sb) );
na02s01 TIMEBOOST_cell_16754 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(g64154_sb), .o(TIMEBOOST_net_3634) );
na02s04 TIMEBOOST_cell_45762 ( .a(TIMEBOOST_net_15119), .b(FE_OFN1327_n_13547), .o(TIMEBOOST_net_14953) );
na02s01 TIMEBOOST_cell_16755 ( .a(TIMEBOOST_net_3634), .b(g64154_db), .o(n_4011) );
in01s01 g61718_u0 ( .a(FE_OFN2081_n_8176), .o(g61718_sb) );
no02f04 TIMEBOOST_cell_10132 ( .a(FE_RN_159_0), .b(FE_RN_160_0), .o(TIMEBOOST_net_1633) );
na02s01 TIMEBOOST_cell_17811 ( .a(TIMEBOOST_net_4162), .b(g61755_sb), .o(n_8304) );
na02f02 TIMEBOOST_cell_22555 ( .a(TIMEBOOST_net_6534), .b(FE_OFN1733_n_16317), .o(n_12663) );
in01s01 g61719_u0 ( .a(FE_OFN704_n_8069), .o(g61719_sb) );
na02m02 TIMEBOOST_cell_15821 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_2__Q), .b(TIMEBOOST_net_3167), .o(n_9118) );
na02s01 TIMEBOOST_cell_9234 ( .a(pci_target_unit_fifos_pcir_data_in_188), .b(g65695_sb), .o(TIMEBOOST_net_1184) );
in01s01 TIMEBOOST_cell_32850 ( .a(TIMEBOOST_net_10351), .o(TIMEBOOST_net_10330) );
in01s01 g61720_u0 ( .a(FE_OFN2084_n_8407), .o(g61720_sb) );
na02s01 TIMEBOOST_cell_18115 ( .a(TIMEBOOST_net_4314), .b(g63560_db), .o(n_4114) );
na02s01 TIMEBOOST_cell_40513 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__Q), .b(wishbone_slave_unit_pcim_sm_data_in_663), .o(TIMEBOOST_net_12495) );
na02s01 TIMEBOOST_cell_39426 ( .a(TIMEBOOST_net_11951), .b(FE_OFN237_n_9118), .o(n_9043) );
in01s01 g61721_u0 ( .a(FE_OFN717_n_8176), .o(g61721_sb) );
na02s01 TIMEBOOST_cell_18117 ( .a(TIMEBOOST_net_4315), .b(g63562_db), .o(n_4112) );
na02s01 TIMEBOOST_cell_9238 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(g65701_sb), .o(TIMEBOOST_net_1186) );
na02s01 TIMEBOOST_cell_18119 ( .a(TIMEBOOST_net_4316), .b(g63574_db), .o(n_4107) );
in01s01 g61722_u0 ( .a(FE_OFN2081_n_8176), .o(g61722_sb) );
na02m02 TIMEBOOST_cell_39411 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_409), .b(g54144_sb), .o(TIMEBOOST_net_11944) );
na02m02 TIMEBOOST_cell_44379 ( .a(n_9136), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__Q), .o(TIMEBOOST_net_14428) );
na02s03 TIMEBOOST_cell_45428 ( .a(TIMEBOOST_net_14952), .b(g53920_sb), .o(n_13524) );
in01s01 g61723_u0 ( .a(FE_OFN713_n_8140), .o(g61723_sb) );
na02s01 TIMEBOOST_cell_18121 ( .a(TIMEBOOST_net_4317), .b(FE_OFN262_n_9851), .o(n_9813) );
na02s01 TIMEBOOST_cell_9240 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(g65703_sb), .o(TIMEBOOST_net_1187) );
in01s01 g61724_u0 ( .a(FE_OFN717_n_8176), .o(g61724_sb) );
na02f02 TIMEBOOST_cell_38787 ( .a(n_9594), .b(g57331_sb), .o(TIMEBOOST_net_11632) );
na02s01 TIMEBOOST_cell_9242 ( .a(pci_target_unit_fifos_pcir_data_in_185), .b(g65706_sb), .o(TIMEBOOST_net_1188) );
na02s01 TIMEBOOST_cell_40485 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__Q), .b(wishbone_slave_unit_pcim_sm_data_in_665), .o(TIMEBOOST_net_12481) );
in01s01 g61725_u0 ( .a(FE_OFN1812_n_7845), .o(g61725_sb) );
na03s02 TIMEBOOST_cell_37779 ( .a(g65839_da), .b(g65839_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__Q), .o(TIMEBOOST_net_11128) );
na02s01 TIMEBOOST_cell_36404 ( .a(TIMEBOOST_net_10440), .b(g65776_db), .o(n_2191) );
na02s01 TIMEBOOST_cell_36406 ( .a(TIMEBOOST_net_10441), .b(g58108_sb), .o(TIMEBOOST_net_361) );
in01s01 g61726_u0 ( .a(n_8069), .o(g61726_sb) );
na02s01 TIMEBOOST_cell_42794 ( .a(TIMEBOOST_net_13635), .b(g63564_db), .o(n_4598) );
na02s01 TIMEBOOST_cell_45058 ( .a(TIMEBOOST_net_14767), .b(FE_OFN1687_n_9528), .o(TIMEBOOST_net_11190) );
na03s02 TIMEBOOST_cell_42795 ( .a(n_18), .b(FE_OFN1628_n_4438), .c(n_4470), .o(TIMEBOOST_net_13636) );
in01s01 g61727_u0 ( .a(FE_OFN2257_n_8060), .o(g61727_sb) );
na02s01 TIMEBOOST_cell_39332 ( .a(TIMEBOOST_net_11904), .b(g64229_db), .o(n_3943) );
na02s01 TIMEBOOST_cell_40539 ( .a(TIMEBOOST_net_994), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_3__Q), .o(TIMEBOOST_net_12508) );
na02s01 TIMEBOOST_cell_38232 ( .a(TIMEBOOST_net_11354), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_4576) );
in01s01 g61728_u0 ( .a(FE_OFN713_n_8140), .o(g61728_sb) );
na02s01 TIMEBOOST_cell_41738 ( .a(TIMEBOOST_net_13107), .b(g65324_db), .o(n_3559) );
na02s01 TIMEBOOST_cell_9246 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(g65687_sb), .o(TIMEBOOST_net_1190) );
na03s02 TIMEBOOST_cell_43309 ( .a(n_3573), .b(FE_OFN1202_n_4090), .c(n_15), .o(TIMEBOOST_net_13893) );
in01s01 g61729_u0 ( .a(FE_OFN713_n_8140), .o(g61729_sb) );
na02s02 TIMEBOOST_cell_38234 ( .a(TIMEBOOST_net_11355), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_4678) );
na02s01 TIMEBOOST_cell_40467 ( .a(wishbone_slave_unit_fifos_outGreyCount_2_), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q), .o(TIMEBOOST_net_12472) );
na02s01 TIMEBOOST_cell_39252 ( .a(TIMEBOOST_net_11864), .b(g58427_sb), .o(TIMEBOOST_net_432) );
in01s01 g61730_u0 ( .a(FE_OFN2256_n_8060), .o(g61730_sb) );
na02f02 TIMEBOOST_cell_41136 ( .a(TIMEBOOST_net_12806), .b(g57305_sb), .o(n_11446) );
na02s01 TIMEBOOST_cell_44956 ( .a(TIMEBOOST_net_14716), .b(g58096_db), .o(n_9080) );
na02s01 TIMEBOOST_cell_18561 ( .a(TIMEBOOST_net_4537), .b(g63182_sb), .o(n_4945) );
in01s01 g61731_u0 ( .a(FE_OFN701_n_7845), .o(g61731_sb) );
na02s02 TIMEBOOST_cell_18563 ( .a(TIMEBOOST_net_4538), .b(g63434_sb), .o(n_4930) );
na02s01 TIMEBOOST_cell_9252 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(g65677_sb), .o(TIMEBOOST_net_1193) );
na02f02 TIMEBOOST_cell_38978 ( .a(TIMEBOOST_net_11727), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10714) );
in01s01 g61732_u0 ( .a(n_8119), .o(g61732_sb) );
na02s01 TIMEBOOST_cell_9074 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__Q), .o(TIMEBOOST_net_1104) );
na02s01 g61732_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__Q), .b(n_8119), .o(g61732_db) );
in01s01 g61733_u0 ( .a(FE_OFN2212_n_8407), .o(g61733_sb) );
na02s02 TIMEBOOST_cell_39820 ( .a(TIMEBOOST_net_12148), .b(g62348_sb), .o(n_6903) );
na02s02 TIMEBOOST_cell_17825 ( .a(TIMEBOOST_net_4169), .b(g62009_sb), .o(n_7877) );
na02f02 TIMEBOOST_cell_39490 ( .a(TIMEBOOST_net_11983), .b(n_17027), .o(TIMEBOOST_net_612) );
in01s01 g61734_u0 ( .a(n_8069), .o(g61734_sb) );
na02s01 TIMEBOOST_cell_9122 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__Q), .b(g65958_sb), .o(TIMEBOOST_net_1128) );
na02s01 g61734_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__Q), .b(n_8069), .o(g61734_db) );
na02s01 TIMEBOOST_cell_9123 ( .a(TIMEBOOST_net_1128), .b(g65958_db), .o(n_2164) );
in01s01 g61735_u0 ( .a(n_8232), .o(g61735_sb) );
na02s01 TIMEBOOST_cell_44859 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q), .b(FE_OFN1650_n_9428), .o(TIMEBOOST_net_14668) );
na02s01 g61735_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__Q), .b(n_8232), .o(g61735_db) );
na02f02 TIMEBOOST_cell_43706 ( .a(TIMEBOOST_net_14091), .b(FE_OFN1349_n_8567), .o(TIMEBOOST_net_13313) );
in01s01 g61736_u0 ( .a(n_8069), .o(g61736_sb) );
na02s01 TIMEBOOST_cell_9126 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__Q), .b(g65960_sb), .o(TIMEBOOST_net_1130) );
na02s01 g61736_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__Q), .b(n_8069), .o(g61736_db) );
na02s01 TIMEBOOST_cell_9127 ( .a(TIMEBOOST_net_1130), .b(g65960_db), .o(n_2162) );
in01s01 g61737_u0 ( .a(FE_OFN719_n_8060), .o(g61737_sb) );
na02m02 TIMEBOOST_cell_38979 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_24__Q), .o(TIMEBOOST_net_11728) );
na02s02 TIMEBOOST_cell_39822 ( .a(TIMEBOOST_net_12149), .b(g62953_sb), .o(n_5975) );
na02s02 TIMEBOOST_cell_38236 ( .a(TIMEBOOST_net_11356), .b(FE_OFN1129_g64577_p), .o(TIMEBOOST_net_4562) );
in01s01 g61738_u0 ( .a(n_8272), .o(g61738_sb) );
na02m02 TIMEBOOST_cell_43965 ( .a(n_9563), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__Q), .o(TIMEBOOST_net_14221) );
na02s01 g61738_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__Q), .b(n_8272), .o(g61738_db) );
na02f02 TIMEBOOST_cell_43966 ( .a(TIMEBOOST_net_14221), .b(FE_OFN1397_n_8567), .o(TIMEBOOST_net_12983) );
in01s01 g61739_u0 ( .a(FE_OFN714_n_8140), .o(g61739_sb) );
na03s02 TIMEBOOST_cell_39413 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__Q), .b(FE_OFN702_n_7845), .c(g61900_sb), .o(TIMEBOOST_net_11945) );
na03s01 TIMEBOOST_cell_34135 ( .a(n_3972), .b(g62843_sb), .c(g62843_db), .o(n_5285) );
na02f02 TIMEBOOST_cell_42294 ( .a(TIMEBOOST_net_13385), .b(g57447_sb), .o(n_10349) );
in01s01 g61740_u0 ( .a(n_8069), .o(g61740_sb) );
na02s01 g61740_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__Q), .b(n_8069), .o(g61740_db) );
na02s01 TIMEBOOST_cell_41885 ( .a(FE_OFN237_n_9118), .b(g57936_sb), .o(TIMEBOOST_net_13181) );
in01s01 g61741_u0 ( .a(n_8232), .o(g61741_sb) );
na02s01 TIMEBOOST_cell_17220 ( .a(n_4493), .b(FE_OFN1643_n_4671), .o(TIMEBOOST_net_3867) );
na02s01 TIMEBOOST_cell_45146 ( .a(TIMEBOOST_net_14811), .b(g57903_db), .o(n_9223) );
na02s02 TIMEBOOST_cell_17221 ( .a(TIMEBOOST_net_3867), .b(g65402_da), .o(n_4236) );
in01s01 g61742_u0 ( .a(n_8119), .o(g61742_sb) );
na02s02 TIMEBOOST_cell_9134 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__Q), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_1134) );
na02s01 g61742_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__Q), .b(n_8119), .o(g61742_db) );
na02s02 TIMEBOOST_cell_43116 ( .a(TIMEBOOST_net_13796), .b(FE_OFN1197_n_4090), .o(TIMEBOOST_net_12096) );
in01s01 g61743_u0 ( .a(n_8407), .o(g61743_sb) );
na02s02 TIMEBOOST_cell_9136 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__Q), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_1135) );
na02s01 g61743_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__Q), .b(n_8407), .o(g61743_db) );
na02s02 TIMEBOOST_cell_9137 ( .a(TIMEBOOST_net_1135), .b(g57795_sb), .o(TIMEBOOST_net_925) );
in01s01 g61744_u0 ( .a(FE_OFN720_n_8060), .o(g61744_sb) );
na02f02 TIMEBOOST_cell_39144 ( .a(FE_OCPN1866_n_12377), .b(TIMEBOOST_net_11810), .o(n_12604) );
na02f02 TIMEBOOST_cell_39069 ( .a(FE_OFN1775_n_13800), .b(TIMEBOOST_net_10152), .o(TIMEBOOST_net_11773) );
na02s02 TIMEBOOST_cell_20672 ( .a(FE_OFN1186_n_3476), .b(configuration_pci_err_cs_bit10), .o(TIMEBOOST_net_5593) );
in01s01 g61745_u0 ( .a(FE_OFN716_n_8176), .o(g61745_sb) );
na02m02 TIMEBOOST_cell_38744 ( .a(TIMEBOOST_net_11610), .b(g53915_sb), .o(n_13527) );
na03s02 TIMEBOOST_cell_34137 ( .a(n_4019), .b(g62799_sb), .c(g62799_db), .o(n_5386) );
in01s01 g61746_u0 ( .a(n_8232), .o(g61746_sb) );
na02s01 TIMEBOOST_cell_44957 ( .a(FE_OFN213_n_9124), .b(g57919_sb), .o(TIMEBOOST_net_14717) );
na02s01 g61746_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__Q), .b(n_8232), .o(g61746_db) );
na02s01 TIMEBOOST_cell_39824 ( .a(TIMEBOOST_net_12150), .b(g62945_sb), .o(n_5991) );
in01s01 g61747_u0 ( .a(FE_OFN712_n_8140), .o(g61747_sb) );
na02s02 TIMEBOOST_cell_38238 ( .a(TIMEBOOST_net_11357), .b(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_4671) );
na02s01 TIMEBOOST_cell_40533 ( .a(TIMEBOOST_net_1825), .b(FE_OFN1082_n_13221), .o(TIMEBOOST_net_12505) );
na02s01 TIMEBOOST_cell_18845 ( .a(TIMEBOOST_net_4679), .b(g63070_sb), .o(n_5110) );
in01s01 g61748_u0 ( .a(n_8232), .o(g61748_sb) );
na02s01 TIMEBOOST_cell_9138 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__Q), .o(TIMEBOOST_net_1136) );
na02s01 g61748_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__Q), .b(n_8232), .o(g61748_db) );
na02s01 TIMEBOOST_cell_9139 ( .a(TIMEBOOST_net_1136), .b(n_4730), .o(TIMEBOOST_net_174) );
in01s01 g61749_u0 ( .a(n_8069), .o(g61749_sb) );
na02s01 TIMEBOOST_cell_45091 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__Q), .b(FE_OFN523_n_9428), .o(TIMEBOOST_net_14784) );
na02s01 g61749_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__Q), .b(n_8069), .o(g61749_db) );
na02s02 TIMEBOOST_cell_39826 ( .a(TIMEBOOST_net_12151), .b(g62606_sb), .o(n_6340) );
in01s01 g61750_u0 ( .a(FE_OFN717_n_8176), .o(g61750_sb) );
na02s02 TIMEBOOST_cell_38240 ( .a(TIMEBOOST_net_11358), .b(FE_OFN1129_g64577_p), .o(TIMEBOOST_net_4683) );
na02s01 TIMEBOOST_cell_9256 ( .a(pci_target_unit_fifos_pcir_data_in_178), .b(g65685_sb), .o(TIMEBOOST_net_1195) );
na02s02 TIMEBOOST_cell_38242 ( .a(TIMEBOOST_net_11359), .b(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_4542) );
in01s01 g61751_u0 ( .a(FE_OFN2081_n_8176), .o(g61751_sb) );
na02m02 TIMEBOOST_cell_43707 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__Q), .b(n_9886), .o(TIMEBOOST_net_14092) );
na02f02 TIMEBOOST_cell_41648 ( .a(FE_OFN1436_n_9372), .b(TIMEBOOST_net_13062), .o(TIMEBOOST_net_11658) );
na02s01 TIMEBOOST_cell_15797 ( .a(TIMEBOOST_net_3155), .b(g67049_sb), .o(n_1274) );
in01s01 g61752_u0 ( .a(n_8272), .o(g61752_sb) );
na02s01 TIMEBOOST_cell_18849 ( .a(TIMEBOOST_net_4681), .b(g63098_sb), .o(n_5058) );
na02s01 g61752_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__Q), .b(n_8272), .o(g61752_db) );
na02s01 TIMEBOOST_cell_18851 ( .a(TIMEBOOST_net_4682), .b(g63140_sb), .o(n_4968) );
in01s01 g61753_u0 ( .a(FE_OFN2257_n_8060), .o(g61753_sb) );
na02s01 TIMEBOOST_cell_18853 ( .a(TIMEBOOST_net_4683), .b(g63143_sb), .o(n_4961) );
na02s01 TIMEBOOST_cell_9258 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(g65686_sb), .o(TIMEBOOST_net_1196) );
na02s01 TIMEBOOST_cell_18855 ( .a(TIMEBOOST_net_4684), .b(g63170_sb), .o(n_4953) );
in01s01 g61754_u0 ( .a(FE_OFN704_n_8069), .o(g61754_sb) );
na02s01 TIMEBOOST_cell_18857 ( .a(TIMEBOOST_net_4685), .b(g63075_sb), .o(n_5100) );
na02s01 TIMEBOOST_cell_9260 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(g65689_sb), .o(TIMEBOOST_net_1197) );
na02s02 TIMEBOOST_cell_18859 ( .a(TIMEBOOST_net_4686), .b(g63121_sb), .o(n_5014) );
in01s01 g61755_u0 ( .a(FE_OFN704_n_8069), .o(g61755_sb) );
na02s01 TIMEBOOST_cell_37202 ( .a(TIMEBOOST_net_10839), .b(g58108_sb), .o(TIMEBOOST_net_9342) );
na02f02 TIMEBOOST_cell_38913 ( .a(n_3332), .b(wbu_addr_in_273), .o(TIMEBOOST_net_11695) );
na02s02 TIMEBOOST_cell_44833 ( .a(FE_OFN640_n_4669), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__Q), .o(TIMEBOOST_net_14655) );
in01s01 g61756_u0 ( .a(FE_OFN719_n_8060), .o(g61756_sb) );
na03s02 TIMEBOOST_cell_38241 ( .a(g64320_da), .b(g64320_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__Q), .o(TIMEBOOST_net_11359) );
na02s02 TIMEBOOST_cell_41774 ( .a(TIMEBOOST_net_13125), .b(g58349_db), .o(n_9472) );
na02s01 TIMEBOOST_cell_39418 ( .a(TIMEBOOST_net_11947), .b(g61896_db), .o(n_8034) );
in01s01 g61757_u0 ( .a(FE_OFN2257_n_8060), .o(g61757_sb) );
na02s02 TIMEBOOST_cell_38244 ( .a(TIMEBOOST_net_11360), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_4498) );
na02f02 TIMEBOOST_cell_39063 ( .a(TIMEBOOST_net_10145), .b(FE_OFN1770_n_14054), .o(TIMEBOOST_net_11770) );
na02s02 TIMEBOOST_cell_18865 ( .a(TIMEBOOST_net_4689), .b(g62813_sb), .o(n_5351) );
in01s01 g61758_u0 ( .a(FE_OFN2084_n_8407), .o(g61758_sb) );
na02s02 TIMEBOOST_cell_38246 ( .a(TIMEBOOST_net_11361), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_4702) );
na02f02 TIMEBOOST_cell_39065 ( .a(TIMEBOOST_net_10141), .b(FE_OFN1770_n_14054), .o(TIMEBOOST_net_11771) );
na02s02 TIMEBOOST_cell_38248 ( .a(TIMEBOOST_net_11362), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_4497) );
in01s01 g61759_u0 ( .a(FE_OFN717_n_8176), .o(g61759_sb) );
na02s01 TIMEBOOST_cell_18571 ( .a(TIMEBOOST_net_4542), .b(g63113_sb), .o(n_5029) );
na02s02 TIMEBOOST_cell_9268 ( .a(n_2284), .b(n_12179), .o(TIMEBOOST_net_1201) );
na03s02 TIMEBOOST_cell_34138 ( .a(n_4027), .b(g62780_sb), .c(g62780_db), .o(n_5431) );
in01s01 g61760_u0 ( .a(FE_OFN2084_n_8407), .o(g61760_sb) );
na02s02 TIMEBOOST_cell_38250 ( .a(TIMEBOOST_net_11363), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_4508) );
na02s01 TIMEBOOST_cell_9270 ( .a(n_2284), .b(n_657), .o(TIMEBOOST_net_1202) );
na02s02 TIMEBOOST_cell_18873 ( .a(TIMEBOOST_net_4693), .b(g62722_sb), .o(n_5539) );
in01s01 g61761_u0 ( .a(FE_OFN714_n_8140), .o(g61761_sb) );
na02f02 TIMEBOOST_cell_43708 ( .a(TIMEBOOST_net_14092), .b(FE_OFN1349_n_8567), .o(TIMEBOOST_net_13314) );
na02s01 TIMEBOOST_cell_15798 ( .a(parchk_pci_ad_reg_in_1215), .b(g67075_db), .o(TIMEBOOST_net_3156) );
na02s01 TIMEBOOST_cell_15859 ( .a(TIMEBOOST_net_3186), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_394), .o(TIMEBOOST_net_65) );
in01s01 g61762_u0 ( .a(FE_OFN719_n_8060), .o(g61762_sb) );
na02f02 TIMEBOOST_cell_39071 ( .a(FE_OFN1775_n_13800), .b(TIMEBOOST_net_10150), .o(TIMEBOOST_net_11774) );
na02f02 TIMEBOOST_cell_38980 ( .a(TIMEBOOST_net_11728), .b(FE_OFN2156_n_16439), .o(TIMEBOOST_net_10713) );
na02s02 TIMEBOOST_cell_38252 ( .a(TIMEBOOST_net_11364), .b(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_4628) );
in01s01 g61763_u0 ( .a(FE_OFN2256_n_8060), .o(g61763_sb) );
na02s02 TIMEBOOST_cell_41959 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__Q), .b(g58345_sb), .o(TIMEBOOST_net_13218) );
na02f02 TIMEBOOST_cell_39067 ( .a(FE_OFN1771_n_14054), .b(TIMEBOOST_net_10137), .o(TIMEBOOST_net_11772) );
na02s01 TIMEBOOST_cell_38254 ( .a(TIMEBOOST_net_11365), .b(FE_OFN1127_g64577_p), .o(TIMEBOOST_net_4657) );
in01s01 g61764_u0 ( .a(n_8140), .o(g61764_sb) );
na02s01 TIMEBOOST_cell_43095 ( .a(n_2181), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__Q), .o(TIMEBOOST_net_13786) );
na02s01 g61764_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__Q), .b(n_8140), .o(g61764_db) );
na02s01 TIMEBOOST_cell_17187 ( .a(TIMEBOOST_net_3850), .b(g65354_db), .o(n_3539) );
in01s01 g61765_u0 ( .a(n_8119), .o(g61765_sb) );
na02f02 TIMEBOOST_cell_40934 ( .a(TIMEBOOST_net_12705), .b(g57051_sb), .o(n_10509) );
na02s01 g61765_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__Q), .b(n_8119), .o(g61765_db) );
na02s01 TIMEBOOST_cell_39828 ( .a(TIMEBOOST_net_12152), .b(g62763_sb), .o(n_6117) );
in01s01 g61766_u0 ( .a(FE_OFN2257_n_8060), .o(g61766_sb) );
na02s01 TIMEBOOST_cell_18579 ( .a(TIMEBOOST_net_4546), .b(g63059_sb), .o(n_5132) );
na02s01 g61766_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__Q), .b(FE_OFN2257_n_8060), .o(g61766_db) );
in01s01 TIMEBOOST_cell_32840 ( .a(TIMEBOOST_net_10341), .o(wbs_dat_i_26_) );
in01s01 g61767_u0 ( .a(n_8119), .o(g61767_sb) );
na02s01 TIMEBOOST_cell_30774 ( .a(pci_target_unit_del_sync_bc_in_201), .b(n_2520), .o(TIMEBOOST_net_9298) );
na02s01 g61767_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__Q), .b(n_8119), .o(g61767_db) );
na02s01 TIMEBOOST_cell_44958 ( .a(TIMEBOOST_net_14717), .b(g57919_db), .o(n_9134) );
in01s01 g61768_u0 ( .a(n_8272), .o(g61768_sb) );
na02s01 TIMEBOOST_cell_9872 ( .a(wishbone_slave_unit_pci_initiator_if_current_byte_address), .b(FE_OFN2072_n_15978), .o(TIMEBOOST_net_1503) );
na02s01 g61768_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__Q), .b(n_8272), .o(g61768_db) );
na02s01 TIMEBOOST_cell_9873 ( .a(TIMEBOOST_net_1503), .b(g53946_sb), .o(TIMEBOOST_net_883) );
in01s01 g61769_u0 ( .a(FE_OFN714_n_8140), .o(g61769_sb) );
na02m02 TIMEBOOST_cell_10140 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__Q), .b(n_504), .o(TIMEBOOST_net_1637) );
na02m02 TIMEBOOST_cell_30784 ( .a(n_2428), .b(n_2228), .o(TIMEBOOST_net_9303) );
in01s01 g61770_u0 ( .a(FE_OFN707_n_8119), .o(g61770_sb) );
na02s02 TIMEBOOST_cell_43082 ( .a(TIMEBOOST_net_13779), .b(FE_OFN1244_n_4092), .o(TIMEBOOST_net_12135) );
na02m04 TIMEBOOST_cell_39037 ( .a(wbs_wbb3_2_wbb2_dat_o_i_113), .b(wbs_dat_o_14_), .o(TIMEBOOST_net_11757) );
na03s02 TIMEBOOST_cell_33464 ( .a(n_4442), .b(g64871_sb), .c(g64871_db), .o(n_4423) );
in01s01 g61771_u0 ( .a(n_8119), .o(g61771_sb) );
na02f02 TIMEBOOST_cell_44380 ( .a(TIMEBOOST_net_14428), .b(FE_OFN1391_n_8567), .o(TIMEBOOST_net_12723) );
na02s01 g61771_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__Q), .b(n_8119), .o(g61771_db) );
na02f02 TIMEBOOST_cell_38810 ( .a(TIMEBOOST_net_11643), .b(FE_OFN1428_n_8567), .o(n_11289) );
in01s01 g61772_u0 ( .a(n_8232), .o(g61772_sb) );
na02s02 TIMEBOOST_cell_43620 ( .a(TIMEBOOST_net_14048), .b(FE_OFN1315_n_6624), .o(TIMEBOOST_net_12249) );
na02s01 g61772_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__Q), .b(n_8232), .o(g61772_db) );
na02s01 TIMEBOOST_cell_42688 ( .a(TIMEBOOST_net_13582), .b(g57928_db), .o(n_9133) );
in01s01 g61773_u0 ( .a(FE_OFN699_n_7845), .o(g61773_sb) );
na02m02 TIMEBOOST_cell_32508 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__16__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__16__Q), .o(TIMEBOOST_net_10165) );
na02m02 TIMEBOOST_cell_43967 ( .a(n_9482), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__Q), .o(TIMEBOOST_net_14222) );
na02f02 TIMEBOOST_cell_41530 ( .a(TIMEBOOST_net_13003), .b(g57544_sb), .o(n_11200) );
in01s01 g61774_u0 ( .a(FE_OFN702_n_7845), .o(g61774_sb) );
na02s02 TIMEBOOST_cell_38256 ( .a(TIMEBOOST_net_11366), .b(FE_OFN1140_g64577_p), .o(TIMEBOOST_net_4615) );
na02s01 TIMEBOOST_cell_9278 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__Q), .b(g65425_sb), .o(TIMEBOOST_net_1206) );
na02f02 TIMEBOOST_cell_22073 ( .a(n_14027), .b(TIMEBOOST_net_6293), .o(n_16211) );
in01s01 g61775_u0 ( .a(n_8407), .o(g61775_sb) );
na02s01 TIMEBOOST_cell_42654 ( .a(TIMEBOOST_net_13565), .b(g64992_db), .o(n_3645) );
na02s01 g61775_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__Q), .b(n_8407), .o(g61775_db) );
na02s01 TIMEBOOST_cell_43368 ( .a(TIMEBOOST_net_13922), .b(n_6287), .o(TIMEBOOST_net_11581) );
na02s02 TIMEBOOST_cell_42704 ( .a(TIMEBOOST_net_13590), .b(g58005_db), .o(n_9790) );
na02s01 g61776_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__Q), .b(n_7102), .o(g61776_db) );
na02s02 TIMEBOOST_cell_43415 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__Q), .b(n_4330), .o(TIMEBOOST_net_13946) );
in01s01 g61777_u0 ( .a(n_8232), .o(g61777_sb) );
na02f02 TIMEBOOST_cell_40936 ( .a(TIMEBOOST_net_12706), .b(g57400_sb), .o(n_10368) );
na02s01 g61777_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__Q), .b(n_8232), .o(g61777_db) );
na02s01 TIMEBOOST_cell_42895 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__Q), .b(FE_OFN572_n_9502), .o(TIMEBOOST_net_13686) );
in01s01 g61778_u0 ( .a(FE_OFN719_n_8060), .o(g61778_sb) );
na02m02 TIMEBOOST_cell_38868 ( .a(TIMEBOOST_net_11672), .b(g58484_sb), .o(n_9353) );
na02s02 TIMEBOOST_cell_38258 ( .a(TIMEBOOST_net_11367), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_4631) );
na02s01 TIMEBOOST_cell_19015 ( .a(TIMEBOOST_net_4764), .b(g58331_db), .o(n_9214) );
in01s01 g61779_u0 ( .a(n_8119), .o(g61779_sb) );
na02m02 TIMEBOOST_cell_40937 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__Q), .b(n_9504), .o(TIMEBOOST_net_12707) );
na02s01 g61779_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__Q), .b(n_8119), .o(g61779_db) );
na02s01 TIMEBOOST_cell_39830 ( .a(TIMEBOOST_net_12153), .b(g62588_sb), .o(n_6374) );
in01s01 g61780_u0 ( .a(FE_OFN2084_n_8407), .o(g61780_sb) );
na02s02 TIMEBOOST_cell_38260 ( .a(TIMEBOOST_net_11368), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_4486) );
na02s01 TIMEBOOST_cell_9280 ( .a(n_1450), .b(pciu_pciif_stop_reg_in), .o(TIMEBOOST_net_1207) );
na02s02 TIMEBOOST_cell_39832 ( .a(TIMEBOOST_net_12154), .b(g62457_sb), .o(n_6682) );
in01s01 g61781_u0 ( .a(n_8272), .o(g61781_sb) );
na02s01 TIMEBOOST_cell_17572 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_2__Q), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_4043) );
na02s01 g61781_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__Q), .b(n_8272), .o(g61781_db) );
na02m01 TIMEBOOST_cell_17573 ( .a(TIMEBOOST_net_4043), .b(n_13221), .o(TIMEBOOST_net_511) );
in01s01 g61782_u0 ( .a(FE_OFN720_n_8060), .o(g61782_sb) );
na02s01 TIMEBOOST_cell_37740 ( .a(TIMEBOOST_net_11108), .b(g61824_sb), .o(n_8139) );
na02s02 TIMEBOOST_cell_43621 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__Q), .b(n_4265), .o(TIMEBOOST_net_14049) );
na02s01 TIMEBOOST_cell_37204 ( .a(TIMEBOOST_net_10840), .b(g65674_db), .o(n_2213) );
in01s01 g61783_u0 ( .a(n_8232), .o(g61783_sb) );
na02f02 TIMEBOOST_cell_40938 ( .a(TIMEBOOST_net_12707), .b(g57444_sb), .o(TIMEBOOST_net_11643) );
na02s01 g61783_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__Q), .b(n_8232), .o(g61783_db) );
na02s01 TIMEBOOST_cell_44959 ( .a(FE_OFN213_n_9124), .b(g58233_sb), .o(TIMEBOOST_net_14718) );
in01s01 g61784_u0 ( .a(FE_OFN713_n_8140), .o(g61784_sb) );
na02s01 TIMEBOOST_cell_42880 ( .a(TIMEBOOST_net_13678), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_11160) );
na02s01 TIMEBOOST_cell_9282 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(g65873_sb), .o(TIMEBOOST_net_1208) );
na04s02 TIMEBOOST_cell_34193 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__Q), .b(FE_OFN1666_n_9477), .c(FE_OFN262_n_9851), .d(g58350_sb), .o(n_9471) );
in01s01 g61785_u0 ( .a(FE_OFN709_n_8232), .o(g61785_sb) );
na02f02 TIMEBOOST_cell_39133 ( .a(TIMEBOOST_net_10169), .b(FE_OFN1606_n_13997), .o(TIMEBOOST_net_11805) );
na02s01 TIMEBOOST_cell_42689 ( .a(n_3770), .b(g65001_sb), .o(TIMEBOOST_net_13583) );
na02s04 TIMEBOOST_cell_45430 ( .a(TIMEBOOST_net_14953), .b(g53926_sb), .o(n_13519) );
in01s01 g61786_u0 ( .a(FE_OFN2081_n_8176), .o(g61786_sb) );
na02s02 TIMEBOOST_cell_45042 ( .a(TIMEBOOST_net_14759), .b(FE_OFN720_n_8060), .o(TIMEBOOST_net_11251) );
na02s02 TIMEBOOST_cell_45696 ( .a(TIMEBOOST_net_15086), .b(FE_OFN1284_n_4097), .o(TIMEBOOST_net_13249) );
na02s02 TIMEBOOST_cell_32011 ( .a(TIMEBOOST_net_9916), .b(FE_OFN1185_n_3476), .o(TIMEBOOST_net_4898) );
in01s01 g61787_u0 ( .a(FE_OFN706_n_8119), .o(g61787_sb) );
na02m02 TIMEBOOST_cell_10146 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__Q), .b(n_504), .o(TIMEBOOST_net_1640) );
na02f02 TIMEBOOST_cell_40940 ( .a(TIMEBOOST_net_12708), .b(g57483_sb), .o(n_10334) );
na02f02 TIMEBOOST_cell_41618 ( .a(FE_OFN1441_n_9372), .b(TIMEBOOST_net_13047), .o(TIMEBOOST_net_11669) );
in01s01 g61788_u0 ( .a(FE_OFN2084_n_8407), .o(g61788_sb) );
na03s03 TIMEBOOST_cell_45431 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__Q), .b(n_13228), .c(FE_OFN1332_n_13547), .o(TIMEBOOST_net_14954) );
na02f01 TIMEBOOST_cell_9284 ( .a(n_15755), .b(wbu_map_in_132), .o(TIMEBOOST_net_1209) );
na04s02 TIMEBOOST_cell_34194 ( .a(g64358_da), .b(g64358_db), .c(g63179_sb), .d(g63179_db), .o(n_7112) );
in01s01 g61789_u0 ( .a(FE_OFN707_n_8119), .o(g61789_sb) );
na02f02 TIMEBOOST_cell_42296 ( .a(TIMEBOOST_net_13386), .b(g57361_sb), .o(n_11385) );
na02m02 TIMEBOOST_cell_9286 ( .a(n_1442), .b(n_2914), .o(TIMEBOOST_net_1210) );
na04s02 TIMEBOOST_cell_34196 ( .a(g63570_da), .b(g63570_db), .c(g61965_sb), .d(g61965_db), .o(n_6946) );
in01s01 g61790_u0 ( .a(FE_OFN706_n_8119), .o(g61790_sb) );
na02s02 TIMEBOOST_cell_45059 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__Q), .b(FE_OFN1666_n_9477), .o(TIMEBOOST_net_14768) );
na02s03 TIMEBOOST_cell_45432 ( .a(TIMEBOOST_net_14954), .b(g53910_sb), .o(n_13531) );
na02m02 TIMEBOOST_cell_41619 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_9__Q), .b(n_9825), .o(TIMEBOOST_net_13048) );
in01s01 g61791_u0 ( .a(FE_OFN2257_n_8060), .o(g61791_sb) );
na02s02 TIMEBOOST_cell_43117 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__Q), .b(n_4346), .o(TIMEBOOST_net_13797) );
na02m06 TIMEBOOST_cell_9288 ( .a(n_2078), .b(n_1742), .o(TIMEBOOST_net_1211) );
na02s02 TIMEBOOST_cell_42559 ( .a(n_2705), .b(n_1480), .o(TIMEBOOST_net_13518) );
in01s01 g61792_u0 ( .a(FE_OFN717_n_8176), .o(g61792_sb) );
no02f04 TIMEBOOST_cell_22415 ( .a(TIMEBOOST_net_6464), .b(FE_RN_810_0), .o(n_14261) );
na02s01 TIMEBOOST_cell_9290 ( .a(FE_OFN197_n_2683), .b(FE_OFN992_n_2373), .o(TIMEBOOST_net_1212) );
na02s02 TIMEBOOST_cell_43118 ( .a(TIMEBOOST_net_13797), .b(FE_OFN1289_n_4098), .o(TIMEBOOST_net_12098) );
in01s01 g61793_u0 ( .a(FE_OFN2081_n_8176), .o(g61793_sb) );
na02s01 TIMEBOOST_cell_39334 ( .a(TIMEBOOST_net_11905), .b(g64243_db), .o(n_3929) );
na02s02 TIMEBOOST_cell_45663 ( .a(TIMEBOOST_net_9805), .b(FE_OFN1170_n_5592), .o(TIMEBOOST_net_15070) );
na04s02 TIMEBOOST_cell_34200 ( .a(g64261_da), .b(g64261_db), .c(g63047_sb), .d(g63047_db), .o(n_5158) );
in01s01 g61794_u0 ( .a(FE_OFN716_n_8176), .o(g61794_sb) );
na02f02 TIMEBOOST_cell_45035 ( .a(TIMEBOOST_net_9630), .b(FE_OFN1150_n_13249), .o(TIMEBOOST_net_14756) );
na02s01 TIMEBOOST_cell_42632 ( .a(TIMEBOOST_net_13554), .b(g58255_db), .o(n_9041) );
na02s01 TIMEBOOST_cell_32010 ( .a(configuration_pci_err_data_512), .b(wbm_dat_o_11_), .o(TIMEBOOST_net_9916) );
in01s01 g61795_u0 ( .a(FE_OFN710_n_8232), .o(g61795_sb) );
na02s02 TIMEBOOST_cell_37742 ( .a(TIMEBOOST_net_11109), .b(FE_OFN1670_n_9477), .o(TIMEBOOST_net_4335) );
na02s01 TIMEBOOST_cell_9294 ( .a(pci_target_unit_fifos_pcir_data_in_167), .b(g65750_sb), .o(TIMEBOOST_net_1214) );
na02s02 TIMEBOOST_cell_38262 ( .a(TIMEBOOST_net_11369), .b(n_14839), .o(g52404_db) );
in01s01 g61796_u0 ( .a(n_8176), .o(g61796_sb) );
na02s01 g61796_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__Q), .b(n_8176), .o(g61796_db) );
na02s02 TIMEBOOST_cell_39415 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_61), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_11946) );
in01s01 g61797_u0 ( .a(n_8140), .o(g61797_sb) );
na02s02 TIMEBOOST_cell_32009 ( .a(TIMEBOOST_net_9915), .b(FE_OFN1183_n_3476), .o(TIMEBOOST_net_4897) );
na02s01 g61797_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__Q), .b(n_8140), .o(g61797_db) );
na02f02 TIMEBOOST_cell_38870 ( .a(TIMEBOOST_net_11673), .b(g58462_sb), .o(n_9391) );
in01s01 g61798_u0 ( .a(n_8232), .o(g61798_sb) );
na02f02 TIMEBOOST_cell_41574 ( .a(TIMEBOOST_net_13025), .b(g57194_sb), .o(n_11559) );
na02s01 g61798_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__Q), .b(n_8232), .o(g61798_db) );
na02f02 TIMEBOOST_cell_44226 ( .a(TIMEBOOST_net_14351), .b(FE_OFN1388_n_8567), .o(TIMEBOOST_net_12766) );
in01s01 g61799_u0 ( .a(FE_OFN701_n_7845), .o(g61799_sb) );
na02s02 TIMEBOOST_cell_37544 ( .a(TIMEBOOST_net_11010), .b(FE_OFN704_n_8069), .o(TIMEBOOST_net_4162) );
na02s01 TIMEBOOST_cell_9296 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(g65755_sb), .o(TIMEBOOST_net_1215) );
na02f02 TIMEBOOST_cell_44318 ( .a(TIMEBOOST_net_14397), .b(FE_OFN1376_n_8567), .o(TIMEBOOST_net_12307) );
in01s01 g61800_u0 ( .a(FE_OFN699_n_7845), .o(g61800_sb) );
na02s01 TIMEBOOST_cell_42759 ( .a(g64176_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__Q), .o(TIMEBOOST_net_13618) );
na02s01 TIMEBOOST_cell_9298 ( .a(pci_target_unit_fifos_pcir_data_in_165), .b(g65756_sb), .o(TIMEBOOST_net_1216) );
na02f02 TIMEBOOST_cell_43000 ( .a(TIMEBOOST_net_13738), .b(n_3373), .o(TIMEBOOST_net_617) );
in01s01 g61801_u0 ( .a(n_8069), .o(g61801_sb) );
na02s02 TIMEBOOST_cell_43541 ( .a(n_4903), .b(n_323), .o(TIMEBOOST_net_14009) );
na02s02 TIMEBOOST_cell_43510 ( .a(TIMEBOOST_net_13993), .b(FE_OFN1230_n_6391), .o(TIMEBOOST_net_12626) );
na02s02 TIMEBOOST_cell_39834 ( .a(TIMEBOOST_net_12155), .b(g62919_sb), .o(n_6041) );
in01s01 g61802_u0 ( .a(FE_OFN716_n_8176), .o(g61802_sb) );
na02s01 TIMEBOOST_cell_42723 ( .a(g64225_db), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__Q), .o(TIMEBOOST_net_13600) );
na02f02 TIMEBOOST_cell_40986 ( .a(TIMEBOOST_net_12731), .b(g57077_sb), .o(n_11666) );
na02s02 TIMEBOOST_cell_43239 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__Q), .b(n_4485), .o(TIMEBOOST_net_13858) );
in01s01 g61803_u0 ( .a(FE_OFN714_n_8140), .o(g61803_sb) );
na02m02 TIMEBOOST_cell_43709 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__Q), .b(n_9713), .o(TIMEBOOST_net_14093) );
na02s04 TIMEBOOST_cell_45434 ( .a(TIMEBOOST_net_14955), .b(g53905_sb), .o(n_13536) );
na02f02 TIMEBOOST_cell_40942 ( .a(TIMEBOOST_net_12709), .b(g57363_sb), .o(n_11384) );
in01s01 g61804_u0 ( .a(n_8140), .o(g61804_sb) );
na02f04 TIMEBOOST_cell_45844 ( .a(TIMEBOOST_net_15160), .b(n_11118), .o(n_12550) );
na02s02 TIMEBOOST_cell_45187 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__Q), .b(n_4439), .o(TIMEBOOST_net_14832) );
in01s01 g61805_u0 ( .a(FE_OFN714_n_8140), .o(g61805_sb) );
na02s02 TIMEBOOST_cell_43416 ( .a(TIMEBOOST_net_13946), .b(n_6319), .o(TIMEBOOST_net_12172) );
na02s03 TIMEBOOST_cell_45436 ( .a(TIMEBOOST_net_14956), .b(g53927_sb), .o(n_13518) );
in01s01 g61806_u0 ( .a(FE_OFN714_n_8140), .o(g61806_sb) );
na02s02 TIMEBOOST_cell_43369 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__Q), .b(n_4334), .o(TIMEBOOST_net_13923) );
na02s03 TIMEBOOST_cell_45438 ( .a(TIMEBOOST_net_14957), .b(g53932_sb), .o(n_13513) );
in01s01 g61807_u0 ( .a(n_8272), .o(g61807_sb) );
in01s01 TIMEBOOST_cell_45882 ( .a(TIMEBOOST_net_15188), .o(TIMEBOOST_net_15189) );
na02s01 g61807_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__Q), .b(n_8272), .o(g61807_db) );
na02f02 TIMEBOOST_cell_41600 ( .a(FE_OFN1437_n_9372), .b(TIMEBOOST_net_13038), .o(TIMEBOOST_net_11671) );
in01s01 g61808_u0 ( .a(n_8176), .o(g61808_sb) );
na02s01 TIMEBOOST_cell_40369 ( .a(TIMEBOOST_net_990), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__Q), .o(TIMEBOOST_net_12423) );
na02s02 TIMEBOOST_cell_40792 ( .a(TIMEBOOST_net_12634), .b(g62532_sb), .o(n_6509) );
in01s01 g61809_u0 ( .a(FE_OFN2258_n_8060), .o(g61809_sb) );
na02s02 TIMEBOOST_cell_37546 ( .a(TIMEBOOST_net_11011), .b(FE_OFN712_n_8140), .o(TIMEBOOST_net_4168) );
na02s01 g61809_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__Q), .b(FE_OFN2258_n_8060), .o(g61809_db) );
na04s02 TIMEBOOST_cell_34202 ( .a(g64269_da), .b(g64269_db), .c(g63056_sb), .d(g63056_db), .o(n_5138) );
in01s01 g61810_u0 ( .a(n_8069), .o(g61810_sb) );
na02s01 TIMEBOOST_cell_39167 ( .a(TIMEBOOST_net_1079), .b(n_2299), .o(TIMEBOOST_net_11822) );
na02s01 g61810_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__Q), .b(n_8069), .o(g61810_db) );
na02f02 TIMEBOOST_cell_42386 ( .a(TIMEBOOST_net_13431), .b(g57232_sb), .o(n_11523) );
in01s01 g61811_u0 ( .a(FE_OFN716_n_8176), .o(g61811_sb) );
na02s02 TIMEBOOST_cell_42724 ( .a(TIMEBOOST_net_13600), .b(g64225_da), .o(TIMEBOOST_net_10972) );
na02f02 TIMEBOOST_cell_40944 ( .a(TIMEBOOST_net_12710), .b(g57257_sb), .o(n_11496) );
na02f02 TIMEBOOST_cell_43710 ( .a(TIMEBOOST_net_14093), .b(FE_OFN1349_n_8567), .o(TIMEBOOST_net_13415) );
in01s01 g61812_u0 ( .a(n_8176), .o(g61812_sb) );
na02s02 TIMEBOOST_cell_43417 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__Q), .b(n_4234), .o(TIMEBOOST_net_13947) );
na02s01 TIMEBOOST_cell_39553 ( .a(configuration_wb_err_addr_533), .b(n_2960), .o(TIMEBOOST_net_12015) );
na02s02 TIMEBOOST_cell_39836 ( .a(TIMEBOOST_net_12156), .b(g62973_sb), .o(n_5936) );
in01s01 g61813_u0 ( .a(FE_OFN710_n_8232), .o(g61813_sb) );
na03s02 TIMEBOOST_cell_6701 ( .a(FE_OFN268_n_9880), .b(g58068_sb), .c(g58068_db), .o(n_9724) );
na02f06 TIMEBOOST_cell_44777 ( .a(n_2000), .b(n_1535), .o(TIMEBOOST_net_14627) );
in01s01 g61814_u0 ( .a(FE_OFN709_n_8232), .o(g61814_sb) );
na02m02 TIMEBOOST_cell_10150 ( .a(n_691), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__Q), .o(TIMEBOOST_net_1642) );
no04m10 TIMEBOOST_cell_15376 ( .a(parchk_pci_ad_out_in_1168), .b(parchk_pci_ad_out_in), .c(FE_RN_797_0), .d(FE_RN_798_0), .o(n_584) );
in01s01 g61815_u0 ( .a(FE_OFN720_n_8060), .o(g61815_sb) );
na02s02 TIMEBOOST_cell_20670 ( .a(FE_OFN1186_n_3476), .b(configuration_pci_err_cs_bit9), .o(TIMEBOOST_net_5592) );
na02s02 TIMEBOOST_cell_38264 ( .a(TIMEBOOST_net_11370), .b(n_8757), .o(TIMEBOOST_net_535) );
na02s02 TIMEBOOST_cell_38266 ( .a(TIMEBOOST_net_11371), .b(FE_OFN1173_n_5592), .o(n_5623) );
in01s01 g61816_u0 ( .a(FE_OFN706_n_8119), .o(g61816_sb) );
na02s03 TIMEBOOST_cell_45440 ( .a(TIMEBOOST_net_14958), .b(g53917_sb), .o(n_13525) );
na02f02 TIMEBOOST_cell_44450 ( .a(TIMEBOOST_net_14463), .b(g57047_sb), .o(n_11687) );
na03s02 TIMEBOOST_cell_34204 ( .a(n_3827), .b(FE_OFN1138_g64577_p), .c(g63127_db), .o(n_4999) );
in01s01 g61817_u0 ( .a(FE_OFN1812_n_7845), .o(g61817_sb) );
na02s01 TIMEBOOST_cell_18863 ( .a(TIMEBOOST_net_4688), .b(g63046_sb), .o(n_5161) );
na02s01 TIMEBOOST_cell_36408 ( .a(TIMEBOOST_net_10442), .b(g65847_db), .o(n_1655) );
na02s01 TIMEBOOST_cell_36410 ( .a(TIMEBOOST_net_10443), .b(g58108_sb), .o(TIMEBOOST_net_291) );
in01s01 g61818_u0 ( .a(FE_OFN701_n_7845), .o(g61818_sb) );
na02s02 TIMEBOOST_cell_42058 ( .a(TIMEBOOST_net_13267), .b(g62567_sb), .o(n_6423) );
na02s01 TIMEBOOST_cell_40449 ( .a(conf_wb_err_addr_in_957), .b(configuration_wb_err_addr_548), .o(TIMEBOOST_net_12463) );
na02s01 TIMEBOOST_cell_42091 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q), .b(n_3787), .o(TIMEBOOST_net_13284) );
in01s01 g61819_u0 ( .a(FE_OFN2084_n_8407), .o(g61819_sb) );
na02s01 TIMEBOOST_cell_9304 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(g65790_sb), .o(TIMEBOOST_net_1219) );
na03s02 TIMEBOOST_cell_34206 ( .a(TIMEBOOST_net_861), .b(g61982_db), .c(g63609_da), .o(n_7155) );
in01s01 g61820_u0 ( .a(n_8140), .o(g61820_sb) );
na02s01 TIMEBOOST_cell_8996 ( .a(wbu_addr_in_274), .b(g58770_sb), .o(TIMEBOOST_net_1065) );
na02s02 TIMEBOOST_cell_45060 ( .a(TIMEBOOST_net_14768), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_11205) );
na02s02 TIMEBOOST_cell_39838 ( .a(TIMEBOOST_net_12157), .b(g62396_sb), .o(n_7388) );
in01s01 g61821_u0 ( .a(FE_OFN2081_n_8176), .o(g61821_sb) );
na02m02 TIMEBOOST_cell_10152 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__Q), .b(g53892_sb), .o(TIMEBOOST_net_1643) );
na02s02 TIMEBOOST_cell_43240 ( .a(TIMEBOOST_net_13858), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_12072) );
in01s01 g61822_u0 ( .a(FE_OFN2212_n_8407), .o(g61822_sb) );
na02s02 TIMEBOOST_cell_39840 ( .a(TIMEBOOST_net_12158), .b(g62992_sb), .o(n_5898) );
na03s02 TIMEBOOST_cell_37851 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__Q), .b(FE_OFN532_n_9823), .c(FE_OFN266_n_9884), .o(TIMEBOOST_net_11164) );
no02m02 TIMEBOOST_cell_19016 ( .a(FE_RN_559_0), .b(FE_OFN969_n_13784), .o(TIMEBOOST_net_4765) );
in01s01 g61823_u0 ( .a(FE_OFN712_n_8140), .o(g61823_sb) );
na03s02 TIMEBOOST_cell_34207 ( .a(TIMEBOOST_net_860), .b(g61978_db), .c(g63606_da), .o(n_7163) );
na02s01 TIMEBOOST_cell_39476 ( .a(TIMEBOOST_net_11976), .b(FE_OFN1174_n_5592), .o(n_5569) );
in01s01 g61824_u0 ( .a(FE_OFN712_n_8140), .o(g61824_sb) );
in01s01 TIMEBOOST_cell_32839 ( .a(TIMEBOOST_net_10340), .o(TIMEBOOST_net_10339) );
na02s01 TIMEBOOST_cell_40551 ( .a(TIMEBOOST_net_992), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_1__Q), .o(TIMEBOOST_net_12514) );
in01s01 TIMEBOOST_cell_32838 ( .a(TIMEBOOST_net_10339), .o(wbs_dat_i_4_) );
in01s01 g61825_u0 ( .a(FE_OFN2212_n_8407), .o(g61825_sb) );
na03s02 TIMEBOOST_cell_38243 ( .a(TIMEBOOST_net_3984), .b(g64079_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__Q), .o(TIMEBOOST_net_11360) );
na02s01 TIMEBOOST_cell_37419 ( .a(wbu_latency_tim_val_in_244), .b(n_6986), .o(TIMEBOOST_net_10948) );
na02s01 TIMEBOOST_cell_18133 ( .a(TIMEBOOST_net_4323), .b(FE_OFN262_n_9851), .o(n_9775) );
in01s01 g61826_u0 ( .a(FE_OFN2084_n_8407), .o(g61826_sb) );
na02s01 TIMEBOOST_cell_9310 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(g65805_sb), .o(TIMEBOOST_net_1222) );
na02f02 TIMEBOOST_cell_42298 ( .a(TIMEBOOST_net_13387), .b(g57083_sb), .o(n_10493) );
in01s01 g61827_u0 ( .a(FE_OFN719_n_8060), .o(g61827_sb) );
na02s01 TIMEBOOST_cell_38624 ( .a(TIMEBOOST_net_11550), .b(g62657_sb), .o(n_6230) );
na02f02 TIMEBOOST_cell_44170 ( .a(TIMEBOOST_net_14323), .b(FE_OFN1415_n_8567), .o(TIMEBOOST_net_13394) );
na02s02 TIMEBOOST_cell_17827 ( .a(TIMEBOOST_net_4170), .b(g62013_sb), .o(n_7869) );
in01s01 g61828_u0 ( .a(FE_OFN1812_n_7845), .o(g61828_sb) );
na02s02 TIMEBOOST_cell_18861 ( .a(TIMEBOOST_net_4687), .b(g63072_sb), .o(n_5106) );
na02s01 TIMEBOOST_cell_36412 ( .a(TIMEBOOST_net_10444), .b(g65718_db), .o(n_2197) );
no02f02 TIMEBOOST_cell_36414 ( .a(TIMEBOOST_net_10445), .b(FE_RN_647_0), .o(FE_RN_666_0) );
in01s01 g61829_u0 ( .a(FE_OFN720_n_8060), .o(g61829_sb) );
na02s02 TIMEBOOST_cell_38080 ( .a(TIMEBOOST_net_11278), .b(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_4558) );
na02s02 TIMEBOOST_cell_38670 ( .a(TIMEBOOST_net_11573), .b(g62379_sb), .o(n_6845) );
na02s01 TIMEBOOST_cell_38082 ( .a(TIMEBOOST_net_11279), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_4577) );
in01s01 g61830_u0 ( .a(FE_OFN701_n_7845), .o(g61830_sb) );
na02s02 TIMEBOOST_cell_37548 ( .a(TIMEBOOST_net_11012), .b(g58258_sb), .o(n_9539) );
na02s03 TIMEBOOST_cell_45442 ( .a(TIMEBOOST_net_14959), .b(g53911_sb), .o(n_13530) );
na02f02 TIMEBOOST_cell_36918 ( .a(TIMEBOOST_net_10697), .b(g52595_sb), .o(n_10278) );
na02s01 g61831_u2 ( .a(n_5641), .b(n_692), .o(g61831_db) );
na02s01 TIMEBOOST_cell_18521 ( .a(TIMEBOOST_net_4517), .b(g62825_sb), .o(n_5327) );
no02s02 g61832_u0 ( .a(wbm_adr_o_28_), .b(n_2942), .o(g61832_p) );
ao12s02 g61832_u1 ( .a(g61832_p), .b(wbm_adr_o_28_), .c(n_2942), .o(n_3472) );
no02f02 g61833_u0 ( .a(n_2947), .b(wbu_addr_in_277), .o(g61833_p) );
ao12f02 g61833_u1 ( .a(g61833_p), .b(wbu_addr_in_277), .c(n_2947), .o(n_3471) );
no02m02 g61834_u0 ( .a(n_3142), .b(n_539), .o(g61834_p) );
ao12m02 g61834_u1 ( .a(g61834_p), .b(n_539), .c(n_3142), .o(n_4196) );
in01s01 g61835_u0 ( .a(FE_OFN1118_g64577_p), .o(g61835_sb) );
na02m02 TIMEBOOST_cell_32690 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__Q), .o(TIMEBOOST_net_10256) );
na02m02 TIMEBOOST_cell_43622 ( .a(TIMEBOOST_net_14049), .b(FE_OFN1311_n_6624), .o(TIMEBOOST_net_12244) );
na02f02 TIMEBOOST_cell_32689 ( .a(FE_OFN1761_n_10780), .b(TIMEBOOST_net_10255), .o(TIMEBOOST_net_6516) );
in01s01 g61836_u0 ( .a(FE_OFN1095_g64577_p), .o(g61836_sb) );
na02s02 TIMEBOOST_cell_36850 ( .a(TIMEBOOST_net_10663), .b(g60640_sb), .o(n_5689) );
na02s01 g61836_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__Q), .b(FE_OFN1095_g64577_p), .o(g61836_db) );
na02s02 TIMEBOOST_cell_36852 ( .a(TIMEBOOST_net_10664), .b(g60658_sb), .o(n_5663) );
in01s01 g61837_u0 ( .a(FE_OFN1097_g64577_p), .o(g61837_sb) );
na02s02 TIMEBOOST_cell_36854 ( .a(TIMEBOOST_net_10665), .b(g60667_sb), .o(n_5651) );
na02s01 g61837_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__Q), .b(FE_OFN1097_g64577_p), .o(g61837_db) );
na02f08 TIMEBOOST_cell_36856 ( .a(n_15915), .b(TIMEBOOST_net_10666), .o(n_16322) );
no02m02 g61838_u0 ( .a(n_3318), .b(wbm_adr_o_31_), .o(g61838_p) );
ao12m02 g61838_u1 ( .a(g61838_p), .b(wbm_adr_o_31_), .c(n_3318), .o(n_4688) );
no02m02 g61839_u0 ( .a(FE_OFN2074_n_2723), .b(conf_wb_err_addr_in_969), .o(g61839_p) );
ao12m02 g61839_u1 ( .a(g61839_p), .b(conf_wb_err_addr_in_969), .c(FE_OFN2074_n_2723), .o(n_3344) );
in01s01 g61840_u0 ( .a(FE_OFN1094_g64577_p), .o(g61840_sb) );
na02m02 TIMEBOOST_cell_44381 ( .a(n_9753), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__Q), .o(TIMEBOOST_net_14429) );
na02s01 g61840_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__Q), .b(FE_OFN1094_g64577_p), .o(g61840_db) );
na02f02 TIMEBOOST_cell_22559 ( .a(TIMEBOOST_net_6536), .b(FE_OFN1736_n_16317), .o(n_12613) );
in01s01 g61841_u0 ( .a(FE_OFN1094_g64577_p), .o(g61841_sb) );
na02s01 g61841_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__Q), .b(FE_OFN1094_g64577_p), .o(g61841_db) );
na02s01 TIMEBOOST_cell_30939 ( .a(TIMEBOOST_net_9380), .b(g65004_sb), .o(n_3639) );
in01s01 g61842_u0 ( .a(FE_OFN1095_g64577_p), .o(g61842_sb) );
na03s02 TIMEBOOST_cell_38047 ( .a(g64274_da), .b(g64274_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__15__Q), .o(TIMEBOOST_net_11262) );
na02s01 g61842_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__Q), .b(FE_OFN1095_g64577_p), .o(g61842_db) );
na02s01 TIMEBOOST_cell_38268 ( .a(TIMEBOOST_net_11372), .b(g62140_sb), .o(n_5553) );
in01s02 g61843_u0 ( .a(n_13825), .o(g61843_sb) );
na02s01 TIMEBOOST_cell_18843 ( .a(TIMEBOOST_net_4678), .b(g63068_sb), .o(n_5114) );
na02s01 TIMEBOOST_cell_36416 ( .a(TIMEBOOST_net_10446), .b(g65998_db), .o(n_3118) );
na02s01 TIMEBOOST_cell_36418 ( .a(TIMEBOOST_net_10447), .b(g63590_sb), .o(n_2567) );
na02s02 TIMEBOOST_cell_42959 ( .a(TIMEBOOST_net_331), .b(g61743_sb), .o(TIMEBOOST_net_13718) );
na02s02 TIMEBOOST_cell_39842 ( .a(TIMEBOOST_net_12159), .b(g63009_sb), .o(n_5864) );
no02s01 g61846_u0 ( .a(conf_wb_err_addr_in_950), .b(n_2011), .o(g61846_p) );
ao12s01 g61846_u1 ( .a(g61846_p), .b(conf_wb_err_addr_in_950), .c(n_2011), .o(n_2981) );
in01s01 g61847_u0 ( .a(n_7210), .o(n_7211) );
na02s02 TIMEBOOST_cell_39844 ( .a(TIMEBOOST_net_12160), .b(g62406_sb), .o(n_6788) );
ao22f02 g61849_u0 ( .a(n_3429), .b(n_1041), .c(n_21), .d(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(n_4818) );
no02s02 g61850_u0 ( .a(wbu_addr_in_258), .b(n_2680), .o(g61850_p) );
ao12s02 g61850_u1 ( .a(g61850_p), .b(wbu_addr_in_258), .c(n_2680), .o(n_2740) );
no02m01 g61851_u0 ( .a(wbm_adr_o_9_), .b(n_2738), .o(g61851_p) );
ao12m01 g61851_u1 ( .a(g61851_p), .b(wbm_adr_o_9_), .c(n_2738), .o(n_2739) );
na02s01 TIMEBOOST_cell_40416 ( .a(TIMEBOOST_net_12446), .b(FE_OFN272_n_9828), .o(n_9625) );
oa12s02 g61853_u0 ( .a(n_7733), .b(FE_OFN2079_n_8069), .c(n_8876), .o(n_8501) );
oa22f06 g61854_u0 ( .a(n_5763), .b(n_16763), .c(wishbone_slave_unit_pci_initiator_if_write_req_int), .d(n_2354), .o(n_13547) );
in01m01 g61855_u0 ( .a(FE_OFN1699_n_5751), .o(g61855_sb) );
na02s01 TIMEBOOST_cell_32006 ( .a(configuration_pci_err_addr_478), .b(wbm_adr_o_8_), .o(TIMEBOOST_net_9914) );
na02f02 TIMEBOOST_cell_22371 ( .a(n_13993), .b(TIMEBOOST_net_6442), .o(TIMEBOOST_net_2900) );
no02f04 TIMEBOOST_cell_22416 ( .a(FE_RN_828_0), .b(FE_RN_829_0), .o(TIMEBOOST_net_6465) );
in01s01 g61856_u0 ( .a(FE_OFN1700_n_5751), .o(g61856_sb) );
na02f02 TIMEBOOST_cell_38905 ( .a(n_3140), .b(wbu_addr_in_268), .o(TIMEBOOST_net_11691) );
na02s01 TIMEBOOST_cell_43711 ( .a(g57915_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__Q), .o(TIMEBOOST_net_14094) );
na02s03 TIMEBOOST_cell_45444 ( .a(TIMEBOOST_net_14960), .b(g53909_sb), .o(n_13532) );
no02s01 g61857_u0 ( .a(n_1273), .b(pci_target_unit_wishbone_master_rty_counter_4_), .o(g61857_p) );
ao12m01 g61857_u1 ( .a(g61857_p), .b(pci_target_unit_wishbone_master_rty_counter_4_), .c(n_1273), .o(n_2289) );
in01s01 g61858_u0 ( .a(n_8140), .o(g61858_sb) );
na02f02 TIMEBOOST_cell_38989 ( .a(TIMEBOOST_net_10102), .b(FE_OFN2158_n_16439), .o(TIMEBOOST_net_11733) );
na02s01 g61858_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__Q), .b(n_8140), .o(g61858_db) );
na02f02 TIMEBOOST_cell_38982 ( .a(TIMEBOOST_net_11729), .b(FE_OFN2156_n_16439), .o(TIMEBOOST_net_10721) );
in01s01 g61859_u0 ( .a(n_8119), .o(g61859_sb) );
na02m02 TIMEBOOST_cell_38983 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_10__Q), .o(TIMEBOOST_net_11730) );
na02s01 g61859_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__Q), .b(n_8119), .o(g61859_db) );
na02s02 TIMEBOOST_cell_38270 ( .a(TIMEBOOST_net_11373), .b(FE_OFN1173_n_5592), .o(n_5620) );
in01s01 g61860_u0 ( .a(FE_OFN719_n_8060), .o(g61860_sb) );
na02s02 TIMEBOOST_cell_43586 ( .a(TIMEBOOST_net_14031), .b(FE_OFN1323_n_6436), .o(TIMEBOOST_net_12233) );
na02s02 TIMEBOOST_cell_17829 ( .a(TIMEBOOST_net_4171), .b(g62016_sb), .o(n_7863) );
na02s02 TIMEBOOST_cell_10931 ( .a(TIMEBOOST_net_2032), .b(g58438_sb), .o(n_9201) );
in01s01 g61861_u0 ( .a(FE_OFN702_n_7845), .o(g61861_sb) );
na02f04 TIMEBOOST_cell_39146 ( .a(TIMEBOOST_net_11811), .b(FE_OCPN1865_n_12377), .o(n_12610) );
na02s02 TIMEBOOST_cell_43028 ( .a(TIMEBOOST_net_13752), .b(g63137_sb), .o(n_4975) );
na02s02 TIMEBOOST_cell_18761 ( .a(TIMEBOOST_net_4637), .b(g63093_sb), .o(n_5066) );
in01s01 g61862_u0 ( .a(FE_OFN699_n_7845), .o(g61862_sb) );
na02s01 TIMEBOOST_cell_37749 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__Q), .b(wbs_dat_i_16_), .o(TIMEBOOST_net_11113) );
na02s01 TIMEBOOST_cell_40555 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_1__Q), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_1__Q), .o(TIMEBOOST_net_12516) );
na02m02 TIMEBOOST_cell_38872 ( .a(g58482_sb), .b(TIMEBOOST_net_11674), .o(n_8975) );
in01s01 g61863_u0 ( .a(n_8119), .o(g61863_sb) );
na02s02 TIMEBOOST_cell_38479 ( .a(wbm_adr_o_10_), .b(n_3005), .o(TIMEBOOST_net_11478) );
na02s01 g61863_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__Q), .b(n_8119), .o(g61863_db) );
na02s01 TIMEBOOST_cell_39367 ( .a(TIMEBOOST_net_3841), .b(FE_OFN2113_n_2053), .o(TIMEBOOST_net_11922) );
in01s01 g61864_u0 ( .a(n_8119), .o(g61864_sb) );
na02m02 TIMEBOOST_cell_10316 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_412), .b(n_13447), .o(TIMEBOOST_net_1725) );
na02s01 g61864_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__Q), .b(n_8119), .o(g61864_db) );
na02m02 TIMEBOOST_cell_38874 ( .a(TIMEBOOST_net_11675), .b(g58468_sb), .o(n_9379) );
in01s01 g61865_u0 ( .a(n_8272), .o(g61865_sb) );
na02s01 TIMEBOOST_cell_44960 ( .a(TIMEBOOST_net_14718), .b(g58233_db), .o(n_9046) );
na02s01 g61865_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__Q), .b(n_8272), .o(g61865_db) );
na02s01 TIMEBOOST_cell_38606 ( .a(TIMEBOOST_net_11541), .b(g62375_sb), .o(n_6853) );
in01s01 g61866_u0 ( .a(n_8407), .o(g61866_sb) );
na02s01 TIMEBOOST_cell_18527 ( .a(TIMEBOOST_net_4520), .b(g62839_sb), .o(n_5296) );
na02s01 g61866_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q), .b(n_8407), .o(g61866_db) );
na02f02 TIMEBOOST_cell_39148 ( .a(TIMEBOOST_net_3076), .b(TIMEBOOST_net_11812), .o(n_12637) );
in01s01 g61867_u0 ( .a(FE_OFN712_n_8140), .o(g61867_sb) );
na02s01 TIMEBOOST_cell_39311 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__Q), .b(g65894_sb), .o(TIMEBOOST_net_11894) );
na02m02 TIMEBOOST_cell_43623 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__Q), .b(n_4244), .o(TIMEBOOST_net_14050) );
na02f04 TIMEBOOST_cell_39150 ( .a(TIMEBOOST_net_11813), .b(n_16244), .o(n_16247) );
in01s01 g61868_u0 ( .a(n_8069), .o(g61868_sb) );
na02s01 TIMEBOOST_cell_38608 ( .a(TIMEBOOST_net_11542), .b(g62602_sb), .o(n_6347) );
na02s02 TIMEBOOST_cell_42081 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__Q), .b(n_3745), .o(TIMEBOOST_net_13279) );
na02s01 TIMEBOOST_cell_43712 ( .a(TIMEBOOST_net_14094), .b(TIMEBOOST_net_9744), .o(TIMEBOOST_net_10053) );
in01s01 g61869_u0 ( .a(FE_OFN714_n_8140), .o(g61869_sb) );
na02s02 TIMEBOOST_cell_10190 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__Q), .b(g61943_sb), .o(TIMEBOOST_net_1662) );
na02s02 TIMEBOOST_cell_45213 ( .a(n_3665), .b(n_3666), .o(TIMEBOOST_net_14845) );
na02s02 TIMEBOOST_cell_44422 ( .a(TIMEBOOST_net_14449), .b(FE_OFN1305_n_13124), .o(TIMEBOOST_net_13425) );
in01s01 g61870_u0 ( .a(n_8407), .o(g61870_sb) );
na02s02 TIMEBOOST_cell_18242 ( .a(n_4662), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_7_), .o(TIMEBOOST_net_4378) );
na02s01 g61870_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__Q), .b(n_8407), .o(g61870_db) );
na02s02 TIMEBOOST_cell_18243 ( .a(TIMEBOOST_net_4378), .b(g59092_sb), .o(TIMEBOOST_net_471) );
in01s01 g61871_u0 ( .a(FE_OFN713_n_8140), .o(g61871_sb) );
na02s01 TIMEBOOST_cell_37751 ( .a(g58118_db), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__Q), .o(TIMEBOOST_net_11114) );
in01s01 TIMEBOOST_cell_45867 ( .a(pci_rst_oe_o), .o(TIMEBOOST_net_15174) );
na02s02 TIMEBOOST_cell_38272 ( .a(TIMEBOOST_net_11374), .b(FE_OFN1173_n_5592), .o(n_5614) );
in01s01 g61872_u0 ( .a(FE_OFN716_n_8176), .o(g61872_sb) );
na02s01 TIMEBOOST_cell_37390 ( .a(TIMEBOOST_net_10933), .b(FE_OFN681_n_4460), .o(TIMEBOOST_net_9494) );
na02f04 TIMEBOOST_cell_22235 ( .a(TIMEBOOST_net_6374), .b(FE_OCP_RBN2224_n_16322), .o(n_16547) );
na02s02 TIMEBOOST_cell_32019 ( .a(TIMEBOOST_net_9920), .b(FE_OFN1183_n_3476), .o(TIMEBOOST_net_4902) );
in01s01 g61873_u0 ( .a(FE_OFN701_n_7845), .o(g61873_sb) );
na02m02 TIMEBOOST_cell_19153 ( .a(TIMEBOOST_net_4833), .b(g58261_sb), .o(TIMEBOOST_net_613) );
na02s01 TIMEBOOST_cell_45092 ( .a(TIMEBOOST_net_14784), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_11200) );
na02s02 TIMEBOOST_cell_19155 ( .a(TIMEBOOST_net_4834), .b(g58800_sb), .o(TIMEBOOST_net_588) );
in01s01 g61874_u0 ( .a(FE_OFN717_n_8176), .o(g61874_sb) );
na02s02 TIMEBOOST_cell_38274 ( .a(TIMEBOOST_net_11375), .b(FE_OFN1166_n_5615), .o(n_5567) );
na02m04 TIMEBOOST_cell_39039 ( .a(wbs_wbb3_2_wbb2_dat_o_i_129), .b(wbs_dat_o_30_), .o(TIMEBOOST_net_11758) );
na02s01 TIMEBOOST_cell_39336 ( .a(TIMEBOOST_net_11906), .b(g64230_db), .o(n_3942) );
in01s01 g61875_u0 ( .a(FE_OFN706_n_8119), .o(g61875_sb) );
na02s02 TIMEBOOST_cell_37550 ( .a(TIMEBOOST_net_11013), .b(g58381_sb), .o(n_9450) );
na02s01 TIMEBOOST_cell_31798 ( .a(configuration_wb_err_addr_538), .b(conf_wb_err_addr_in_947), .o(TIMEBOOST_net_9810) );
in01s01 g61876_u0 ( .a(FE_OFN709_n_8232), .o(g61876_sb) );
na02f02 TIMEBOOST_cell_39152 ( .a(TIMEBOOST_net_11814), .b(FE_OFN1566_n_12502), .o(n_12753) );
na02m04 TIMEBOOST_cell_39047 ( .a(wbs_wbb3_2_wbb2_dat_o_i_100), .b(wbs_dat_o_1_), .o(TIMEBOOST_net_11762) );
na02s02 TIMEBOOST_cell_38276 ( .a(TIMEBOOST_net_11376), .b(FE_OFN1166_n_5615), .o(n_5558) );
in01s01 g61877_u0 ( .a(n_8272), .o(g61877_sb) );
na02s01 TIMEBOOST_cell_10336 ( .a(n_3503), .b(n_2308), .o(TIMEBOOST_net_1735) );
na02s01 g61877_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__Q), .b(n_8272), .o(g61877_db) );
na02s01 TIMEBOOST_cell_10337 ( .a(TIMEBOOST_net_1735), .b(n_4743), .o(TIMEBOOST_net_461) );
in01s01 g61878_u0 ( .a(FE_OFN1812_n_7845), .o(g61878_sb) );
na02s02 TIMEBOOST_cell_18833 ( .a(TIMEBOOST_net_4673), .b(g63012_sb), .o(n_5225) );
na02s01 TIMEBOOST_cell_36420 ( .a(TIMEBOOST_net_10448), .b(g65994_sb), .o(n_2372) );
na02s01 TIMEBOOST_cell_36422 ( .a(TIMEBOOST_net_10449), .b(g65994_sb), .o(n_2568) );
in01s01 g61879_u0 ( .a(n_8069), .o(g61879_sb) );
na02s01 TIMEBOOST_cell_44961 ( .a(FE_OFN233_n_9876), .b(g57913_sb), .o(TIMEBOOST_net_14719) );
na02s01 g61879_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__Q), .b(n_8069), .o(g61879_db) );
na02s01 TIMEBOOST_cell_38610 ( .a(TIMEBOOST_net_11543), .b(g63108_sb), .o(n_5854) );
in01s01 g61880_u0 ( .a(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61880_sb) );
na02f02 TIMEBOOST_cell_41138 ( .a(TIMEBOOST_net_12807), .b(g57048_sb), .o(n_10511) );
na02s01 g61880_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61880_db) );
na02m02 TIMEBOOST_cell_32534 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__28__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__28__Q), .o(TIMEBOOST_net_10178) );
in01s01 g61881_u0 ( .a(FE_OFN706_n_8119), .o(g61881_sb) );
na02m02 TIMEBOOST_cell_43805 ( .a(n_9873), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__Q), .o(TIMEBOOST_net_14141) );
na02s02 TIMEBOOST_cell_37552 ( .a(TIMEBOOST_net_11014), .b(g58105_sb), .o(n_9691) );
na02s01 TIMEBOOST_cell_31796 ( .a(configuration_wb_err_data_574), .b(parchk_pci_ad_out_in_1171), .o(TIMEBOOST_net_9809) );
in01s01 g61882_u0 ( .a(FE_OFN707_n_8119), .o(g61882_sb) );
na02f02 TIMEBOOST_cell_22333 ( .a(TIMEBOOST_net_6423), .b(n_10163), .o(n_12159) );
na02m04 TIMEBOOST_cell_39049 ( .a(wbs_wbb3_2_wbb2_dat_o_i_128), .b(wbs_dat_o_29_), .o(TIMEBOOST_net_11763) );
na02m02 TIMEBOOST_cell_43713 ( .a(n_1039), .b(wishbone_slave_unit_fifos_inGreyCount_reg_1__Q), .o(TIMEBOOST_net_14095) );
in01s01 g61883_u0 ( .a(FE_OFN710_n_8232), .o(g61883_sb) );
na02f02 TIMEBOOST_cell_22335 ( .a(TIMEBOOST_net_6424), .b(n_12228), .o(n_15441) );
na02f02 TIMEBOOST_cell_44628 ( .a(TIMEBOOST_net_14552), .b(FE_OFN2187_n_8567), .o(TIMEBOOST_net_13007) );
na03f02 TIMEBOOST_cell_22336 ( .a(n_10010), .b(n_10014), .c(n_10599), .o(TIMEBOOST_net_6425) );
in01s01 g61884_u0 ( .a(FE_OFN2256_n_8060), .o(g61884_sb) );
na02s02 TIMEBOOST_cell_43575 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__31__Q), .b(n_4222), .o(TIMEBOOST_net_14026) );
na02m02 TIMEBOOST_cell_44201 ( .a(n_9508), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__Q), .o(TIMEBOOST_net_14339) );
na02s01 TIMEBOOST_cell_42633 ( .a(FE_OFN250_n_9789), .b(g58195_sb), .o(TIMEBOOST_net_13555) );
in01s01 g61885_u0 ( .a(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61885_sb) );
na02m02 TIMEBOOST_cell_38794 ( .a(TIMEBOOST_net_11635), .b(g54360_sb), .o(n_13082) );
na02s01 g61885_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61885_db) );
na02s02 TIMEBOOST_cell_43370 ( .a(TIMEBOOST_net_13923), .b(n_6645), .o(TIMEBOOST_net_12173) );
in01s01 g61886_u0 ( .a(FE_OFN710_n_8232), .o(g61886_sb) );
na02s02 TIMEBOOST_cell_38278 ( .a(TIMEBOOST_net_11377), .b(FE_OFN1173_n_5592), .o(n_5627) );
na02f02 TIMEBOOST_cell_39057 ( .a(FE_OFN1771_n_14054), .b(TIMEBOOST_net_10146), .o(TIMEBOOST_net_11767) );
na02s02 TIMEBOOST_cell_18779 ( .a(TIMEBOOST_net_4646), .b(g62782_sb), .o(n_5427) );
in01s01 g61887_u0 ( .a(n_8407), .o(g61887_sb) );
na02f02 TIMEBOOST_cell_44244 ( .a(TIMEBOOST_net_14360), .b(FE_OFN1394_n_8567), .o(TIMEBOOST_net_13376) );
na02s01 g61887_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__Q), .b(n_8407), .o(g61887_db) );
na02s01 TIMEBOOST_cell_18637 ( .a(TIMEBOOST_net_4575), .b(g63064_sb), .o(n_5122) );
in01s01 g61888_u0 ( .a(FE_OFN712_n_8140), .o(g61888_sb) );
na02m02 TIMEBOOST_cell_36740 ( .a(TIMEBOOST_net_463), .b(TIMEBOOST_net_10608), .o(TIMEBOOST_net_2412) );
na02f02 TIMEBOOST_cell_39059 ( .a(TIMEBOOST_net_10147), .b(FE_OFN1770_n_14054), .o(TIMEBOOST_net_11768) );
na02s02 TIMEBOOST_cell_36742 ( .a(TIMEBOOST_net_10609), .b(g63095_db), .o(n_5064) );
in01s01 g61889_u0 ( .a(n_8176), .o(g61889_sb) );
na02s02 TIMEBOOST_cell_18831 ( .a(TIMEBOOST_net_4672), .b(g63010_sb), .o(n_5227) );
na02s01 g61889_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__Q), .b(n_8176), .o(g61889_db) );
na02s01 TIMEBOOST_cell_39338 ( .a(TIMEBOOST_net_11907), .b(g64234_db), .o(n_3938) );
in01s01 g61890_u0 ( .a(FE_OFN699_n_7845), .o(g61890_sb) );
na02f02 TIMEBOOST_cell_36972 ( .a(TIMEBOOST_net_10724), .b(g58803_sb), .o(n_8638) );
na02m02 TIMEBOOST_cell_38947 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_20__Q), .o(TIMEBOOST_net_11712) );
na02m02 TIMEBOOST_cell_36744 ( .a(TIMEBOOST_net_337), .b(TIMEBOOST_net_10610), .o(TIMEBOOST_net_4867) );
in01s01 g61891_u0 ( .a(n_8119), .o(g61891_sb) );
na02s01 g61891_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__Q), .b(n_8119), .o(g61891_db) );
na02s01 TIMEBOOST_cell_18795 ( .a(TIMEBOOST_net_4654), .b(g63191_sb), .o(n_4941) );
in01s01 g61892_u0 ( .a(FE_OFN710_n_8232), .o(g61892_sb) );
na02s02 TIMEBOOST_cell_36746 ( .a(TIMEBOOST_net_10611), .b(TIMEBOOST_net_581), .o(n_5644) );
na02s01 TIMEBOOST_cell_9336 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(g64122_sb), .o(TIMEBOOST_net_1235) );
na02f02 TIMEBOOST_cell_42244 ( .a(TIMEBOOST_net_13360), .b(FE_OFN1394_n_8567), .o(TIMEBOOST_net_12312) );
in01s01 g61893_u0 ( .a(n_8272), .o(g61893_sb) );
na03s02 TIMEBOOST_cell_38351 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__15__Q), .b(FE_OFN1134_g64577_p), .c(n_3939), .o(TIMEBOOST_net_11414) );
na02s01 g61893_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__Q), .b(n_8272), .o(g61893_db) );
na02f02 TIMEBOOST_cell_38984 ( .a(TIMEBOOST_net_11730), .b(FE_OFN2153_n_16439), .o(TIMEBOOST_net_10726) );
in01s01 g61894_u0 ( .a(n_8407), .o(g61894_sb) );
na02f06 TIMEBOOST_cell_44778 ( .a(TIMEBOOST_net_14627), .b(n_2298), .o(n_3304) );
na02s01 g61894_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__Q), .b(n_8407), .o(g61894_db) );
na02f02 TIMEBOOST_cell_38986 ( .a(TIMEBOOST_net_11731), .b(g52606_db), .o(n_11865) );
in01s01 g61895_u0 ( .a(n_8119), .o(g61895_sb) );
na02s02 TIMEBOOST_cell_18677 ( .a(TIMEBOOST_net_4595), .b(g63550_sb), .o(n_4607) );
na02s01 g61895_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__Q), .b(n_8119), .o(g61895_db) );
na02s02 TIMEBOOST_cell_39360 ( .a(TIMEBOOST_net_11918), .b(g61751_sb), .o(n_8313) );
na02s02 TIMEBOOST_cell_38280 ( .a(TIMEBOOST_net_11378), .b(FE_OFN1173_n_5592), .o(n_5619) );
na02s01 g61896_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__Q), .b(n_8119), .o(g61896_db) );
na02s01 TIMEBOOST_cell_38282 ( .a(TIMEBOOST_net_11379), .b(g62115_sb), .o(n_5581) );
in01s01 g61897_u0 ( .a(n_8176), .o(g61897_sb) );
na02s02 TIMEBOOST_cell_38284 ( .a(TIMEBOOST_net_11380), .b(FE_OFN1166_n_5615), .o(n_5579) );
na02s01 g61897_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__Q), .b(n_8176), .o(g61897_db) );
na02s01 TIMEBOOST_cell_18803 ( .a(TIMEBOOST_net_4658), .b(g63111_sb), .o(n_5033) );
na02s01 TIMEBOOST_cell_18689 ( .a(TIMEBOOST_net_4601), .b(g62819_sb), .o(n_5337) );
na02s01 g61898_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__Q), .b(n_8407), .o(g61898_db) );
na02s02 TIMEBOOST_cell_18805 ( .a(TIMEBOOST_net_4659), .b(g63061_sb), .o(n_5128) );
in01s01 g61899_u0 ( .a(n_8407), .o(g61899_sb) );
na02f02 TIMEBOOST_cell_38988 ( .a(TIMEBOOST_net_11732), .b(g58819_sb), .o(n_8622) );
na02s01 g61899_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__Q), .b(n_8407), .o(g61899_db) );
na02s01 TIMEBOOST_cell_18807 ( .a(TIMEBOOST_net_4660), .b(g63019_sb), .o(n_5210) );
in01s01 g61900_u0 ( .a(FE_OFN702_n_7845), .o(g61900_sb) );
na02f02 TIMEBOOST_cell_36952 ( .a(TIMEBOOST_net_10714), .b(g58815_sb), .o(n_8626) );
na02s02 TIMEBOOST_cell_40537 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__Q), .b(g58364_sb), .o(TIMEBOOST_net_12507) );
na02m02 TIMEBOOST_cell_20345 ( .a(TIMEBOOST_net_5429), .b(n_5745), .o(n_7723) );
in01s01 g61901_u0 ( .a(FE_OFN2256_n_8060), .o(g61901_sb) );
na02s01 TIMEBOOST_cell_39350 ( .a(TIMEBOOST_net_11913), .b(g64308_db), .o(n_3867) );
na03s02 TIMEBOOST_cell_39329 ( .a(TIMEBOOST_net_3760), .b(g65727_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__Q), .o(TIMEBOOST_net_11903) );
na02s02 TIMEBOOST_cell_20349 ( .a(TIMEBOOST_net_5431), .b(g59796_db), .o(n_7621) );
in01s01 g61902_u0 ( .a(FE_OFN1812_n_7845), .o(g61902_sb) );
na03s02 TIMEBOOST_cell_37781 ( .a(g65842_da), .b(g65842_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__Q), .o(TIMEBOOST_net_11129) );
na02s01 TIMEBOOST_cell_36424 ( .a(TIMEBOOST_net_10450), .b(g65096_sb), .o(TIMEBOOST_net_218) );
na02s01 TIMEBOOST_cell_36426 ( .a(TIMEBOOST_net_10451), .b(n_3780), .o(n_3697) );
in01s01 g61903_u0 ( .a(n_8272), .o(g61903_sb) );
na02s01 TIMEBOOST_cell_18617 ( .a(TIMEBOOST_net_4565), .b(g62765_sb), .o(n_5465) );
na02s01 g61903_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__Q), .b(n_8272), .o(g61903_db) );
na02f02 TIMEBOOST_cell_44731 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__Q), .b(FE_OFN1749_n_12004), .o(TIMEBOOST_net_14604) );
in01s01 g61904_u0 ( .a(n_8232), .o(g61904_sb) );
na02s02 TIMEBOOST_cell_38286 ( .a(TIMEBOOST_net_11381), .b(g62020_sb), .o(n_7855) );
na02s01 g61904_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__Q), .b(n_8232), .o(g61904_db) );
na02s01 TIMEBOOST_cell_18809 ( .a(TIMEBOOST_net_4661), .b(g62779_sb), .o(n_5433) );
in01s01 g61905_u0 ( .a(FE_OFN706_n_8119), .o(g61905_sb) );
na02s01 TIMEBOOST_cell_18621 ( .a(TIMEBOOST_net_4567), .b(g62778_sb), .o(n_5435) );
na02s02 TIMEBOOST_cell_37554 ( .a(TIMEBOOST_net_11015), .b(g58380_sb), .o(n_9008) );
na02s01 TIMEBOOST_cell_31794 ( .a(configuration_wb_err_data_581), .b(parchk_pci_ad_out_in_1178), .o(TIMEBOOST_net_9808) );
in01s01 g61906_u0 ( .a(FE_OFN707_n_8119), .o(g61906_sb) );
na03s02 TIMEBOOST_cell_36801 ( .a(g64239_da), .b(g64239_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__Q), .o(TIMEBOOST_net_10639) );
na02m02 TIMEBOOST_cell_45795 ( .a(n_9515), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__Q), .o(TIMEBOOST_net_15136) );
na03s02 TIMEBOOST_cell_36763 ( .a(TIMEBOOST_net_4263), .b(g64112_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__16__Q), .o(TIMEBOOST_net_10620) );
in01s01 g61907_u0 ( .a(FE_OFN2212_n_8407), .o(g61907_sb) );
na02s02 TIMEBOOST_cell_38084 ( .a(TIMEBOOST_net_11280), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_4506) );
na02s01 g61907_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__Q), .b(FE_OFN2212_n_8407), .o(g61907_db) );
na02s02 TIMEBOOST_cell_38086 ( .a(TIMEBOOST_net_11281), .b(FE_OFN1126_g64577_p), .o(TIMEBOOST_net_4538) );
in01s01 g61908_u0 ( .a(FE_OFN709_n_8232), .o(g61908_sb) );
na02s01 TIMEBOOST_cell_18625 ( .a(TIMEBOOST_net_4569), .b(g62775_sb), .o(n_5444) );
na02s02 TIMEBOOST_cell_37556 ( .a(TIMEBOOST_net_11016), .b(g58231_sb), .o(n_9559) );
na02s02 TIMEBOOST_cell_42560 ( .a(TIMEBOOST_net_13518), .b(n_1379), .o(TIMEBOOST_net_196) );
in01s01 g61909_u0 ( .a(n_8272), .o(g61909_sb) );
na02s02 TIMEBOOST_cell_38288 ( .a(TIMEBOOST_net_11382), .b(g61878_sb), .o(n_8073) );
na02s01 g61909_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__Q), .b(n_8272), .o(g61909_db) );
na02f02 TIMEBOOST_cell_39154 ( .a(TIMEBOOST_net_3110), .b(TIMEBOOST_net_11815), .o(n_12600) );
in01s01 g61910_u0 ( .a(FE_OFN2081_n_8176), .o(g61910_sb) );
na02s01 TIMEBOOST_cell_10580 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__Q), .b(g65400_sb), .o(TIMEBOOST_net_1857) );
na02s01 TIMEBOOST_cell_31792 ( .a(parchk_pci_ad_out_in_1176), .b(configuration_wb_err_data_579), .o(TIMEBOOST_net_9807) );
na02s02 TIMEBOOST_cell_41960 ( .a(TIMEBOOST_net_13218), .b(g58345_db), .o(n_9475) );
in01s01 g61911_u0 ( .a(FE_OFN701_n_7845), .o(g61911_sb) );
na02s02 TIMEBOOST_cell_20355 ( .a(TIMEBOOST_net_5434), .b(FE_OFN1312_n_6624), .o(TIMEBOOST_net_2477) );
na02f02 TIMEBOOST_cell_45796 ( .a(TIMEBOOST_net_15136), .b(FE_OFN1383_n_8567), .o(TIMEBOOST_net_14578) );
no02f04 TIMEBOOST_cell_20063 ( .a(FE_RN_211_0), .b(TIMEBOOST_net_5288), .o(TIMEBOOST_net_2899) );
in01s01 g61912_u0 ( .a(FE_OFN2257_n_8060), .o(g61912_sb) );
na02m02 TIMEBOOST_cell_20367 ( .a(TIMEBOOST_net_5440), .b(FE_OFN1312_n_6624), .o(TIMEBOOST_net_2446) );
na02s01 g61912_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__Q), .b(FE_OFN2257_n_8060), .o(g61912_db) );
no02f02 TIMEBOOST_cell_22364 ( .a(TIMEBOOST_net_2300), .b(FE_RN_362_0), .o(TIMEBOOST_net_6439) );
in01s01 g61913_u0 ( .a(FE_OFN709_n_8232), .o(g61913_sb) );
na02s01 TIMEBOOST_cell_39203 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__Q), .b(n_8119), .o(TIMEBOOST_net_11840) );
na02s01 TIMEBOOST_cell_45664 ( .a(TIMEBOOST_net_15070), .b(g62120_sb), .o(n_5576) );
in01s01 TIMEBOOST_cell_45926 ( .a(TIMEBOOST_net_15232), .o(TIMEBOOST_net_15233) );
in01s01 g61914_u0 ( .a(FE_OFN709_n_8232), .o(g61914_sb) );
na02f02 TIMEBOOST_cell_38990 ( .a(TIMEBOOST_net_11733), .b(g58811_sb), .o(n_8630) );
na02f02 TIMEBOOST_cell_41542 ( .a(TIMEBOOST_net_13009), .b(g57581_sb), .o(n_11169) );
na02f02 TIMEBOOST_cell_42300 ( .a(TIMEBOOST_net_13388), .b(g57411_sb), .o(n_10365) );
in01s01 g61915_u0 ( .a(FE_OFN704_n_8069), .o(g61915_sb) );
na02m02 TIMEBOOST_cell_42245 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__Q), .b(n_9579), .o(TIMEBOOST_net_13361) );
na02f02 TIMEBOOST_cell_38992 ( .a(TIMEBOOST_net_11734), .b(g58809_sb), .o(n_8632) );
na03s02 TIMEBOOST_cell_36771 ( .a(TIMEBOOST_net_4273), .b(g64080_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__12__Q), .o(TIMEBOOST_net_10624) );
in01s01 g61916_u0 ( .a(FE_OFN704_n_8069), .o(g61916_sb) );
na02s02 TIMEBOOST_cell_20363 ( .a(TIMEBOOST_net_5438), .b(FE_OFN1312_n_6624), .o(TIMEBOOST_net_2431) );
na02s01 TIMEBOOST_cell_9348 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__Q), .b(n_4677), .o(TIMEBOOST_net_1241) );
na03s02 TIMEBOOST_cell_36749 ( .a(g65681_da), .b(g65681_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__Q), .o(TIMEBOOST_net_10613) );
in01s01 g61917_u0 ( .a(FE_OFN1812_n_7845), .o(g61917_sb) );
na03s02 TIMEBOOST_cell_37783 ( .a(g65825_da), .b(g65825_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__Q), .o(TIMEBOOST_net_11130) );
na02f06 TIMEBOOST_cell_36428 ( .a(TIMEBOOST_net_10452), .b(FE_OFN1026_n_16760), .o(FE_RN_838_0) );
na02s02 TIMEBOOST_cell_36430 ( .a(TIMEBOOST_net_10453), .b(n_1169), .o(n_2233) );
in01s01 g61918_u0 ( .a(n_8407), .o(g61918_sb) );
na02s02 TIMEBOOST_cell_18823 ( .a(TIMEBOOST_net_4668), .b(g59373_sb), .o(n_7687) );
na02s01 g61918_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__Q), .b(n_8407), .o(g61918_db) );
na02s01 TIMEBOOST_cell_18811 ( .a(TIMEBOOST_net_4662), .b(g63114_sb), .o(n_5027) );
in01s01 g61919_u0 ( .a(FE_OFN714_n_8140), .o(g61919_sb) );
na03s02 TIMEBOOST_cell_10586 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__Q), .b(FE_OFN1112_g64577_p), .c(n_3909), .o(TIMEBOOST_net_1860) );
na02s02 TIMEBOOST_cell_45665 ( .a(TIMEBOOST_net_862), .b(g61981_db), .o(TIMEBOOST_net_15071) );
na02s02 TIMEBOOST_cell_45754 ( .a(TIMEBOOST_net_15115), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_13244) );
na02s01 TIMEBOOST_cell_42796 ( .a(TIMEBOOST_net_13636), .b(g64850_sb), .o(n_4434) );
na02s02 TIMEBOOST_cell_16798 ( .a(n_3774), .b(g65056_sb), .o(TIMEBOOST_net_3656) );
in01s01 g61921_u0 ( .a(FE_OFN716_n_8176), .o(g61921_sb) );
na02s01 TIMEBOOST_cell_39428 ( .a(TIMEBOOST_net_11952), .b(g61997_sb), .o(n_7901) );
na02s01 TIMEBOOST_cell_18114 ( .a(g63560_sb), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_), .o(TIMEBOOST_net_4314) );
na02s01 TIMEBOOST_cell_37785 ( .a(g64226_da), .b(g64226_db), .o(TIMEBOOST_net_11131) );
na02s02 TIMEBOOST_cell_16801 ( .a(TIMEBOOST_net_3657), .b(g65393_db), .o(n_3523) );
na02s01 g61922_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__Q), .b(n_8232), .o(g61922_db) );
na02s01 TIMEBOOST_cell_41868 ( .a(TIMEBOOST_net_13172), .b(g61894_db), .o(n_8039) );
in01s01 g61923_u0 ( .a(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61923_sb) );
na02m02 TIMEBOOST_cell_42189 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__Q), .b(n_9861), .o(TIMEBOOST_net_13333) );
na02s01 g61923_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61923_db) );
na02f02 TIMEBOOST_cell_43968 ( .a(TIMEBOOST_net_14222), .b(FE_OFN1400_n_8567), .o(TIMEBOOST_net_12821) );
in01s01 g61924_u0 ( .a(n_8069), .o(g61924_sb) );
na02s01 TIMEBOOST_cell_41869 ( .a(conf_wb_err_addr_in_963), .b(configuration_wb_err_addr_554), .o(TIMEBOOST_net_13173) );
na02s01 TIMEBOOST_cell_41870 ( .a(TIMEBOOST_net_13173), .b(FE_OFN1170_n_5592), .o(TIMEBOOST_net_12456) );
in01s01 g61925_u0 ( .a(n_8119), .o(g61925_sb) );
na02s01 TIMEBOOST_cell_41871 ( .a(TIMEBOOST_net_978), .b(configuration_wb_err_addr_549), .o(TIMEBOOST_net_13174) );
na02s01 TIMEBOOST_cell_44962 ( .a(TIMEBOOST_net_14719), .b(g57913_db), .o(n_9897) );
na02s01 TIMEBOOST_cell_41872 ( .a(TIMEBOOST_net_13174), .b(FE_OFN1170_n_5592), .o(TIMEBOOST_net_12467) );
in01s01 g61926_u0 ( .a(FE_OFN707_n_8119), .o(g61926_sb) );
na02s01 TIMEBOOST_cell_37482 ( .a(TIMEBOOST_net_10979), .b(g58299_sb), .o(n_9509) );
na02s01 TIMEBOOST_cell_9350 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(g64122_sb), .o(TIMEBOOST_net_1242) );
na02s01 TIMEBOOST_cell_37484 ( .a(TIMEBOOST_net_10980), .b(g65887_db), .o(n_1862) );
in01s01 g61927_u0 ( .a(FE_OFN2256_n_8060), .o(g61927_sb) );
na02s02 TIMEBOOST_cell_37486 ( .a(TIMEBOOST_net_10981), .b(g65357_sb), .o(n_4256) );
na02s01 TIMEBOOST_cell_17200 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__Q), .b(g65348_sb), .o(TIMEBOOST_net_3857) );
na02s01 TIMEBOOST_cell_37488 ( .a(TIMEBOOST_net_10982), .b(FE_OFN1807_n_4501), .o(TIMEBOOST_net_9641) );
na02s01 TIMEBOOST_cell_41873 ( .a(TIMEBOOST_net_980), .b(configuration_wb_err_addr_537), .o(TIMEBOOST_net_13175) );
na02s01 TIMEBOOST_cell_44963 ( .a(FE_OFN221_n_9846), .b(g57926_sb), .o(TIMEBOOST_net_14720) );
na02s01 TIMEBOOST_cell_41874 ( .a(TIMEBOOST_net_13175), .b(FE_OFN1170_n_5592), .o(TIMEBOOST_net_12465) );
in01s01 g61929_u0 ( .a(n_8272), .o(g61929_sb) );
na02s01 TIMEBOOST_cell_41875 ( .a(conf_wb_err_addr_in_965), .b(configuration_wb_err_addr_556), .o(TIMEBOOST_net_13176) );
na02s01 g61929_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__Q), .b(n_8272), .o(g61929_db) );
na02s02 TIMEBOOST_cell_41876 ( .a(TIMEBOOST_net_13176), .b(FE_OFN1170_n_5592), .o(TIMEBOOST_net_12464) );
in01s01 g61930_u0 ( .a(n_8272), .o(g61930_sb) );
na02s01 TIMEBOOST_cell_41877 ( .a(conf_wb_err_addr_in_966), .b(configuration_wb_err_addr_557), .o(TIMEBOOST_net_13177) );
na02s02 TIMEBOOST_cell_42110 ( .a(TIMEBOOST_net_13293), .b(g58448_db), .o(n_9197) );
na02s01 TIMEBOOST_cell_39466 ( .a(TIMEBOOST_net_11971), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_4673) );
in01s01 g61931_u0 ( .a(n_8140), .o(g61931_sb) );
na02s02 TIMEBOOST_cell_41878 ( .a(TIMEBOOST_net_13177), .b(FE_OFN1170_n_5592), .o(TIMEBOOST_net_12468) );
na02s01 TIMEBOOST_cell_40371 ( .a(TIMEBOOST_net_988), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__Q), .o(TIMEBOOST_net_12424) );
na02s02 TIMEBOOST_cell_41879 ( .a(TIMEBOOST_net_4368), .b(g54182_sb), .o(TIMEBOOST_net_13178) );
in01s01 g61932_u0 ( .a(n_8176), .o(g61932_sb) );
na02s02 TIMEBOOST_cell_41880 ( .a(TIMEBOOST_net_13178), .b(g54182_db), .o(n_13431) );
na02s01 TIMEBOOST_cell_41881 ( .a(g62734_sb), .b(g62734_db), .o(TIMEBOOST_net_13179) );
in01s01 g61933_u0 ( .a(n_8232), .o(g61933_sb) );
na02s01 TIMEBOOST_cell_41882 ( .a(TIMEBOOST_net_13179), .b(n_4044), .o(n_5511) );
na02s02 TIMEBOOST_cell_45188 ( .a(TIMEBOOST_net_14832), .b(FE_OFN1268_n_4095), .o(TIMEBOOST_net_12091) );
na02s01 TIMEBOOST_cell_16809 ( .a(TIMEBOOST_net_3661), .b(g64990_db), .o(n_3646) );
in01s01 g61934_u0 ( .a(n_8119), .o(g61934_sb) );
na02s01 TIMEBOOST_cell_44964 ( .a(TIMEBOOST_net_14720), .b(g57926_db), .o(n_9883) );
na02s03 TIMEBOOST_cell_45446 ( .a(TIMEBOOST_net_14961), .b(g53918_sb), .o(n_13469) );
na02s02 TIMEBOOST_cell_16882 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__Q), .b(g64304_sb), .o(TIMEBOOST_net_3698) );
na02s02 TIMEBOOST_cell_43418 ( .a(TIMEBOOST_net_13947), .b(n_6645), .o(TIMEBOOST_net_12193) );
in01s01 g61936_u0 ( .a(FE_OFN1812_n_7845), .o(g61936_sb) );
na02s01 TIMEBOOST_cell_18813 ( .a(TIMEBOOST_net_4663), .b(g63062_sb), .o(n_5126) );
na02s01 TIMEBOOST_cell_36432 ( .a(TIMEBOOST_net_10454), .b(g65713_db), .o(n_1612) );
na02s01 TIMEBOOST_cell_36434 ( .a(TIMEBOOST_net_10455), .b(g65782_db), .o(n_1650) );
in01s01 g61937_u0 ( .a(FE_OFN716_n_8176), .o(g61937_sb) );
na02m02 TIMEBOOST_cell_10154 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__Q), .b(n_13447), .o(TIMEBOOST_net_1644) );
na02m02 TIMEBOOST_cell_42301 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__31__Q), .b(n_9729), .o(TIMEBOOST_net_13389) );
na02f02 TIMEBOOST_cell_42302 ( .a(TIMEBOOST_net_13389), .b(g57198_sb), .o(TIMEBOOST_net_11639) );
na02s01 TIMEBOOST_cell_16883 ( .a(TIMEBOOST_net_3698), .b(g64304_db), .o(n_3871) );
na02s01 TIMEBOOST_cell_45147 ( .a(FE_OFN201_n_9230), .b(g58415_sb), .o(TIMEBOOST_net_14812) );
na02s01 TIMEBOOST_cell_43044 ( .a(TIMEBOOST_net_13760), .b(g58400_sb), .o(n_9208) );
in01s01 g61939_u0 ( .a(n_8272), .o(g61939_sb) );
na02s01 TIMEBOOST_cell_44965 ( .a(g58123_sb), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_14721) );
na02s01 g61939_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__Q), .b(n_8272), .o(g61939_db) );
na02s02 TIMEBOOST_cell_39846 ( .a(TIMEBOOST_net_12161), .b(g62623_sb), .o(n_6311) );
in01s01 g61940_u0 ( .a(FE_OFN713_n_8140), .o(g61940_sb) );
na02s02 TIMEBOOST_cell_18801 ( .a(TIMEBOOST_net_4657), .b(g63054_sb), .o(n_7122) );
na02m02 TIMEBOOST_cell_44171 ( .a(n_9014), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__Q), .o(TIMEBOOST_net_14324) );
na02s02 TIMEBOOST_cell_37743 ( .a(FE_OFN252_n_9868), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__Q), .o(TIMEBOOST_net_11110) );
in01s01 g61941_u0 ( .a(FE_OFN2212_n_8407), .o(g61941_sb) );
na02s01 TIMEBOOST_cell_38554 ( .a(TIMEBOOST_net_11515), .b(g62032_sb), .o(n_7783) );
na02s01 TIMEBOOST_cell_38746 ( .a(TIMEBOOST_net_11611), .b(g53913_sb), .o(n_13528) );
na02f02 TIMEBOOST_cell_38994 ( .a(TIMEBOOST_net_11735), .b(g58835_sb), .o(n_8602) );
in01s01 g61942_u0 ( .a(FE_OFN2257_n_8060), .o(g61942_sb) );
na02f02 TIMEBOOST_cell_38876 ( .a(TIMEBOOST_net_11676), .b(g58481_sb), .o(n_8977) );
na02s01 TIMEBOOST_cell_18116 ( .a(g63562_sb), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_), .o(TIMEBOOST_net_4315) );
na02m02 TIMEBOOST_cell_39477 ( .a(FE_OFN1149_n_13249), .b(TIMEBOOST_net_9658), .o(TIMEBOOST_net_11977) );
in01s03 g61943_u0 ( .a(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61943_sb) );
na02s01 TIMEBOOST_cell_22302 ( .a(g52461_da), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_6408) );
na02s01 g61943_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61943_db) );
na02s01 TIMEBOOST_cell_22306 ( .a(g52463_da), .b(FE_OFN1022_n_11877), .o(TIMEBOOST_net_6410) );
in01s01 g61944_u0 ( .a(FE_OFN709_n_8232), .o(g61944_sb) );
na02s02 TIMEBOOST_cell_10156 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__Q), .b(FE_OFN2059_n_13447), .o(TIMEBOOST_net_1645) );
na02s02 TIMEBOOST_cell_45447 ( .a(n_3522), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q), .o(TIMEBOOST_net_14962) );
na02s01 TIMEBOOST_cell_41948 ( .a(TIMEBOOST_net_13212), .b(g58277_db), .o(n_9525) );
in01s01 g61945_u0 ( .a(FE_OFN2257_n_8060), .o(g61945_sb) );
na02s01 TIMEBOOST_cell_37745 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__Q), .b(wbs_dat_i_10_), .o(TIMEBOOST_net_11111) );
na02s01 TIMEBOOST_cell_18118 ( .a(g63574_sb), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_), .o(TIMEBOOST_net_4316) );
na02s01 TIMEBOOST_cell_40382 ( .a(TIMEBOOST_net_12429), .b(g65391_db), .o(n_4241) );
in01s01 g61946_u0 ( .a(FE_OFN710_n_8232), .o(g61946_sb) );
na02s01 TIMEBOOST_cell_37490 ( .a(TIMEBOOST_net_10983), .b(g65834_sb), .o(TIMEBOOST_net_332) );
na02s01 TIMEBOOST_cell_17122 ( .a(pci_target_unit_del_sync_addr_in_219), .b(parchk_pci_ad_reg_in_1220), .o(TIMEBOOST_net_3818) );
na02s02 TIMEBOOST_cell_37744 ( .a(TIMEBOOST_net_11110), .b(FE_OFN1670_n_9477), .o(TIMEBOOST_net_4350) );
in01s01 g61947_u0 ( .a(FE_OFN2257_n_8060), .o(g61947_sb) );
na02s01 TIMEBOOST_cell_37492 ( .a(TIMEBOOST_net_10984), .b(g65831_sb), .o(TIMEBOOST_net_329) );
na03s02 TIMEBOOST_cell_40621 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__Q), .b(n_3698), .c(FE_OFN1208_n_6356), .o(TIMEBOOST_net_12549) );
na02f02 TIMEBOOST_cell_37077 ( .a(FE_OCP_RBN1998_n_13971), .b(TIMEBOOST_net_10237), .o(TIMEBOOST_net_10777) );
in01s01 g61948_u0 ( .a(FE_OFN709_n_8232), .o(g61948_sb) );
na02s02 TIMEBOOST_cell_40384 ( .a(TIMEBOOST_net_12430), .b(g64831_sb), .o(n_4449) );
na02f02 TIMEBOOST_cell_41628 ( .a(FE_OFN1441_n_9372), .b(TIMEBOOST_net_13052), .o(TIMEBOOST_net_11679) );
na02s02 TIMEBOOST_cell_39406 ( .a(TIMEBOOST_net_11941), .b(g58158_sb), .o(n_9631) );
in01s01 g61949_u0 ( .a(n_8272), .o(g61949_sb) );
na02s01 TIMEBOOST_cell_45093 ( .a(g64316_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__Q), .o(TIMEBOOST_net_14785) );
na02s01 g61949_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__Q), .b(n_8272), .o(g61949_db) );
na02s01 TIMEBOOST_cell_42916 ( .a(TIMEBOOST_net_13696), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_11182) );
in01s01 g61950_u0 ( .a(FE_OFN2081_n_8176), .o(g61950_sb) );
na02s02 TIMEBOOST_cell_38290 ( .a(TIMEBOOST_net_11383), .b(g61902_sb), .o(n_8019) );
na02s02 TIMEBOOST_cell_37392 ( .a(TIMEBOOST_net_10934), .b(FE_OFN2072_n_15978), .o(TIMEBOOST_net_9854) );
na02s02 TIMEBOOST_cell_38292 ( .a(TIMEBOOST_net_11384), .b(g61917_sb), .o(n_7987) );
in01s01 g61951_u0 ( .a(FE_OFN710_n_8232), .o(g61951_sb) );
na02s01 TIMEBOOST_cell_37494 ( .a(TIMEBOOST_net_10985), .b(g65846_sb), .o(TIMEBOOST_net_334) );
na02f04 TIMEBOOST_cell_44773 ( .a(TIMEBOOST_net_3225), .b(TIMEBOOST_net_3252), .o(TIMEBOOST_net_14625) );
na02s01 TIMEBOOST_cell_37496 ( .a(TIMEBOOST_net_10986), .b(g65833_sb), .o(TIMEBOOST_net_331) );
in01s01 g61952_u0 ( .a(FE_OFN707_n_8119), .o(g61952_sb) );
na02s02 TIMEBOOST_cell_38294 ( .a(TIMEBOOST_net_11385), .b(g61828_sb), .o(n_8130) );
na02s01 TIMEBOOST_cell_39365 ( .a(TIMEBOOST_net_3861), .b(FE_OFN2113_n_2053), .o(TIMEBOOST_net_11921) );
na02s01 TIMEBOOST_cell_37213 ( .a(parchk_pci_ad_reg_in_1216), .b(pci_target_unit_del_sync_addr_in_215), .o(TIMEBOOST_net_10845) );
na02s02 TIMEBOOST_cell_22281 ( .a(n_10278), .b(TIMEBOOST_net_6397), .o(n_11878) );
na02s01 g61953_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__Q), .b(n_7102), .o(g61953_db) );
na03f02 TIMEBOOST_cell_36090 ( .a(FE_OFN1565_n_12502), .b(TIMEBOOST_net_10190), .c(n_12313), .o(n_12726) );
in01s01 g61954_u0 ( .a(FE_OFN707_n_8119), .o(g61954_sb) );
na02m02 TIMEBOOST_cell_10158 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__Q), .b(FE_OFN2059_n_13447), .o(TIMEBOOST_net_1646) );
na02f02 TIMEBOOST_cell_41570 ( .a(TIMEBOOST_net_13023), .b(g57119_sb), .o(n_11626) );
na02s02 TIMEBOOST_cell_43241 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__Q), .b(n_3653), .o(TIMEBOOST_net_13859) );
in01s01 g61955_u0 ( .a(FE_OFN1094_g64577_p), .o(g61955_sb) );
na02s01 TIMEBOOST_cell_30940 ( .a(n_3744), .b(g65060_sb), .o(TIMEBOOST_net_9381) );
na02s01 TIMEBOOST_cell_42690 ( .a(TIMEBOOST_net_13583), .b(g65001_db), .o(n_3640) );
na02s01 TIMEBOOST_cell_30941 ( .a(TIMEBOOST_net_9381), .b(g65060_db), .o(n_3613) );
in01s01 g61956_u0 ( .a(FE_OFN1097_g64577_p), .o(g61956_sb) );
na02s01 TIMEBOOST_cell_36536 ( .a(TIMEBOOST_net_10506), .b(g65767_sb), .o(TIMEBOOST_net_273) );
na02s01 g61956_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__1__Q), .b(FE_OFN1097_g64577_p), .o(g61956_db) );
na02s01 TIMEBOOST_cell_36538 ( .a(TIMEBOOST_net_10507), .b(g65749_sb), .o(TIMEBOOST_net_271) );
in01s01 g61957_u0 ( .a(FE_OFN1095_g64577_p), .o(g61957_sb) );
na02f02 TIMEBOOST_cell_36858 ( .a(TIMEBOOST_net_10667), .b(n_16162), .o(TIMEBOOST_net_9984) );
na02s01 g61957_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__Q), .b(FE_OFN1095_g64577_p), .o(g61957_db) );
na02s01 TIMEBOOST_cell_36860 ( .a(TIMEBOOST_net_10668), .b(g61743_db), .o(n_8331) );
in01s01 g61958_u0 ( .a(FE_OFN1094_g64577_p), .o(g61958_sb) );
na02f02 TIMEBOOST_cell_42190 ( .a(TIMEBOOST_net_13333), .b(FE_OFN1425_n_8567), .o(TIMEBOOST_net_12285) );
na02s02 TIMEBOOST_cell_30943 ( .a(TIMEBOOST_net_9382), .b(g65070_sb), .o(n_3606) );
in01s01 g61959_u0 ( .a(FE_OFN1097_g64577_p), .o(g61959_sb) );
na02m02 TIMEBOOST_cell_36862 ( .a(TIMEBOOST_net_10669), .b(TIMEBOOST_net_608), .o(n_14845) );
na02s01 g61959_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q), .b(FE_OFN1097_g64577_p), .o(g61959_db) );
na02s01 TIMEBOOST_cell_36864 ( .a(TIMEBOOST_net_10670), .b(g63124_db), .o(n_5006) );
na02s01 TIMEBOOST_cell_17815 ( .a(TIMEBOOST_net_4164), .b(g61793_sb), .o(n_8213) );
na02s01 g61960_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61960_db) );
in01s01 g61961_u0 ( .a(FE_OFN1094_g64577_p), .o(g61961_sb) );
na02s02 TIMEBOOST_cell_30944 ( .a(n_3752), .b(g65050_sb), .o(TIMEBOOST_net_9383) );
na02s01 g61961_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__Q), .b(FE_OFN1095_g64577_p), .o(g61961_db) );
na02s02 TIMEBOOST_cell_30945 ( .a(TIMEBOOST_net_9383), .b(g65050_db), .o(n_3620) );
in01s01 g61962_u0 ( .a(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61962_sb) );
na02s01 TIMEBOOST_cell_44879 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__Q), .b(g65896_sb), .o(TIMEBOOST_net_14678) );
na02s01 g61962_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61962_db) );
na02m02 TIMEBOOST_cell_43969 ( .a(n_9445), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__Q), .o(TIMEBOOST_net_14223) );
in01s01 g61963_u0 ( .a(FE_OFN1095_g64577_p), .o(g61963_sb) );
na02s02 TIMEBOOST_cell_19137 ( .a(TIMEBOOST_net_4825), .b(g59231_sb), .o(TIMEBOOST_net_590) );
na02s01 g61963_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__Q), .b(FE_OFN1095_g64577_p), .o(g61963_db) );
na02s02 TIMEBOOST_cell_44423 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_795), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_30__Q), .o(TIMEBOOST_net_14450) );
na02s02 TIMEBOOST_cell_38748 ( .a(TIMEBOOST_net_11612), .b(g53916_sb), .o(n_13526) );
na02s01 g61964_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61964_db) );
na02s02 TIMEBOOST_cell_38296 ( .a(TIMEBOOST_net_11386), .b(g61817_sb), .o(n_8157) );
in01s01 g61965_u0 ( .a(FE_OFN1095_g64577_p), .o(g61965_sb) );
na02s01 TIMEBOOST_cell_36866 ( .a(TIMEBOOST_net_10671), .b(g61775_db), .o(n_8258) );
na02s01 g61965_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__Q), .b(FE_OFN1095_g64577_p), .o(g61965_db) );
na02s01 TIMEBOOST_cell_36868 ( .a(TIMEBOOST_net_10672), .b(g61771_db), .o(n_8267) );
na02s02 TIMEBOOST_cell_38298 ( .a(TIMEBOOST_net_11387), .b(g61725_sb), .o(n_8371) );
na02s01 g61966_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61966_db) );
no02f06 TIMEBOOST_cell_16372 ( .a(FE_RN_9_0), .b(n_15456), .o(TIMEBOOST_net_3443) );
na02s02 TIMEBOOST_cell_38300 ( .a(TIMEBOOST_net_11388), .b(g61714_sb), .o(n_8397) );
na02s01 g61967_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61967_db) );
na02f06 TIMEBOOST_cell_36836 ( .a(TIMEBOOST_net_10656), .b(g75162_db), .o(n_16534) );
na02s02 TIMEBOOST_cell_43242 ( .a(TIMEBOOST_net_13859), .b(FE_OFN1253_n_4143), .o(TIMEBOOST_net_12043) );
na02s01 g61968_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61968_db) );
na02f02 TIMEBOOST_cell_44522 ( .a(TIMEBOOST_net_14499), .b(FE_OFN2179_n_8567), .o(TIMEBOOST_net_12999) );
na02s01 TIMEBOOST_cell_37250 ( .a(TIMEBOOST_net_10863), .b(FE_OFN665_n_4495), .o(TIMEBOOST_net_9382) );
na02s01 g61969_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61969_db) );
na02s02 TIMEBOOST_cell_18633 ( .a(TIMEBOOST_net_4573), .b(g63079_sb), .o(n_5094) );
na02s02 TIMEBOOST_cell_38302 ( .a(TIMEBOOST_net_11389), .b(g61936_sb), .o(n_7951) );
na02s01 g61970_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61970_db) );
na02s02 TIMEBOOST_cell_43419 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__Q), .b(n_3620), .o(TIMEBOOST_net_13948) );
na02s01 g61971_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61971_db) );
na02f02 TIMEBOOST_cell_43970 ( .a(TIMEBOOST_net_14223), .b(FE_OFN1391_n_8567), .o(TIMEBOOST_net_12702) );
na02s01 TIMEBOOST_cell_36436 ( .a(TIMEBOOST_net_10456), .b(g65760_db), .o(n_1603) );
na02s01 g61972_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61972_db) );
na02s02 TIMEBOOST_cell_19305 ( .a(TIMEBOOST_net_4909), .b(g60662_sb), .o(n_5657) );
na02f02 TIMEBOOST_cell_22319 ( .a(TIMEBOOST_net_6416), .b(FE_OFN1748_n_12004), .o(n_12512) );
na02s01 g61973_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61973_db) );
na02f02 TIMEBOOST_cell_43806 ( .a(TIMEBOOST_net_14141), .b(FE_OFN1392_n_8567), .o(TIMEBOOST_net_12960) );
na02s02 TIMEBOOST_cell_43511 ( .a(n_4372), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__Q), .o(TIMEBOOST_net_13994) );
na02s01 g61974_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61974_db) );
na03s02 TIMEBOOST_cell_38091 ( .a(TIMEBOOST_net_3471), .b(g64334_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__Q), .o(TIMEBOOST_net_11284) );
na02f02 TIMEBOOST_cell_43714 ( .a(TIMEBOOST_net_14095), .b(n_9144), .o(TIMEBOOST_net_13373) );
na02s01 g61975_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61975_db) );
na02f02 TIMEBOOST_cell_22321 ( .a(TIMEBOOST_net_6417), .b(FE_OFN1748_n_12004), .o(n_12669) );
na02s01 TIMEBOOST_cell_36438 ( .a(TIMEBOOST_net_10457), .b(g64172_db), .o(n_3993) );
na02s01 g61976_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61976_db) );
na02s02 TIMEBOOST_cell_19307 ( .a(TIMEBOOST_net_4910), .b(g60665_sb), .o(n_5654) );
na02s01 TIMEBOOST_cell_18911 ( .a(TIMEBOOST_net_4712), .b(g63133_sb), .o(n_4984) );
na02s01 g61977_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61977_db) );
na02m02 TIMEBOOST_cell_43759 ( .a(n_9418), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__Q), .o(TIMEBOOST_net_14118) );
na02s01 TIMEBOOST_cell_36324 ( .a(TIMEBOOST_net_10400), .b(g65951_db), .o(n_2168) );
na02s01 g61978_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61978_db) );
na02s02 TIMEBOOST_cell_19309 ( .a(TIMEBOOST_net_4911), .b(g60609_sb), .o(n_4845) );
na02s02 TIMEBOOST_cell_43243 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__Q), .b(n_3594), .o(TIMEBOOST_net_13860) );
na02s01 g61979_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61979_db) );
na02f02 TIMEBOOST_cell_22337 ( .a(TIMEBOOST_net_6425), .b(n_10596), .o(n_12141) );
na03f02 TIMEBOOST_cell_22338 ( .a(n_9260), .b(n_10023), .c(n_10026), .o(TIMEBOOST_net_6426) );
na02s01 g61980_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61980_db) );
na02f02 TIMEBOOST_cell_22339 ( .a(TIMEBOOST_net_6426), .b(n_10614), .o(n_12144) );
na02s01 TIMEBOOST_cell_36326 ( .a(TIMEBOOST_net_10401), .b(g67051_sb), .o(n_1444) );
na02s01 g61981_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61981_db) );
na02s02 TIMEBOOST_cell_19313 ( .a(TIMEBOOST_net_4913), .b(g60673_sb), .o(n_5646) );
na02s01 TIMEBOOST_cell_36328 ( .a(TIMEBOOST_net_10402), .b(g65961_db), .o(n_2161) );
na02s01 g61982_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61982_db) );
na02s02 TIMEBOOST_cell_19311 ( .a(TIMEBOOST_net_4912), .b(g60668_sb), .o(n_5650) );
na03f02 TIMEBOOST_cell_22340 ( .a(n_9315), .b(n_9319), .c(n_10188), .o(TIMEBOOST_net_6427) );
na02s01 g61983_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61983_db) );
na02f02 TIMEBOOST_cell_22341 ( .a(TIMEBOOST_net_6427), .b(n_10183), .o(n_12161) );
na02f02 TIMEBOOST_cell_38996 ( .a(TIMEBOOST_net_11736), .b(g58824_sb), .o(n_8617) );
na02s01 g61984_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61984_db) );
na02s01 TIMEBOOST_cell_43244 ( .a(TIMEBOOST_net_13860), .b(FE_OFN1208_n_6356), .o(TIMEBOOST_net_12113) );
na03f02 TIMEBOOST_cell_22342 ( .a(n_10102), .b(n_9290), .c(n_9293), .o(TIMEBOOST_net_6428) );
na02s01 g61985_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61985_db) );
na02f02 TIMEBOOST_cell_22343 ( .a(TIMEBOOST_net_6428), .b(n_10944), .o(n_12153) );
na02s02 TIMEBOOST_cell_38304 ( .a(TIMEBOOST_net_11390), .b(n_5743), .o(n_7722) );
na02s01 g61986_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61986_db) );
na02s01 TIMEBOOST_cell_43310 ( .a(TIMEBOOST_net_13893), .b(g63145_sb), .o(n_5850) );
na03f02 TIMEBOOST_cell_22344 ( .a(n_10066), .b(n_9272), .c(n_9271), .o(TIMEBOOST_net_6429) );
na02s01 g61987_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61987_db) );
na02m02 TIMEBOOST_cell_42191 ( .a(n_9406), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__Q), .o(TIMEBOOST_net_13334) );
na02s02 TIMEBOOST_cell_18923 ( .a(TIMEBOOST_net_4718), .b(g62768_sb), .o(n_5458) );
na02s01 g61988_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61988_db) );
na02s02 TIMEBOOST_cell_43420 ( .a(TIMEBOOST_net_13948), .b(n_6431), .o(TIMEBOOST_net_12203) );
na02s01 g61989_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61989_db) );
na02m02 TIMEBOOST_cell_43971 ( .a(n_9048), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q), .o(TIMEBOOST_net_14224) );
in01s01 g61990_u0 ( .a(n_8069), .o(g61990_sb) );
na02s02 TIMEBOOST_cell_39848 ( .a(TIMEBOOST_net_12162), .b(g62941_sb), .o(n_5999) );
na02s02 TIMEBOOST_cell_40367 ( .a(pci_target_unit_fifos_pcir_data_in_163), .b(g65709_sb), .o(TIMEBOOST_net_12422) );
na02s01 TIMEBOOST_cell_16888 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__Q), .o(TIMEBOOST_net_3701) );
in01s01 g61991_u0 ( .a(FE_OFN2212_n_8407), .o(g61991_sb) );
na02s02 TIMEBOOST_cell_38306 ( .a(TIMEBOOST_net_11391), .b(g58357_db), .o(n_9015) );
na02s02 TIMEBOOST_cell_18583 ( .a(TIMEBOOST_net_4548), .b(g63110_sb), .o(n_5036) );
na02s02 TIMEBOOST_cell_18585 ( .a(TIMEBOOST_net_4549), .b(g59370_sb), .o(n_7694) );
in01s01 g61992_u0 ( .a(n_8069), .o(g61992_sb) );
na02f02 TIMEBOOST_cell_44634 ( .a(TIMEBOOST_net_14555), .b(FE_OFN2173_n_8567), .o(TIMEBOOST_net_13488) );
na02s02 TIMEBOOST_cell_45189 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q), .b(n_4481), .o(TIMEBOOST_net_14833) );
na02s01 TIMEBOOST_cell_45148 ( .a(TIMEBOOST_net_14812), .b(g58415_db), .o(n_9203) );
in01s01 g61993_u0 ( .a(FE_OFN699_n_7845), .o(g61993_sb) );
na02s02 TIMEBOOST_cell_10554 ( .a(pci_cbe_o_2_), .b(n_14389), .o(TIMEBOOST_net_1844) );
na02s01 TIMEBOOST_cell_17392 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__Q), .b(g64245_sb), .o(TIMEBOOST_net_3953) );
na02s01 TIMEBOOST_cell_37452 ( .a(TIMEBOOST_net_10964), .b(FE_OFN775_n_15366), .o(TIMEBOOST_net_10563) );
in01s01 g61994_u0 ( .a(n_8272), .o(g61994_sb) );
na02s01 TIMEBOOST_cell_16890 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__Q), .o(TIMEBOOST_net_3702) );
na02s01 g61994_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__Q), .b(n_8272), .o(g61994_db) );
na03f04 TIMEBOOST_cell_36076 ( .a(FE_OFN1601_n_13995), .b(TIMEBOOST_net_10158), .c(FE_OFN1605_n_13997), .o(FE_RN_893_0) );
in01s01 g61995_u0 ( .a(FE_OFN702_n_7845), .o(g61995_sb) );
na02s02 TIMEBOOST_cell_37394 ( .a(TIMEBOOST_net_10935), .b(g65434_sb), .o(n_4220) );
na03f02 TIMEBOOST_cell_2003 ( .a(g52401_db), .b(g52401_sb), .c(n_3483), .o(n_14818) );
na02s01 TIMEBOOST_cell_41804 ( .a(TIMEBOOST_net_13140), .b(g62029_sb), .o(n_7838) );
na02f02 TIMEBOOST_cell_44202 ( .a(TIMEBOOST_net_14339), .b(FE_OFN1382_n_8567), .o(TIMEBOOST_net_12771) );
na02s01 g61996_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__Q), .b(n_8232), .o(g61996_db) );
na03s02 TIMEBOOST_cell_40357 ( .a(n_4488), .b(g64988_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__Q), .o(TIMEBOOST_net_12417) );
in01s01 g61997_u0 ( .a(n_8119), .o(g61997_sb) );
na02s02 TIMEBOOST_cell_42677 ( .a(g64905_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__Q), .o(TIMEBOOST_net_13577) );
na02f02 TIMEBOOST_cell_40051 ( .a(n_9425), .b(g57565_sb), .o(TIMEBOOST_net_12264) );
na02s01 TIMEBOOST_cell_39850 ( .a(TIMEBOOST_net_12163), .b(g62601_sb), .o(n_6348) );
in01s01 g61998_u0 ( .a(FE_OFN699_n_7845), .o(g61998_sb) );
na02s01 TIMEBOOST_cell_18725 ( .a(TIMEBOOST_net_4619), .b(g63034_sb), .o(n_5179) );
na02s01 TIMEBOOST_cell_17396 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__Q), .b(g64251_sb), .o(TIMEBOOST_net_3955) );
na02s02 TIMEBOOST_cell_18727 ( .a(TIMEBOOST_net_4620), .b(g62855_sb), .o(n_5258) );
in01s01 g61999_u0 ( .a(n_8232), .o(g61999_sb) );
na02s02 TIMEBOOST_cell_45149 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__Q), .b(n_2455), .o(TIMEBOOST_net_14813) );
na02s01 TIMEBOOST_cell_16824 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__Q), .b(g65311_sb), .o(TIMEBOOST_net_3669) );
na02f02 g61_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__Q), .o(n_15537) );
in01s01 g62000_u0 ( .a(FE_OFN2258_n_8060), .o(g62000_sb) );
na02s01 TIMEBOOST_cell_18729 ( .a(TIMEBOOST_net_4621), .b(g62856_sb), .o(n_5255) );
na02s01 TIMEBOOST_cell_45061 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__Q), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_14769) );
na02m02 TIMEBOOST_cell_38308 ( .a(FE_OCPN1911_FE_OFN1152_n_13249), .b(TIMEBOOST_net_11392), .o(TIMEBOOST_net_4752) );
in01s01 g62001_u0 ( .a(FE_OFN717_n_8176), .o(g62001_sb) );
na02s01 TIMEBOOST_cell_38310 ( .a(TIMEBOOST_net_11393), .b(g58396_db), .o(n_9005) );
na02s01 TIMEBOOST_cell_17420 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__Q), .b(g60687_sb), .o(TIMEBOOST_net_3967) );
na02s01 TIMEBOOST_cell_18735 ( .a(TIMEBOOST_net_4624), .b(g62826_sb), .o(n_5325) );
in01s01 g62002_u0 ( .a(FE_OFN702_n_7845), .o(g62002_sb) );
na02s02 TIMEBOOST_cell_18737 ( .a(TIMEBOOST_net_4625), .b(g62762_sb), .o(n_5470) );
na02s01 TIMEBOOST_cell_17398 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__Q), .b(g64259_sb), .o(TIMEBOOST_net_3956) );
na02s01 TIMEBOOST_cell_18739 ( .a(TIMEBOOST_net_4626), .b(g63119_sb), .o(n_5018) );
in01s01 g62003_u0 ( .a(n_8232), .o(g62003_sb) );
na02s01 TIMEBOOST_cell_39303 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__Q), .b(g65838_sb), .o(TIMEBOOST_net_11890) );
na02s02 TIMEBOOST_cell_45150 ( .a(TIMEBOOST_net_14813), .b(FE_OFN1252_n_4143), .o(TIMEBOOST_net_12067) );
na02s01 TIMEBOOST_cell_39852 ( .a(TIMEBOOST_net_12164), .b(g62971_sb), .o(n_5940) );
na02s01 TIMEBOOST_cell_40301 ( .a(n_4452), .b(g65052_sb), .o(TIMEBOOST_net_12389) );
na02s01 TIMEBOOST_cell_16902 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__Q), .b(g64282_sb), .o(TIMEBOOST_net_3708) );
in01s01 g62005_u0 ( .a(FE_OFN712_n_8140), .o(g62005_sb) );
na02s02 TIMEBOOST_cell_18875 ( .a(TIMEBOOST_net_4694), .b(g62725_sb), .o(n_5531) );
na02s01 TIMEBOOST_cell_17400 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__Q), .b(g64252_sb), .o(TIMEBOOST_net_3957) );
na02s01 TIMEBOOST_cell_38312 ( .a(TIMEBOOST_net_11394), .b(g63553_sb), .o(n_4924) );
in01s01 g62006_u0 ( .a(FE_OFN706_n_8119), .o(g62006_sb) );
na02m02 TIMEBOOST_cell_10160 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__Q), .b(n_13447), .o(TIMEBOOST_net_1647) );
na02s01 TIMEBOOST_cell_42948 ( .a(TIMEBOOST_net_13712), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_11937) );
na02s02 TIMEBOOST_cell_43025 ( .a(n_3954), .b(g62864_sb), .o(TIMEBOOST_net_13751) );
in01s01 g62007_u0 ( .a(n_8069), .o(g62007_sb) );
na02s02 TIMEBOOST_cell_36540 ( .a(TIMEBOOST_net_10508), .b(g64924_sb), .o(TIMEBOOST_net_9605) );
na02s01 TIMEBOOST_cell_36542 ( .a(TIMEBOOST_net_10509), .b(g65696_sb), .o(TIMEBOOST_net_267) );
na02s02 TIMEBOOST_cell_9269 ( .a(TIMEBOOST_net_1201), .b(n_13820), .o(TIMEBOOST_net_604) );
na02s01 g62008_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__Q), .b(n_8407), .o(g62008_db) );
na02f02 TIMEBOOST_cell_38998 ( .a(TIMEBOOST_net_11737), .b(g58820_sb), .o(n_8621) );
in01s01 g62009_u0 ( .a(FE_OFN713_n_8140), .o(g62009_sb) );
na02s01 TIMEBOOST_cell_18879 ( .a(TIMEBOOST_net_4696), .b(g62742_sb), .o(n_5495) );
na02s01 TIMEBOOST_cell_17402 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__Q), .b(g64341_sb), .o(TIMEBOOST_net_3958) );
na02s01 TIMEBOOST_cell_38314 ( .a(TIMEBOOST_net_11395), .b(g63152_sb), .o(n_4959) );
in01s01 g62010_u0 ( .a(FE_OFN706_n_8119), .o(g62010_sb) );
na02s01 TIMEBOOST_cell_42725 ( .a(g65942_db), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__Q), .o(TIMEBOOST_net_13601) );
na02s01 TIMEBOOST_cell_39254 ( .a(TIMEBOOST_net_11865), .b(g58383_db), .o(n_9448) );
na02f02 TIMEBOOST_cell_44294 ( .a(TIMEBOOST_net_14385), .b(FE_OFN1419_n_8567), .o(TIMEBOOST_net_12864) );
in01s01 g62011_u0 ( .a(FE_OFN704_n_8069), .o(g62011_sb) );
na02s01 TIMEBOOST_cell_38316 ( .a(TIMEBOOST_net_11396), .b(g63557_sb), .o(n_4920) );
na02s02 TIMEBOOST_cell_37396 ( .a(TIMEBOOST_net_10936), .b(TIMEBOOST_net_3437), .o(TIMEBOOST_net_5434) );
na02s02 TIMEBOOST_cell_38318 ( .a(TIMEBOOST_net_11397), .b(g62830_sb), .o(n_5315) );
in01s01 g62012_u0 ( .a(FE_OFN712_n_8140), .o(g62012_sb) );
na02s01 TIMEBOOST_cell_18741 ( .a(TIMEBOOST_net_4627), .b(g62752_sb), .o(n_5476) );
na02s02 TIMEBOOST_cell_43602 ( .a(TIMEBOOST_net_14039), .b(FE_OFN1250_n_4093), .o(TIMEBOOST_net_12574) );
na02s01 TIMEBOOST_cell_18743 ( .a(TIMEBOOST_net_4628), .b(g62767_sb), .o(n_5461) );
in01s01 g62013_u0 ( .a(FE_OFN712_n_8140), .o(g62013_sb) );
na02s01 TIMEBOOST_cell_18887 ( .a(TIMEBOOST_net_4700), .b(g62764_sb), .o(n_5467) );
na02s01 TIMEBOOST_cell_17404 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__Q), .b(g64342_sb), .o(TIMEBOOST_net_3959) );
na02f02 TIMEBOOST_cell_18889 ( .a(TIMEBOOST_net_4701), .b(g54318_db), .o(n_13290) );
in01s01 g62014_u0 ( .a(FE_OFN2084_n_8407), .o(g62014_sb) );
na02s02 TIMEBOOST_cell_18891 ( .a(TIMEBOOST_net_4702), .b(g62766_sb), .o(n_5463) );
na02s02 TIMEBOOST_cell_39854 ( .a(TIMEBOOST_net_12165), .b(g62533_sb), .o(n_6506) );
na02s02 TIMEBOOST_cell_38320 ( .a(TIMEBOOST_net_11398), .b(g62790_sb), .o(n_5409) );
in01s01 g62015_u0 ( .a(FE_OFN709_n_8232), .o(g62015_sb) );
na02m02 TIMEBOOST_cell_10162 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__Q), .b(n_13447), .o(TIMEBOOST_net_1648) );
na02s01 TIMEBOOST_cell_17279 ( .a(TIMEBOOST_net_3896), .b(g65427_da), .o(n_3508) );
na03s01 TIMEBOOST_cell_624 ( .a(n_4594), .b(g61959_sb), .c(g61959_db), .o(n_6953) );
in01s01 g62016_u0 ( .a(FE_OFN712_n_8140), .o(g62016_sb) );
na02s01 TIMEBOOST_cell_38322 ( .a(TIMEBOOST_net_11399), .b(g63136_sb), .o(n_4978) );
na02s01 TIMEBOOST_cell_17406 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__Q), .b(g64260_sb), .o(TIMEBOOST_net_3960) );
na02s02 TIMEBOOST_cell_18897 ( .a(TIMEBOOST_net_4705), .b(g62817_sb), .o(n_5342) );
in01s01 g62017_u0 ( .a(FE_OFN2212_n_8407), .o(g62017_sb) );
na02s02 TIMEBOOST_cell_38324 ( .a(TIMEBOOST_net_11400), .b(g63041_sb), .o(n_5168) );
na02s01 TIMEBOOST_cell_44880 ( .a(TIMEBOOST_net_14678), .b(g65896_db), .o(n_1858) );
na02f02 TIMEBOOST_cell_10941 ( .a(TIMEBOOST_net_2037), .b(g54320_da), .o(n_13287) );
in01s01 g62018_u0 ( .a(FE_OFN2084_n_8407), .o(g62018_sb) );
na02s01 TIMEBOOST_cell_39386 ( .a(TIMEBOOST_net_11931), .b(g62773_sb), .o(TIMEBOOST_net_9746) );
na03s02 TIMEBOOST_cell_39197 ( .a(n_8884), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_18__Q), .c(g58776_sb), .o(TIMEBOOST_net_11837) );
na02s01 TIMEBOOST_cell_18747 ( .a(TIMEBOOST_net_4630), .b(g63109_sb), .o(n_5038) );
in01s01 g62019_u0 ( .a(FE_OFN2212_n_8407), .o(g62019_sb) );
na02m02 TIMEBOOST_cell_42828 ( .a(TIMEBOOST_net_13652), .b(n_3027), .o(TIMEBOOST_net_340) );
na02s01 TIMEBOOST_cell_17199 ( .a(TIMEBOOST_net_3856), .b(g65365_db), .o(n_3534) );
in01s01 TIMEBOOST_cell_45905 ( .a(wbm_dat_i_12_), .o(TIMEBOOST_net_15212) );
in01s01 g62020_u0 ( .a(FE_OFN1812_n_7845), .o(g62020_sb) );
na03s02 TIMEBOOST_cell_37699 ( .a(n_2213), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__Q), .c(FE_OFN716_n_8176), .o(TIMEBOOST_net_11088) );
na02s01 TIMEBOOST_cell_36440 ( .a(TIMEBOOST_net_10458), .b(g58078_sb), .o(TIMEBOOST_net_9769) );
na02s01 TIMEBOOST_cell_36442 ( .a(TIMEBOOST_net_10459), .b(g63537_db), .o(n_4618) );
na02s01 TIMEBOOST_cell_16961 ( .a(TIMEBOOST_net_3737), .b(g65222_sb), .o(n_2665) );
na02s01 g62021_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g62021_db) );
na02s02 TIMEBOOST_cell_43421 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__Q), .b(n_3635), .o(TIMEBOOST_net_13949) );
in01s01 g62022_u0 ( .a(FE_OFN699_n_7845), .o(g62022_sb) );
na02s02 TIMEBOOST_cell_38326 ( .a(TIMEBOOST_net_11401), .b(g63080_sb), .o(n_5092) );
na02s01 TIMEBOOST_cell_17408 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__Q), .b(g64256_sb), .o(TIMEBOOST_net_3961) );
na02s01 TIMEBOOST_cell_38328 ( .a(TIMEBOOST_net_11402), .b(g63014_sb), .o(n_5221) );
in01s01 g62023_u0 ( .a(FE_OFN719_n_8060), .o(g62023_sb) );
na02s02 TIMEBOOST_cell_38672 ( .a(TIMEBOOST_net_11574), .b(g62619_sb), .o(n_6321) );
na02f02 TIMEBOOST_cell_39000 ( .a(TIMEBOOST_net_11738), .b(g58805_sb), .o(n_8636) );
na02f02 TIMEBOOST_cell_39002 ( .a(TIMEBOOST_net_11739), .b(g58816_sb), .o(n_8625) );
in01s01 g62024_u0 ( .a(FE_OFN720_n_8060), .o(g62024_sb) );
na02s02 TIMEBOOST_cell_38088 ( .a(TIMEBOOST_net_11282), .b(FE_OFN1126_g64577_p), .o(TIMEBOOST_net_4549) );
na02m02 TIMEBOOST_cell_43624 ( .a(TIMEBOOST_net_14050), .b(FE_OFN1311_n_6624), .o(TIMEBOOST_net_12235) );
na02s01 TIMEBOOST_cell_37925 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__Q), .o(TIMEBOOST_net_11201) );
in01s01 g62025_u0 ( .a(FE_OFN701_n_7845), .o(g62025_sb) );
na02m02 TIMEBOOST_cell_44245 ( .a(n_9744), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q), .o(TIMEBOOST_net_14361) );
na02s01 g62025_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__Q), .b(FE_OFN701_n_7845), .o(g62025_db) );
in01s01 TIMEBOOST_cell_32849 ( .a(TIMEBOOST_net_10350), .o(TIMEBOOST_net_10349) );
in01s01 g62026_u0 ( .a(FE_OFN720_n_8060), .o(g62026_sb) );
na02s01 TIMEBOOST_cell_38076 ( .a(TIMEBOOST_net_11276), .b(FE_OFN1139_g64577_p), .o(TIMEBOOST_net_4593) );
na02f02 TIMEBOOST_cell_38812 ( .a(TIMEBOOST_net_11644), .b(g57471_sb), .o(n_10342) );
na02s02 TIMEBOOST_cell_38072 ( .a(TIMEBOOST_net_11274), .b(FE_OFN2106_g64577_p), .o(TIMEBOOST_net_4676) );
in01s01 g62027_u0 ( .a(FE_OFN699_n_7845), .o(g62027_sb) );
na02s01 TIMEBOOST_cell_18787 ( .a(TIMEBOOST_net_4650), .b(g63033_sb), .o(n_5181) );
na02s02 TIMEBOOST_cell_17410 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__Q), .b(g64263_sb), .o(TIMEBOOST_net_3962) );
na02s01 TIMEBOOST_cell_38330 ( .a(TIMEBOOST_net_11403), .b(g63026_sb), .o(n_5194) );
in01s01 g62028_u0 ( .a(FE_OFN702_n_7845), .o(g62028_sb) );
no02s02 TIMEBOOST_cell_41700 ( .a(TIMEBOOST_net_13088), .b(n_1666), .o(TIMEBOOST_net_10822) );
na02s01 TIMEBOOST_cell_17412 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q), .b(g64250_sb), .o(TIMEBOOST_net_3963) );
na02s02 TIMEBOOST_cell_45151 ( .a(n_3582), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__Q), .o(TIMEBOOST_net_14814) );
in01s01 g62029_u0 ( .a(FE_OFN702_n_7845), .o(g62029_sb) );
na02f02 TIMEBOOST_cell_41140 ( .a(TIMEBOOST_net_12808), .b(g57587_sb), .o(n_10290) );
na02f02 TIMEBOOST_cell_44172 ( .a(TIMEBOOST_net_14324), .b(FE_OFN1413_n_8567), .o(TIMEBOOST_net_13395) );
no02f02 TIMEBOOST_cell_22069 ( .a(TIMEBOOST_net_6291), .b(n_7824), .o(g53077_p) );
in01s01 g62030_u0 ( .a(FE_OFN1700_n_5751), .o(g62030_sb) );
na03s02 TIMEBOOST_cell_37787 ( .a(g65901_da), .b(g65901_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__Q), .o(TIMEBOOST_net_11132) );
na02s02 TIMEBOOST_cell_16959 ( .a(TIMEBOOST_net_3736), .b(g65218_sb), .o(n_2669) );
na02s02 TIMEBOOST_cell_16957 ( .a(TIMEBOOST_net_3735), .b(g65228_sb), .o(n_2659) );
in01s02 g62031_u0 ( .a(FE_OFN1145_n_15261), .o(g62031_sb) );
na02s02 TIMEBOOST_cell_3311 ( .a(TIMEBOOST_net_235), .b(n_4465), .o(n_4419) );
na02s02 TIMEBOOST_cell_43396 ( .a(TIMEBOOST_net_13936), .b(n_6319), .o(TIMEBOOST_net_12180) );
na02s01 TIMEBOOST_cell_37678 ( .a(TIMEBOOST_net_11077), .b(g61739_sb), .o(n_8339) );
in01s01 g62032_u0 ( .a(FE_OFN1300_n_5763), .o(g62032_sb) );
na02s01 TIMEBOOST_cell_18783 ( .a(TIMEBOOST_net_4648), .b(g63024_sb), .o(n_5198) );
na02s02 TIMEBOOST_cell_16955 ( .a(TIMEBOOST_net_3734), .b(g65223_sb), .o(n_2664) );
na02s02 TIMEBOOST_cell_43607 ( .a(n_4918), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__Q), .o(TIMEBOOST_net_14042) );
in01s02 g62033_u0 ( .a(FE_OFN1143_n_15261), .o(g62033_sb) );
na02s02 TIMEBOOST_cell_38332 ( .a(TIMEBOOST_net_11404), .b(g63083_sb), .o(n_5088) );
na02m02 TIMEBOOST_cell_44173 ( .a(n_9507), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__Q), .o(TIMEBOOST_net_14325) );
na02s01 TIMEBOOST_cell_42678 ( .a(TIMEBOOST_net_13577), .b(n_4447), .o(TIMEBOOST_net_12392) );
in01s01 g62034_u0 ( .a(FE_OFN1302_n_5763), .o(g62034_sb) );
na02m02 TIMEBOOST_cell_41591 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_27__Q), .b(FE_OFN233_n_9876), .o(TIMEBOOST_net_13034) );
na02s02 TIMEBOOST_cell_39256 ( .a(TIMEBOOST_net_11866), .b(g58444_db), .o(n_9409) );
na02s02 TIMEBOOST_cell_45448 ( .a(TIMEBOOST_net_14962), .b(FE_OFN1231_n_6391), .o(TIMEBOOST_net_13288) );
in01s01 g62035_u0 ( .a(FE_OFN1301_n_5763), .o(g62035_sb) );
na02f02 TIMEBOOST_cell_42304 ( .a(TIMEBOOST_net_13390), .b(g57501_sb), .o(n_11236) );
na03s02 TIMEBOOST_cell_36765 ( .a(g64106_da), .b(g64106_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__Q), .o(TIMEBOOST_net_10621) );
na02f02 TIMEBOOST_cell_41582 ( .a(TIMEBOOST_net_13029), .b(g57433_sb), .o(n_10823) );
in01s01 g62036_u0 ( .a(FE_OFN1301_n_5763), .o(g62036_sb) );
na03s01 TIMEBOOST_cell_37713 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__Q), .b(FE_OFN702_n_7845), .c(n_2209), .o(TIMEBOOST_net_11095) );
na02f02 TIMEBOOST_cell_43972 ( .a(TIMEBOOST_net_14224), .b(FE_OFN1382_n_8567), .o(TIMEBOOST_net_12809) );
na02f02 TIMEBOOST_cell_44336 ( .a(TIMEBOOST_net_14406), .b(FE_OFN1404_n_8567), .o(TIMEBOOST_net_12686) );
in01s01 g62037_u0 ( .a(FE_OFN1301_n_5763), .o(g62037_sb) );
na02s02 TIMEBOOST_cell_43494 ( .a(TIMEBOOST_net_13985), .b(FE_OFN1234_n_6391), .o(TIMEBOOST_net_12204) );
na02s01 TIMEBOOST_cell_39319 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__Q), .b(g65874_sb), .o(TIMEBOOST_net_11898) );
na02s01 TIMEBOOST_cell_2852 ( .a(pci_target_unit_wishbone_master_burst_chopped), .b(n_1183), .o(TIMEBOOST_net_6) );
in01s01 g62038_u0 ( .a(FE_OFN1302_n_5763), .o(g62038_sb) );
na02s01 TIMEBOOST_cell_2853 ( .a(TIMEBOOST_net_6), .b(n_898), .o(n_1185) );
na02s04 TIMEBOOST_cell_45819 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_19__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_784), .o(TIMEBOOST_net_15148) );
na02s01 TIMEBOOST_cell_2854 ( .a(pci_target_unit_wishbone_master_first_wb_data_access), .b(n_705), .o(TIMEBOOST_net_7) );
in01s01 g62039_u0 ( .a(FE_OFN1302_n_5763), .o(g62039_sb) );
na02s01 TIMEBOOST_cell_2855 ( .a(TIMEBOOST_net_7), .b(n_1183), .o(n_2027) );
na02s01 TIMEBOOST_cell_37767 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__Q), .b(wbs_dat_i_2_), .o(TIMEBOOST_net_11122) );
no02s01 TIMEBOOST_cell_2856 ( .a(n_23), .b(wbs_bte_i_1_), .o(TIMEBOOST_net_8) );
in01s01 g62040_u0 ( .a(FE_OFN1302_n_5763), .o(g62040_sb) );
no02s01 TIMEBOOST_cell_2857 ( .a(TIMEBOOST_net_8), .b(n_748), .o(g64630_BP) );
na02s01 TIMEBOOST_cell_37769 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__Q), .b(wbs_dat_i_13_), .o(TIMEBOOST_net_11123) );
na02s02 TIMEBOOST_cell_43504 ( .a(TIMEBOOST_net_13990), .b(FE_OFN1231_n_6391), .o(TIMEBOOST_net_12623) );
in01s01 g62041_u0 ( .a(FE_OFN1301_n_5763), .o(g62041_sb) );
na02s01 TIMEBOOST_cell_45449 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q), .b(TIMEBOOST_net_899), .o(TIMEBOOST_net_14963) );
na03s02 TIMEBOOST_cell_36767 ( .a(g64105_da), .b(g64105_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__Q), .o(TIMEBOOST_net_10622) );
na02f02 TIMEBOOST_cell_44694 ( .a(TIMEBOOST_net_14585), .b(TIMEBOOST_net_6264), .o(n_9236) );
in01s01 g62042_u0 ( .a(FE_OFN1302_n_5763), .o(g62042_sb) );
na02s01 TIMEBOOST_cell_41994 ( .a(TIMEBOOST_net_13235), .b(g62543_sb), .o(n_6480) );
na02f02 TIMEBOOST_cell_44174 ( .a(TIMEBOOST_net_14325), .b(FE_OFN1413_n_8567), .o(TIMEBOOST_net_13396) );
na02s01 TIMEBOOST_cell_2862 ( .a(n_705), .b(pci_target_unit_wishbone_master_rty_counter_0_), .o(TIMEBOOST_net_11) );
in01s01 g62043_u0 ( .a(FE_OFN1299_n_5763), .o(g62043_sb) );
na02s01 TIMEBOOST_cell_39301 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__Q), .b(g65890_sb), .o(TIMEBOOST_net_11889) );
no02f04 TIMEBOOST_cell_22417 ( .a(FE_RN_827_0), .b(TIMEBOOST_net_6465), .o(n_14402) );
na02s01 TIMEBOOST_cell_30857 ( .a(TIMEBOOST_net_9339), .b(g65889_db), .o(n_1860) );
in01s01 g62044_u0 ( .a(FE_OFN1300_n_5763), .o(g62044_sb) );
na03s02 TIMEBOOST_cell_39473 ( .a(TIMEBOOST_net_3953), .b(g64245_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__Q), .o(TIMEBOOST_net_11975) );
na02s02 TIMEBOOST_cell_43371 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__Q), .b(n_4156), .o(TIMEBOOST_net_13924) );
na02s02 TIMEBOOST_cell_16953 ( .a(TIMEBOOST_net_3733), .b(g65219_sb), .o(n_2668) );
in01s01 g62045_u0 ( .a(FE_OFN1302_n_5763), .o(g62045_sb) );
na02s01 TIMEBOOST_cell_2863 ( .a(TIMEBOOST_net_11), .b(pci_target_unit_wishbone_master_reset_rty_cnt), .o(n_8678) );
na03s02 TIMEBOOST_cell_37717 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__Q), .b(FE_OFN704_n_8069), .c(n_2200), .o(TIMEBOOST_net_11097) );
na02s01 TIMEBOOST_cell_2864 ( .a(pci_target_unit_del_sync_comp_done_reg_main), .b(n_1816), .o(TIMEBOOST_net_12) );
in01s01 g62046_u0 ( .a(FE_OFN1299_n_5763), .o(g62046_sb) );
na02s01 TIMEBOOST_cell_18749 ( .a(TIMEBOOST_net_4631), .b(g63032_sb), .o(n_5183) );
na02s02 TIMEBOOST_cell_30917 ( .a(TIMEBOOST_net_9369), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_3727) );
na02s01 TIMEBOOST_cell_43245 ( .a(n_4469), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__Q), .o(TIMEBOOST_net_13861) );
in01s01 g62047_u0 ( .a(FE_OFN1302_n_5763), .o(g62047_sb) );
na02s01 TIMEBOOST_cell_2865 ( .a(TIMEBOOST_net_12), .b(n_1817), .o(n_2468) );
na02s01 TIMEBOOST_cell_18745 ( .a(TIMEBOOST_net_4629), .b(g63028_sb), .o(n_5190) );
na02s01 TIMEBOOST_cell_45062 ( .a(TIMEBOOST_net_14769), .b(FE_OFN531_n_9823), .o(TIMEBOOST_net_11162) );
in01s01 g62048_u0 ( .a(FE_OFN1301_n_5763), .o(g62048_sb) );
na02f02 TIMEBOOST_cell_39004 ( .a(TIMEBOOST_net_11740), .b(g52533_sb), .o(n_13686) );
na03s02 TIMEBOOST_cell_38207 ( .a(TIMEBOOST_net_4071), .b(g64322_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__Q), .o(TIMEBOOST_net_11342) );
na03s02 TIMEBOOST_cell_40303 ( .a(n_4482), .b(g64890_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__Q), .o(TIMEBOOST_net_12390) );
in01s01 g62049_u0 ( .a(FE_OFN1301_n_5763), .o(g62049_sb) );
na02s02 TIMEBOOST_cell_39856 ( .a(TIMEBOOST_net_12166), .b(g62363_sb), .o(n_6875) );
na02s02 TIMEBOOST_cell_38439 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__Q), .b(FE_OFN201_n_9230), .o(TIMEBOOST_net_11458) );
na02s01 TIMEBOOST_cell_38334 ( .a(TIMEBOOST_net_11405), .b(g63088_sb), .o(n_5078) );
in01s01 g62050_u0 ( .a(FE_OFN1301_n_5763), .o(g62050_sb) );
na02s01 TIMEBOOST_cell_18485 ( .a(TIMEBOOST_net_4499), .b(g62740_sb), .o(n_5499) );
na03s02 TIMEBOOST_cell_38429 ( .a(n_3867), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__12__Q), .c(FE_OFN2106_g64577_p), .o(TIMEBOOST_net_11453) );
na02s02 TIMEBOOST_cell_43471 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__Q), .b(n_1852), .o(TIMEBOOST_net_13974) );
in01s01 g62051_u0 ( .a(FE_OFN1299_n_5763), .o(g62051_sb) );
na02s01 TIMEBOOST_cell_18733 ( .a(TIMEBOOST_net_4623), .b(g63084_sb), .o(n_5086) );
na02s01 TIMEBOOST_cell_9342 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(g64197_sb), .o(TIMEBOOST_net_1238) );
in01s01 TIMEBOOST_cell_32855 ( .a(TIMEBOOST_net_10356), .o(TIMEBOOST_net_10355) );
in01s01 g62052_u0 ( .a(FE_OFN1301_n_5763), .o(g62052_sb) );
na02s02 TIMEBOOST_cell_38336 ( .a(TIMEBOOST_net_11406), .b(g63049_sb), .o(n_5153) );
na02s01 TIMEBOOST_cell_19064 ( .a(configuration_pci_err_data_504), .b(wbm_dat_o_3_), .o(TIMEBOOST_net_4789) );
na02s01 TIMEBOOST_cell_38338 ( .a(TIMEBOOST_net_11407), .b(g62837_sb), .o(n_7128) );
in01s01 g62053_u0 ( .a(FE_OFN1302_n_5763), .o(g62053_sb) );
na03s02 TIMEBOOST_cell_42691 ( .a(FE_OFN225_n_9122), .b(g58182_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__Q), .o(TIMEBOOST_net_13584) );
na03s02 TIMEBOOST_cell_37719 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__Q), .b(FE_OFN713_n_8140), .c(n_2187), .o(TIMEBOOST_net_11098) );
na02f02 TIMEBOOST_cell_37805 ( .a(TIMEBOOST_net_9679), .b(g54335_sb), .o(TIMEBOOST_net_11141) );
in01s01 g62054_u0 ( .a(FE_OFN1302_n_5763), .o(g62054_sb) );
na02s01 TIMEBOOST_cell_18577 ( .a(TIMEBOOST_net_4545), .b(g63022_sb), .o(n_5203) );
na02s01 TIMEBOOST_cell_16951 ( .a(TIMEBOOST_net_3732), .b(g65231_sb), .o(n_2656) );
na02s01 TIMEBOOST_cell_42597 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__Q), .b(FE_OFN950_n_2055), .o(TIMEBOOST_net_13537) );
in01s01 g62055_u0 ( .a(FE_OFN1299_n_5763), .o(g62055_sb) );
na02s01 TIMEBOOST_cell_18575 ( .a(TIMEBOOST_net_4544), .b(g63021_sb), .o(n_5205) );
na02s01 TIMEBOOST_cell_30947 ( .a(TIMEBOOST_net_9384), .b(g65086_sb), .o(n_3599) );
na02s02 TIMEBOOST_cell_16949 ( .a(TIMEBOOST_net_3731), .b(g65226_sb), .o(n_2661) );
in01s01 g62056_u0 ( .a(FE_OFN1301_n_5763), .o(g62056_sb) );
na02s01 TIMEBOOST_cell_42712 ( .a(TIMEBOOST_net_13594), .b(g65748_db), .o(n_1606) );
na02s01 TIMEBOOST_cell_19066 ( .a(configuration_pci_err_data_506), .b(wbm_dat_o_5_), .o(TIMEBOOST_net_4790) );
na02f02 TIMEBOOST_cell_42306 ( .a(TIMEBOOST_net_13391), .b(g57431_sb), .o(n_11303) );
in01s01 g62057_u0 ( .a(FE_OFN1302_n_5763), .o(g62057_sb) );
na02f02 TIMEBOOST_cell_44735 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__Q), .b(FE_OFN1583_n_12306), .o(TIMEBOOST_net_14606) );
na02s02 TIMEBOOST_cell_43422 ( .a(TIMEBOOST_net_13949), .b(n_6554), .o(TIMEBOOST_net_12206) );
in01s01 g62058_u0 ( .a(FE_OFN2079_n_8069), .o(g62058_sb) );
na02s02 TIMEBOOST_cell_18753 ( .a(TIMEBOOST_net_4633), .b(g62781_sb), .o(n_5429) );
na02s01 TIMEBOOST_cell_37398 ( .a(TIMEBOOST_net_10937), .b(g61930_sb), .o(n_7963) );
na02s01 TIMEBOOST_cell_38340 ( .a(TIMEBOOST_net_11408), .b(g62801_sb), .o(n_5380) );
in01s01 g62059_u0 ( .a(FE_OFN1299_n_5763), .o(g62059_sb) );
na02s01 TIMEBOOST_cell_45450 ( .a(TIMEBOOST_net_14963), .b(g58634_sb), .o(TIMEBOOST_net_14075) );
na03s02 TIMEBOOST_cell_38217 ( .a(g64191_da), .b(g64191_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q), .o(TIMEBOOST_net_11347) );
na02s10 TIMEBOOST_cell_2880 ( .a(conf_wb_err_addr_in_950), .b(conf_wb_err_addr_in_947), .o(TIMEBOOST_net_20) );
in01s01 g62060_u0 ( .a(FE_OFN1301_n_5763), .o(g62060_sb) );
na02m08 TIMEBOOST_cell_2881 ( .a(n_1165), .b(TIMEBOOST_net_20), .o(n_1972) );
na02s02 TIMEBOOST_cell_43587 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__Q), .b(n_4297), .o(TIMEBOOST_net_14032) );
na02s10 TIMEBOOST_cell_2882 ( .a(wbm_adr_o_3_), .b(wbm_adr_o_4_), .o(TIMEBOOST_net_21) );
in01s01 g62061_u0 ( .a(FE_OFN1300_n_5763), .o(g62061_sb) );
na02m02 TIMEBOOST_cell_44315 ( .a(n_9404), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__Q), .o(TIMEBOOST_net_14396) );
na02s02 TIMEBOOST_cell_3415 ( .a(TIMEBOOST_net_287), .b(FE_OFN215_n_9856), .o(n_9683) );
na02f02 TIMEBOOST_cell_44382 ( .a(TIMEBOOST_net_14429), .b(FE_OFN1400_n_8567), .o(TIMEBOOST_net_12724) );
in01s01 g62062_u0 ( .a(FE_OFN1300_n_5763), .o(g62062_sb) );
na03s02 TIMEBOOST_cell_37723 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__Q), .b(FE_OFN717_n_8176), .c(n_2201), .o(TIMEBOOST_net_11100) );
na02f02 TIMEBOOST_cell_22435 ( .a(TIMEBOOST_net_6474), .b(FE_OFN1752_n_12086), .o(n_12766) );
in01s01 g62063_u0 ( .a(FE_OFN1301_n_5763), .o(g62063_sb) );
na02m06 TIMEBOOST_cell_2883 ( .a(n_562), .b(TIMEBOOST_net_21), .o(n_1477) );
na02f02 TIMEBOOST_cell_44664 ( .a(TIMEBOOST_net_14570), .b(FE_OFN1417_n_8567), .o(TIMEBOOST_net_12790) );
na02s08 TIMEBOOST_cell_2884 ( .a(conf_wb_err_addr_in_955), .b(conf_wb_err_addr_in_954), .o(TIMEBOOST_net_22) );
in01s01 g62064_u0 ( .a(FE_OFN1302_n_5763), .o(g62064_sb) );
na02s02 TIMEBOOST_cell_43552 ( .a(TIMEBOOST_net_14014), .b(FE_OFN1310_n_6624), .o(TIMEBOOST_net_12214) );
na02m02 TIMEBOOST_cell_44383 ( .a(n_9818), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__Q), .o(TIMEBOOST_net_14430) );
na02f02 TIMEBOOST_cell_41654 ( .a(FE_OFN1436_n_9372), .b(TIMEBOOST_net_13065), .o(TIMEBOOST_net_11659) );
in01s01 g62065_u0 ( .a(FE_OFN1301_n_5763), .o(g62065_sb) );
na02m04 TIMEBOOST_cell_2885 ( .a(n_913), .b(TIMEBOOST_net_22), .o(n_2750) );
na02s01 TIMEBOOST_cell_39369 ( .a(TIMEBOOST_net_9578), .b(FE_OFN2113_n_2053), .o(TIMEBOOST_net_11923) );
na02s01 TIMEBOOST_cell_2886 ( .a(wbm_adr_o_29_), .b(wbm_adr_o_30_), .o(TIMEBOOST_net_23) );
in01s01 g62066_u0 ( .a(FE_OFN2079_n_8069), .o(g62066_sb) );
na02m02 TIMEBOOST_cell_10164 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__Q), .b(FE_OFN2059_n_13447), .o(TIMEBOOST_net_1649) );
na02s01 TIMEBOOST_cell_40514 ( .a(TIMEBOOST_net_12495), .b(FE_OFN1300_n_5763), .o(TIMEBOOST_net_11505) );
na02f02 TIMEBOOST_cell_38878 ( .a(TIMEBOOST_net_11677), .b(g58479_sb), .o(n_9358) );
in01m01 g62067_u0 ( .a(FE_OFN1700_n_5751), .o(g62067_sb) );
na02s02 TIMEBOOST_cell_18709 ( .a(TIMEBOOST_net_4611), .b(g63071_sb), .o(n_5108) );
na02f02 TIMEBOOST_cell_42192 ( .a(TIMEBOOST_net_13334), .b(FE_OFN1388_n_8567), .o(TIMEBOOST_net_12286) );
na02m02 TIMEBOOST_cell_42193 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__Q), .b(n_9446), .o(TIMEBOOST_net_13335) );
in01s01 g62068_u0 ( .a(FE_OFN1699_n_5751), .o(g62068_sb) );
na03s02 TIMEBOOST_cell_43311 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__Q), .b(n_3735), .c(FE_OFN1264_n_4095), .o(TIMEBOOST_net_13894) );
na02s01 TIMEBOOST_cell_19032 ( .a(wishbone_slave_unit_pcim_sm_data_in_656), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__Q), .o(TIMEBOOST_net_4773) );
na02s01 TIMEBOOST_cell_44794 ( .a(TIMEBOOST_net_14635), .b(g64819_db), .o(n_3740) );
in01s01 g62069_u0 ( .a(FE_OFN2079_n_8069), .o(g62069_sb) );
na02s02 TIMEBOOST_cell_10166 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__Q), .b(n_13447), .o(TIMEBOOST_net_1650) );
na02f02 TIMEBOOST_cell_42308 ( .a(TIMEBOOST_net_13392), .b(g57216_sb), .o(n_11542) );
na02s02 TIMEBOOST_cell_45451 ( .a(n_826), .b(TIMEBOOST_net_900), .o(TIMEBOOST_net_14964) );
in01s01 g62070_u0 ( .a(FE_OFN2079_n_8069), .o(g62070_sb) );
na02m02 TIMEBOOST_cell_10168 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__Q), .b(n_504), .o(TIMEBOOST_net_1651) );
na02m02 TIMEBOOST_cell_44295 ( .a(n_9661), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__Q), .o(TIMEBOOST_net_14386) );
na02f02 TIMEBOOST_cell_42310 ( .a(TIMEBOOST_net_13393), .b(g57072_sb), .o(n_10497) );
in01s01 g62071_u0 ( .a(FE_OFN2079_n_8069), .o(g62071_sb) );
na02s01 TIMEBOOST_cell_18525 ( .a(TIMEBOOST_net_4519), .b(g62838_sb), .o(n_5298) );
na02s02 TIMEBOOST_cell_45452 ( .a(TIMEBOOST_net_14964), .b(g58635_sb), .o(TIMEBOOST_net_14076) );
na02m02 TIMEBOOST_cell_37747 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__Q), .b(n_13447), .o(TIMEBOOST_net_11112) );
in01s01 g62072_u0 ( .a(n_5633), .o(g62072_sb) );
na02s01 TIMEBOOST_cell_44966 ( .a(TIMEBOOST_net_14721), .b(g58134_db), .o(n_9071) );
na02s01 TIMEBOOST_cell_9144 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__Q), .o(TIMEBOOST_net_1139) );
in01s01 TIMEBOOST_cell_32848 ( .a(TIMEBOOST_net_10349), .o(wbs_dat_i_18_) );
in01s01 g62073_u0 ( .a(FE_OFN1174_n_5592), .o(g62073_sb) );
na02s01 TIMEBOOST_cell_19875 ( .a(TIMEBOOST_net_5194), .b(g62986_sb), .o(n_5910) );
na02s02 TIMEBOOST_cell_39388 ( .a(TIMEBOOST_net_11932), .b(g57996_sb), .o(n_9798) );
na03m02 TIMEBOOST_cell_39409 ( .a(TIMEBOOST_net_505), .b(g63533_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__Q), .o(TIMEBOOST_net_11943) );
in01s01 g62074_u0 ( .a(FE_OFN1170_n_5592), .o(g62074_sb) );
na02s01 TIMEBOOST_cell_38630 ( .a(TIMEBOOST_net_11553), .b(g59113_sb), .o(n_8703) );
na02f02 TIMEBOOST_cell_42312 ( .a(TIMEBOOST_net_13394), .b(g57125_sb), .o(n_11620) );
in01s01 g62075_u0 ( .a(FE_OFN1163_n_5615), .o(g62075_sb) );
na02s02 TIMEBOOST_cell_37558 ( .a(TIMEBOOST_net_11017), .b(g52636_db), .o(n_14755) );
na02s01 TIMEBOOST_cell_38556 ( .a(TIMEBOOST_net_11516), .b(g62050_sb), .o(n_7760) );
na02s02 TIMEBOOST_cell_36748 ( .a(TIMEBOOST_net_10612), .b(FE_OFN1129_g64577_p), .o(TIMEBOOST_net_4510) );
in01s01 g62076_u0 ( .a(FE_OFN1174_n_5592), .o(g62076_sb) );
na02s02 TIMEBOOST_cell_45453 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_1__Q), .b(TIMEBOOST_net_896), .o(TIMEBOOST_net_14965) );
na03s02 TIMEBOOST_cell_38255 ( .a(g64247_da), .b(g64247_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__21__Q), .o(TIMEBOOST_net_11366) );
na02m02 TIMEBOOST_cell_11729 ( .a(TIMEBOOST_net_2431), .b(g62948_sb), .o(n_5985) );
in01s01 g62077_u0 ( .a(n_5633), .o(g62077_sb) );
na02s01 TIMEBOOST_cell_41740 ( .a(TIMEBOOST_net_13108), .b(g65059_db), .o(n_3614) );
na02s01 TIMEBOOST_cell_9146 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__Q), .o(TIMEBOOST_net_1140) );
na02m02 TIMEBOOST_cell_32506 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__Q), .o(TIMEBOOST_net_10164) );
in01s01 g62078_u0 ( .a(n_5633), .o(g62078_sb) );
na02f02 TIMEBOOST_cell_41142 ( .a(TIMEBOOST_net_12809), .b(g57368_sb), .o(n_10381) );
na02s01 TIMEBOOST_cell_17232 ( .a(n_4482), .b(FE_OFN654_n_4508), .o(TIMEBOOST_net_3873) );
na02f02 TIMEBOOST_cell_44384 ( .a(TIMEBOOST_net_14430), .b(FE_OFN1415_n_8567), .o(TIMEBOOST_net_12758) );
in01s01 g62079_u0 ( .a(FE_OFN1163_n_5615), .o(g62079_sb) );
na02s02 TIMEBOOST_cell_36750 ( .a(TIMEBOOST_net_10613), .b(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_4553) );
na02s01 TIMEBOOST_cell_38309 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__Q), .b(g58396_sb), .o(TIMEBOOST_net_11393) );
na02s01 TIMEBOOST_cell_44845 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__Q), .b(g65413_sb), .o(TIMEBOOST_net_14661) );
in01s02 g62080_u0 ( .a(FE_OFN1169_n_5592), .o(g62080_sb) );
na02s02 TIMEBOOST_cell_39390 ( .a(TIMEBOOST_net_11933), .b(FE_OFN272_n_9828), .o(n_9662) );
na02s02 TIMEBOOST_cell_39858 ( .a(TIMEBOOST_net_12167), .b(g62679_sb), .o(n_6181) );
na02s02 TIMEBOOST_cell_39392 ( .a(TIMEBOOST_net_11934), .b(FE_OFN270_n_9836), .o(n_9414) );
in01s01 g62081_u0 ( .a(FE_OFN1169_n_5592), .o(g62081_sb) );
na02s01 TIMEBOOST_cell_39306 ( .a(TIMEBOOST_net_11891), .b(g65836_db), .o(n_1883) );
na02s02 TIMEBOOST_cell_38342 ( .a(TIMEBOOST_net_11409), .b(g62809_sb), .o(n_5361) );
na02s01 TIMEBOOST_cell_44846 ( .a(TIMEBOOST_net_14661), .b(g65413_db), .o(n_3514) );
in01s02 g62082_u0 ( .a(FE_OFN1173_n_5592), .o(g62082_sb) );
na02s01 TIMEBOOST_cell_18705 ( .a(TIMEBOOST_net_4609), .b(g63023_sb), .o(n_5200) );
na02f02 TIMEBOOST_cell_38796 ( .a(TIMEBOOST_net_11636), .b(n_2865), .o(TIMEBOOST_net_6032) );
na02f04 TIMEBOOST_cell_37154 ( .a(n_12962), .b(TIMEBOOST_net_10815), .o(n_13143) );
in01s01 g62083_u0 ( .a(FE_OFN1173_n_5592), .o(g62083_sb) );
na02s01 TIMEBOOST_cell_18569 ( .a(TIMEBOOST_net_4541), .b(g63055_sb), .o(n_5140) );
na02f02 TIMEBOOST_cell_39156 ( .a(n_12250), .b(TIMEBOOST_net_11816), .o(n_12678) );
na02s02 TIMEBOOST_cell_36752 ( .a(TIMEBOOST_net_10614), .b(FE_OFN1128_g64577_p), .o(TIMEBOOST_net_4523) );
in01s01 g62084_u0 ( .a(FE_OFN1165_n_5615), .o(g62084_sb) );
na02s02 TIMEBOOST_cell_18699 ( .a(TIMEBOOST_net_4606), .b(g62759_sb), .o(n_5472) );
na02s02 TIMEBOOST_cell_36754 ( .a(TIMEBOOST_net_10615), .b(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_4684) );
na02m02 TIMEBOOST_cell_39158 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_397), .b(TIMEBOOST_net_11817), .o(TIMEBOOST_net_9631) );
in01s02 g62085_u0 ( .a(FE_OFN1173_n_5592), .o(g62085_sb) );
na02s01 TIMEBOOST_cell_18697 ( .a(TIMEBOOST_net_4605), .b(g62847_sb), .o(n_5277) );
na02s01 TIMEBOOST_cell_36544 ( .a(TIMEBOOST_net_10510), .b(g65741_db), .o(n_1930) );
no02f06 TIMEBOOST_cell_20383 ( .a(TIMEBOOST_net_5448), .b(FE_RN_154_0), .o(n_4699) );
in01s01 g62086_u0 ( .a(FE_OFN1173_n_5592), .o(g62086_sb) );
na02s01 TIMEBOOST_cell_39289 ( .a(pci_target_unit_fifos_pcir_data_in_164), .b(g65771_sb), .o(TIMEBOOST_net_11883) );
na02s01 TIMEBOOST_cell_36545 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__Q), .b(n_4460), .o(TIMEBOOST_net_10511) );
na02s02 TIMEBOOST_cell_36756 ( .a(TIMEBOOST_net_10616), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_4718) );
in01s02 g62087_u0 ( .a(FE_OFN1173_n_5592), .o(g62087_sb) );
na02f02 TIMEBOOST_cell_44736 ( .a(TIMEBOOST_net_14606), .b(n_12024), .o(n_17036) );
na02s02 TIMEBOOST_cell_36758 ( .a(TIMEBOOST_net_10617), .b(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_4616) );
na02s01 TIMEBOOST_cell_36708 ( .a(TIMEBOOST_net_10592), .b(g61904_db), .o(n_8014) );
in01s02 g62088_u0 ( .a(FE_OFN1173_n_5592), .o(g62088_sb) );
na02s01 TIMEBOOST_cell_39291 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(g65735_sb), .o(TIMEBOOST_net_11884) );
na02s02 TIMEBOOST_cell_36710 ( .a(TIMEBOOST_net_10593), .b(g63589_sb), .o(n_4779) );
na02m02 TIMEBOOST_cell_38880 ( .a(TIMEBOOST_net_11678), .b(g58477_sb), .o(n_8979) );
in01s01 g62089_u0 ( .a(FE_OFN1164_n_5615), .o(g62089_sb) );
na03s02 TIMEBOOST_cell_37703 ( .a(n_1877), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__Q), .c(FE_OFN709_n_8232), .o(TIMEBOOST_net_11090) );
na02s01 TIMEBOOST_cell_36276 ( .a(TIMEBOOST_net_10376), .b(FE_OFN988_n_574), .o(n_1647) );
na02s01 TIMEBOOST_cell_36546 ( .a(TIMEBOOST_net_10511), .b(n_4470), .o(TIMEBOOST_net_3566) );
in01s01 g62090_u0 ( .a(n_5633), .o(g62090_sb) );
in01s01 TIMEBOOST_cell_32837 ( .a(TIMEBOOST_net_10338), .o(TIMEBOOST_net_10337) );
na02f02 TIMEBOOST_cell_38917 ( .a(n_3133), .b(wbu_addr_in_264), .o(TIMEBOOST_net_11697) );
in01s01 TIMEBOOST_cell_32836 ( .a(TIMEBOOST_net_10337), .o(wbs_dat_i_24_) );
in01s02 g62091_u0 ( .a(FE_OFN1164_n_5615), .o(g62091_sb) );
na02m02 TIMEBOOST_cell_37560 ( .a(TIMEBOOST_net_11018), .b(g52625_db), .o(n_14681) );
na02s02 TIMEBOOST_cell_38344 ( .a(TIMEBOOST_net_11410), .b(g62788_sb), .o(n_5414) );
na02s02 TIMEBOOST_cell_39308 ( .a(TIMEBOOST_net_11892), .b(g58287_db), .o(n_9516) );
in01s02 g62092_u0 ( .a(FE_OFN1173_n_5592), .o(g62092_sb) );
na03s02 TIMEBOOST_cell_39439 ( .a(g64103_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__Q), .c(FE_OFN877_g64577_p), .o(TIMEBOOST_net_11958) );
na02s02 TIMEBOOST_cell_36548 ( .a(TIMEBOOST_net_10512), .b(g64826_db), .o(n_4455) );
na02s01 TIMEBOOST_cell_36550 ( .a(TIMEBOOST_net_10513), .b(g64755_db), .o(n_4500) );
in01s01 g62093_u0 ( .a(FE_OFN1168_n_5592), .o(g62093_sb) );
na02s01 TIMEBOOST_cell_37403 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__Q), .b(g58442_sb), .o(TIMEBOOST_net_10940) );
na02s02 TIMEBOOST_cell_39860 ( .a(TIMEBOOST_net_12168), .b(g63029_sb), .o(n_5860) );
na02m02 TIMEBOOST_cell_42349 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__Q), .b(n_9875), .o(TIMEBOOST_net_13413) );
in01s01 g62094_u0 ( .a(n_5633), .o(g62094_sb) );
na02s02 TIMEBOOST_cell_43083 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__Q), .b(n_4492), .o(TIMEBOOST_net_13780) );
na02m04 TIMEBOOST_cell_39043 ( .a(wbs_wbb3_2_wbb2_dat_o_i_110), .b(wbs_dat_o_11_), .o(TIMEBOOST_net_11760) );
na02f02 TIMEBOOST_cell_44712 ( .a(TIMEBOOST_net_14594), .b(n_11921), .o(n_12640) );
in01s01 g62095_u0 ( .a(n_5633), .o(g62095_sb) );
na02f02 TIMEBOOST_cell_44660 ( .a(TIMEBOOST_net_14568), .b(FE_OFN2182_n_8567), .o(TIMEBOOST_net_13016) );
na02m02 TIMEBOOST_cell_39347 ( .a(pci_target_unit_pcit_if_strd_addr_in_693), .b(g52652_sb), .o(TIMEBOOST_net_11912) );
na02s01 TIMEBOOST_cell_15824 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_83), .b(FE_OFN2119_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3169) );
in01s01 g62096_u0 ( .a(FE_OFN1168_n_5592), .o(g62096_sb) );
na02s02 TIMEBOOST_cell_37562 ( .a(TIMEBOOST_net_11019), .b(g52639_db), .o(n_14751) );
na02m02 TIMEBOOST_cell_38830 ( .a(TIMEBOOST_net_11653), .b(g58483_sb), .o(n_8973) );
na02s02 TIMEBOOST_cell_37564 ( .a(TIMEBOOST_net_11020), .b(g52638_db), .o(n_14753) );
in01s01 g62097_u0 ( .a(FE_OFN1168_n_5592), .o(g62097_sb) );
na02f02 TIMEBOOST_cell_42350 ( .a(TIMEBOOST_net_13413), .b(FE_OFN2171_n_8567), .o(TIMEBOOST_net_12331) );
in01s01 TIMEBOOST_cell_45927 ( .a(wbm_dat_i_22_), .o(TIMEBOOST_net_15234) );
na02s02 TIMEBOOST_cell_19907 ( .a(TIMEBOOST_net_5210), .b(g63150_sb), .o(n_5840) );
in01s01 g62098_u0 ( .a(FE_OFN1168_n_5592), .o(g62098_sb) );
na02s01 TIMEBOOST_cell_37566 ( .a(TIMEBOOST_net_11021), .b(g65893_db), .o(n_2590) );
na02s01 TIMEBOOST_cell_38346 ( .a(TIMEBOOST_net_11411), .b(g63437_sb), .o(n_4928) );
na02s02 TIMEBOOST_cell_37910 ( .a(TIMEBOOST_net_11193), .b(g58309_sb), .o(n_9501) );
in01s01 g62099_u0 ( .a(FE_OFN1163_n_5615), .o(g62099_sb) );
na02m02 TIMEBOOST_cell_11759 ( .a(TIMEBOOST_net_2446), .b(g62961_sb), .o(n_5960) );
na02s02 TIMEBOOST_cell_44834 ( .a(TIMEBOOST_net_14655), .b(n_4470), .o(TIMEBOOST_net_10908) );
na03m02 TIMEBOOST_cell_41715 ( .a(g58769_sb), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_11__Q), .c(n_8884), .o(TIMEBOOST_net_13096) );
in01s01 g62100_u0 ( .a(FE_OFN1168_n_5592), .o(g62100_sb) );
na02s02 TIMEBOOST_cell_43072 ( .a(TIMEBOOST_net_13774), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_12029) );
na03s02 TIMEBOOST_cell_38327 ( .a(n_3943), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__12__Q), .c(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_11402) );
na02s01 TIMEBOOST_cell_36552 ( .a(TIMEBOOST_net_10514), .b(g64748_db), .o(n_4506) );
in01s01 g62101_u0 ( .a(n_5633), .o(g62101_sb) );
na02s01 TIMEBOOST_cell_16300 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__13__Q), .o(TIMEBOOST_net_3407) );
na02s01 TIMEBOOST_cell_16945 ( .a(TIMEBOOST_net_3729), .b(g65243_sb), .o(n_2639) );
na02m02 TIMEBOOST_cell_44241 ( .a(n_9794), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__Q), .o(TIMEBOOST_net_14359) );
in01s01 g62102_u0 ( .a(FE_OFN1164_n_5615), .o(g62102_sb) );
na02s02 TIMEBOOST_cell_43073 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__Q), .b(n_3688), .o(TIMEBOOST_net_13775) );
na02s02 TIMEBOOST_cell_38674 ( .a(TIMEBOOST_net_11575), .b(g63186_sb), .o(n_5780) );
na02s01 TIMEBOOST_cell_37568 ( .a(TIMEBOOST_net_11022), .b(g58254_sb), .o(n_9042) );
in01s02 g62103_u0 ( .a(FE_OFN1164_n_5615), .o(g62103_sb) );
na02s01 TIMEBOOST_cell_37978 ( .a(TIMEBOOST_net_11227), .b(n_4728), .o(n_7125) );
na03s02 TIMEBOOST_cell_38329 ( .a(n_3929), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__Q), .c(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_11403) );
na02s01 TIMEBOOST_cell_37980 ( .a(TIMEBOOST_net_11228), .b(g54184_db), .o(n_13359) );
in01s01 g62104_u0 ( .a(FE_OFN1163_n_5615), .o(g62104_sb) );
na03m02 TIMEBOOST_cell_34221 ( .a(TIMEBOOST_net_4338), .b(g54158_sb), .c(g53891_db), .o(n_13555) );
na02s02 TIMEBOOST_cell_38676 ( .a(TIMEBOOST_net_11576), .b(g62540_sb), .o(n_6488) );
na02s01 TIMEBOOST_cell_43123 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__Q), .b(n_3628), .o(TIMEBOOST_net_13800) );
in01s01 g62105_u0 ( .a(FE_OFN1174_n_5592), .o(g62105_sb) );
na02s01 TIMEBOOST_cell_37400 ( .a(TIMEBOOST_net_10938), .b(g61741_sb), .o(n_8335) );
na02s02 TIMEBOOST_cell_37746 ( .a(TIMEBOOST_net_11111), .b(FE_OFN2022_n_4778), .o(TIMEBOOST_net_10605) );
na02s01 TIMEBOOST_cell_39296 ( .a(TIMEBOOST_net_11886), .b(g65972_sb), .o(n_2152) );
in01s01 g62106_u0 ( .a(n_5633), .o(g62106_sb) );
na03s02 TIMEBOOST_cell_871 ( .a(n_4612), .b(g61697_sb), .c(g61697_db), .o(n_6980) );
na02s01 TIMEBOOST_cell_17240 ( .a(n_4488), .b(FE_OFN652_n_4508), .o(TIMEBOOST_net_3877) );
in01s01 TIMEBOOST_cell_32844 ( .a(TIMEBOOST_net_10345), .o(wbs_dat_i_25_) );
in01s01 g62107_u0 ( .a(FE_OFN1174_n_5592), .o(g62107_sb) );
na02s01 TIMEBOOST_cell_37402 ( .a(TIMEBOOST_net_10939), .b(g58454_db), .o(n_8990) );
in01s01 TIMEBOOST_cell_45928 ( .a(TIMEBOOST_net_15234), .o(TIMEBOOST_net_15235) );
na02s01 TIMEBOOST_cell_37404 ( .a(TIMEBOOST_net_10940), .b(g58442_db), .o(n_8993) );
in01s01 g62108_u0 ( .a(FE_OFN1174_n_5592), .o(g62108_sb) );
na02s01 TIMEBOOST_cell_37406 ( .a(TIMEBOOST_net_10941), .b(g58336_db), .o(n_9020) );
in01s01 TIMEBOOST_cell_45929 ( .a(wbm_dat_i_23_), .o(TIMEBOOST_net_15236) );
na02s01 TIMEBOOST_cell_37408 ( .a(TIMEBOOST_net_10942), .b(g58451_db), .o(n_8991) );
in01s01 g62109_u0 ( .a(FE_OFN1169_n_5592), .o(g62109_sb) );
na02s01 TIMEBOOST_cell_37410 ( .a(TIMEBOOST_net_10943), .b(g65788_db), .o(n_1597) );
na02f02 TIMEBOOST_cell_37748 ( .a(TIMEBOOST_net_11112), .b(FE_OFN1148_n_13249), .o(TIMEBOOST_net_4414) );
na02s01 TIMEBOOST_cell_37412 ( .a(TIMEBOOST_net_10944), .b(g65211_db), .o(n_2677) );
in01s01 g62110_u0 ( .a(FE_OFN1165_n_5615), .o(g62110_sb) );
na02f02 TIMEBOOST_cell_39115 ( .a(TIMEBOOST_net_10160), .b(FE_OFN1606_n_13997), .o(TIMEBOOST_net_11796) );
na02s02 TIMEBOOST_cell_36554 ( .a(TIMEBOOST_net_10515), .b(g58391_db), .o(n_9441) );
na02s01 TIMEBOOST_cell_36556 ( .a(TIMEBOOST_net_10516), .b(g64786_db), .o(n_3765) );
in01s01 g62111_u0 ( .a(n_5633), .o(g62111_sb) );
na03s02 TIMEBOOST_cell_34259 ( .a(TIMEBOOST_net_9816), .b(FE_OFN1174_n_5592), .c(g62076_sb), .o(n_5635) );
na02s01 g62111_u2 ( .a(configuration_wb_err_addr_542), .b(n_5633), .o(g62111_db) );
na02s01 TIMEBOOST_cell_38348 ( .a(TIMEBOOST_net_11412), .b(g63169_sb), .o(n_4955) );
in01s01 g62112_u0 ( .a(FE_OFN1171_n_5592), .o(g62112_sb) );
na02s01 TIMEBOOST_cell_37414 ( .a(TIMEBOOST_net_10945), .b(g65225_db), .o(n_2662) );
na02s01 TIMEBOOST_cell_37416 ( .a(TIMEBOOST_net_10946), .b(g65786_sb), .o(n_1598) );
in01s01 g62113_u0 ( .a(FE_OFN1170_n_5592), .o(g62113_sb) );
na02s01 TIMEBOOST_cell_42767 ( .a(TIMEBOOST_net_3895), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__Q), .o(TIMEBOOST_net_13622) );
na02s01 TIMEBOOST_cell_38558 ( .a(TIMEBOOST_net_11517), .b(g62035_sb), .o(n_7781) );
na02m02 TIMEBOOST_cell_37252 ( .a(TIMEBOOST_net_10864), .b(g58778_sb), .o(n_9884) );
in01s01 g62114_u0 ( .a(n_5633), .o(g62114_sb) );
in01s01 TIMEBOOST_cell_32843 ( .a(TIMEBOOST_net_10344), .o(TIMEBOOST_net_10343) );
na02s01 g62114_u2 ( .a(configuration_wb_err_addr_545), .b(n_5633), .o(g62114_db) );
na03s02 TIMEBOOST_cell_876 ( .a(n_4072), .b(g62811_sb), .c(g62811_db), .o(n_5356) );
in01s01 g62115_u0 ( .a(FE_OFN1166_n_5615), .o(g62115_sb) );
na02s01 TIMEBOOST_cell_16065 ( .a(TIMEBOOST_net_3289), .b(g65860_db), .o(n_1579) );
na02s01 TIMEBOOST_cell_36558 ( .a(TIMEBOOST_net_10517), .b(g64171_db), .o(n_3994) );
na02f02 TIMEBOOST_cell_41677 ( .a(n_14895), .b(n_13484), .o(TIMEBOOST_net_13077) );
in01s01 g62116_u0 ( .a(n_5633), .o(g62116_sb) );
na03s02 TIMEBOOST_cell_877 ( .a(n_3949), .b(g62859_sb), .c(g62859_db), .o(n_5248) );
na02s01 g62116_u2 ( .a(configuration_wb_err_addr_547), .b(n_5633), .o(g62116_db) );
na02m02 TIMEBOOST_cell_44271 ( .a(n_9206), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__Q), .o(TIMEBOOST_net_14374) );
in01s01 g62117_u0 ( .a(FE_OFN1166_n_5615), .o(g62117_sb) );
na02s01 TIMEBOOST_cell_36560 ( .a(TIMEBOOST_net_10518), .b(g65312_sb), .o(n_3568) );
na02s01 TIMEBOOST_cell_36562 ( .a(TIMEBOOST_net_10519), .b(g64160_db), .o(n_4005) );
in01s01 g62118_u0 ( .a(FE_OFN1171_n_5592), .o(g62118_sb) );
na02s01 TIMEBOOST_cell_36564 ( .a(TIMEBOOST_net_10520), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_3650) );
na02s01 TIMEBOOST_cell_36566 ( .a(TIMEBOOST_net_10521), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_3648) );
in01s01 g62119_u0 ( .a(n_5633), .o(g62119_sb) );
na03s02 TIMEBOOST_cell_6552 ( .a(n_4645), .b(g64873_sb), .c(g64873_db), .o(n_4422) );
na02s01 g62119_u2 ( .a(configuration_wb_err_addr_550), .b(n_5633), .o(g62119_db) );
na02f08 TIMEBOOST_cell_44781 ( .a(n_1519), .b(n_763), .o(TIMEBOOST_net_14629) );
in01s01 g62120_u0 ( .a(FE_OFN1170_n_5592), .o(g62120_sb) );
na03s02 TIMEBOOST_cell_37709 ( .a(n_1907), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__Q), .c(FE_OFN716_n_8176), .o(TIMEBOOST_net_11093) );
na02s01 TIMEBOOST_cell_36568 ( .a(TIMEBOOST_net_10522), .b(g58402_sb), .o(TIMEBOOST_net_9568) );
na02s01 TIMEBOOST_cell_36570 ( .a(TIMEBOOST_net_10523), .b(g65822_db), .o(n_1894) );
in01s01 g62121_u0 ( .a(FE_OFN1171_n_5592), .o(g62121_sb) );
na02s02 TIMEBOOST_cell_37570 ( .a(TIMEBOOST_net_11023), .b(g58242_sb), .o(n_9549) );
na02m02 TIMEBOOST_cell_44175 ( .a(n_8991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__Q), .o(TIMEBOOST_net_14326) );
na02s02 TIMEBOOST_cell_39408 ( .a(TIMEBOOST_net_11942), .b(FE_OFN270_n_9836), .o(n_9569) );
in01s01 g62122_u0 ( .a(FE_OFN1172_n_5592), .o(g62122_sb) );
in01s01 TIMEBOOST_cell_45906 ( .a(TIMEBOOST_net_15212), .o(TIMEBOOST_net_15213) );
na02s02 TIMEBOOST_cell_37750 ( .a(TIMEBOOST_net_11113), .b(FE_OFN2022_n_4778), .o(TIMEBOOST_net_10601) );
na02s02 TIMEBOOST_cell_38750 ( .a(TIMEBOOST_net_11613), .b(g53901_sb), .o(n_13540) );
in01s01 g62123_u0 ( .a(FE_OFN1171_n_5592), .o(g62123_sb) );
na03s02 TIMEBOOST_cell_37711 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__Q), .b(FE_OFN2084_n_8407), .c(n_1604), .o(TIMEBOOST_net_11094) );
na02s01 TIMEBOOST_cell_36572 ( .a(TIMEBOOST_net_10524), .b(g64224_db), .o(n_4518) );
na02s01 TIMEBOOST_cell_36574 ( .a(TIMEBOOST_net_10525), .b(g65954_db), .o(n_1844) );
in01s01 g62124_u0 ( .a(n_5633), .o(g62124_sb) );
na02s01 TIMEBOOST_cell_39258 ( .a(TIMEBOOST_net_11867), .b(g64130_db), .o(n_4032) );
na02m04 TIMEBOOST_cell_39045 ( .a(wbs_wbb3_2_wbb2_dat_o_i_109), .b(wbs_dat_o_10_), .o(TIMEBOOST_net_11761) );
na02f08 TIMEBOOST_cell_44782 ( .a(TIMEBOOST_net_14629), .b(n_16539), .o(n_16540) );
in01s01 g62125_u0 ( .a(FE_OFN1170_n_5592), .o(g62125_sb) );
na02f02 TIMEBOOST_cell_39119 ( .a(TIMEBOOST_net_10171), .b(FE_OCPN2219_n_13997), .o(TIMEBOOST_net_11798) );
na02s01 TIMEBOOST_cell_36576 ( .a(TIMEBOOST_net_10526), .b(g65230_db), .o(n_2657) );
na02s01 TIMEBOOST_cell_36578 ( .a(TIMEBOOST_net_10527), .b(g60603_sb), .o(TIMEBOOST_net_9837) );
in01s01 g62126_u0 ( .a(FE_OFN1170_n_5592), .o(g62126_sb) );
na02s01 TIMEBOOST_cell_18553 ( .a(TIMEBOOST_net_4533), .b(g63037_sb), .o(n_5174) );
na02s01 TIMEBOOST_cell_36580 ( .a(TIMEBOOST_net_10528), .b(g62008_db), .o(n_7879) );
na02f02 TIMEBOOST_cell_41678 ( .a(TIMEBOOST_net_13077), .b(n_14829), .o(n_14893) );
in01s01 g62127_u0 ( .a(FE_OFN1172_n_5592), .o(g62127_sb) );
na02f02 TIMEBOOST_cell_41679 ( .a(n_14895), .b(n_13488), .o(TIMEBOOST_net_13078) );
na02f02 TIMEBOOST_cell_39147 ( .a(FE_OFN1552_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__Q), .o(TIMEBOOST_net_11812) );
na02m02 TIMEBOOST_cell_11821 ( .a(TIMEBOOST_net_2477), .b(g62599_sb), .o(n_6353) );
in01s01 g62128_u0 ( .a(FE_OFN1171_n_5592), .o(g62128_sb) );
na02s02 TIMEBOOST_cell_37870 ( .a(TIMEBOOST_net_11173), .b(g58032_sb), .o(n_9754) );
na02s02 TIMEBOOST_cell_43588 ( .a(TIMEBOOST_net_14032), .b(FE_OFN1285_n_4097), .o(TIMEBOOST_net_12047) );
na02s02 TIMEBOOST_cell_37872 ( .a(TIMEBOOST_net_11174), .b(g58178_sb), .o(n_9610) );
in01s01 g62129_u0 ( .a(FE_OFN1166_n_5615), .o(g62129_sb) );
na02s02 TIMEBOOST_cell_18631 ( .a(TIMEBOOST_net_4572), .b(g63082_sb), .o(n_7119) );
na02s02 TIMEBOOST_cell_36582 ( .a(TIMEBOOST_net_10529), .b(n_16748), .o(TIMEBOOST_net_4178) );
na02s01 TIMEBOOST_cell_36584 ( .a(TIMEBOOST_net_10530), .b(g63586_sb), .o(n_4101) );
in01s01 g62130_u0 ( .a(FE_OFN1171_n_5592), .o(g62130_sb) );
na02s02 TIMEBOOST_cell_37874 ( .a(TIMEBOOST_net_11175), .b(g57961_sb), .o(n_9843) );
na02m02 TIMEBOOST_cell_43589 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__Q), .b(n_3705), .o(TIMEBOOST_net_14033) );
na02s01 TIMEBOOST_cell_37860 ( .a(TIMEBOOST_net_11168), .b(g58280_sb), .o(n_9522) );
in01s01 g62131_u0 ( .a(FE_OFN1171_n_5592), .o(g62131_sb) );
na02f02 TIMEBOOST_cell_36920 ( .a(TIMEBOOST_net_10698), .b(g52598_sb), .o(n_10275) );
na02s01 TIMEBOOST_cell_39337 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q), .b(g64234_sb), .o(TIMEBOOST_net_11907) );
na02s01 TIMEBOOST_cell_36444 ( .a(TIMEBOOST_net_10460), .b(g64199_db), .o(n_3970) );
in01s01 g62132_u0 ( .a(n_5633), .o(g62132_sb) );
na02s01 TIMEBOOST_cell_43066 ( .a(TIMEBOOST_net_13771), .b(FE_OFN1293_n_4098), .o(TIMEBOOST_net_12024) );
na02s01 TIMEBOOST_cell_17244 ( .a(n_4444), .b(FE_OFN652_n_4508), .o(TIMEBOOST_net_3879) );
na02s01 TIMEBOOST_cell_37992 ( .a(TIMEBOOST_net_11234), .b(TIMEBOOST_net_9714), .o(n_5084) );
in01s01 g62133_u0 ( .a(n_5633), .o(g62133_sb) );
na02s02 TIMEBOOST_cell_38350 ( .a(TIMEBOOST_net_11413), .b(g63392_sb), .o(n_4134) );
na02s01 TIMEBOOST_cell_17246 ( .a(n_4470), .b(FE_OFN651_n_4508), .o(TIMEBOOST_net_3880) );
na02s02 TIMEBOOST_cell_37886 ( .a(TIMEBOOST_net_11181), .b(g58192_sb), .o(n_9592) );
in01s01 g62134_u0 ( .a(n_5633), .o(g62134_sb) );
in01s01 TIMEBOOST_cell_32842 ( .a(TIMEBOOST_net_10343), .o(wbs_dat_i_2_) );
na02s01 TIMEBOOST_cell_39195 ( .a(TIMEBOOST_net_3334), .b(FE_OFN1003_n_2047), .o(TIMEBOOST_net_11836) );
na02s01 TIMEBOOST_cell_30864 ( .a(pci_target_unit_pcit_if_strd_addr_in_690), .b(n_2544), .o(TIMEBOOST_net_9343) );
in01s01 g62135_u0 ( .a(FE_OFN1166_n_5615), .o(g62135_sb) );
na02s01 TIMEBOOST_cell_18551 ( .a(TIMEBOOST_net_4532), .b(g63030_sb), .o(n_5188) );
na02s01 TIMEBOOST_cell_36586 ( .a(TIMEBOOST_net_10531), .b(g63586_sb), .o(n_4102) );
na02s01 TIMEBOOST_cell_36588 ( .a(TIMEBOOST_net_10532), .b(g63584_sb), .o(n_4104) );
in01s01 g62136_u0 ( .a(FE_OFN1171_n_5592), .o(g62136_sb) );
na03s02 TIMEBOOST_cell_37773 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__Q), .b(FE_OFN709_n_8232), .c(n_1580), .o(TIMEBOOST_net_11125) );
na02s01 TIMEBOOST_cell_36590 ( .a(TIMEBOOST_net_10533), .b(g63584_sb), .o(n_4103) );
na02s01 TIMEBOOST_cell_36592 ( .a(TIMEBOOST_net_10534), .b(g63582_db), .o(n_4106) );
in01s01 g62137_u0 ( .a(FE_OFN1171_n_5592), .o(g62137_sb) );
na02s01 TIMEBOOST_cell_36446 ( .a(TIMEBOOST_net_10461), .b(g65778_db), .o(n_1600) );
na02f02 TIMEBOOST_cell_38832 ( .a(TIMEBOOST_net_11654), .b(g58455_sb), .o(n_9402) );
na02s01 TIMEBOOST_cell_36448 ( .a(TIMEBOOST_net_10462), .b(g65795_db), .o(n_1592) );
in01s01 g62138_u0 ( .a(FE_OFN1170_n_5592), .o(g62138_sb) );
na03s02 TIMEBOOST_cell_37775 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__Q), .b(FE_OFN2081_n_8176), .c(n_1564), .o(TIMEBOOST_net_11126) );
no02f04 TIMEBOOST_cell_36594 ( .a(TIMEBOOST_net_10535), .b(FE_RN_151_0), .o(n_2939) );
na02s01 TIMEBOOST_cell_36596 ( .a(TIMEBOOST_net_10536), .b(TIMEBOOST_net_4052), .o(n_4105) );
in01s01 g62139_u0 ( .a(FE_OFN1171_n_5592), .o(g62139_sb) );
na02s01 TIMEBOOST_cell_37862 ( .a(TIMEBOOST_net_11169), .b(g58273_sb), .o(n_9527) );
na02m02 TIMEBOOST_cell_43590 ( .a(TIMEBOOST_net_14033), .b(FE_OFN1323_n_6436), .o(TIMEBOOST_net_12248) );
na02s02 TIMEBOOST_cell_37864 ( .a(TIMEBOOST_net_11170), .b(g58394_sb), .o(n_9439) );
in01s01 g62140_u0 ( .a(FE_OFN1166_n_5615), .o(g62140_sb) );
na03f02 TIMEBOOST_cell_21816 ( .a(n_3062), .b(n_2913), .c(n_2836), .o(TIMEBOOST_net_6165) );
na02s02 TIMEBOOST_cell_36598 ( .a(TIMEBOOST_net_10537), .b(FE_OFN2079_n_8069), .o(TIMEBOOST_net_4115) );
na02s02 TIMEBOOST_cell_36600 ( .a(TIMEBOOST_net_10538), .b(n_3126), .o(TIMEBOOST_net_4079) );
in01s01 g62141_u0 ( .a(FE_OFN1174_n_5592), .o(g62141_sb) );
na02s02 g52441_u2 ( .a(n_14680), .b(n_14839), .o(g52441_db) );
na02f02 TIMEBOOST_cell_39153 ( .a(n_12313), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__Q), .o(TIMEBOOST_net_11815) );
na02s02 TIMEBOOST_cell_37856 ( .a(TIMEBOOST_net_11166), .b(g57957_sb), .o(n_9848) );
in01m01 g62143_u0 ( .a(n_2035), .o(n_2281) );
in01s01 g62144_u0 ( .a(n_1694), .o(n_1695) );
in01s01 g62145_u0 ( .a(n_1692), .o(n_1693) );
na02m06 g62193_u0 ( .a(n_15931), .b(n_1698), .o(n_7427) );
na02f06 g62194_u0 ( .a(n_15931), .b(n_2044), .o(n_7420) );
na02f08 g62195_u0 ( .a(n_15931), .b(n_1061), .o(n_7410) );
na02f02 g62196_u0 ( .a(n_7466), .b(FE_OCPN1854_n_2071), .o(n_7437) );
oa12s02 g62197_u0 ( .a(configuration_wb_err_cs_bit8), .b(n_3282), .c(n_8440), .o(n_7743) );
na02m08 g62198_u0 ( .a(FE_OFN1158_n_15325), .b(n_1061), .o(n_7015) );
na02m02 g62199_u0 ( .a(n_7809), .b(FE_OCPN1854_n_2071), .o(n_7810) );
na02f02 g62200_u0 ( .a(n_7803), .b(FE_OCPN1854_n_2071), .o(n_7804) );
oa12s02 g62201_u0 ( .a(configuration_isr_bit_2975), .b(n_3800), .c(n_8440), .o(n_7742) );
na02s08 g62202_u0 ( .a(n_7466), .b(n_1698), .o(n_7467) );
oa12s02 g62203_u0 ( .a(configuration_status_bit8), .b(n_3257), .c(n_8440), .o(n_7740) );
oa12s01 g62204_u0 ( .a(configuration_status_bit_322), .b(n_3256), .c(n_8440), .o(n_7739) );
na02f08 g62205_u0 ( .a(n_16916), .b(n_1698), .o(n_7283) );
na02f06 g62207_u0 ( .a(n_16916), .b(n_2044), .o(n_7273) );
na02s08 g62208_u0 ( .a(FE_OFN1159_n_15325), .b(n_1698), .o(n_7012) );
na02s08 g62209_u0 ( .a(FE_OFN1159_n_15325), .b(n_2044), .o(n_7007) );
na02f08 g62210_u0 ( .a(n_16916), .b(n_1061), .o(n_7293) );
oa12s02 g62211_u0 ( .a(configuration_status_bit_435), .b(n_3255), .c(n_8440), .o(n_7738) );
oa12s02 g62212_u0 ( .a(configuration_status_bit_379), .b(n_3258), .c(n_8440), .o(n_7737) );
oa12s02 g62213_u0 ( .a(configuration_status_bit_351), .b(n_3262), .c(n_8440), .o(n_7735) );
oa12s02 g62214_u0 ( .a(configuration_status_bit_407), .b(n_3254), .c(n_8440), .o(n_7734) );
na02f02 g62215_u0 ( .a(n_7795), .b(FE_OCPN1854_n_2071), .o(n_7796) );
no02f06 g62217_u0 ( .a(n_4686), .b(n_4685), .o(n_4853) );
in01f01 g62218_u0 ( .a(n_4815), .o(n_4816) );
no02f04 g62219_u0 ( .a(n_2708), .b(n_4685), .o(g62219_p) );
in01f04 g62219_u1 ( .a(g62219_p), .o(n_4815) );
na02f04 g62220_u0 ( .a(n_1390), .b(n_2680), .o(g62220_p) );
in01f04 g62220_u1 ( .a(g62220_p), .o(n_2970) );
na02m02 g62221_u0 ( .a(n_2738), .b(n_2463), .o(g62221_p) );
in01m02 g62221_u1 ( .a(g62221_p), .o(n_2873) );
na02f01 g62222_u0 ( .a(FE_OCP_RBN2222_n_15347), .b(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(n_6944) );
na02f02 g62223_u0 ( .a(wishbone_slave_unit_wishbone_slave_do_del_request), .b(FE_OCP_RBN2220_n_15347), .o(g62223_p) );
in01f02 g62223_u1 ( .a(g62223_p), .o(n_4814) );
in01s01 TIMEBOOST_cell_32835 ( .a(TIMEBOOST_net_10336), .o(TIMEBOOST_net_10335) );
na02s02 g62225_u0 ( .a(FE_OFN1169_n_5592), .b(configuration_wb_err_cs_bit9), .o(n_4813) );
na02s02 TIMEBOOST_cell_40418 ( .a(TIMEBOOST_net_12447), .b(FE_OFN272_n_9828), .o(n_9704) );
na02f03 g62254_u0 ( .a(n_3342), .b(n_3341), .o(g62254_p) );
in01f03 g62254_u1 ( .a(g62254_p), .o(n_3476) );
oa12f02 g62258_u0 ( .a(n_4123), .b(n_2972), .c(n_2127), .o(n_4812) );
na02s02 g62259_u0 ( .a(FE_OFN2079_n_8069), .b(n_8876), .o(n_7733) );
no02s02 g62260_u0 ( .a(n_2721), .b(FE_OFN778_n_4152), .o(n_3162) );
ao12s01 g62261_u0 ( .a(configuration_sync_pci_err_cs_8_del_bit_reg_Q), .b(n_4721), .c(n_4743), .o(n_7574) );
na02m02 g62262_u0 ( .a(n_3436), .b(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(n_7078) );
na02s02 g62263_u0 ( .a(FE_OFN2079_n_8069), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_), .o(n_7731) );
na02m02 g62264_u0 ( .a(n_2461), .b(n_2680), .o(g62264_p) );
in01f02 g62264_u1 ( .a(g62264_p), .o(n_2462) );
na02s02 g62265_u0 ( .a(FE_OFN1171_n_5592), .b(configuration_wb_err_addr), .o(n_4811) );
no02m06 g62267_u0 ( .a(n_7398), .b(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(n_7725) );
na02f06 TIMEBOOST_cell_41934 ( .a(g54237_sb), .b(TIMEBOOST_net_13205), .o(n_13651) );
na02m02 g62273_u0 ( .a(n_1111), .b(n_13825), .o(n_6942) );
na02s02 g62274_u0 ( .a(wishbone_slave_unit_pcim_sm_be_in_558), .b(n_13825), .o(n_6941) );
na02m02 g62275_u0 ( .a(wishbone_slave_unit_pcim_sm_be_in_559), .b(n_13825), .o(n_6940) );
in01m01 g62277_u0 ( .a(n_2460), .o(n_2735) );
no02m04 g62278_u0 ( .a(n_2011), .b(n_1639), .o(n_2460) );
no02f02 g62279_u0 ( .a(n_2940), .b(FE_OFN1142_n_15261), .o(n_3339) );
na02s02 TIMEBOOST_cell_45223 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__Q), .b(n_4279), .o(TIMEBOOST_net_14850) );
no02m02 g62281_u0 ( .a(FE_OFN1144_n_15261), .b(n_2941), .o(n_3338) );
no02m02 g62282_u0 ( .a(n_3136), .b(FE_OFN1145_n_15261), .o(n_3468) );
ao12s01 g62283_u0 ( .a(configuration_sync_isr_2_del_bit_reg_Q), .b(n_3799), .c(n_4743), .o(n_7571) );
na02s01 TIMEBOOST_cell_38352 ( .a(TIMEBOOST_net_11414), .b(g63017_sb), .o(n_5214) );
na02m02 g62285_u0 ( .a(n_3160), .b(wishbone_slave_unit_pcim_if_del_we_in), .o(g62285_p) );
in01m02 g62285_u1 ( .a(g62285_p), .o(n_3391) );
no02m01 g62286_u0 ( .a(FE_OFN1172_n_5592), .b(n_16763), .o(n_4809) );
na03s01 TIMEBOOST_cell_34153 ( .a(n_4011), .b(g62807_sb), .c(g62807_db), .o(n_5366) );
no02s02 g62288_u0 ( .a(n_2943), .b(n_692), .o(n_3337) );
no02f01 g62289_u0 ( .a(n_16163), .b(pci_target_unit_wishbone_master_retried), .o(TIMEBOOST_net_3148) );
no02s02 g62290_u0 ( .a(n_2010), .b(FE_OFN778_n_4152), .o(n_2980) );
na02s02 TIMEBOOST_cell_39862 ( .a(TIMEBOOST_net_12169), .b(g62614_sb), .o(n_6329) );
na02s01 g62293_u0 ( .a(n_7350), .b(n_7569), .o(n_8503) );
na02f08 g62294_u0 ( .a(n_15920), .b(n_15347), .o(n_15014) );
in01s01 TIMEBOOST_cell_45875 ( .a(n_7174), .o(TIMEBOOST_net_15182) );
na02f02 TIMEBOOST_cell_42314 ( .a(TIMEBOOST_net_13395), .b(g57502_sb), .o(n_10327) );
na02m02 TIMEBOOST_cell_45454 ( .a(TIMEBOOST_net_14965), .b(g58631_sb), .o(TIMEBOOST_net_14077) );
na02f02 TIMEBOOST_cell_42316 ( .a(TIMEBOOST_net_13396), .b(g57441_sb), .o(n_11295) );
na02s02 TIMEBOOST_cell_45455 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_0__Q), .b(TIMEBOOST_net_895), .o(TIMEBOOST_net_14966) );
na02s02 TIMEBOOST_cell_41702 ( .a(TIMEBOOST_net_13089), .b(n_8832), .o(n_9228) );
na02f04 TIMEBOOST_cell_44779 ( .a(n_16388), .b(n_16393), .o(TIMEBOOST_net_14628) );
na02f02 TIMEBOOST_cell_22345 ( .a(TIMEBOOST_net_6429), .b(n_10641), .o(n_12147) );
na02f02 TIMEBOOST_cell_44267 ( .a(n_9659), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__Q), .o(TIMEBOOST_net_14372) );
na02s01 TIMEBOOST_cell_44870 ( .a(TIMEBOOST_net_14673), .b(g58315_sb), .o(TIMEBOOST_net_12443) );
na02s01 TIMEBOOST_cell_44783 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__Q), .b(FE_OFN575_n_9902), .o(TIMEBOOST_net_14630) );
na02f02 TIMEBOOST_cell_44248 ( .a(TIMEBOOST_net_14362), .b(FE_OFN1373_n_8567), .o(TIMEBOOST_net_13403) );
na02s01 TIMEBOOST_cell_30918 ( .a(pci_target_unit_pcit_if_strd_addr_in), .b(n_2671), .o(TIMEBOOST_net_9370) );
na02f02 TIMEBOOST_cell_42318 ( .a(TIMEBOOST_net_13397), .b(g57564_sb), .o(n_10297) );
na02s01 TIMEBOOST_cell_42960 ( .a(TIMEBOOST_net_13718), .b(g61898_db), .o(n_8030) );
na02f02 g62312_u0 ( .a(n_1970), .b(n_2738), .o(g62312_p) );
in01m02 g62312_u1 ( .a(g62312_p), .o(n_2456) );
na03f02 TIMEBOOST_cell_22346 ( .a(n_10057), .b(n_9270), .c(n_9269), .o(TIMEBOOST_net_6430) );
ao22f02 g62314_u0 ( .a(n_2264), .b(n_2727), .c(n_2711), .d(n_2430), .o(n_4197) );
oa12s01 g62316_u0 ( .a(n_5545), .b(n_5546), .c(pci_target_unit_fifos_pciw_inTransactionCount_1_), .o(n_5548) );
oa12s01 g62317_u0 ( .a(n_5545), .b(pci_target_unit_fifos_inGreyCount_0_), .c(n_5546), .o(n_5547) );
no02m02 g62318_u0 ( .a(n_1557), .b(n_4680), .o(g62318_p) );
in01m02 g62318_u1 ( .a(g62318_p), .o(n_4681) );
na02m01 g62319_u0 ( .a(n_3450), .b(n_4718), .o(g62319_p) );
in01s01 g62319_u1 ( .a(g62319_p), .o(n_4679) );
ao12f02 g62320_u0 ( .a(n_2956), .b(n_1445), .c(FE_OCP_RBN2239_g74749_p), .o(n_4165) );
ao12s01 g62321_u0 ( .a(n_3157), .b(n_1335), .c(wbm_rty_i), .o(n_3159) );
ao12s01 g62322_u0 ( .a(n_1714), .b(n_1226), .c(wishbone_slave_unit_pci_initiator_sm_latency_timer_3_), .o(n_2034) );
na02s01 TIMEBOOST_cell_37269 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(g65675_sb), .o(TIMEBOOST_net_10873) );
oa12s01 g62325_u0 ( .a(n_7136), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_0_), .c(FE_OFN1192_n_6935), .o(n_7137) );
in01s01 g62326_u0 ( .a(FE_OFN1192_n_6935), .o(g62326_sb) );
na02s02 TIMEBOOST_cell_3045 ( .a(TIMEBOOST_net_102), .b(n_2236), .o(n_2706) );
na02s01 g62326_u2 ( .a(n_1510), .b(FE_OFN1192_n_6935), .o(g62326_db) );
na03f02 TIMEBOOST_cell_36093 ( .a(n_12224), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__Q), .c(n_12010), .o(n_12652) );
ao12m01 g62327_u0 ( .a(n_3157), .b(n_2291), .c(wbm_rty_i), .o(n_3158) );
ao12m01 g62328_u0 ( .a(n_3157), .b(n_2396), .c(wbm_rty_i), .o(n_3156) );
ao12f01 g62329_u0 ( .a(n_1808), .b(n_4675), .c(n_4674), .o(n_4896) );
in01m01 g62330_u0 ( .a(n_7400), .o(n_7135) );
no02m02 g62331_u0 ( .a(n_4793), .b(n_3811), .o(n_7400) );
oa12f02 g62332_u0 ( .a(n_1099), .b(n_2728), .c(n_2959), .o(n_3333) );
in01s01 g62333_u0 ( .a(FE_OFN1269_n_4095), .o(g62333_sb) );
na02f02 TIMEBOOST_cell_44176 ( .a(TIMEBOOST_net_14326), .b(FE_OFN1370_n_8567), .o(TIMEBOOST_net_13397) );
na02f02 TIMEBOOST_cell_42194 ( .a(TIMEBOOST_net_13335), .b(FE_OFN1388_n_8567), .o(TIMEBOOST_net_12289) );
na02m02 TIMEBOOST_cell_42195 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__Q), .b(n_9598), .o(TIMEBOOST_net_13336) );
in01s01 g62334_u0 ( .a(FE_OFN1269_n_4095), .o(g62334_sb) );
na02s01 TIMEBOOST_cell_37243 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__Q), .b(n_3755), .o(TIMEBOOST_net_10860) );
na02s01 TIMEBOOST_cell_43312 ( .a(TIMEBOOST_net_13894), .b(g62684_sb), .o(n_6171) );
na02m02 TIMEBOOST_cell_43579 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__Q), .b(n_4246), .o(TIMEBOOST_net_14028) );
in01s01 g62335_u0 ( .a(FE_OFN1275_n_4096), .o(g62335_sb) );
na02m04 TIMEBOOST_cell_3047 ( .a(n_2229), .b(TIMEBOOST_net_103), .o(n_2230) );
na03s02 TIMEBOOST_cell_37777 ( .a(g65869_da), .b(g65869_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__Q), .o(TIMEBOOST_net_11127) );
na02s06 TIMEBOOST_cell_3048 ( .a(n_1824), .b(n_373), .o(TIMEBOOST_net_104) );
in01s01 g62336_u0 ( .a(FE_OFN1257_n_4143), .o(g62336_sb) );
na02s01 TIMEBOOST_cell_37245 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__Q), .b(n_3749), .o(TIMEBOOST_net_10861) );
na02f02 TIMEBOOST_cell_43716 ( .a(TIMEBOOST_net_14096), .b(g57421_sb), .o(n_11316) );
na03s02 TIMEBOOST_cell_43313 ( .a(n_4673), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__Q), .c(g62942_sb), .o(TIMEBOOST_net_13895) );
in01s01 g62337_u0 ( .a(FE_OFN1231_n_6391), .o(g62337_sb) );
na02s02 TIMEBOOST_cell_3581 ( .a(TIMEBOOST_net_370), .b(FE_OFN262_n_9851), .o(n_9647) );
na03f04 TIMEBOOST_cell_37149 ( .a(n_11818), .b(n_11956), .c(n_11957), .o(TIMEBOOST_net_10813) );
na02s01 TIMEBOOST_cell_15793 ( .a(TIMEBOOST_net_3153), .b(g67042_sb), .o(n_1272) );
in01s01 g62338_u0 ( .a(FE_OFN1231_n_6391), .o(g62338_sb) );
na02m02 TIMEBOOST_cell_43973 ( .a(n_9826), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__Q), .o(TIMEBOOST_net_14225) );
na02f02 TIMEBOOST_cell_37143 ( .a(n_14253), .b(n_14440), .o(TIMEBOOST_net_10810) );
in01s01 g62339_u0 ( .a(FE_OFN2064_n_6391), .o(g62339_sb) );
na02f02 TIMEBOOST_cell_37145 ( .a(n_14255), .b(n_14442), .o(TIMEBOOST_net_10811) );
na02s01 TIMEBOOST_cell_42747 ( .a(g65378_da), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__Q), .o(TIMEBOOST_net_13612) );
na02s01 TIMEBOOST_cell_3444 ( .a(FE_OFN207_n_9865), .b(g58106_sb), .o(TIMEBOOST_net_302) );
in01s01 g62340_u0 ( .a(FE_OFN1275_n_4096), .o(g62340_sb) );
na02m03 TIMEBOOST_cell_3049 ( .a(TIMEBOOST_net_104), .b(n_8498), .o(n_2678) );
na02m02 TIMEBOOST_cell_3999 ( .a(TIMEBOOST_net_579), .b(n_3131), .o(n_4192) );
na02m02 TIMEBOOST_cell_45456 ( .a(TIMEBOOST_net_14966), .b(g58630_sb), .o(TIMEBOOST_net_14078) );
in01s01 g62341_u0 ( .a(FE_OFN1295_n_4098), .o(g62341_sb) );
na02s01 TIMEBOOST_cell_37247 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__Q), .b(wishbone_slave_unit_fifos_wbr_control_in), .o(TIMEBOOST_net_10862) );
na02s02 TIMEBOOST_cell_42726 ( .a(TIMEBOOST_net_13601), .b(g65942_da), .o(TIMEBOOST_net_10973) );
na02s01 g57797_u1 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .b(g57797_sb), .o(g57797_da) );
in01s01 g62342_u0 ( .a(FE_OFN1259_n_4143), .o(g62342_sb) );
na02s02 TIMEBOOST_cell_37187 ( .a(g57795_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_2_), .o(TIMEBOOST_net_10832) );
na02s02 TIMEBOOST_cell_45750 ( .a(TIMEBOOST_net_15113), .b(FE_OFN1194_n_6935), .o(TIMEBOOST_net_13247) );
na02m02 TIMEBOOST_cell_42102 ( .a(TIMEBOOST_net_13289), .b(n_7618), .o(TIMEBOOST_net_11597) );
in01s01 g62343_u0 ( .a(FE_OFN1219_n_6886), .o(g62343_sb) );
na02m02 TIMEBOOST_cell_37189 ( .a(n_2458), .b(n_2475), .o(TIMEBOOST_net_10833) );
na02s02 TIMEBOOST_cell_41691 ( .a(n_707), .b(n_378), .o(TIMEBOOST_net_13084) );
na02m02 TIMEBOOST_cell_44277 ( .a(n_9542), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__Q), .o(TIMEBOOST_net_14377) );
in01s01 g62344_u0 ( .a(FE_OFN1275_n_4096), .o(g62344_sb) );
na02m02 TIMEBOOST_cell_41716 ( .a(TIMEBOOST_net_13096), .b(wbu_addr_in_260), .o(n_9860) );
na02f02 TIMEBOOST_cell_44316 ( .a(TIMEBOOST_net_14396), .b(FE_OFN1376_n_8567), .o(TIMEBOOST_net_12282) );
na02s01 TIMEBOOST_cell_3052 ( .a(n_2411), .b(wbm_adr_o_2_), .o(TIMEBOOST_net_106) );
in01s02 g62345_u0 ( .a(FE_OFN1311_n_6624), .o(g62345_sb) );
na03s02 TIMEBOOST_cell_38259 ( .a(TIMEBOOST_net_3981), .b(g64183_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q), .o(TIMEBOOST_net_11368) );
na02s01 TIMEBOOST_cell_43246 ( .a(TIMEBOOST_net_13861), .b(FE_OFN1275_n_4096), .o(TIMEBOOST_net_12551) );
na02s02 TIMEBOOST_cell_39864 ( .a(TIMEBOOST_net_12170), .b(g62978_sb), .o(n_5926) );
in01s01 g62346_u0 ( .a(FE_OFN1231_n_6391), .o(g62346_sb) );
na02m02 TIMEBOOST_cell_44385 ( .a(n_9091), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__Q), .o(TIMEBOOST_net_14431) );
na02f02 TIMEBOOST_cell_37133 ( .a(FE_RN_89_0), .b(n_10644), .o(TIMEBOOST_net_10805) );
na02s02 TIMEBOOST_cell_38354 ( .a(TIMEBOOST_net_11415), .b(g62841_sb), .o(n_5290) );
in01s01 g62347_u0 ( .a(FE_OFN1219_n_6886), .o(g62347_sb) );
no02f04 TIMEBOOST_cell_42562 ( .a(TIMEBOOST_net_13519), .b(FE_RN_638_0), .o(TIMEBOOST_net_130) );
na02s01 TIMEBOOST_cell_16016 ( .a(FE_OFN2094_n_2520), .b(g66419_db), .o(TIMEBOOST_net_3265) );
na02f04 TIMEBOOST_cell_44768 ( .a(TIMEBOOST_net_14622), .b(FE_RN_270_0), .o(TIMEBOOST_net_1096) );
in01s01 g62348_u0 ( .a(n_6319), .o(g62348_sb) );
na02f02 TIMEBOOST_cell_37147 ( .a(n_14511), .b(n_14429), .o(TIMEBOOST_net_10812) );
na02s01 TIMEBOOST_cell_39201 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__Q), .b(n_8119), .o(TIMEBOOST_net_11839) );
no02f08 TIMEBOOST_cell_3346 ( .a(FE_OCPN1843_n_16033), .b(n_15999), .o(TIMEBOOST_net_253) );
in01s01 g62349_u0 ( .a(FE_OFN1269_n_4095), .o(g62349_sb) );
na02s01 TIMEBOOST_cell_37191 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(g65711_sb), .o(TIMEBOOST_net_10834) );
na02s02 TIMEBOOST_cell_42103 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__Q), .b(n_3632), .o(TIMEBOOST_net_13290) );
na02s02 TIMEBOOST_cell_42104 ( .a(TIMEBOOST_net_13290), .b(FE_OFN1317_n_6624), .o(TIMEBOOST_net_11590) );
in01s01 g62350_u0 ( .a(FE_OFN1278_n_4097), .o(g62350_sb) );
na02s01 TIMEBOOST_cell_37193 ( .a(pci_target_unit_fifos_pcir_data_in_167), .b(g65775_sb), .o(TIMEBOOST_net_10835) );
na02s01 TIMEBOOST_cell_16061 ( .a(TIMEBOOST_net_3287), .b(g65867_db), .o(n_1577) );
na02s02 TIMEBOOST_cell_43247 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q), .b(n_4376), .o(TIMEBOOST_net_13862) );
in01s02 g62351_u0 ( .a(FE_OFN1322_n_6436), .o(g62351_sb) );
na02s02 TIMEBOOST_cell_43314 ( .a(TIMEBOOST_net_13895), .b(FE_OFN1225_n_6391), .o(n_5997) );
na02s02 TIMEBOOST_cell_43372 ( .a(TIMEBOOST_net_13924), .b(n_6319), .o(TIMEBOOST_net_12174) );
na02s01 TIMEBOOST_cell_31244 ( .a(n_4442), .b(g65014_sb), .o(TIMEBOOST_net_9533) );
in01s01 g62352_u0 ( .a(FE_OFN1250_n_4093), .o(g62352_sb) );
na02s02 TIMEBOOST_cell_3053 ( .a(TIMEBOOST_net_106), .b(n_1975), .o(n_2934) );
na02s02 TIMEBOOST_cell_18619 ( .a(TIMEBOOST_net_4566), .b(g62771_sb), .o(n_5452) );
no02s01 TIMEBOOST_cell_3054 ( .a(n_1460), .b(n_169), .o(TIMEBOOST_net_107) );
in01s01 g62353_u0 ( .a(FE_OFN1261_n_4143), .o(g62353_sb) );
na02s01 TIMEBOOST_cell_37195 ( .a(pci_target_unit_fifos_pcir_data_in_173), .b(g65678_sb), .o(TIMEBOOST_net_10836) );
na02m02 TIMEBOOST_cell_43717 ( .a(n_9044), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__Q), .o(TIMEBOOST_net_14097) );
na02f02 TIMEBOOST_cell_44334 ( .a(TIMEBOOST_net_14405), .b(FE_OFN1377_n_8567), .o(TIMEBOOST_net_12737) );
in01s01 g62354_u0 ( .a(FE_OFN1261_n_4143), .o(g62354_sb) );
na02m02 TIMEBOOST_cell_37197 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_3_), .o(TIMEBOOST_net_10837) );
na03s01 TIMEBOOST_cell_33543 ( .a(n_1908), .b(g61748_sb), .c(g61748_db), .o(n_8321) );
na02s01 TIMEBOOST_cell_45220 ( .a(TIMEBOOST_net_14848), .b(FE_OFN1218_n_6886), .o(TIMEBOOST_net_12112) );
in01s01 g62355_u0 ( .a(FE_OFN1232_n_6391), .o(g62355_sb) );
na03f04 TIMEBOOST_cell_37129 ( .a(n_11716), .b(n_10527), .c(n_10859), .o(TIMEBOOST_net_10803) );
na02s01 TIMEBOOST_cell_3445 ( .a(TIMEBOOST_net_302), .b(g58106_db), .o(n_9689) );
na02s01 TIMEBOOST_cell_15895 ( .a(TIMEBOOST_net_3204), .b(g56933_sb), .o(TIMEBOOST_net_897) );
in01s01 g62356_u0 ( .a(FE_OFN1218_n_6886), .o(g62356_sb) );
na02s01 TIMEBOOST_cell_37199 ( .a(pci_target_unit_fifos_pcir_data_in_187), .b(g65698_sb), .o(TIMEBOOST_net_10838) );
na02f02 TIMEBOOST_cell_42150 ( .a(TIMEBOOST_net_13313), .b(g57353_sb), .o(n_11394) );
na03s01 TIMEBOOST_cell_33542 ( .a(n_1914), .b(g61742_sb), .c(g61742_db), .o(n_8333) );
in01s01 g62357_u0 ( .a(FE_OFN1284_n_4097), .o(g62357_sb) );
na02s01 TIMEBOOST_cell_37753 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__Q), .b(wbs_dat_i_24_), .o(TIMEBOOST_net_11115) );
in01s01 g62358_u0 ( .a(FE_OFN1273_n_4096), .o(g62358_sb) );
na02m02 TIMEBOOST_cell_32688 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__Q), .o(TIMEBOOST_net_10255) );
no03f06 TIMEBOOST_cell_37169 ( .a(FE_RN_677_0), .b(n_376), .c(n_2844), .o(TIMEBOOST_net_10823) );
na02f02 TIMEBOOST_cell_41496 ( .a(TIMEBOOST_net_12986), .b(g57486_sb), .o(n_11251) );
in01s01 g62359_u0 ( .a(FE_OFN1216_n_4151), .o(g62359_sb) );
na02f04 TIMEBOOST_cell_11924 ( .a(n_16325), .b(FE_RN_592_0), .o(TIMEBOOST_net_2529) );
na03s01 TIMEBOOST_cell_33541 ( .a(TIMEBOOST_net_267), .b(g61765_sb), .c(g61765_db), .o(n_8281) );
na03s02 TIMEBOOST_cell_43315 ( .a(n_4434), .b(FE_OFN1274_n_4096), .c(n_18), .o(TIMEBOOST_net_13896) );
in01s01 g62360_u0 ( .a(FE_OFN1282_n_4097), .o(g62360_sb) );
na02s01 TIMEBOOST_cell_37755 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__Q), .b(wbs_dat_i_22_), .o(TIMEBOOST_net_11116) );
na02f02 TIMEBOOST_cell_41670 ( .a(TIMEBOOST_net_13073), .b(FE_OFN1768_n_14054), .o(n_14508) );
na02f02 TIMEBOOST_cell_44310 ( .a(TIMEBOOST_net_14393), .b(FE_OFN1412_n_8567), .o(TIMEBOOST_net_12738) );
in01s01 g62361_u0 ( .a(FE_OFN1246_n_4093), .o(g62361_sb) );
na02m02 TIMEBOOST_cell_39160 ( .a(g58780_db), .b(TIMEBOOST_net_11818), .o(n_9844) );
na02f02 TIMEBOOST_cell_42476 ( .a(TIMEBOOST_net_13476), .b(g57505_sb), .o(n_10817) );
na02s01 TIMEBOOST_cell_45666 ( .a(TIMEBOOST_net_15071), .b(g63617_da), .o(n_7157) );
in01s01 g62362_u0 ( .a(FE_OFN1274_n_4096), .o(g62362_sb) );
no02f06 TIMEBOOST_cell_3059 ( .a(TIMEBOOST_net_109), .b(n_16286), .o(n_16288) );
na02f02 TIMEBOOST_cell_37139 ( .a(FE_RN_137_0), .b(n_10907), .o(TIMEBOOST_net_10808) );
na02s02 TIMEBOOST_cell_43248 ( .a(TIMEBOOST_net_13862), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_12042) );
in01s01 g62363_u0 ( .a(n_6431), .o(g62363_sb) );
na03s02 TIMEBOOST_cell_37771 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__Q), .b(FE_OFN716_n_8176), .c(n_1587), .o(TIMEBOOST_net_11124) );
no02f20 TIMEBOOST_cell_3347 ( .a(TIMEBOOST_net_253), .b(FE_RN_149_0), .o(n_16810) );
na02f02 TIMEBOOST_cell_3348 ( .a(n_1358), .b(conf_wb_err_addr_in_943), .o(TIMEBOOST_net_254) );
in01s01 g62364_u0 ( .a(FE_OFN1258_n_4143), .o(g62364_sb) );
na02s02 TIMEBOOST_cell_39866 ( .a(TIMEBOOST_net_12171), .b(g62911_sb), .o(n_6056) );
na02f02 TIMEBOOST_cell_44232 ( .a(TIMEBOOST_net_14354), .b(FE_OFN1424_n_8567), .o(TIMEBOOST_net_13402) );
na02s01 TIMEBOOST_cell_43132 ( .a(TIMEBOOST_net_13804), .b(FE_OFN1265_n_4095), .o(TIMEBOOST_net_12128) );
in01s01 g62365_u0 ( .a(FE_OFN1222_n_6391), .o(g62365_sb) );
na02f02 TIMEBOOST_cell_32687 ( .a(FE_OFN1762_n_10780), .b(TIMEBOOST_net_10254), .o(TIMEBOOST_net_6515) );
na03s02 TIMEBOOST_cell_37727 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__Q), .b(FE_OFN717_n_8176), .c(n_1933), .o(TIMEBOOST_net_11102) );
na02s01 TIMEBOOST_cell_3062 ( .a(n_1089), .b(parchk_pci_par_en_in), .o(TIMEBOOST_net_111) );
in01s01 g62366_u0 ( .a(FE_OFN1192_n_6935), .o(g62366_sb) );
na02s01 TIMEBOOST_cell_3063 ( .a(TIMEBOOST_net_111), .b(n_12855), .o(n_13332) );
na02s01 g62366_u2 ( .a(n_3765), .b(FE_OFN1192_n_6935), .o(g62366_db) );
in01s01 g62367_u0 ( .a(FE_OFN2063_n_6391), .o(g62367_sb) );
na03f04 TIMEBOOST_cell_37093 ( .a(n_10672), .b(n_10096), .c(n_10675), .o(TIMEBOOST_net_10785) );
na02f02 TIMEBOOST_cell_43974 ( .a(TIMEBOOST_net_14225), .b(FE_OFN1425_n_8567), .o(TIMEBOOST_net_12907) );
na03s02 TIMEBOOST_cell_34794 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__Q), .b(g62925_sb), .c(g62925_db), .o(n_6031) );
in01s01 g62368_u0 ( .a(n_6287), .o(g62368_sb) );
na02f02 TIMEBOOST_cell_37095 ( .a(FE_RN_35_0), .b(n_10974), .o(TIMEBOOST_net_10786) );
na02f02 TIMEBOOST_cell_3349 ( .a(TIMEBOOST_net_254), .b(n_2397), .o(n_2266) );
na02m02 TIMEBOOST_cell_32686 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__Q), .o(TIMEBOOST_net_10254) );
in01s01 g62369_u0 ( .a(FE_OFN1293_n_4098), .o(g62369_sb) );
na02s02 TIMEBOOST_cell_45152 ( .a(TIMEBOOST_net_14814), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_13230) );
na02s01 TIMEBOOST_cell_43133 ( .a(n_4296), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__Q), .o(TIMEBOOST_net_13805) );
na02s02 TIMEBOOST_cell_42603 ( .a(n_3764), .b(g65016_sb), .o(TIMEBOOST_net_13540) );
in01s01 g62370_u0 ( .a(FE_OFN1230_n_6391), .o(g62370_sb) );
in01s01 TIMEBOOST_cell_45907 ( .a(wbm_dat_i_13_), .o(TIMEBOOST_net_15214) );
na02s01 TIMEBOOST_cell_44967 ( .a(FE_OFN215_n_9856), .b(g57920_sb), .o(TIMEBOOST_net_14722) );
na02s01 TIMEBOOST_cell_31051 ( .a(TIMEBOOST_net_9436), .b(g64964_db), .o(n_4375) );
in01s01 g62371_u0 ( .a(FE_OFN1194_n_6935), .o(g62371_sb) );
na02s01 TIMEBOOST_cell_3065 ( .a(TIMEBOOST_net_112), .b(FE_OFN992_n_2373), .o(n_7397) );
na02f06 TIMEBOOST_cell_36835 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_), .b(g75162_sb), .o(TIMEBOOST_net_10656) );
na02s01 TIMEBOOST_cell_3066 ( .a(n_1690), .b(n_1187), .o(TIMEBOOST_net_113) );
in01s01 g62372_u0 ( .a(FE_OFN1284_n_4097), .o(g62372_sb) );
na02s02 TIMEBOOST_cell_3067 ( .a(TIMEBOOST_net_113), .b(n_1438), .o(n_2295) );
na02s01 TIMEBOOST_cell_37757 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__Q), .b(wbs_dat_i_18_), .o(TIMEBOOST_net_11117) );
na02s02 TIMEBOOST_cell_3068 ( .a(n_1689), .b(n_1186), .o(TIMEBOOST_net_114) );
in01s01 g62373_u0 ( .a(FE_OFN1295_n_4098), .o(g62373_sb) );
na02s01 TIMEBOOST_cell_44968 ( .a(TIMEBOOST_net_14722), .b(g57920_db), .o(n_9891) );
na02f04 TIMEBOOST_cell_42585 ( .a(TIMEBOOST_net_3293), .b(n_16391), .o(TIMEBOOST_net_13531) );
na02s02 TIMEBOOST_cell_43134 ( .a(TIMEBOOST_net_13805), .b(FE_OFN1224_n_6391), .o(TIMEBOOST_net_12524) );
in01s01 g62374_u0 ( .a(FE_OFN1207_n_6356), .o(g62374_sb) );
na02s01 TIMEBOOST_cell_42838 ( .a(TIMEBOOST_net_13657), .b(g63597_da), .o(n_7195) );
na02f06 TIMEBOOST_cell_42586 ( .a(TIMEBOOST_net_13531), .b(n_16311), .o(n_16798) );
na02m02 TIMEBOOST_cell_42563 ( .a(FE_OFN2059_n_13447), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__Q), .o(TIMEBOOST_net_13520) );
in01s01 g62375_u0 ( .a(FE_OFN1269_n_4095), .o(g62375_sb) );
na02f02 TIMEBOOST_cell_37099 ( .a(FE_RN_32_0), .b(n_10986), .o(TIMEBOOST_net_10788) );
na02f02 TIMEBOOST_cell_44721 ( .a(TIMEBOOST_net_10177), .b(FE_OCPN2218_n_13997), .o(TIMEBOOST_net_14599) );
in01s01 g62376_u0 ( .a(FE_OFN1261_n_4143), .o(g62376_sb) );
na02f04 TIMEBOOST_cell_42818 ( .a(TIMEBOOST_net_13647), .b(n_7321), .o(TIMEBOOST_net_9882) );
na02s02 TIMEBOOST_cell_42024 ( .a(TIMEBOOST_net_13250), .b(g62507_sb), .o(n_6566) );
na03s02 TIMEBOOST_cell_42025 ( .a(n_4382), .b(FE_OFN1223_n_6391), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__Q), .o(TIMEBOOST_net_13251) );
in01s01 g62377_u0 ( .a(FE_OFN1260_n_4143), .o(g62377_sb) );
na04m02 TIMEBOOST_cell_34388 ( .a(g52394_sb), .b(n_8757), .c(g52632_da), .d(g52632_db), .o(TIMEBOOST_net_5442) );
na02s02 TIMEBOOST_cell_43006 ( .a(TIMEBOOST_net_13741), .b(g63621_da), .o(n_7174) );
in01s01 g62378_u0 ( .a(FE_OFN1231_n_6391), .o(g62378_sb) );
na02s02 TIMEBOOST_cell_43423 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__31__Q), .b(n_4670), .o(TIMEBOOST_net_13950) );
na03f02 TIMEBOOST_cell_36895 ( .a(n_354), .b(FE_OFN1394_n_8567), .c(n_8549), .o(TIMEBOOST_net_10686) );
na03s02 TIMEBOOST_cell_34281 ( .a(TIMEBOOST_net_9806), .b(FE_OFN1173_n_5592), .c(g62083_sb), .o(n_5626) );
in01s01 g62379_u0 ( .a(FE_OFN1230_n_6391), .o(g62379_sb) );
na02s02 TIMEBOOST_cell_39295 ( .a(TIMEBOOST_net_9400), .b(FE_OFN1797_n_2299), .o(TIMEBOOST_net_11886) );
na02s01 TIMEBOOST_cell_3451 ( .a(TIMEBOOST_net_305), .b(n_4450), .o(n_4221) );
na02s02 TIMEBOOST_cell_37994 ( .a(TIMEBOOST_net_11235), .b(g52630_sb), .o(n_14676) );
in01s01 g62380_u0 ( .a(FE_OFN1269_n_4095), .o(g62380_sb) );
no02f02 TIMEBOOST_cell_36891 ( .a(FE_RN_569_0), .b(n_7552), .o(TIMEBOOST_net_10684) );
na02s02 TIMEBOOST_cell_42075 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__Q), .b(n_3784), .o(TIMEBOOST_net_13276) );
na02s02 TIMEBOOST_cell_42088 ( .a(TIMEBOOST_net_13282), .b(n_6554), .o(TIMEBOOST_net_11579) );
in01s01 g62381_u0 ( .a(FE_OFN2064_n_6391), .o(g62381_sb) );
na02s02 TIMEBOOST_cell_36897 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_769), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_4__Q), .o(TIMEBOOST_net_10687) );
na02s02 TIMEBOOST_cell_3453 ( .a(TIMEBOOST_net_306), .b(n_4450), .o(n_4451) );
na02f02 TIMEBOOST_cell_44386 ( .a(TIMEBOOST_net_14431), .b(FE_OFN1412_n_8567), .o(TIMEBOOST_net_12782) );
in01s01 g62382_u0 ( .a(n_6554), .o(g62382_sb) );
na02s02 TIMEBOOST_cell_42774 ( .a(TIMEBOOST_net_13625), .b(g58174_db), .o(n_9061) );
na02s01 TIMEBOOST_cell_3351 ( .a(TIMEBOOST_net_255), .b(g65797_sb), .o(n_1591) );
na02f04 TIMEBOOST_cell_37295 ( .a(TIMEBOOST_net_193), .b(n_2447), .o(TIMEBOOST_net_10886) );
in01s01 g62383_u0 ( .a(FE_OFN1218_n_6886), .o(g62383_sb) );
na02s01 TIMEBOOST_cell_40386 ( .a(TIMEBOOST_net_12431), .b(g64257_db), .o(n_3916) );
na02f02 TIMEBOOST_cell_44229 ( .a(n_9625), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__Q), .o(TIMEBOOST_net_14353) );
na02f02 TIMEBOOST_cell_32588 ( .a(FE_OFN1747_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__Q), .o(TIMEBOOST_net_10205) );
in01s01 g62384_u0 ( .a(FE_OFN1284_n_4097), .o(g62384_sb) );
na02s02 TIMEBOOST_cell_3069 ( .a(TIMEBOOST_net_114), .b(n_1476), .o(n_2275) );
na03s01 TIMEBOOST_cell_38049 ( .a(g64141_da), .b(g64141_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__Q), .o(TIMEBOOST_net_11263) );
na02s02 TIMEBOOST_cell_45063 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__Q), .b(FE_OFN1654_n_9502), .o(TIMEBOOST_net_14770) );
in01s01 g62385_u0 ( .a(FE_OFN1285_n_4097), .o(g62385_sb) );
na02f02 TIMEBOOST_cell_37083 ( .a(FE_OCP_RBN1998_n_13971), .b(TIMEBOOST_net_10236), .o(TIMEBOOST_net_10780) );
na03s02 TIMEBOOST_cell_41995 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__Q), .b(n_4319), .c(FE_OFN1241_n_4092), .o(TIMEBOOST_net_13236) );
in01s01 g62386_u0 ( .a(FE_OFN1261_n_4143), .o(g62386_sb) );
na02f02 TIMEBOOST_cell_37085 ( .a(FE_OCP_RBN1996_n_13971), .b(TIMEBOOST_net_10234), .o(TIMEBOOST_net_10781) );
na03s02 TIMEBOOST_cell_42059 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__Q), .b(n_4370), .c(FE_OFN1249_n_4093), .o(TIMEBOOST_net_13268) );
na02s02 TIMEBOOST_cell_45786 ( .a(TIMEBOOST_net_15131), .b(FE_OFN1812_n_7845), .o(TIMEBOOST_net_11384) );
in01s01 g62387_u0 ( .a(FE_OFN1273_n_4096), .o(g62387_sb) );
na02s02 TIMEBOOST_cell_45457 ( .a(n_982), .b(TIMEBOOST_net_898), .o(TIMEBOOST_net_14967) );
na02s01 TIMEBOOST_cell_37759 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__Q), .b(wbs_dat_i_5_), .o(TIMEBOOST_net_11118) );
no02m01 TIMEBOOST_cell_3072 ( .a(n_2263), .b(wishbone_slave_unit_pcim_sm_be_in_557), .o(TIMEBOOST_net_116) );
in01s01 g62388_u0 ( .a(FE_OFN1213_n_4151), .o(g62388_sb) );
na02f02 TIMEBOOST_cell_37087 ( .a(TIMEBOOST_net_10230), .b(FE_OCP_RBN1997_n_13971), .o(TIMEBOOST_net_10782) );
na02s02 TIMEBOOST_cell_42012 ( .a(TIMEBOOST_net_13244), .b(g62411_sb), .o(n_6776) );
na03s02 TIMEBOOST_cell_42013 ( .a(n_4395), .b(FE_OFN1275_n_4096), .c(n_4394), .o(TIMEBOOST_net_13245) );
in01s01 g62389_u0 ( .a(FE_OFN1212_n_4151), .o(g62389_sb) );
na02s02 TIMEBOOST_cell_37622 ( .a(TIMEBOOST_net_11049), .b(g62010_sb), .o(n_7875) );
na02s01 TIMEBOOST_cell_2887 ( .a(TIMEBOOST_net_23), .b(n_879), .o(n_880) );
na02s01 TIMEBOOST_cell_2888 ( .a(wbm_adr_o_28_), .b(wbm_adr_o_29_), .o(TIMEBOOST_net_24) );
in01s01 g62390_u0 ( .a(FE_OFN1279_n_4097), .o(g62390_sb) );
na02f02 TIMEBOOST_cell_37091 ( .a(FE_OCP_RBN1995_n_13971), .b(TIMEBOOST_net_10232), .o(TIMEBOOST_net_10784) );
na02s01 TIMEBOOST_cell_42014 ( .a(TIMEBOOST_net_13245), .b(g62344_sb), .o(n_6911) );
na02s02 TIMEBOOST_cell_41996 ( .a(TIMEBOOST_net_13236), .b(g62436_sb), .o(n_6724) );
in01s01 g62391_u0 ( .a(FE_OFN1285_n_4097), .o(g62391_sb) );
na02f02 TIMEBOOST_cell_37089 ( .a(FE_OCP_RBN1998_n_13971), .b(TIMEBOOST_net_10229), .o(TIMEBOOST_net_10783) );
na02s02 TIMEBOOST_cell_42060 ( .a(TIMEBOOST_net_13268), .b(g62524_sb), .o(n_6528) );
na02f02 TIMEBOOST_cell_42320 ( .a(TIMEBOOST_net_13398), .b(g57430_sb), .o(n_10359) );
in01s01 g62392_u0 ( .a(FE_OFN1208_n_6356), .o(g62392_sb) );
na02f02 TIMEBOOST_cell_37063 ( .a(FE_RN_188_0), .b(n_10890), .o(TIMEBOOST_net_10770) );
na02s02 TIMEBOOST_cell_45458 ( .a(TIMEBOOST_net_14967), .b(g58633_sb), .o(TIMEBOOST_net_14079) );
in01s01 g62393_u0 ( .a(FE_OFN1250_n_4093), .o(g62393_sb) );
na02m02 TIMEBOOST_cell_43975 ( .a(n_9466), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__Q), .o(TIMEBOOST_net_14226) );
na02s02 TIMEBOOST_cell_38612 ( .a(TIMEBOOST_net_11544), .b(g62888_sb), .o(n_6101) );
na02f02 TIMEBOOST_cell_41022 ( .a(TIMEBOOST_net_12749), .b(g57419_sb), .o(n_11320) );
in01s01 g62394_u0 ( .a(FE_OFN1275_n_4096), .o(g62394_sb) );
na02s01 TIMEBOOST_cell_3075 ( .a(TIMEBOOST_net_117), .b(g65810_sb), .o(n_2186) );
na02s01 TIMEBOOST_cell_37761 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__Q), .b(wbs_dat_i_6_), .o(TIMEBOOST_net_11119) );
na02f02 TIMEBOOST_cell_32685 ( .a(FE_OFN1761_n_10780), .b(TIMEBOOST_net_10253), .o(TIMEBOOST_net_6513) );
in01s02 g62395_u0 ( .a(FE_OFN1316_n_6624), .o(g62395_sb) );
na03m02 TIMEBOOST_cell_34807 ( .a(TIMEBOOST_net_5442), .b(n_3486), .c(TIMEBOOST_net_587), .o(n_14803) );
na02f02 TIMEBOOST_cell_43976 ( .a(TIMEBOOST_net_14226), .b(FE_OFN1424_n_8567), .o(TIMEBOOST_net_13377) );
na02s02 TIMEBOOST_cell_40726 ( .a(TIMEBOOST_net_12601), .b(g62638_sb), .o(n_6273) );
in01s01 g62396_u0 ( .a(n_6431), .o(g62396_sb) );
na02f02 TIMEBOOST_cell_37065 ( .a(n_13987), .b(TIMEBOOST_net_10223), .o(TIMEBOOST_net_10771) );
na02f01 TIMEBOOST_cell_3353 ( .a(n_15014), .b(TIMEBOOST_net_256), .o(n_5742) );
na02s01 TIMEBOOST_cell_3354 ( .a(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .b(FE_OCPN1875_n_14526), .o(TIMEBOOST_net_257) );
in01s01 g62397_u0 ( .a(FE_OFN1214_n_4151), .o(g62397_sb) );
na02f02 TIMEBOOST_cell_37069 ( .a(n_13987), .b(TIMEBOOST_net_10224), .o(TIMEBOOST_net_10773) );
na03s02 TIMEBOOST_cell_42061 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__Q), .b(n_3655), .c(FE_OFN1249_n_4093), .o(TIMEBOOST_net_13269) );
na02s02 TIMEBOOST_cell_42727 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__Q), .b(FE_OFN569_n_9528), .o(TIMEBOOST_net_13602) );
in01s01 g62398_u0 ( .a(FE_OFN1260_n_4143), .o(g62398_sb) );
na02s02 TIMEBOOST_cell_42775 ( .a(FE_OFN1687_n_9528), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__Q), .o(TIMEBOOST_net_13626) );
na02s01 TIMEBOOST_cell_43373 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__Q), .b(n_4263), .o(TIMEBOOST_net_13925) );
na02s02 TIMEBOOST_cell_41998 ( .a(TIMEBOOST_net_13237), .b(g63151_sb), .o(n_5838) );
in01s01 g62399_u0 ( .a(FE_OFN1193_n_6935), .o(g62399_sb) );
na02s01 TIMEBOOST_cell_3077 ( .a(TIMEBOOST_net_118), .b(g65835_sb), .o(n_2185) );
na02s01 TIMEBOOST_cell_37763 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__Q), .b(wbs_dat_i_26_), .o(TIMEBOOST_net_11120) );
na02s02 TIMEBOOST_cell_45459 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_2__Q), .b(TIMEBOOST_net_897), .o(TIMEBOOST_net_14968) );
in01s01 g62400_u0 ( .a(n_6645), .o(g62400_sb) );
na02f02 TIMEBOOST_cell_36899 ( .a(FE_RN_570_0), .b(FE_RN_572_0), .o(TIMEBOOST_net_10688) );
na02m01 TIMEBOOST_cell_3355 ( .a(n_15014), .b(TIMEBOOST_net_257), .o(n_7329) );
na02f02 TIMEBOOST_cell_3356 ( .a(n_16021), .b(n_15055), .o(TIMEBOOST_net_258) );
in01s01 g62401_u0 ( .a(FE_OFN1313_n_6624), .o(g62401_sb) );
na02f02 TIMEBOOST_cell_42196 ( .a(TIMEBOOST_net_13336), .b(FE_OFN1419_n_8567), .o(TIMEBOOST_net_12288) );
na02m02 TIMEBOOST_cell_42239 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__Q), .b(n_9500), .o(TIMEBOOST_net_13358) );
na02f02 TIMEBOOST_cell_44306 ( .a(TIMEBOOST_net_14391), .b(FE_OFN1408_n_8567), .o(TIMEBOOST_net_13407) );
in01s01 g62402_u0 ( .a(FE_OFN1236_n_6391), .o(g62402_sb) );
na02m02 TIMEBOOST_cell_42819 ( .a(pci_target_unit_pcit_if_strd_addr_in_689), .b(g52648_sb), .o(TIMEBOOST_net_13648) );
na02m04 TIMEBOOST_cell_3455 ( .a(n_3132), .b(TIMEBOOST_net_307), .o(n_3142) );
na02s02 TIMEBOOST_cell_21977 ( .a(n_10139), .b(TIMEBOOST_net_6245), .o(n_11853) );
in01s01 g62403_u0 ( .a(FE_OFN1232_n_6391), .o(g62403_sb) );
na02s02 TIMEBOOST_cell_42776 ( .a(TIMEBOOST_net_13626), .b(FE_OFN254_n_9825), .o(TIMEBOOST_net_10990) );
na02s01 TIMEBOOST_cell_3457 ( .a(TIMEBOOST_net_308), .b(n_4450), .o(n_4503) );
na04f04 TIMEBOOST_cell_36223 ( .a(n_13972), .b(n_14556), .c(n_14454), .d(n_13857), .o(n_14601) );
in01s01 g62404_u0 ( .a(n_6319), .o(g62404_sb) );
na02m02 TIMEBOOST_cell_42820 ( .a(TIMEBOOST_net_13648), .b(g52648_db), .o(n_14740) );
na02f02 TIMEBOOST_cell_3357 ( .a(n_15014), .b(TIMEBOOST_net_258), .o(n_15446) );
na02s01 TIMEBOOST_cell_45743 ( .a(n_1937), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__Q), .o(TIMEBOOST_net_15110) );
in01s01 g62405_u0 ( .a(FE_OFN1219_n_6886), .o(g62405_sb) );
na02m02 TIMEBOOST_cell_42821 ( .a(pci_target_unit_pcit_if_strd_addr_in_694), .b(g52653_sb), .o(TIMEBOOST_net_13649) );
na03s02 TIMEBOOST_cell_41999 ( .a(n_6), .b(n_4433), .c(FE_OFN369_n_4092), .o(TIMEBOOST_net_13238) );
na02m02 TIMEBOOST_cell_42197 ( .a(n_9580), .b(FE_RN_484_0), .o(TIMEBOOST_net_13337) );
in01s01 g62406_u0 ( .a(FE_OFN1235_n_6391), .o(g62406_sb) );
na02s01 TIMEBOOST_cell_42694 ( .a(TIMEBOOST_net_13585), .b(g58333_sb), .o(TIMEBOOST_net_10970) );
na02m04 TIMEBOOST_cell_3459 ( .a(n_3378), .b(TIMEBOOST_net_309), .o(n_8750) );
na02m02 TIMEBOOST_cell_40872 ( .a(TIMEBOOST_net_12674), .b(FE_OFN1331_n_13547), .o(TIMEBOOST_net_11625) );
in01s02 g62407_u0 ( .a(FE_OFN1310_n_6624), .o(g62407_sb) );
na02f02 TIMEBOOST_cell_41088 ( .a(TIMEBOOST_net_12782), .b(g57196_sb), .o(n_10446) );
na03s02 TIMEBOOST_cell_33755 ( .a(FE_OFN221_n_9846), .b(g57989_sb), .c(g57989_db), .o(n_9807) );
na02s01 TIMEBOOST_cell_40402 ( .a(g63619_da), .b(TIMEBOOST_net_12439), .o(n_7200) );
in01s02 g62408_u0 ( .a(FE_OFN1310_n_6624), .o(g62408_sb) );
na03s02 TIMEBOOST_cell_38381 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__Q), .b(FE_OFN1115_g64577_p), .c(n_4068), .o(TIMEBOOST_net_11429) );
na02f02 TIMEBOOST_cell_44751 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q), .b(FE_OCPN1825_n_12030), .o(TIMEBOOST_net_14614) );
na02s01 TIMEBOOST_cell_38039 ( .a(n_2174), .b(g61735_sb), .o(TIMEBOOST_net_11258) );
in01s01 g62409_u0 ( .a(FE_OFN1234_n_6391), .o(g62409_sb) );
na02s01 TIMEBOOST_cell_41739 ( .a(n_3761), .b(g65059_sb), .o(TIMEBOOST_net_13108) );
na03s02 TIMEBOOST_cell_40689 ( .a(n_4298), .b(FE_OFN1215_n_4151), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__Q), .o(TIMEBOOST_net_12583) );
na03f02 TIMEBOOST_cell_3462 ( .a(FE_RN_631_0), .b(FE_RN_641_0), .c(FE_RN_666_0), .o(TIMEBOOST_net_311) );
in01s01 g62410_u0 ( .a(FE_OFN1270_n_4095), .o(g62410_sb) );
na02m02 TIMEBOOST_cell_42822 ( .a(TIMEBOOST_net_13649), .b(g52653_db), .o(n_14733) );
na02s01 TIMEBOOST_cell_43249 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__Q), .b(n_3570), .o(TIMEBOOST_net_13863) );
na02s02 TIMEBOOST_cell_41990 ( .a(TIMEBOOST_net_13233), .b(g63001_sb), .o(n_5880) );
in01s01 g62411_u0 ( .a(FE_OFN1272_n_4096), .o(g62411_sb) );
na02s01 TIMEBOOST_cell_3079 ( .a(TIMEBOOST_net_119), .b(g65907_sb), .o(n_2151) );
na02s02 TIMEBOOST_cell_18653 ( .a(TIMEBOOST_net_4583), .b(g63142_sb), .o(n_4963) );
na02s02 TIMEBOOST_cell_42634 ( .a(TIMEBOOST_net_13555), .b(g58195_db), .o(n_9591) );
in01s01 g62412_u0 ( .a(FE_OFN1202_n_4090), .o(g62412_sb) );
na02s02 TIMEBOOST_cell_40728 ( .a(TIMEBOOST_net_12602), .b(g63011_sb), .o(n_5862) );
na02f02 TIMEBOOST_cell_44695 ( .a(n_973), .b(n_14971), .o(TIMEBOOST_net_14586) );
na02f02 TIMEBOOST_cell_44674 ( .a(TIMEBOOST_net_14575), .b(g57528_sb), .o(n_11213) );
in01s01 g62413_u0 ( .a(FE_OFN1253_n_4143), .o(g62413_sb) );
na02f02 TIMEBOOST_cell_36903 ( .a(n_3366), .b(n_3228), .o(TIMEBOOST_net_10690) );
na02m02 TIMEBOOST_cell_43576 ( .a(TIMEBOOST_net_14026), .b(FE_OFN1323_n_6436), .o(TIMEBOOST_net_12215) );
na02s01 TIMEBOOST_cell_42030 ( .a(TIMEBOOST_net_13253), .b(g62609_sb), .o(n_6335) );
in01s01 g62414_u0 ( .a(FE_OFN1214_n_4151), .o(g62414_sb) );
na02s01 TIMEBOOST_cell_42612 ( .a(TIMEBOOST_net_13544), .b(g58034_db), .o(n_9097) );
na02s01 TIMEBOOST_cell_42000 ( .a(TIMEBOOST_net_13238), .b(g62506_sb), .o(n_6567) );
na02s02 TIMEBOOST_cell_41807 ( .a(n_4482), .b(g64870_db), .o(TIMEBOOST_net_13142) );
in01s01 g62415_u0 ( .a(FE_OFN1219_n_6886), .o(g62415_sb) );
na02s01 TIMEBOOST_cell_42613 ( .a(FE_OFN217_n_9889), .b(g57984_sb), .o(TIMEBOOST_net_13545) );
na02s02 TIMEBOOST_cell_43374 ( .a(TIMEBOOST_net_13925), .b(n_6287), .o(TIMEBOOST_net_12178) );
na02s02 TIMEBOOST_cell_43577 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__Q), .b(n_4416), .o(TIMEBOOST_net_14027) );
in01s02 g62416_u0 ( .a(FE_OFN1316_n_6624), .o(g62416_sb) );
na03s02 TIMEBOOST_cell_39363 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__Q), .b(FE_OFN717_n_8176), .c(n_1897), .o(TIMEBOOST_net_11920) );
na02s01 TIMEBOOST_cell_42748 ( .a(TIMEBOOST_net_13612), .b(TIMEBOOST_net_3877), .o(TIMEBOOST_net_4796) );
na02s01 TIMEBOOST_cell_36330 ( .a(TIMEBOOST_net_10403), .b(g65959_db), .o(n_2163) );
in01s01 g62417_u0 ( .a(FE_OFN1253_n_4143), .o(g62417_sb) );
na02f08 TIMEBOOST_cell_36855 ( .a(n_16524), .b(FE_OCPN1823_n_16560), .o(TIMEBOOST_net_10666) );
na02s01 TIMEBOOST_cell_42062 ( .a(TIMEBOOST_net_13269), .b(g62531_sb), .o(n_6512) );
na03s02 TIMEBOOST_cell_42001 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__Q), .b(n_4467), .c(FE_OFN1219_n_6886), .o(TIMEBOOST_net_13239) );
in01s01 g62418_u0 ( .a(FE_OFN1241_n_4092), .o(g62418_sb) );
na02f02 TIMEBOOST_cell_36857 ( .a(TIMEBOOST_net_208), .b(FE_OCP_RBN2004_FE_OFN1026_n_16760), .o(TIMEBOOST_net_10667) );
na02m02 TIMEBOOST_cell_44227 ( .a(n_9635), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__Q), .o(TIMEBOOST_net_14352) );
na02s02 TIMEBOOST_cell_42002 ( .a(TIMEBOOST_net_13239), .b(g62415_sb), .o(n_6768) );
in01s01 g62419_u0 ( .a(FE_OFN1243_n_4092), .o(g62419_sb) );
na02s01 TIMEBOOST_cell_36859 ( .a(n_1954), .b(g61743_sb), .o(TIMEBOOST_net_10668) );
na02f02 TIMEBOOST_cell_44696 ( .a(TIMEBOOST_net_14586), .b(TIMEBOOST_net_6265), .o(n_9235) );
na02m02 TIMEBOOST_cell_32684 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__31__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__31__Q), .o(TIMEBOOST_net_10253) );
in01s01 g62420_u0 ( .a(FE_OFN1268_n_4095), .o(g62420_sb) );
na03m02 TIMEBOOST_cell_36861 ( .a(g52447_db), .b(n_4209), .c(g52447_sb), .o(TIMEBOOST_net_10669) );
na02m02 TIMEBOOST_cell_42120 ( .a(TIMEBOOST_net_13298), .b(FE_OFN1315_n_6624), .o(TIMEBOOST_net_11589) );
na02m02 TIMEBOOST_cell_41601 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_8__Q), .b(FE_OFN252_n_9868), .o(TIMEBOOST_net_13039) );
in01s01 g62421_u0 ( .a(n_6554), .o(g62421_sb) );
na02s01 TIMEBOOST_cell_36453 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(g65717_sb), .o(TIMEBOOST_net_10465) );
na02s01 TIMEBOOST_cell_3359 ( .a(TIMEBOOST_net_259), .b(n_3437), .o(n_4591) );
na02m02 TIMEBOOST_cell_45460 ( .a(TIMEBOOST_net_14968), .b(g58632_sb), .o(TIMEBOOST_net_14080) );
in01s01 g62422_u0 ( .a(FE_OFN1244_n_4092), .o(g62422_sb) );
na02s02 TIMEBOOST_cell_36863 ( .a(n_3848), .b(g63124_sb), .o(TIMEBOOST_net_10670) );
na02f02 TIMEBOOST_cell_41602 ( .a(FE_OFN1437_n_9372), .b(TIMEBOOST_net_13039), .o(TIMEBOOST_net_11681) );
na02m02 TIMEBOOST_cell_41603 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_7__Q), .b(FE_OFN250_n_9789), .o(TIMEBOOST_net_13040) );
in01s01 g62423_u0 ( .a(FE_OFN1224_n_6391), .o(g62423_sb) );
na02f02 TIMEBOOST_cell_3083 ( .a(TIMEBOOST_net_121), .b(n_15922), .o(n_15927) );
na02s01 TIMEBOOST_cell_37765 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__Q), .b(wbs_dat_i_4_), .o(TIMEBOOST_net_11121) );
na03f02 TIMEBOOST_cell_3084 ( .a(FE_RN_613_0), .b(FE_RN_615_0), .c(FE_RN_618_0), .o(TIMEBOOST_net_122) );
in01s01 g62424_u0 ( .a(FE_OFN1252_n_4143), .o(g62424_sb) );
na02s01 TIMEBOOST_cell_36865 ( .a(TIMEBOOST_net_266), .b(g61775_sb), .o(TIMEBOOST_net_10671) );
na03s02 TIMEBOOST_cell_34262 ( .a(TIMEBOOST_net_9813), .b(FE_OFN1174_n_5592), .c(g62107_sb), .o(n_5593) );
na02f02 TIMEBOOST_cell_32683 ( .a(FE_OFN1760_n_10780), .b(TIMEBOOST_net_10252), .o(TIMEBOOST_net_6511) );
in01s02 g62425_u0 ( .a(FE_OFN1311_n_6624), .o(g62425_sb) );
na02s02 TIMEBOOST_cell_37982 ( .a(TIMEBOOST_net_11229), .b(g54175_db), .o(n_13218) );
na02s02 TIMEBOOST_cell_43591 ( .a(n_7373), .b(n_4907), .o(TIMEBOOST_net_14034) );
na02s01 TIMEBOOST_cell_9081 ( .a(TIMEBOOST_net_1107), .b(n_4725), .o(TIMEBOOST_net_161) );
in01s01 g62426_u0 ( .a(FE_OFN1223_n_6391), .o(g62426_sb) );
na02f02 TIMEBOOST_cell_3085 ( .a(TIMEBOOST_net_122), .b(FE_RN_611_0), .o(FE_RN_619_0) );
in01s01 TIMEBOOST_cell_45868 ( .a(TIMEBOOST_net_15174), .o(TIMEBOOST_net_15175) );
na03s01 TIMEBOOST_cell_34248 ( .a(TIMEBOOST_net_9798), .b(FE_OFN1165_n_5615), .c(g62089_sb), .o(n_5618) );
in01s02 g62427_u0 ( .a(FE_OFN1316_n_6624), .o(g62427_sb) );
na02s01 TIMEBOOST_cell_36332 ( .a(TIMEBOOST_net_10404), .b(g65907_sb), .o(n_2174) );
na02s01 TIMEBOOST_cell_42971 ( .a(n_2308), .b(n_3108), .o(TIMEBOOST_net_13724) );
na02s01 TIMEBOOST_cell_40516 ( .a(TIMEBOOST_net_12496), .b(FE_OFN1301_n_5763), .o(TIMEBOOST_net_11504) );
in01s01 g62428_u0 ( .a(FE_OFN1224_n_6391), .o(g62428_sb) );
na03s02 TIMEBOOST_cell_34249 ( .a(TIMEBOOST_net_9797), .b(FE_OFN1174_n_5592), .c(g62141_sb), .o(n_5552) );
in01s01 TIMEBOOST_cell_45908 ( .a(TIMEBOOST_net_15214), .o(TIMEBOOST_net_15215) );
na02m02 TIMEBOOST_cell_32682 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__Q), .o(TIMEBOOST_net_10252) );
in01s01 g62429_u0 ( .a(FE_OFN1219_n_6886), .o(g62429_sb) );
na02s01 TIMEBOOST_cell_36867 ( .a(TIMEBOOST_net_268), .b(g61771_sb), .o(TIMEBOOST_net_10672) );
na02s01 TIMEBOOST_cell_45697 ( .a(n_3697), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__Q), .o(TIMEBOOST_net_15087) );
na02f02 TIMEBOOST_cell_44387 ( .a(n_9041), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__Q), .o(TIMEBOOST_net_14432) );
in01s01 g62430_u0 ( .a(FE_OFN1269_n_4095), .o(g62430_sb) );
na02s01 TIMEBOOST_cell_36869 ( .a(TIMEBOOST_net_270), .b(g61796_sb), .o(TIMEBOOST_net_10673) );
na02f02 TIMEBOOST_cell_43718 ( .a(TIMEBOOST_net_14097), .b(FE_OFN1381_n_8567), .o(TIMEBOOST_net_12842) );
na02m02 TIMEBOOST_cell_42564 ( .a(TIMEBOOST_net_13520), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_386), .o(TIMEBOOST_net_9851) );
in01s01 g62431_u0 ( .a(FE_OFN2063_n_6391), .o(g62431_sb) );
na03s02 TIMEBOOST_cell_36751 ( .a(g65252_da), .b(g65252_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__Q), .o(TIMEBOOST_net_10614) );
na02f02 TIMEBOOST_cell_3463 ( .a(TIMEBOOST_net_311), .b(FE_RN_702_0), .o(FE_RN_703_0) );
in01s01 g62432_u0 ( .a(FE_OFN1235_n_6391), .o(g62432_sb) );
na02s01 TIMEBOOST_cell_36389 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__Q), .b(g65923_sb), .o(TIMEBOOST_net_10433) );
na02m02 TIMEBOOST_cell_32388 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_30__Q), .o(TIMEBOOST_net_10105) );
na02s01 TIMEBOOST_cell_18487 ( .a(TIMEBOOST_net_4500), .b(g62741_sb), .o(n_5497) );
in01s01 g62433_u0 ( .a(FE_OFN1313_n_6624), .o(g62433_sb) );
na02m02 TIMEBOOST_cell_39354 ( .a(FE_OFN1150_n_13249), .b(TIMEBOOST_net_11915), .o(TIMEBOOST_net_4287) );
na02s02 TIMEBOOST_cell_3729 ( .a(TIMEBOOST_net_444), .b(FE_OFN264_n_9849), .o(n_9850) );
na02s01 TIMEBOOST_cell_40517 ( .a(wishbone_slave_unit_pcim_sm_data_in_659), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__Q), .o(TIMEBOOST_net_12497) );
in01s01 g62434_u0 ( .a(n_6554), .o(g62434_sb) );
na02s01 TIMEBOOST_cell_36445 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(g65778_sb), .o(TIMEBOOST_net_10461) );
na02f01 TIMEBOOST_cell_3361 ( .a(TIMEBOOST_net_260), .b(n_3335), .o(n_3498) );
na03f02 TIMEBOOST_cell_36095 ( .a(n_10634), .b(FE_RN_474_0), .c(n_12574), .o(n_12836) );
in01s01 g62435_u0 ( .a(n_6645), .o(g62435_sb) );
na02s01 TIMEBOOST_cell_36379 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__Q), .b(g65853_sb), .o(TIMEBOOST_net_10428) );
na02s02 TIMEBOOST_cell_44416 ( .a(TIMEBOOST_net_14446), .b(FE_OFN1306_n_13124), .o(TIMEBOOST_net_13420) );
na02s02 TIMEBOOST_cell_3364 ( .a(n_2426), .b(n_2433), .o(TIMEBOOST_net_262) );
in01s01 g62436_u0 ( .a(FE_OFN1241_n_4092), .o(g62436_sb) );
na02s01 TIMEBOOST_cell_36871 ( .a(TIMEBOOST_net_272), .b(g61779_sb), .o(TIMEBOOST_net_10674) );
na02m04 TIMEBOOST_cell_31878 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_385), .b(TIMEBOOST_net_1820), .o(TIMEBOOST_net_9850) );
na02m02 TIMEBOOST_cell_32504 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__13__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__13__Q), .o(TIMEBOOST_net_10163) );
in01s01 g62437_u0 ( .a(FE_OFN1283_n_4097), .o(g62437_sb) );
na02s01 TIMEBOOST_cell_36873 ( .a(TIMEBOOST_net_274), .b(g61767_sb), .o(TIMEBOOST_net_10675) );
na02m02 TIMEBOOST_cell_42565 ( .a(n_8884), .b(wbu_addr_in_250), .o(TIMEBOOST_net_13521) );
na02f02 TIMEBOOST_cell_32681 ( .a(FE_OFN1760_n_10780), .b(TIMEBOOST_net_10251), .o(TIMEBOOST_net_6510) );
in01s01 g62438_u0 ( .a(FE_OFN1241_n_4092), .o(g62438_sb) );
na02s01 TIMEBOOST_cell_36875 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__Q), .b(g58297_sb), .o(TIMEBOOST_net_10676) );
na02s02 TIMEBOOST_cell_41701 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_33__Q), .b(FE_OFN2054_n_8831), .o(TIMEBOOST_net_13089) );
na02m02 TIMEBOOST_cell_44242 ( .a(TIMEBOOST_net_14359), .b(FE_OFN1401_n_8567), .o(TIMEBOOST_net_12792) );
in01s02 g62439_u0 ( .a(FE_OFN1310_n_6624), .o(g62439_sb) );
na02s01 TIMEBOOST_cell_36252 ( .a(TIMEBOOST_net_10364), .b(FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_1008) );
na03s02 TIMEBOOST_cell_40691 ( .a(n_4312), .b(n_4313), .c(FE_OFN1246_n_4093), .o(TIMEBOOST_net_12584) );
na02s01 TIMEBOOST_cell_40518 ( .a(TIMEBOOST_net_12497), .b(FE_OFN1301_n_5763), .o(TIMEBOOST_net_11516) );
in01s01 g62440_u0 ( .a(FE_OFN1278_n_4097), .o(g62440_sb) );
na02s03 TIMEBOOST_cell_3089 ( .a(TIMEBOOST_net_124), .b(g58773_sb), .o(n_9856) );
na03s02 TIMEBOOST_cell_37593 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__Q), .b(FE_OFN2256_n_8060), .c(n_2193), .o(TIMEBOOST_net_11035) );
na02f02 TIMEBOOST_cell_42322 ( .a(TIMEBOOST_net_13399), .b(g57166_sb), .o(n_10459) );
in01s01 g62441_u0 ( .a(FE_OFN2064_n_6391), .o(g62441_sb) );
na02s01 TIMEBOOST_cell_36449 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__Q), .b(FE_OFN575_n_9902), .o(TIMEBOOST_net_10463) );
na02s02 TIMEBOOST_cell_3467 ( .a(TIMEBOOST_net_313), .b(n_3337), .o(n_4080) );
na02s01 TIMEBOOST_cell_40520 ( .a(TIMEBOOST_net_12498), .b(FE_OFN1299_n_5763), .o(TIMEBOOST_net_11519) );
in01s01 g62442_u0 ( .a(FE_OFN1261_n_4143), .o(g62442_sb) );
no02f04 TIMEBOOST_cell_36877 ( .a(FE_RN_396_0), .b(FE_OFN1710_n_4868), .o(TIMEBOOST_net_10677) );
na02s01 TIMEBOOST_cell_42598 ( .a(TIMEBOOST_net_13537), .b(g61705_sb), .o(TIMEBOOST_net_10991) );
na02s02 TIMEBOOST_cell_45461 ( .a(TIMEBOOST_net_4796), .b(FE_OFN1200_n_4090), .o(TIMEBOOST_net_14969) );
in01s01 g62443_u0 ( .a(FE_OFN1247_n_4093), .o(g62443_sb) );
na02s02 TIMEBOOST_cell_42711 ( .a(pci_target_unit_fifos_pcir_data_in), .b(g65748_sb), .o(TIMEBOOST_net_13594) );
na03s02 TIMEBOOST_cell_13817 ( .a(FE_OFN235_n_9834), .b(g58188_sb), .c(g58188_db), .o(n_9596) );
na03s02 TIMEBOOST_cell_33247 ( .a(FE_OFN227_n_9841), .b(g57993_sb), .c(g57993_db), .o(n_9802) );
in01s02 g62444_u0 ( .a(FE_OFN1323_n_6436), .o(g62444_sb) );
na02m02 TIMEBOOST_cell_43977 ( .a(n_9039), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__Q), .o(TIMEBOOST_net_14227) );
na02f02 TIMEBOOST_cell_43978 ( .a(TIMEBOOST_net_14227), .b(FE_OFN1377_n_8567), .o(TIMEBOOST_net_12964) );
na02s02 TIMEBOOST_cell_32214 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_772), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_7__Q), .o(TIMEBOOST_net_10018) );
in01s01 g62445_u0 ( .a(FE_OFN1212_n_4151), .o(g62445_sb) );
na02s02 TIMEBOOST_cell_36881 ( .a(n_1904), .b(g61858_sb), .o(TIMEBOOST_net_10679) );
na02s02 TIMEBOOST_cell_39868 ( .a(TIMEBOOST_net_12172), .b(g62475_sb), .o(n_6639) );
na02s02 TIMEBOOST_cell_45094 ( .a(TIMEBOOST_net_14785), .b(g64316_da), .o(TIMEBOOST_net_11332) );
in01s02 g62446_u0 ( .a(FE_OFN1311_n_6624), .o(g62446_sb) );
na02m02 TIMEBOOST_cell_44523 ( .a(n_9220), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__Q), .o(TIMEBOOST_net_14500) );
na02m02 TIMEBOOST_cell_43979 ( .a(n_9434), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q), .o(TIMEBOOST_net_14228) );
na02s01 TIMEBOOST_cell_42823 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__Q), .b(g65317_sb), .o(TIMEBOOST_net_13650) );
in01s01 g62447_u0 ( .a(n_6431), .o(g62447_sb) );
na02f02 TIMEBOOST_cell_43980 ( .a(TIMEBOOST_net_14228), .b(FE_OFN1409_n_8567), .o(TIMEBOOST_net_12978) );
na02s02 TIMEBOOST_cell_36883 ( .a(n_1858), .b(g61859_sb), .o(TIMEBOOST_net_10680) );
na02m02 TIMEBOOST_cell_38882 ( .a(TIMEBOOST_net_11679), .b(g58473_sb), .o(n_9371) );
in01s01 g62448_u0 ( .a(FE_OFN1215_n_4151), .o(g62448_sb) );
na02f06 TIMEBOOST_cell_36887 ( .a(TIMEBOOST_net_893), .b(n_16438), .o(TIMEBOOST_net_10682) );
na02s01 TIMEBOOST_cell_38356 ( .a(TIMEBOOST_net_11416), .b(g62829_sb), .o(n_5318) );
no02f06 TIMEBOOST_cell_20069 ( .a(TIMEBOOST_net_5291), .b(FE_RN_124_0), .o(TIMEBOOST_net_944) );
in01s01 g62449_u0 ( .a(FE_OFN1293_n_4098), .o(g62449_sb) );
na02s02 TIMEBOOST_cell_36885 ( .a(n_1902), .b(g61863_sb), .o(TIMEBOOST_net_10681) );
na02s02 TIMEBOOST_cell_39870 ( .a(TIMEBOOST_net_12173), .b(g62472_sb), .o(n_6647) );
na03s02 TIMEBOOST_cell_34282 ( .a(TIMEBOOST_net_4178), .b(g52629_sb), .c(n_8757), .o(g52443_db) );
in01s01 g62450_u0 ( .a(FE_OFN1222_n_6391), .o(g62450_sb) );
na02s02 TIMEBOOST_cell_3091 ( .a(TIMEBOOST_net_125), .b(g58788_sb), .o(n_9834) );
na03s01 TIMEBOOST_cell_37681 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q), .b(FE_OFN699_n_7845), .c(n_2151), .o(TIMEBOOST_net_11079) );
na03s02 TIMEBOOST_cell_41971 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__Q), .b(n_3583), .c(FE_OFN1214_n_4151), .o(TIMEBOOST_net_13224) );
in01s02 g62451_u0 ( .a(FE_OFN1317_n_6624), .o(g62451_sb) );
na02f02 TIMEBOOST_cell_43981 ( .a(n_9084), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__Q), .o(TIMEBOOST_net_14229) );
na02f02 TIMEBOOST_cell_44258 ( .a(TIMEBOOST_net_14367), .b(FE_OFN1400_n_8567), .o(TIMEBOOST_net_12890) );
na03s02 TIMEBOOST_cell_34795 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__Q), .b(g63154_sb), .c(g63154_db), .o(n_5833) );
in01s01 g62452_u0 ( .a(FE_OFN1285_n_4097), .o(g62452_sb) );
na02m02 g52447_u2 ( .a(n_14839), .b(n_14750), .o(g52447_db) );
na02s01 TIMEBOOST_cell_41897 ( .a(configuration_wb_err_addr_553), .b(conf_wb_err_addr_in_962), .o(TIMEBOOST_net_13187) );
in01s01 g62453_u0 ( .a(FE_OFN1319_n_6436), .o(g62453_sb) );
na02f02 TIMEBOOST_cell_43982 ( .a(TIMEBOOST_net_14229), .b(FE_OFN1397_n_8567), .o(TIMEBOOST_net_12954) );
na02s01 TIMEBOOST_cell_36254 ( .a(TIMEBOOST_net_10365), .b(wishbone_slave_unit_pci_initiator_if_read_count_3_), .o(TIMEBOOST_net_259) );
na02f02 TIMEBOOST_cell_36922 ( .a(TIMEBOOST_net_10699), .b(g52601_sb), .o(n_10263) );
in01s01 g62454_u0 ( .a(FE_OFN1208_n_6356), .o(g62454_sb) );
na02m02 TIMEBOOST_cell_44337 ( .a(n_9757), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__Q), .o(TIMEBOOST_net_14407) );
na02s01 TIMEBOOST_cell_38358 ( .a(TIMEBOOST_net_11417), .b(g63018_sb), .o(n_5212) );
na02s01 TIMEBOOST_cell_42797 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(g64091_sb), .o(TIMEBOOST_net_13637) );
in01s01 g62455_u0 ( .a(FE_OFN1232_n_6391), .o(g62455_sb) );
na02m04 TIMEBOOST_cell_20634 ( .a(FE_RN_578_0), .b(FE_OFN1946_n_13784), .o(TIMEBOOST_net_5574) );
na02s01 TIMEBOOST_cell_18615 ( .a(TIMEBOOST_net_4564), .b(g63103_sb), .o(n_5048) );
na02s01 TIMEBOOST_cell_40522 ( .a(TIMEBOOST_net_12499), .b(FE_OFN1299_n_5763), .o(TIMEBOOST_net_11518) );
in01s01 g62456_u0 ( .a(FE_OFN1193_n_6935), .o(g62456_sb) );
na02s01 TIMEBOOST_cell_3093 ( .a(TIMEBOOST_net_126), .b(g58798_sb), .o(n_9825) );
na03s02 TIMEBOOST_cell_37683 ( .a(n_2192), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__Q), .c(FE_OFN2081_n_8176), .o(TIMEBOOST_net_11080) );
na02f02 TIMEBOOST_cell_44222 ( .a(TIMEBOOST_net_14349), .b(FE_OFN1413_n_8567), .o(TIMEBOOST_net_12854) );
in01s01 g62457_u0 ( .a(FE_OFN2063_n_6391), .o(g62457_sb) );
na02s01 TIMEBOOST_cell_36381 ( .a(n_2651), .b(g65999_db), .o(TIMEBOOST_net_10429) );
no02m02 TIMEBOOST_cell_3471 ( .a(TIMEBOOST_net_315), .b(n_7715), .o(g59232_p) );
na02s02 TIMEBOOST_cell_9003 ( .a(TIMEBOOST_net_1068), .b(n_294), .o(n_13548) );
in01s01 g62458_u0 ( .a(FE_OFN1212_n_4151), .o(g62458_sb) );
na02f06 TIMEBOOST_cell_36833 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_), .b(g75160_sb), .o(TIMEBOOST_net_10655) );
na03f02 TIMEBOOST_cell_2511 ( .a(n_9852), .b(g57078_sb), .c(g57078_db), .o(n_11665) );
na02s02 TIMEBOOST_cell_45667 ( .a(TIMEBOOST_net_859), .b(g61976_db), .o(TIMEBOOST_net_15072) );
in01s01 g62459_u0 ( .a(FE_OFN1285_n_4097), .o(g62459_sb) );
na02s02 TIMEBOOST_cell_36811 ( .a(n_3839), .b(g63036_sb), .o(TIMEBOOST_net_10644) );
na03f02 TIMEBOOST_cell_2513 ( .a(n_9109), .b(g57117_sb), .c(g57117_db), .o(n_10477) );
na03f02 TIMEBOOST_cell_2514 ( .a(n_9785), .b(g57140_sb), .c(g57140_db), .o(n_11609) );
in01s01 g62460_u0 ( .a(FE_OFN1225_n_6391), .o(g62460_sb) );
na02f02 TIMEBOOST_cell_3095 ( .a(TIMEBOOST_net_127), .b(n_2378), .o(n_4680) );
na03s02 TIMEBOOST_cell_37625 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__Q), .b(FE_OFN707_n_8119), .c(n_1931), .o(TIMEBOOST_net_11051) );
na02m02 TIMEBOOST_cell_32680 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__Q), .o(TIMEBOOST_net_10251) );
in01s01 g62461_u0 ( .a(FE_OFN1232_n_6391), .o(g62461_sb) );
na02s02 TIMEBOOST_cell_36813 ( .a(n_4005), .b(g62833_db), .o(TIMEBOOST_net_10645) );
na02s01 TIMEBOOST_cell_3473 ( .a(TIMEBOOST_net_316), .b(g64255_sb), .o(n_3918) );
na02s01 TIMEBOOST_cell_43316 ( .a(TIMEBOOST_net_13896), .b(g62500_sb), .o(n_6582) );
in01s01 g62462_u0 ( .a(FE_OFN1204_n_4090), .o(g62462_sb) );
in01s01 TIMEBOOST_cell_45938 ( .a(TIMEBOOST_net_15244), .o(TIMEBOOST_net_15245) );
na02s01 TIMEBOOST_cell_42026 ( .a(TIMEBOOST_net_13251), .b(g62649_sb), .o(n_6249) );
na03s02 TIMEBOOST_cell_41981 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__17__Q), .b(n_4503), .c(FE_OFN1261_n_4143), .o(TIMEBOOST_net_13229) );
in01s01 g62463_u0 ( .a(FE_OFN1294_n_4098), .o(g62463_sb) );
na02s01 TIMEBOOST_cell_36823 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_384), .b(g53947_da), .o(TIMEBOOST_net_10650) );
na03f02 TIMEBOOST_cell_2515 ( .a(n_9101), .b(g57153_sb), .c(g57153_db), .o(n_10463) );
na02s02 TIMEBOOST_cell_20085 ( .a(TIMEBOOST_net_5299), .b(g62966_sb), .o(n_5950) );
in01s01 g62464_u0 ( .a(FE_OFN1213_n_4151), .o(g62464_sb) );
na02f02 TIMEBOOST_cell_37067 ( .a(n_13987), .b(TIMEBOOST_net_10222), .o(TIMEBOOST_net_10772) );
na02f02 TIMEBOOST_cell_41604 ( .a(FE_OFN1440_n_9372), .b(TIMEBOOST_net_13040), .o(TIMEBOOST_net_11672) );
na02f02 TIMEBOOST_cell_39006 ( .a(TIMEBOOST_net_11741), .b(g52531_sb), .o(n_13792) );
in01s01 g62465_u0 ( .a(FE_OFN1235_n_6391), .o(g62465_sb) );
na02s01 TIMEBOOST_cell_36439 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__Q), .b(FE_OFN577_n_9902), .o(TIMEBOOST_net_10458) );
na02s01 TIMEBOOST_cell_3475 ( .a(TIMEBOOST_net_317), .b(g65905_sb), .o(n_3207) );
na02s03 TIMEBOOST_cell_3476 ( .a(pci_target_unit_del_sync_comp_cycle_count_14_), .b(pci_target_unit_del_sync_comp_cycle_count_15_), .o(TIMEBOOST_net_318) );
in01s01 g62466_u0 ( .a(FE_OFN1219_n_6886), .o(g62466_sb) );
na02f02 TIMEBOOST_cell_37071 ( .a(n_13987), .b(TIMEBOOST_net_10225), .o(TIMEBOOST_net_10774) );
na02m02 TIMEBOOST_cell_44665 ( .a(n_9226), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__Q), .o(TIMEBOOST_net_14571) );
in01s01 g62467_u0 ( .a(FE_OFN1260_n_4143), .o(g62467_sb) );
na02f02 TIMEBOOST_cell_36815 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_796), .b(g54321_sb), .o(TIMEBOOST_net_10646) );
na02s01 TIMEBOOST_cell_38548 ( .a(TIMEBOOST_net_11512), .b(g62062_sb), .o(n_7747) );
na02s01 TIMEBOOST_cell_43250 ( .a(TIMEBOOST_net_13863), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_11546) );
in01s01 g62468_u0 ( .a(FE_OFN1193_n_6935), .o(g62468_sb) );
no02f02 TIMEBOOST_cell_3097 ( .a(TIMEBOOST_net_128), .b(FE_RN_682_0), .o(FE_RN_683_0) );
na02s01 g62468_u2 ( .a(n_3729), .b(n_6935), .o(g62468_db) );
na02s02 TIMEBOOST_cell_45462 ( .a(TIMEBOOST_net_14969), .b(g63094_sb), .o(n_5856) );
in01s01 g62469_u0 ( .a(FE_OFN2064_n_6391), .o(g62469_sb) );
na02f02 TIMEBOOST_cell_37107 ( .a(FE_RN_143_0), .b(n_10865), .o(TIMEBOOST_net_10792) );
na02s02 TIMEBOOST_cell_3477 ( .a(TIMEBOOST_net_318), .b(n_3025), .o(n_3463) );
na02s03 TIMEBOOST_cell_3478 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__Q), .o(TIMEBOOST_net_319) );
in01s01 g62470_u0 ( .a(FE_OFN1208_n_6356), .o(g62470_sb) );
na02f02 TIMEBOOST_cell_37057 ( .a(TIMEBOOST_net_10128), .b(n_13891), .o(TIMEBOOST_net_10767) );
na02m02 TIMEBOOST_cell_39162 ( .a(TIMEBOOST_net_11819), .b(wbu_addr_in_256), .o(n_9789) );
na02m02 TIMEBOOST_cell_43983 ( .a(n_9668), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__Q), .o(TIMEBOOST_net_14230) );
in01s01 g62471_u0 ( .a(FE_OFN1261_n_4143), .o(g62471_sb) );
na02s01 TIMEBOOST_cell_36817 ( .a(n_1567), .b(g61939_sb), .o(TIMEBOOST_net_10647) );
na03s02 TIMEBOOST_cell_36837 ( .a(TIMEBOOST_net_4082), .b(g65389_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__Q), .o(TIMEBOOST_net_10657) );
na02s01 TIMEBOOST_cell_36256 ( .a(TIMEBOOST_net_10366), .b(n_550), .o(n_1382) );
in01s01 g62472_u0 ( .a(n_6645), .o(g62472_sb) );
na02s02 TIMEBOOST_cell_36819 ( .a(wishbone_slave_unit_pcim_if_wbw_cbe_in_417), .b(g53944_da), .o(TIMEBOOST_net_10648) );
na02m02 TIMEBOOST_cell_3365 ( .a(TIMEBOOST_net_262), .b(n_2441), .o(n_2434) );
na02f02 TIMEBOOST_cell_41518 ( .a(TIMEBOOST_net_12997), .b(g57567_sb), .o(n_11186) );
in01s01 g62473_u0 ( .a(FE_OFN1234_n_6391), .o(g62473_sb) );
na02s01 TIMEBOOST_cell_36829 ( .a(n_4399), .b(g62607_sb), .o(TIMEBOOST_net_10653) );
na02m04 TIMEBOOST_cell_3479 ( .a(TIMEBOOST_net_319), .b(n_3074), .o(n_3462) );
na02f01 TIMEBOOST_cell_3480 ( .a(n_16485), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q), .o(TIMEBOOST_net_320) );
in01s01 g62474_u0 ( .a(FE_OFN1275_n_4096), .o(g62474_sb) );
no02f02 TIMEBOOST_cell_3099 ( .a(TIMEBOOST_net_129), .b(FE_RN_689_0), .o(FE_RN_691_0) );
na03s02 TIMEBOOST_cell_37627 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__Q), .b(FE_OFN707_n_8119), .c(n_1932), .o(TIMEBOOST_net_11052) );
na02s01 TIMEBOOST_cell_42635 ( .a(n_3761), .b(g65018_sb), .o(TIMEBOOST_net_13556) );
in01s01 g62475_u0 ( .a(n_6319), .o(g62475_sb) );
na02s01 TIMEBOOST_cell_42599 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(g65684_sb), .o(TIMEBOOST_net_13538) );
na02s01 TIMEBOOST_cell_16109 ( .a(TIMEBOOST_net_3311), .b(g65697_sb), .o(n_2204) );
in01s01 g62476_u0 ( .a(FE_OFN1206_n_6356), .o(g62476_sb) );
no02f02 TIMEBOOST_cell_3101 ( .a(TIMEBOOST_net_130), .b(FE_RN_636_0), .o(FE_RN_641_0) );
na03s02 TIMEBOOST_cell_37629 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__Q), .b(FE_OFN713_n_8140), .c(n_1947), .o(TIMEBOOST_net_11053) );
na02s01 TIMEBOOST_cell_45668 ( .a(TIMEBOOST_net_15072), .b(g63604_da), .o(n_7168) );
in01s02 g62477_u0 ( .a(FE_OFN1311_n_6624), .o(g62477_sb) );
na02s02 TIMEBOOST_cell_43424 ( .a(TIMEBOOST_net_13950), .b(n_6232), .o(TIMEBOOST_net_12190) );
na02s01 TIMEBOOST_cell_37984 ( .a(TIMEBOOST_net_11230), .b(g63025_db), .o(n_5196) );
na02f02 TIMEBOOST_cell_45463 ( .a(n_7329), .b(TIMEBOOST_net_600), .o(TIMEBOOST_net_14970) );
in01s01 g62478_u0 ( .a(n_6232), .o(g62478_sb) );
na02s02 TIMEBOOST_cell_36827 ( .a(wishbone_slave_unit_pcim_if_wbw_cbe_in_416), .b(g53943_da), .o(TIMEBOOST_net_10652) );
na02s01 TIMEBOOST_cell_39872 ( .a(TIMEBOOST_net_12174), .b(g62979_sb), .o(n_5924) );
no02m02 TIMEBOOST_cell_3370 ( .a(n_15929), .b(n_15924), .o(TIMEBOOST_net_265) );
in01s01 g62479_u0 ( .a(FE_OFN1222_n_6391), .o(g62479_sb) );
na02f02 TIMEBOOST_cell_3103 ( .a(TIMEBOOST_net_131), .b(n_2238), .o(n_2954) );
na02s03 TIMEBOOST_cell_3104 ( .a(n_2244), .b(wbu_addr_in_251), .o(TIMEBOOST_net_132) );
in01s01 g62480_u0 ( .a(FE_OFN1222_n_6391), .o(g62480_sb) );
na02m04 TIMEBOOST_cell_3105 ( .a(TIMEBOOST_net_132), .b(n_1362), .o(n_2716) );
na03s02 TIMEBOOST_cell_37633 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__Q), .b(FE_OFN702_n_7845), .c(n_1920), .o(TIMEBOOST_net_11055) );
na02s02 TIMEBOOST_cell_3106 ( .a(n_2244), .b(n_2225), .o(TIMEBOOST_net_133) );
in01s02 g62481_u0 ( .a(FE_OFN1317_n_6624), .o(g62481_sb) );
na02f02 TIMEBOOST_cell_12678 ( .a(n_13903), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__Q), .o(TIMEBOOST_net_2906) );
na02f02 TIMEBOOST_cell_43984 ( .a(TIMEBOOST_net_14230), .b(FE_OFN1374_n_8567), .o(TIMEBOOST_net_12921) );
na02f02 TIMEBOOST_cell_37813 ( .a(g54333_sb), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_777), .o(TIMEBOOST_net_11145) );
in01s01 g62482_u0 ( .a(FE_OFN1288_n_4098), .o(g62482_sb) );
na02s02 TIMEBOOST_cell_36805 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_66), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_10641) );
na02s01 TIMEBOOST_cell_43251 ( .a(n_4295), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__Q), .o(TIMEBOOST_net_13864) );
na02f02 TIMEBOOST_cell_44388 ( .a(TIMEBOOST_net_14432), .b(FE_OFN1405_n_8567), .o(TIMEBOOST_net_12762) );
in01s01 g62483_u0 ( .a(FE_OFN1293_n_4098), .o(g62483_sb) );
na02s02 TIMEBOOST_cell_37164 ( .a(TIMEBOOST_net_10820), .b(TIMEBOOST_net_19), .o(n_5769) );
na02m02 TIMEBOOST_cell_43985 ( .a(n_9058), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__Q), .o(TIMEBOOST_net_14231) );
na02m02 TIMEBOOST_cell_44233 ( .a(n_9224), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__Q), .o(TIMEBOOST_net_14355) );
in01s02 g62484_u0 ( .a(FE_OFN1317_n_6624), .o(g62484_sb) );
na02f02 TIMEBOOST_cell_43986 ( .a(TIMEBOOST_net_14231), .b(FE_OFN1368_n_8567), .o(TIMEBOOST_net_12920) );
na02s01 TIMEBOOST_cell_43425 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__Q), .b(n_4437), .o(TIMEBOOST_net_13951) );
na02s01 TIMEBOOST_cell_15794 ( .a(parchk_pci_ad_reg_in_1235), .b(g67050_db), .o(TIMEBOOST_net_3154) );
in01s01 g62485_u0 ( .a(FE_OFN1258_n_4143), .o(g62485_sb) );
na02s02 TIMEBOOST_cell_36821 ( .a(wishbone_slave_unit_pcim_if_wbw_cbe_in), .b(g53945_da), .o(TIMEBOOST_net_10649) );
na02s01 TIMEBOOST_cell_42656 ( .a(TIMEBOOST_net_13566), .b(FE_OFN2108_n_2047), .o(TIMEBOOST_net_11888) );
na02s02 TIMEBOOST_cell_43516 ( .a(TIMEBOOST_net_13996), .b(FE_OFN1235_n_6391), .o(TIMEBOOST_net_12147) );
in01s02 g62486_u0 ( .a(FE_OFN1317_n_6624), .o(g62486_sb) );
na02s02 TIMEBOOST_cell_16971 ( .a(TIMEBOOST_net_3742), .b(g65247_sb), .o(n_2635) );
na02m02 TIMEBOOST_cell_43987 ( .a(n_9475), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__Q), .o(TIMEBOOST_net_14232) );
na04s02 TIMEBOOST_cell_34237 ( .a(g63566_da), .b(g63566_db), .c(g61963_sb), .d(g61963_db), .o(n_6948) );
in01s01 g62487_u0 ( .a(FE_OFN1268_n_4095), .o(g62487_sb) );
na02s02 TIMEBOOST_cell_37166 ( .a(TIMEBOOST_net_10821), .b(n_1993), .o(TIMEBOOST_net_136) );
na02s02 TIMEBOOST_cell_42982 ( .a(TIMEBOOST_net_13729), .b(g61822_sb), .o(n_8144) );
na02s02 TIMEBOOST_cell_43426 ( .a(TIMEBOOST_net_13951), .b(n_6232), .o(TIMEBOOST_net_11572) );
in01s01 g62488_u0 ( .a(FE_OFN1294_n_4098), .o(g62488_sb) );
na02s02 TIMEBOOST_cell_36825 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in), .b(TIMEBOOST_net_883), .o(TIMEBOOST_net_10651) );
na02s02 TIMEBOOST_cell_38360 ( .a(TIMEBOOST_net_11418), .b(g62795_sb), .o(n_5396) );
na02s02 TIMEBOOST_cell_39874 ( .a(TIMEBOOST_net_12175), .b(g62644_sb), .o(n_6261) );
in01s01 g62489_u0 ( .a(FE_OFN1193_n_6935), .o(g62489_sb) );
na02f02 TIMEBOOST_cell_3107 ( .a(TIMEBOOST_net_133), .b(n_2243), .o(n_2712) );
na03s02 TIMEBOOST_cell_37635 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__Q), .b(FE_OFN699_n_7845), .c(n_1928), .o(TIMEBOOST_net_11056) );
na02s01 TIMEBOOST_cell_31243 ( .a(TIMEBOOST_net_9532), .b(g64955_sb), .o(n_3663) );
in01s01 g62490_u0 ( .a(FE_OFN1248_n_4093), .o(g62490_sb) );
na02m04 TIMEBOOST_cell_3109 ( .a(TIMEBOOST_net_134), .b(n_2238), .o(n_2714) );
na02s04 TIMEBOOST_cell_45820 ( .a(TIMEBOOST_net_15148), .b(FE_OFN2135_n_13124), .o(TIMEBOOST_net_14990) );
in01s01 g62491_u0 ( .a(n_6232), .o(g62491_sb) );
na02s01 TIMEBOOST_cell_17745 ( .a(TIMEBOOST_net_4129), .b(g61937_sb), .o(n_7949) );
no02m04 TIMEBOOST_cell_3371 ( .a(n_15324), .b(TIMEBOOST_net_265), .o(n_15325) );
na02s01 TIMEBOOST_cell_42636 ( .a(TIMEBOOST_net_13556), .b(g65018_db), .o(n_3633) );
in01s01 g62492_u0 ( .a(FE_OFN1241_n_4092), .o(g62492_sb) );
na03s02 TIMEBOOST_cell_36783 ( .a(g64367_da), .b(g64367_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__Q), .o(TIMEBOOST_net_10630) );
na02s02 TIMEBOOST_cell_40702 ( .a(TIMEBOOST_net_12589), .b(g62340_sb), .o(n_6919) );
na02s01 TIMEBOOST_cell_44881 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__Q), .b(g65809_sb), .o(TIMEBOOST_net_14679) );
in01s01 g62493_u0 ( .a(n_6554), .o(g62493_sb) );
na02f02 TIMEBOOST_cell_37061 ( .a(FE_RN_230_0), .b(n_10885), .o(TIMEBOOST_net_10769) );
na02m02 TIMEBOOST_cell_10170 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__Q), .b(n_13447), .o(TIMEBOOST_net_1652) );
na02f08 TIMEBOOST_cell_15899 ( .a(TIMEBOOST_net_3206), .b(output_backup_trdy_out_reg_Q), .o(n_1192) );
in01s01 g62494_u0 ( .a(FE_OFN1276_n_4096), .o(g62494_sb) );
na02s01 TIMEBOOST_cell_3111 ( .a(TIMEBOOST_net_135), .b(n_2708), .o(n_2709) );
na02m04 TIMEBOOST_cell_45821 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_785), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_20__Q), .o(TIMEBOOST_net_15149) );
na02s01 TIMEBOOST_cell_43252 ( .a(TIMEBOOST_net_13864), .b(FE_OFN1250_n_4093), .o(TIMEBOOST_net_12525) );
in01s01 g62495_u0 ( .a(n_6287), .o(g62495_sb) );
na02s02 TIMEBOOST_cell_3591 ( .a(TIMEBOOST_net_375), .b(FE_OFN268_n_9880), .o(n_9639) );
na02f02 TIMEBOOST_cell_12642 ( .a(FE_OFN1771_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__Q), .o(TIMEBOOST_net_2888) );
na02f02 TIMEBOOST_cell_42520 ( .a(TIMEBOOST_net_13498), .b(g57594_sb), .o(n_11159) );
in01s01 g62496_u0 ( .a(FE_OFN1249_n_4093), .o(g62496_sb) );
na02f02 TIMEBOOST_cell_37053 ( .a(TIMEBOOST_net_10124), .b(n_13891), .o(TIMEBOOST_net_10765) );
na02s01 TIMEBOOST_cell_44857 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__Q), .b(FE_OFN1657_n_9502), .o(TIMEBOOST_net_14667) );
na03f02 TIMEBOOST_cell_2540 ( .a(n_9004), .b(g57543_sb), .c(g57543_db), .o(n_10310) );
in01s01 g62497_u0 ( .a(FE_OFN1249_n_4093), .o(g62497_sb) );
na02f02 TIMEBOOST_cell_37037 ( .a(FE_OFN1771_n_14054), .b(TIMEBOOST_net_10143), .o(TIMEBOOST_net_10757) );
na02s02 TIMEBOOST_cell_39876 ( .a(TIMEBOOST_net_12176), .b(g62926_sb), .o(n_6029) );
na02s02 TIMEBOOST_cell_45669 ( .a(TIMEBOOST_net_858), .b(g61972_db), .o(TIMEBOOST_net_15073) );
in01s01 g62498_u0 ( .a(FE_OFN1313_n_6624), .o(g62498_sb) );
na02s02 TIMEBOOST_cell_16969 ( .a(TIMEBOOST_net_3741), .b(g65237_sb), .o(n_2646) );
na02f02 TIMEBOOST_cell_43988 ( .a(TIMEBOOST_net_14232), .b(FE_OFN1415_n_8567), .o(TIMEBOOST_net_12955) );
na02f02 TIMEBOOST_cell_41320 ( .a(TIMEBOOST_net_12898), .b(g57149_sb), .o(n_11601) );
in01s01 g62499_u0 ( .a(FE_OFN1253_n_4143), .o(g62499_sb) );
na02f02 TIMEBOOST_cell_37039 ( .a(FE_OFN1771_n_14054), .b(TIMEBOOST_net_10138), .o(TIMEBOOST_net_10758) );
na02f02 TIMEBOOST_cell_44524 ( .a(TIMEBOOST_net_14500), .b(FE_OFN2174_n_8567), .o(TIMEBOOST_net_13456) );
na02m02 TIMEBOOST_cell_43989 ( .a(n_9732), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q), .o(TIMEBOOST_net_14233) );
in01s01 g62500_u0 ( .a(FE_OFN1274_n_4096), .o(g62500_sb) );
na02s02 TIMEBOOST_cell_3113 ( .a(TIMEBOOST_net_136), .b(n_1630), .o(n_1994) );
na03s02 TIMEBOOST_cell_37641 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__Q), .b(FE_OFN710_n_8232), .c(n_1867), .o(TIMEBOOST_net_11059) );
na03f02 TIMEBOOST_cell_36094 ( .a(FE_OFN1746_n_12004), .b(TIMEBOOST_net_10200), .c(n_12010), .o(n_12521) );
in01s01 g62501_u0 ( .a(FE_OFN1310_n_6624), .o(g62501_sb) );
na02f02 TIMEBOOST_cell_43990 ( .a(TIMEBOOST_net_14233), .b(FE_OFN1385_n_8567), .o(TIMEBOOST_net_12883) );
na02f02 TIMEBOOST_cell_44210 ( .a(TIMEBOOST_net_14343), .b(FE_OFN1405_n_8567), .o(TIMEBOOST_net_12986) );
na02s02 TIMEBOOST_cell_44434 ( .a(TIMEBOOST_net_14455), .b(FE_OFN1305_n_13124), .o(TIMEBOOST_net_13416) );
in01s01 g62502_u0 ( .a(FE_OFN1295_n_4098), .o(g62502_sb) );
na02f02 TIMEBOOST_cell_37041 ( .a(TIMEBOOST_net_10125), .b(n_13891), .o(TIMEBOOST_net_10759) );
na02s02 TIMEBOOST_cell_39878 ( .a(TIMEBOOST_net_12177), .b(g62654_sb), .o(n_6235) );
na02s02 TIMEBOOST_cell_39880 ( .a(TIMEBOOST_net_12178), .b(g62964_sb), .o(n_5954) );
in01s01 g62503_u0 ( .a(FE_OFN1250_n_4093), .o(g62503_sb) );
na02m01 TIMEBOOST_cell_3115 ( .a(TIMEBOOST_net_137), .b(n_1813), .o(n_4720) );
na03s02 TIMEBOOST_cell_37643 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__Q), .b(FE_OFN717_n_8176), .c(n_1917), .o(TIMEBOOST_net_11060) );
na02s01 TIMEBOOST_cell_43253 ( .a(n_4351), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__Q), .o(TIMEBOOST_net_13865) );
in01s02 g62504_u0 ( .a(FE_OFN1322_n_6436), .o(g62504_sb) );
na02m02 TIMEBOOST_cell_43991 ( .a(n_9538), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__Q), .o(TIMEBOOST_net_14234) );
na02s02 TIMEBOOST_cell_42824 ( .a(TIMEBOOST_net_13650), .b(g65317_db), .o(n_3565) );
na03m02 TIMEBOOST_cell_3754 ( .a(n_2929), .b(n_2411), .c(n_1227), .o(TIMEBOOST_net_457) );
in01s01 g62505_u0 ( .a(FE_OFN1268_n_4095), .o(g62505_sb) );
na02f02 TIMEBOOST_cell_37043 ( .a(FE_OFN1775_n_13800), .b(TIMEBOOST_net_10149), .o(TIMEBOOST_net_10760) );
na02s01 TIMEBOOST_cell_38054 ( .a(TIMEBOOST_net_11265), .b(FE_OFN1135_g64577_p), .o(TIMEBOOST_net_4621) );
in01s01 g62506_u0 ( .a(FE_OFN369_n_4092), .o(g62506_sb) );
na02f02 TIMEBOOST_cell_37045 ( .a(FE_OFN1775_n_13800), .b(TIMEBOOST_net_10148), .o(TIMEBOOST_net_10761) );
na02f02 TIMEBOOST_cell_43992 ( .a(TIMEBOOST_net_14234), .b(FE_OFN1422_n_8567), .o(TIMEBOOST_net_12956) );
na02m02 TIMEBOOST_cell_43993 ( .a(n_9000), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__Q), .o(TIMEBOOST_net_14235) );
in01s01 g62507_u0 ( .a(FE_OFN1223_n_6391), .o(g62507_sb) );
na02m04 TIMEBOOST_cell_3117 ( .a(TIMEBOOST_net_138), .b(n_2769), .o(n_3008) );
na03s02 TIMEBOOST_cell_37645 ( .a(n_1717), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__Q), .c(FE_OFN2081_n_8176), .o(TIMEBOOST_net_11061) );
na02m02 TIMEBOOST_cell_3118 ( .a(n_2281), .b(n_3007), .o(TIMEBOOST_net_139) );
in01s01 g62508_u0 ( .a(FE_OFN1243_n_4092), .o(g62508_sb) );
na02s02 TIMEBOOST_cell_42839 ( .a(g65862_db), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__Q), .o(TIMEBOOST_net_13658) );
na02f02 TIMEBOOST_cell_43994 ( .a(TIMEBOOST_net_14235), .b(FE_OFN1377_n_8567), .o(TIMEBOOST_net_12969) );
na02f02 TIMEBOOST_cell_42198 ( .a(TIMEBOOST_net_13337), .b(FE_OFN1389_n_8567), .o(TIMEBOOST_net_12287) );
in01s01 g62509_u0 ( .a(FE_OFN1243_n_4092), .o(g62509_sb) );
na02s02 TIMEBOOST_cell_42840 ( .a(TIMEBOOST_net_13658), .b(g65862_da), .o(TIMEBOOST_net_11929) );
na02s02 TIMEBOOST_cell_41912 ( .a(TIMEBOOST_net_13194), .b(g58344_db), .o(n_9018) );
na02m02 TIMEBOOST_cell_42199 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__Q), .b(n_9496), .o(TIMEBOOST_net_13338) );
in01s01 g62510_u0 ( .a(FE_OFN1270_n_4095), .o(g62510_sb) );
na02f06 TIMEBOOST_cell_36999 ( .a(n_16967), .b(n_16205), .o(TIMEBOOST_net_10738) );
na02f02 TIMEBOOST_cell_41234 ( .a(TIMEBOOST_net_12855), .b(g57165_sb), .o(n_10836) );
in01s01 g62511_u0 ( .a(n_6554), .o(g62511_sb) );
na02s02 TIMEBOOST_cell_42841 ( .a(g65914_db), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__Q), .o(TIMEBOOST_net_13659) );
na02s02 TIMEBOOST_cell_45199 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__Q), .b(n_3566), .o(TIMEBOOST_net_14838) );
na02s02 TIMEBOOST_cell_40730 ( .a(TIMEBOOST_net_12603), .b(g63148_sb), .o(n_5844) );
in01s01 g62512_u0 ( .a(FE_OFN1222_n_6391), .o(g62512_sb) );
na02m04 TIMEBOOST_cell_3119 ( .a(n_1973), .b(TIMEBOOST_net_139), .o(n_2492) );
na03s02 TIMEBOOST_cell_37647 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__Q), .b(FE_OFN2256_n_8060), .c(n_1919), .o(TIMEBOOST_net_11062) );
na02f02 TIMEBOOST_cell_45464 ( .a(TIMEBOOST_net_14970), .b(n_7508), .o(TIMEBOOST_net_11628) );
in01s01 g62513_u0 ( .a(FE_OFN1222_n_6391), .o(g62513_sb) );
na02s01 TIMEBOOST_cell_3121 ( .a(TIMEBOOST_net_140), .b(g65857_sb), .o(n_1581) );
na02s02 TIMEBOOST_cell_43553 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__Q), .b(n_3534), .o(TIMEBOOST_net_14015) );
na02s01 TIMEBOOST_cell_42637 ( .a(FE_OFN245_n_9114), .b(g58193_sb), .o(TIMEBOOST_net_13557) );
in01s01 g62514_u0 ( .a(FE_OFN1244_n_4092), .o(g62514_sb) );
na02s02 TIMEBOOST_cell_42842 ( .a(TIMEBOOST_net_13659), .b(g65914_da), .o(TIMEBOOST_net_11930) );
na02f02 TIMEBOOST_cell_42324 ( .a(TIMEBOOST_net_13400), .b(g57337_sb), .o(n_11415) );
na02f02 TIMEBOOST_cell_42260 ( .a(TIMEBOOST_net_13368), .b(FE_OFN1417_n_8567), .o(TIMEBOOST_net_12335) );
in01s01 g62515_u0 ( .a(FE_OFN1226_n_6391), .o(g62515_sb) );
na02s01 TIMEBOOST_cell_3123 ( .a(TIMEBOOST_net_141), .b(g65863_sb), .o(n_1578) );
na02s02 TIMEBOOST_cell_39882 ( .a(TIMEBOOST_net_12179), .b(g62553_sb), .o(n_6458) );
na02m02 TIMEBOOST_cell_32678 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__Q), .o(TIMEBOOST_net_10250) );
in01s01 g62516_u0 ( .a(FE_OFN1222_n_6391), .o(g62516_sb) );
na02s02 TIMEBOOST_cell_40732 ( .a(TIMEBOOST_net_12604), .b(g62616_sb), .o(n_6325) );
na03s02 TIMEBOOST_cell_37651 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__Q), .b(FE_OFN2084_n_8407), .c(n_2060), .o(TIMEBOOST_net_11064) );
na03m02 TIMEBOOST_cell_45465 ( .a(g52398_db), .b(g52398_sb), .c(n_3331), .o(TIMEBOOST_net_14971) );
in01s01 g62517_u0 ( .a(FE_OFN1224_n_6391), .o(g62517_sb) );
na02s01 TIMEBOOST_cell_3127 ( .a(TIMEBOOST_net_143), .b(g65857_sb), .o(n_1648) );
na02f02 TIMEBOOST_cell_44737 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__Q), .b(FE_OFN1583_n_12306), .o(TIMEBOOST_net_14607) );
na02f02 TIMEBOOST_cell_44740 ( .a(TIMEBOOST_net_14608), .b(n_11934), .o(n_12653) );
in01s02 g62518_u0 ( .a(FE_OFN1314_n_6624), .o(g62518_sb) );
na02s02 TIMEBOOST_cell_43427 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__Q), .b(n_3676), .o(TIMEBOOST_net_13952) );
na02m04 TIMEBOOST_cell_3755 ( .a(n_2931), .b(TIMEBOOST_net_457), .o(n_3324) );
na02m02 TIMEBOOST_cell_3756 ( .a(n_1986), .b(n_2929), .o(TIMEBOOST_net_458) );
in01s01 g62519_u0 ( .a(FE_OFN1317_n_6624), .o(g62519_sb) );
na02s02 TIMEBOOST_cell_16967 ( .a(TIMEBOOST_net_3740), .b(g65229_sb), .o(n_2658) );
na02m02 TIMEBOOST_cell_3757 ( .a(TIMEBOOST_net_458), .b(n_2931), .o(n_2930) );
na02f02 TIMEBOOST_cell_22351 ( .a(TIMEBOOST_net_6432), .b(n_10173), .o(n_12160) );
in01s02 g62520_u0 ( .a(FE_OFN1316_n_6624), .o(g62520_sb) );
na02s02 TIMEBOOST_cell_43428 ( .a(TIMEBOOST_net_13952), .b(n_6431), .o(TIMEBOOST_net_12189) );
na02f02 TIMEBOOST_cell_3759 ( .a(TIMEBOOST_net_459), .b(FE_RN_704_0), .o(FE_RN_705_0) );
na02s01 TIMEBOOST_cell_3760 ( .a(n_4869), .b(n_15856), .o(TIMEBOOST_net_460) );
in01s01 g62521_u0 ( .a(FE_OFN1260_n_4143), .o(g62521_sb) );
na02s01 TIMEBOOST_cell_42843 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__Q), .b(n_2198), .o(TIMEBOOST_net_13660) );
na02f02 TIMEBOOST_cell_44608 ( .a(TIMEBOOST_net_14542), .b(FE_OFN2169_n_8567), .o(TIMEBOOST_net_13478) );
na02f02 TIMEBOOST_cell_13045 ( .a(TIMEBOOST_net_3089), .b(n_11996), .o(n_12517) );
in01s01 g62522_u0 ( .a(FE_OFN1260_n_4143), .o(g62522_sb) );
na02s01 TIMEBOOST_cell_42844 ( .a(TIMEBOOST_net_13660), .b(FE_OFN720_n_8060), .o(TIMEBOOST_net_11254) );
na02f02 TIMEBOOST_cell_41418 ( .a(TIMEBOOST_net_12947), .b(g57574_sb), .o(n_11177) );
na03s02 TIMEBOOST_cell_43317 ( .a(n_3529), .b(FE_OFN1278_n_4097), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__Q), .o(TIMEBOOST_net_13897) );
in01s01 g62523_u0 ( .a(FE_OFN1314_n_6624), .o(g62523_sb) );
na02s02 TIMEBOOST_cell_43429 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__Q), .b(n_4236), .o(TIMEBOOST_net_13953) );
na02f02 TIMEBOOST_cell_3761 ( .a(n_4818), .b(TIMEBOOST_net_460), .o(n_7538) );
na02m02 TIMEBOOST_cell_45466 ( .a(TIMEBOOST_net_14971), .b(TIMEBOOST_net_591), .o(n_14822) );
in01s01 g62524_u0 ( .a(FE_OFN1249_n_4093), .o(g62524_sb) );
na02s01 TIMEBOOST_cell_42845 ( .a(n_1664), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__Q), .o(TIMEBOOST_net_13661) );
na02s01 TIMEBOOST_cell_42749 ( .a(FE_OFN215_n_9856), .b(g58175_sb), .o(TIMEBOOST_net_13613) );
in01s01 g62525_u0 ( .a(FE_OFN1248_n_4093), .o(g62525_sb) );
na02m02 TIMEBOOST_cell_3129 ( .a(TIMEBOOST_net_144), .b(n_2260), .o(n_2429) );
na03s02 TIMEBOOST_cell_37655 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__Q), .b(FE_OFN2257_n_8060), .c(n_2207), .o(TIMEBOOST_net_11066) );
na02s01 TIMEBOOST_cell_30880 ( .a(pci_target_unit_pcit_if_strd_addr_in_689), .b(n_2526), .o(TIMEBOOST_net_9351) );
in01s01 g62526_u0 ( .a(FE_OFN1278_n_4097), .o(g62526_sb) );
na02s04 TIMEBOOST_cell_3131 ( .a(TIMEBOOST_net_145), .b(n_2236), .o(n_2948) );
na03s02 TIMEBOOST_cell_43011 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__Q), .b(FE_OFN1120_g64577_p), .c(g62774_sb), .o(TIMEBOOST_net_13744) );
in01s01 g62527_u0 ( .a(FE_OFN1282_n_4097), .o(g62527_sb) );
na02s02 TIMEBOOST_cell_42846 ( .a(TIMEBOOST_net_13661), .b(FE_OFN719_n_8060), .o(TIMEBOOST_net_11249) );
na02f02 TIMEBOOST_cell_42326 ( .a(TIMEBOOST_net_13401), .b(g57429_sb), .o(n_11305) );
in01s01 g62528_u0 ( .a(FE_OFN1219_n_6886), .o(g62528_sb) );
na02m02 TIMEBOOST_cell_3133 ( .a(TIMEBOOST_net_146), .b(n_1799), .o(n_2876) );
na03s02 TIMEBOOST_cell_37659 ( .a(n_1593), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__Q), .c(FE_OFN714_n_8140), .o(TIMEBOOST_net_11068) );
na02f08 TIMEBOOST_cell_3134 ( .a(n_16516), .b(n_16501), .o(TIMEBOOST_net_147) );
in01s01 g62529_u0 ( .a(FE_OFN1231_n_6391), .o(g62529_sb) );
na02f02 TIMEBOOST_cell_42478 ( .a(TIMEBOOST_net_13477), .b(g57271_sb), .o(n_10416) );
na02s01 TIMEBOOST_cell_42847 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__Q), .b(n_2212), .o(TIMEBOOST_net_13662) );
na02s01 TIMEBOOST_cell_40519 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__Q), .b(wishbone_slave_unit_pcim_sm_data_in_646), .o(TIMEBOOST_net_12498) );
in01s01 g62530_u0 ( .a(FE_OFN1250_n_4093), .o(g62530_sb) );
na02f04 TIMEBOOST_cell_3135 ( .a(n_16499), .b(TIMEBOOST_net_147), .o(n_16503) );
in01s01 TIMEBOOST_cell_45873 ( .a(n_11849), .o(TIMEBOOST_net_15180) );
na03f02 TIMEBOOST_cell_36139 ( .a(n_11013), .b(FE_RN_98_0), .c(n_12591), .o(n_12853) );
in01s01 g62531_u0 ( .a(FE_OFN1249_n_4093), .o(g62531_sb) );
na02s01 TIMEBOOST_cell_42848 ( .a(TIMEBOOST_net_13662), .b(FE_OFN720_n_8060), .o(TIMEBOOST_net_11250) );
na02m02 TIMEBOOST_cell_41605 ( .a(wbu_sel_in_312), .b(wishbone_slave_unit_fifos_wbr_be_in_264), .o(TIMEBOOST_net_13041) );
na02f02 TIMEBOOST_cell_41576 ( .a(TIMEBOOST_net_13026), .b(g57469_sb), .o(n_10820) );
in01s01 g62532_u0 ( .a(FE_OFN1233_n_6391), .o(g62532_sb) );
na02s01 TIMEBOOST_cell_36791 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__Q), .b(g62729_sb), .o(TIMEBOOST_net_10634) );
na02f02 TIMEBOOST_cell_3481 ( .a(TIMEBOOST_net_320), .b(n_13221), .o(g59331_p) );
na02s01 TIMEBOOST_cell_3482 ( .a(FE_OFN2093_n_2301), .b(FE_OCPN1838_n_1238), .o(TIMEBOOST_net_321) );
in01s01 g62533_u0 ( .a(FE_OFN1230_n_6391), .o(g62533_sb) );
na03s02 TIMEBOOST_cell_36787 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__Q), .b(FE_OFN1129_g64577_p), .c(n_4033), .o(TIMEBOOST_net_10632) );
na02s01 TIMEBOOST_cell_3483 ( .a(TIMEBOOST_net_321), .b(n_2725), .o(n_3363) );
na02s02 TIMEBOOST_cell_45095 ( .a(n_1978), .b(wishbone_slave_unit_pcim_sm_be_in_557), .o(TIMEBOOST_net_14786) );
in01s01 g62534_u0 ( .a(FE_OFN2064_n_6391), .o(g62534_sb) );
na02s01 TIMEBOOST_cell_37254 ( .a(TIMEBOOST_net_10865), .b(FE_OFN1626_n_4438), .o(TIMEBOOST_net_9403) );
na02f02 TIMEBOOST_cell_3485 ( .a(TIMEBOOST_net_322), .b(n_4897), .o(n_7322) );
na02f02 TIMEBOOST_cell_44208 ( .a(TIMEBOOST_net_14342), .b(FE_OFN1374_n_8567), .o(TIMEBOOST_net_12987) );
in01s01 g62535_u0 ( .a(FE_OFN1315_n_6624), .o(g62535_sb) );
na02s01 TIMEBOOST_cell_16991 ( .a(TIMEBOOST_net_3752), .b(g65220_sb), .o(n_2667) );
na02s02 TIMEBOOST_cell_3763 ( .a(TIMEBOOST_net_461), .b(n_3107), .o(n_8476) );
na02m01 TIMEBOOST_cell_3764 ( .a(g52624_db), .b(n_14837), .o(TIMEBOOST_net_462) );
in01s01 g62536_u0 ( .a(FE_OFN1261_n_4143), .o(g62536_sb) );
na02f02 TIMEBOOST_cell_41544 ( .a(TIMEBOOST_net_13010), .b(g57367_sb), .o(n_10383) );
na03s02 TIMEBOOST_cell_41961 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__Q), .b(n_4339), .c(FE_OFN1264_n_4095), .o(TIMEBOOST_net_13219) );
in01s01 g62537_u0 ( .a(FE_OFN1258_n_4143), .o(g62537_sb) );
na03s02 TIMEBOOST_cell_36793 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__21__Q), .b(FE_OFN1140_g64577_p), .c(g62777_sb), .o(TIMEBOOST_net_10635) );
na02s01 TIMEBOOST_cell_43254 ( .a(TIMEBOOST_net_13865), .b(FE_OFN1225_n_6391), .o(TIMEBOOST_net_12526) );
na02s02 TIMEBOOST_cell_42604 ( .a(TIMEBOOST_net_13540), .b(g65016_db), .o(n_3634) );
in01s01 g62538_u0 ( .a(FE_OFN1283_n_4097), .o(g62538_sb) );
na03s02 TIMEBOOST_cell_36795 ( .a(g64267_da), .b(g64267_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__Q), .o(TIMEBOOST_net_10636) );
na02f02 TIMEBOOST_cell_41290 ( .a(TIMEBOOST_net_12883), .b(g57195_sb), .o(n_11557) );
na02f02 TIMEBOOST_cell_41242 ( .a(TIMEBOOST_net_12859), .b(g57128_sb), .o(n_11617) );
in01s01 g62539_u0 ( .a(FE_OFN1284_n_4097), .o(g62539_sb) );
na02s02 TIMEBOOST_cell_40704 ( .a(TIMEBOOST_net_12590), .b(g63167_sb), .o(n_5804) );
na02s02 TIMEBOOST_cell_18235 ( .a(TIMEBOOST_net_4374), .b(g61940_sb), .o(n_7943) );
no02m06 TIMEBOOST_cell_3138 ( .a(FE_RN_603_0), .b(FE_RN_604_0), .o(TIMEBOOST_net_149) );
in01s01 g62540_u0 ( .a(n_6645), .o(g62540_sb) );
na02s01 TIMEBOOST_cell_45720 ( .a(TIMEBOOST_net_15098), .b(g62999_sb), .o(n_5884) );
na02s01 TIMEBOOST_cell_39207 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__Q), .b(n_8407), .o(TIMEBOOST_net_11842) );
na02f02 TIMEBOOST_cell_44342 ( .a(TIMEBOOST_net_14409), .b(FE_OFN1409_n_8567), .o(TIMEBOOST_net_12728) );
in01s01 g62541_u0 ( .a(FE_OFN1219_n_6886), .o(g62541_sb) );
na03s02 TIMEBOOST_cell_36797 ( .a(g60686_da), .b(g60686_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__Q), .o(TIMEBOOST_net_10637) );
na02f02 TIMEBOOST_cell_41238 ( .a(TIMEBOOST_net_12857), .b(g57321_sb), .o(n_11429) );
na02m02 TIMEBOOST_cell_45467 ( .a(n_7711), .b(TIMEBOOST_net_703), .o(TIMEBOOST_net_14972) );
in01s01 g62542_u0 ( .a(FE_OFN1242_n_4092), .o(g62542_sb) );
na03s02 TIMEBOOST_cell_36799 ( .a(g64310_da), .b(g64310_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__Q), .o(TIMEBOOST_net_10638) );
na02f02 TIMEBOOST_cell_45468 ( .a(TIMEBOOST_net_14972), .b(n_13747), .o(TIMEBOOST_net_12679) );
na02m02 TIMEBOOST_cell_41606 ( .a(FE_OFN1438_n_9372), .b(TIMEBOOST_net_13041), .o(TIMEBOOST_net_11666) );
in01s01 g62543_u0 ( .a(FE_OFN1284_n_4097), .o(g62543_sb) );
no02f04 TIMEBOOST_cell_3139 ( .a(TIMEBOOST_net_149), .b(FE_RN_605_0), .o(FE_RN_606_0) );
na03s02 TIMEBOOST_cell_37663 ( .a(n_1881), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__Q), .c(FE_OFN706_n_8119), .o(TIMEBOOST_net_11070) );
na03f02 TIMEBOOST_cell_36138 ( .a(n_14545), .b(n_14513), .c(n_14431), .o(n_14590) );
in01s01 g62544_u0 ( .a(FE_OFN1274_n_4096), .o(g62544_sb) );
na02m02 TIMEBOOST_cell_3141 ( .a(n_2558), .b(TIMEBOOST_net_150), .o(n_4778) );
na03s02 TIMEBOOST_cell_37665 ( .a(n_1589), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__Q), .c(FE_OFN2081_n_8176), .o(TIMEBOOST_net_11071) );
na02s02 TIMEBOOST_cell_42638 ( .a(TIMEBOOST_net_13557), .b(g58193_db), .o(n_9057) );
in01m01 g62545_u0 ( .a(FE_OFN1274_n_4096), .o(g62545_sb) );
no02f02 TIMEBOOST_cell_3143 ( .a(TIMEBOOST_net_151), .b(FE_RN_626_0), .o(FE_RN_631_0) );
na02s02 TIMEBOOST_cell_18233 ( .a(TIMEBOOST_net_4373), .b(g61952_sb), .o(n_7921) );
na02f02 TIMEBOOST_cell_41322 ( .a(TIMEBOOST_net_12899), .b(g57167_sb), .o(n_11586) );
in01s01 g62546_u0 ( .a(FE_OFN1244_n_4092), .o(g62546_sb) );
na03s02 TIMEBOOST_cell_36777 ( .a(g64278_da), .b(g64278_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__Q), .o(TIMEBOOST_net_10627) );
na02s02 TIMEBOOST_cell_43084 ( .a(TIMEBOOST_net_13780), .b(FE_OFN1293_n_4098), .o(TIMEBOOST_net_12212) );
na03f02 TIMEBOOST_cell_43085 ( .a(TIMEBOOST_net_557), .b(FE_OFN2069_n_15978), .c(n_4204), .o(TIMEBOOST_net_13781) );
in01s01 g62547_u0 ( .a(FE_OFN1312_n_6624), .o(g62547_sb) );
na02s02 TIMEBOOST_cell_43430 ( .a(TIMEBOOST_net_13953), .b(n_6431), .o(TIMEBOOST_net_12185) );
na03s02 TIMEBOOST_cell_38225 ( .a(g64324_da), .b(g64324_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__Q), .o(TIMEBOOST_net_11351) );
na02m01 TIMEBOOST_cell_3766 ( .a(g52643_db), .b(n_14837), .o(TIMEBOOST_net_463) );
in01s01 g62548_u0 ( .a(FE_OFN1243_n_4092), .o(g62548_sb) );
na02f02 TIMEBOOST_cell_42246 ( .a(TIMEBOOST_net_13361), .b(FE_OFN1374_n_8567), .o(TIMEBOOST_net_12317) );
na02s01 TIMEBOOST_cell_45670 ( .a(TIMEBOOST_net_15073), .b(g63591_da), .o(n_7180) );
na02m02 TIMEBOOST_cell_44655 ( .a(n_9225), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__Q), .o(TIMEBOOST_net_14566) );
in01s01 g62549_u0 ( .a(FE_OFN1244_n_4092), .o(g62549_sb) );
na02s02 TIMEBOOST_cell_36741 ( .a(n_3890), .b(g63095_sb), .o(TIMEBOOST_net_10609) );
na02s01 TIMEBOOST_cell_41982 ( .a(TIMEBOOST_net_13229), .b(g62376_sb), .o(n_6851) );
na02m02 TIMEBOOST_cell_45671 ( .a(TIMEBOOST_net_515), .b(g53939_sb), .o(TIMEBOOST_net_15074) );
in01s01 g62550_u0 ( .a(FE_OFN2063_n_6391), .o(g62550_sb) );
na02s01 TIMEBOOST_cell_36401 ( .a(pci_target_unit_fifos_pcir_data_in_175), .b(g65688_sb), .o(TIMEBOOST_net_10439) );
no02f02 TIMEBOOST_cell_3487 ( .a(TIMEBOOST_net_323), .b(FE_RN_703_0), .o(FE_RN_704_0) );
na02f04 TIMEBOOST_cell_3488 ( .a(n_16451), .b(FE_OCPN1875_n_14526), .o(TIMEBOOST_net_324) );
in01s01 g62551_u0 ( .a(FE_OFN1224_n_6391), .o(g62551_sb) );
na02s01 TIMEBOOST_cell_45469 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__Q), .b(FE_OFN1094_g64577_p), .o(TIMEBOOST_net_14973) );
na03s02 TIMEBOOST_cell_37667 ( .a(n_1594), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__Q), .c(FE_OFN709_n_8232), .o(TIMEBOOST_net_11072) );
na02m02 TIMEBOOST_cell_32676 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__Q), .o(TIMEBOOST_net_10249) );
in01s01 g62552_u0 ( .a(FE_OFN1224_n_6391), .o(g62552_sb) );
na02s01 TIMEBOOST_cell_42639 ( .a(FE_OFN245_n_9114), .b(g57973_sb), .o(TIMEBOOST_net_13558) );
na03s01 TIMEBOOST_cell_37669 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__Q), .b(FE_OFN702_n_7845), .c(n_2186), .o(TIMEBOOST_net_11073) );
na02s01 TIMEBOOST_cell_17961 ( .a(TIMEBOOST_net_4237), .b(g65384_da), .o(n_4656) );
in01s01 g62553_u0 ( .a(FE_OFN1232_n_6391), .o(g62553_sb) );
na02s01 TIMEBOOST_cell_36451 ( .a(pci_target_unit_fifos_pciw_cbe_in), .b(g64138_sb), .o(TIMEBOOST_net_10464) );
na02f04 TIMEBOOST_cell_3489 ( .a(TIMEBOOST_net_324), .b(n_16452), .o(n_16455) );
na02s02 TIMEBOOST_cell_17512 ( .a(pci_target_unit_fifos_pciw_addr_data_in_130), .b(g64208_sb), .o(TIMEBOOST_net_4013) );
in01s01 g62554_u0 ( .a(FE_OFN1268_n_4095), .o(g62554_sb) );
na02f02 TIMEBOOST_cell_37047 ( .a(FE_OFN1775_n_13800), .b(TIMEBOOST_net_10153), .o(TIMEBOOST_net_10762) );
na02s02 TIMEBOOST_cell_41978 ( .a(TIMEBOOST_net_13227), .b(g62489_sb), .o(n_6607) );
na02s02 TIMEBOOST_cell_43318 ( .a(TIMEBOOST_net_13897), .b(g62910_sb), .o(n_6058) );
in01s01 g62555_u0 ( .a(FE_OFN1270_n_4095), .o(g62555_sb) );
na02m02 TIMEBOOST_cell_36743 ( .a(n_3493), .b(g53897_sb), .o(TIMEBOOST_net_10610) );
na02m02 TIMEBOOST_cell_43995 ( .a(n_9494), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__Q), .o(TIMEBOOST_net_14236) );
na02f02 TIMEBOOST_cell_45755 ( .a(TIMEBOOST_net_9567), .b(FE_OFN1063_n_15808), .o(TIMEBOOST_net_15116) );
in01s01 g62556_u0 ( .a(FE_OFN1248_n_4093), .o(g62556_sb) );
na02s02 TIMEBOOST_cell_40852 ( .a(TIMEBOOST_net_12664), .b(FE_OFN1330_n_13547), .o(TIMEBOOST_net_11620) );
na03s02 TIMEBOOST_cell_37671 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__Q), .b(FE_OFN713_n_8140), .c(n_2189), .o(TIMEBOOST_net_11074) );
na02f02 TIMEBOOST_cell_32675 ( .a(FE_OFN1759_n_10780), .b(TIMEBOOST_net_10248), .o(TIMEBOOST_net_6501) );
in01s01 g62557_u0 ( .a(FE_OFN1274_n_4096), .o(g62557_sb) );
na02s01 TIMEBOOST_cell_3151 ( .a(TIMEBOOST_net_155), .b(g60689_sb), .o(n_3815) );
na03s02 TIMEBOOST_cell_37673 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__Q), .b(FE_OFN710_n_8232), .c(n_1865), .o(TIMEBOOST_net_11075) );
na02s01 TIMEBOOST_cell_45012 ( .a(TIMEBOOST_net_14744), .b(FE_OFN714_n_8140), .o(TIMEBOOST_net_11069) );
in01s02 g62558_u0 ( .a(FE_OFN1323_n_6436), .o(g62558_sb) );
na02s02 TIMEBOOST_cell_16965 ( .a(TIMEBOOST_net_3739), .b(g65227_sb), .o(n_2660) );
na03s02 TIMEBOOST_cell_18788 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__Q), .b(FE_OFN1122_g64577_p), .c(n_4060), .o(TIMEBOOST_net_4651) );
na02s02 TIMEBOOST_cell_39884 ( .a(TIMEBOOST_net_12180), .b(g62990_sb), .o(n_5902) );
in01s01 g62559_u0 ( .a(FE_OFN1212_n_4151), .o(g62559_sb) );
na02s01 TIMEBOOST_cell_15810 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_5_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_2_), .o(TIMEBOOST_net_3162) );
na02s02 TIMEBOOST_cell_38362 ( .a(TIMEBOOST_net_11419), .b(g63076_sb), .o(n_5098) );
in01s01 g62560_u0 ( .a(FE_OFN1323_n_6436), .o(g62560_sb) );
na02f02 TIMEBOOST_cell_43996 ( .a(TIMEBOOST_net_14236), .b(FE_OFN1376_n_8567), .o(TIMEBOOST_net_12882) );
na02s02 TIMEBOOST_cell_38263 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_72), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_11370) );
na02s02 TIMEBOOST_cell_3770 ( .a(n_2872), .b(n_2596), .o(TIMEBOOST_net_465) );
in01s01 g62561_u0 ( .a(FE_OFN1323_n_6436), .o(g62561_sb) );
na02m02 TIMEBOOST_cell_43997 ( .a(n_9135), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__Q), .o(TIMEBOOST_net_14237) );
na02m02 TIMEBOOST_cell_3771 ( .a(n_2873), .b(TIMEBOOST_net_465), .o(n_2874) );
na02s01 TIMEBOOST_cell_38550 ( .a(TIMEBOOST_net_11513), .b(g62051_sb), .o(n_7759) );
in01s01 g62562_u0 ( .a(FE_OFN1313_n_6624), .o(g62562_sb) );
na02s02 TIMEBOOST_cell_16941 ( .a(TIMEBOOST_net_3727), .b(g65250_sb), .o(n_2632) );
na02f02 TIMEBOOST_cell_3773 ( .a(TIMEBOOST_net_466), .b(g54323_da), .o(g54039_db) );
na02s02 TIMEBOOST_cell_17665 ( .a(TIMEBOOST_net_4089), .b(g65412_db), .o(n_4670) );
in01s01 g62563_u0 ( .a(n_6431), .o(g62563_sb) );
na02s01 TIMEBOOST_cell_36455 ( .a(n_2675), .b(FE_OFN783_n_2678), .o(TIMEBOOST_net_10466) );
na02m02 TIMEBOOST_cell_43813 ( .a(n_9198), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__Q), .o(TIMEBOOST_net_14145) );
na02s01 TIMEBOOST_cell_37572 ( .a(TIMEBOOST_net_11024), .b(g65925_db), .o(n_2586) );
in01s01 g62564_u0 ( .a(FE_OFN1193_n_6935), .o(g62564_sb) );
na02f08 TIMEBOOST_cell_3155 ( .a(TIMEBOOST_net_157), .b(n_4743), .o(n_7498) );
na02s02 TIMEBOOST_cell_43554 ( .a(TIMEBOOST_net_14015), .b(FE_OFN1317_n_6624), .o(TIMEBOOST_net_12253) );
na02s01 TIMEBOOST_cell_45470 ( .a(TIMEBOOST_net_14973), .b(g62733_sb), .o(TIMEBOOST_net_10024) );
in01s01 g62565_u0 ( .a(FE_OFN1193_n_6935), .o(g62565_sb) );
na02f02 TIMEBOOST_cell_44648 ( .a(TIMEBOOST_net_14562), .b(FE_OFN2169_n_8567), .o(TIMEBOOST_net_13485) );
na03f06 TIMEBOOST_cell_32919 ( .a(n_16388), .b(n_16390), .c(n_16389), .o(n_16391) );
in01s01 g62566_u0 ( .a(FE_OFN1285_n_4097), .o(g62566_sb) );
na02s01 TIMEBOOST_cell_42849 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__Q), .b(n_2293), .o(TIMEBOOST_net_13663) );
na02m02 TIMEBOOST_cell_45672 ( .a(TIMEBOOST_net_15074), .b(g54185_da), .o(TIMEBOOST_net_10643) );
na03m02 TIMEBOOST_cell_32917 ( .a(n_1615), .b(TIMEBOOST_net_3213), .c(n_1616), .o(TIMEBOOST_net_9306) );
in01s01 g62567_u0 ( .a(FE_OFN1284_n_4097), .o(g62567_sb) );
na02s02 TIMEBOOST_cell_40734 ( .a(TIMEBOOST_net_12605), .b(g62483_sb), .o(n_6621) );
no02m01 TIMEBOOST_cell_18229 ( .a(TIMEBOOST_net_4371), .b(g61618_BP), .o(g61618_p) );
na02s02 TIMEBOOST_cell_15811 ( .a(TIMEBOOST_net_3162), .b(n_947), .o(TIMEBOOST_net_32) );
in01s01 g62568_u0 ( .a(FE_OFN1295_n_4098), .o(g62568_sb) );
na02s01 TIMEBOOST_cell_17699 ( .a(TIMEBOOST_net_4106), .b(g61800_sb), .o(n_8196) );
na02m02 TIMEBOOST_cell_32674 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__Q), .o(TIMEBOOST_net_10248) );
na02s02 TIMEBOOST_cell_41972 ( .a(TIMEBOOST_net_13224), .b(g62899_sb), .o(n_6079) );
in01s01 g62569_u0 ( .a(FE_OFN1315_n_6624), .o(g62569_sb) );
na02f02 TIMEBOOST_cell_43998 ( .a(TIMEBOOST_net_14237), .b(FE_OFN1397_n_8567), .o(TIMEBOOST_net_12957) );
na02s02 TIMEBOOST_cell_39886 ( .a(TIMEBOOST_net_12181), .b(g62936_sb), .o(n_6009) );
na02f06 TIMEBOOST_cell_3776 ( .a(n_15910), .b(n_15914), .o(TIMEBOOST_net_468) );
in01s01 g62570_u0 ( .a(FE_OFN1234_n_6391), .o(g62570_sb) );
na02s01 TIMEBOOST_cell_36371 ( .a(FE_OFN945_n_2248), .b(g65849_sb), .o(TIMEBOOST_net_10424) );
na02s01 TIMEBOOST_cell_44969 ( .a(g58075_sb), .b(FE_OFN215_n_9856), .o(TIMEBOOST_net_14723) );
in01s01 TIMEBOOST_cell_8843 ( .a(TIMEBOOST_net_979), .o(TIMEBOOST_net_980) );
in01s01 g62571_u0 ( .a(FE_OFN1314_n_6624), .o(g62571_sb) );
na02m02 TIMEBOOST_cell_43999 ( .a(n_9103), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__Q), .o(TIMEBOOST_net_14238) );
na02f08 TIMEBOOST_cell_3777 ( .a(TIMEBOOST_net_468), .b(FE_OCP_RBN2231_FE_RN_390_0), .o(n_15915) );
in01s01 g62572_u0 ( .a(FE_OFN1200_n_4090), .o(g62572_sb) );
na02s01 TIMEBOOST_cell_38056 ( .a(TIMEBOOST_net_11266), .b(FE_OFN1135_g64577_p), .o(TIMEBOOST_net_4521) );
na02f02 TIMEBOOST_cell_41556 ( .a(TIMEBOOST_net_13016), .b(g57059_sb), .o(n_10848) );
na02f02 TIMEBOOST_cell_32673 ( .a(FE_OFN1759_n_10780), .b(TIMEBOOST_net_10247), .o(TIMEBOOST_net_6500) );
in01s01 g62573_u0 ( .a(FE_OFN1196_n_4090), .o(g62573_sb) );
no02f06 TIMEBOOST_cell_20346 ( .a(FE_OFN1706_n_4868), .b(FE_RN_361_0), .o(TIMEBOOST_net_5430) );
na02s02 TIMEBOOST_cell_45673 ( .a(n_4228), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__Q), .o(TIMEBOOST_net_15075) );
na02m02 TIMEBOOST_cell_44389 ( .a(n_9078), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__Q), .o(TIMEBOOST_net_14433) );
in01s01 g62574_u0 ( .a(FE_OFN1193_n_6935), .o(g62574_sb) );
na02s02 TIMEBOOST_cell_20348 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__Q), .b(g59796_sb), .o(TIMEBOOST_net_5431) );
na02f02 TIMEBOOST_cell_41546 ( .a(TIMEBOOST_net_13011), .b(g57154_sb), .o(n_11597) );
na02s02 TIMEBOOST_cell_43492 ( .a(TIMEBOOST_net_13984), .b(FE_OFN1231_n_6391), .o(TIMEBOOST_net_12618) );
in01s01 g62575_u0 ( .a(FE_OFN1192_n_6935), .o(g62575_sb) );
na02s03 TIMEBOOST_cell_15812 ( .a(pci_target_unit_del_sync_comp_cycle_count_10_), .b(pci_target_unit_del_sync_comp_cycle_count_11_), .o(TIMEBOOST_net_3163) );
na02s01 g62575_u2 ( .a(n_4341), .b(n_6935), .o(g62575_db) );
na02s03 TIMEBOOST_cell_15813 ( .a(TIMEBOOST_net_3163), .b(n_937), .o(TIMEBOOST_net_243) );
in01s01 g62576_u0 ( .a(FE_OFN1320_n_6436), .o(g62576_sb) );
na02f02 TIMEBOOST_cell_44000 ( .a(TIMEBOOST_net_14238), .b(FE_OFN1381_n_8567), .o(TIMEBOOST_net_12872) );
na03s02 TIMEBOOST_cell_37607 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__Q), .b(FE_OFN713_n_8140), .c(n_2205), .o(TIMEBOOST_net_11042) );
na02s01 TIMEBOOST_cell_3780 ( .a(n_5757), .b(n_15741), .o(TIMEBOOST_net_470) );
in01s01 g62577_u0 ( .a(FE_OFN1246_n_4093), .o(g62577_sb) );
na02s01 TIMEBOOST_cell_38364 ( .a(TIMEBOOST_net_11420), .b(g63015_sb), .o(n_5218) );
na02s02 TIMEBOOST_cell_45674 ( .a(TIMEBOOST_net_15075), .b(FE_OFN1248_n_4093), .o(TIMEBOOST_net_13303) );
na02f02 TIMEBOOST_cell_41548 ( .a(TIMEBOOST_net_13012), .b(g57446_sb), .o(n_11286) );
in01s01 g62578_u0 ( .a(FE_OFN1208_n_6356), .o(g62578_sb) );
na02s02 TIMEBOOST_cell_39888 ( .a(TIMEBOOST_net_12182), .b(g62402_sb), .o(n_6795) );
na02f02 TIMEBOOST_cell_41494 ( .a(TIMEBOOST_net_12985), .b(g57182_sb), .o(n_11572) );
na02m02 TIMEBOOST_cell_45471 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__Q), .b(n_9882), .o(TIMEBOOST_net_14974) );
in01s01 g62579_u0 ( .a(FE_OFN1208_n_6356), .o(g62579_sb) );
na02s02 TIMEBOOST_cell_39890 ( .a(TIMEBOOST_net_12183), .b(g62677_sb), .o(n_6186) );
na02s01 TIMEBOOST_cell_41947 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__Q), .b(g58277_sb), .o(TIMEBOOST_net_13212) );
na02m02 TIMEBOOST_cell_41946 ( .a(TIMEBOOST_net_13211), .b(TIMEBOOST_net_9881), .o(n_13500) );
in01s01 g62580_u0 ( .a(FE_OFN1222_n_6391), .o(g62580_sb) );
na02s01 TIMEBOOST_cell_15814 ( .a(n_8831), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_29__Q), .o(TIMEBOOST_net_3164) );
na03s02 TIMEBOOST_cell_37605 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN707_n_8119), .c(n_2210), .o(TIMEBOOST_net_11041) );
na02f02 TIMEBOOST_cell_42480 ( .a(TIMEBOOST_net_13478), .b(g57074_sb), .o(n_10495) );
in01s01 g62581_u0 ( .a(FE_OFN1250_n_4093), .o(g62581_sb) );
na02s01 TIMEBOOST_cell_3163 ( .a(TIMEBOOST_net_161), .b(g60689_sb), .o(n_3204) );
na03s02 TIMEBOOST_cell_37601 ( .a(n_1595), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__Q), .c(FE_OFN714_n_8140), .o(TIMEBOOST_net_11039) );
na02s01 TIMEBOOST_cell_3164 ( .a(n_3761), .b(g65069_sb), .o(TIMEBOOST_net_162) );
in01s01 g62582_u0 ( .a(FE_OFN1194_n_6935), .o(g62582_sb) );
na02s01 TIMEBOOST_cell_3165 ( .a(TIMEBOOST_net_162), .b(g65069_db), .o(n_3607) );
na02m02 TIMEBOOST_cell_19047 ( .a(TIMEBOOST_net_4780), .b(n_7317), .o(n_8535) );
na02f02 TIMEBOOST_cell_41144 ( .a(TIMEBOOST_net_12810), .b(g57497_sb), .o(n_10329) );
in01s01 g62583_u0 ( .a(FE_OFN1224_n_6391), .o(g62583_sb) );
na02f02 TIMEBOOST_cell_41498 ( .a(TIMEBOOST_net_12987), .b(g57213_sb), .o(n_11544) );
na02s02 TIMEBOOST_cell_38589 ( .a(TIMEBOOST_net_9956), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_11533) );
na02s02 TIMEBOOST_cell_43145 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__Q), .b(n_4267), .o(TIMEBOOST_net_13811) );
in01s01 g62584_u0 ( .a(FE_OFN1293_n_4098), .o(g62584_sb) );
na03s02 TIMEBOOST_cell_39357 ( .a(n_1946), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__Q), .c(FE_OFN714_n_8140), .o(TIMEBOOST_net_11917) );
na02f02 TIMEBOOST_cell_45472 ( .a(TIMEBOOST_net_14974), .b(FE_OFN1349_n_8567), .o(TIMEBOOST_net_14463) );
na02s02 TIMEBOOST_cell_45746 ( .a(TIMEBOOST_net_15111), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_13243) );
in01s01 g62585_u0 ( .a(FE_OFN1294_n_4098), .o(g62585_sb) );
na02s02 TIMEBOOST_cell_39892 ( .a(TIMEBOOST_net_12184), .b(g62626_sb), .o(n_6303) );
in01s01 TIMEBOOST_cell_32854 ( .a(TIMEBOOST_net_10355), .o(TIMEBOOST_net_10326) );
no03f08 TIMEBOOST_cell_32870 ( .a(FE_RN_754_0), .b(wishbone_slave_unit_pci_initiator_if_del_read_req), .c(n_15859), .o(n_15979) );
in01s01 g62586_u0 ( .a(FE_OFN1213_n_4151), .o(g62586_sb) );
na02s02 TIMEBOOST_cell_39894 ( .a(TIMEBOOST_net_12185), .b(g62939_sb), .o(n_6003) );
na02m02 TIMEBOOST_cell_44639 ( .a(n_9879), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__Q), .o(TIMEBOOST_net_14558) );
na02f02 TIMEBOOST_cell_41504 ( .a(TIMEBOOST_net_12990), .b(g57183_sb), .o(n_11571) );
in01s01 g62587_u0 ( .a(FE_OFN1202_n_4090), .o(g62587_sb) );
na02s01 TIMEBOOST_cell_3169 ( .a(TIMEBOOST_net_164), .b(n_2477), .o(n_2478) );
na03s02 TIMEBOOST_cell_38209 ( .a(TIMEBOOST_net_4016), .b(g64217_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q), .o(TIMEBOOST_net_11343) );
na02s01 TIMEBOOST_cell_17223 ( .a(TIMEBOOST_net_3868), .b(g65322_da), .o(n_4269) );
in01s01 g62588_u0 ( .a(n_6431), .o(g62588_sb) );
na02s01 TIMEBOOST_cell_36457 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__Q), .b(FE_OFN527_n_9899), .o(TIMEBOOST_net_10467) );
na02s01 TIMEBOOST_cell_17168 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__Q), .o(TIMEBOOST_net_3841) );
na02f02 TIMEBOOST_cell_36924 ( .a(TIMEBOOST_net_10700), .b(g52605_sb), .o(n_10237) );
in01s01 g62589_u0 ( .a(FE_OFN1194_n_6935), .o(g62589_sb) );
na02s01 TIMEBOOST_cell_3171 ( .a(TIMEBOOST_net_165), .b(n_5641), .o(n_1978) );
na02s01 TIMEBOOST_cell_41737 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__Q), .b(g65324_sb), .o(TIMEBOOST_net_13107) );
na02s02 TIMEBOOST_cell_31411 ( .a(TIMEBOOST_net_9616), .b(g65015_db), .o(n_3635) );
in01s01 g62590_u0 ( .a(FE_OFN1206_n_6356), .o(g62590_sb) );
na02s02 TIMEBOOST_cell_39164 ( .a(TIMEBOOST_net_11820), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_9852) );
na02m02 TIMEBOOST_cell_45473 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__Q), .b(n_9518), .o(TIMEBOOST_net_14975) );
na02f02 TIMEBOOST_cell_41506 ( .a(TIMEBOOST_net_12991), .b(g57080_sb), .o(n_11662) );
in01s01 g62591_u0 ( .a(FE_OFN1242_n_4092), .o(g62591_sb) );
na02s01 TIMEBOOST_cell_39260 ( .a(TIMEBOOST_net_11868), .b(g64186_db), .o(n_4735) );
na02s02 TIMEBOOST_cell_41956 ( .a(TIMEBOOST_net_13216), .b(g58271_db), .o(n_9530) );
na02s01 TIMEBOOST_cell_16060 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__Q), .b(g65867_sb), .o(TIMEBOOST_net_3287) );
in01s01 g62592_u0 ( .a(FE_OFN1283_n_4097), .o(g62592_sb) );
na02s02 TIMEBOOST_cell_3173 ( .a(TIMEBOOST_net_166), .b(n_2473), .o(n_2474) );
na03s02 TIMEBOOST_cell_43319 ( .a(n_3514), .b(FE_OFN1206_n_6356), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__Q), .o(TIMEBOOST_net_13898) );
na02s01 TIMEBOOST_cell_22294 ( .a(g52478_da), .b(FE_OFN8_n_11877), .o(TIMEBOOST_net_6404) );
in01s02 g62593_u0 ( .a(FE_OFN1311_n_6624), .o(g62593_sb) );
na02s02 TIMEBOOST_cell_17017 ( .a(TIMEBOOST_net_3765), .b(g65248_sb), .o(n_2634) );
na02m02 TIMEBOOST_cell_3781 ( .a(TIMEBOOST_net_470), .b(n_4809), .o(n_5758) );
na02s02 TIMEBOOST_cell_18459 ( .a(TIMEBOOST_net_4486), .b(g62776_sb), .o(n_5441) );
in01s01 g62594_u0 ( .a(FE_OFN1203_n_4090), .o(g62594_sb) );
na02m02 TIMEBOOST_cell_20366 ( .a(n_3509), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__Q), .o(TIMEBOOST_net_5440) );
na02s02 TIMEBOOST_cell_41945 ( .a(TIMEBOOST_net_1835), .b(FE_OFN1083_n_13221), .o(TIMEBOOST_net_13211) );
na03m08 TIMEBOOST_cell_32863 ( .a(pciu_pciif_idsel_reg_in), .b(n_343), .c(n_8511), .o(TIMEBOOST_net_53) );
no02m02 g62595_u0 ( .a(n_2915), .b(conf_wb_err_addr_in_968), .o(g62595_p) );
ao12m02 g62595_u1 ( .a(g62595_p), .b(conf_wb_err_addr_in_968), .c(n_2915), .o(n_3467) );
in01s01 g62596_u0 ( .a(FE_OFN1294_n_4098), .o(g62596_sb) );
no02f04 TIMEBOOST_cell_12665 ( .a(TIMEBOOST_net_2899), .b(n_13348), .o(g53084_p) );
no04f08 TIMEBOOST_cell_32862 ( .a(TIMEBOOST_net_3149), .b(n_544), .c(n_715), .d(conf_wb_err_bc_in_848), .o(TIMEBOOST_net_3230) );
na02f02 TIMEBOOST_cell_41492 ( .a(TIMEBOOST_net_12984), .b(g57180_sb), .o(n_11575) );
in01s01 g62597_u0 ( .a(FE_OFN1207_n_6356), .o(g62597_sb) );
na02s01 TIMEBOOST_cell_39421 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_404), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_11949) );
na02m02 TIMEBOOST_cell_32446 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__Q), .o(TIMEBOOST_net_10134) );
na02s02 TIMEBOOST_cell_45675 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__Q), .b(n_4259), .o(TIMEBOOST_net_15076) );
in01s01 g62598_u0 ( .a(FE_OFN1207_n_6356), .o(g62598_sb) );
na02s02 TIMEBOOST_cell_38366 ( .a(TIMEBOOST_net_11421), .b(g63087_sb), .o(n_5080) );
na02f02 TIMEBOOST_cell_41532 ( .a(TIMEBOOST_net_13004), .b(g57224_sb), .o(n_11532) );
na02m02 TIMEBOOST_cell_41623 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_23__Q), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_13050) );
in01s01 g62599_u0 ( .a(FE_OFN1312_n_6624), .o(g62599_sb) );
na02s02 TIMEBOOST_cell_17015 ( .a(TIMEBOOST_net_3764), .b(g65246_sb), .o(n_2636) );
na03s02 TIMEBOOST_cell_37611 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__Q), .b(FE_OFN701_n_7845), .c(n_1591), .o(TIMEBOOST_net_11044) );
na02s02 TIMEBOOST_cell_16629 ( .a(TIMEBOOST_net_3571), .b(g65417_db), .o(n_3512) );
in01s01 g62600_u0 ( .a(FE_OFN1314_n_6624), .o(g62600_sb) );
na02m02 TIMEBOOST_cell_44001 ( .a(n_9561), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__Q), .o(TIMEBOOST_net_14239) );
na02f08 TIMEBOOST_cell_3785 ( .a(TIMEBOOST_net_472), .b(n_3379), .o(n_7618) );
na02s02 TIMEBOOST_cell_38368 ( .a(TIMEBOOST_net_11422), .b(g63073_sb), .o(n_5104) );
in01s01 g62601_u0 ( .a(FE_OFN1236_n_6391), .o(g62601_sb) );
na02s01 TIMEBOOST_cell_36377 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__Q), .b(g65865_sb), .o(TIMEBOOST_net_10427) );
na02s02 TIMEBOOST_cell_39896 ( .a(TIMEBOOST_net_12186), .b(g63005_sb), .o(n_5872) );
in01s01 TIMEBOOST_cell_8845 ( .a(TIMEBOOST_net_981), .o(TIMEBOOST_net_982) );
in01s01 g62602_u0 ( .a(FE_OFN1218_n_6886), .o(g62602_sb) );
na02m02 TIMEBOOST_cell_44177 ( .a(n_9031), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__Q), .o(TIMEBOOST_net_14327) );
na03s02 TIMEBOOST_cell_14015 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_394), .b(g54203_sb), .c(TIMEBOOST_net_522), .o(g53942_db) );
na02s02 TIMEBOOST_cell_39340 ( .a(TIMEBOOST_net_11908), .b(g65900_sb), .o(n_1571) );
in01s01 g62603_u0 ( .a(FE_OFN1218_n_6886), .o(g62603_sb) );
na03s02 TIMEBOOST_cell_20374 ( .a(TIMEBOOST_net_535), .b(g52637_da), .c(g52446_sb), .o(TIMEBOOST_net_5444) );
na02f02 TIMEBOOST_cell_42352 ( .a(TIMEBOOST_net_13414), .b(g57297_sb), .o(n_11454) );
na02s02 TIMEBOOST_cell_45676 ( .a(TIMEBOOST_net_15076), .b(FE_OFN1214_n_4151), .o(TIMEBOOST_net_12594) );
in01s01 g62604_u0 ( .a(FE_OFN1253_n_4143), .o(g62604_sb) );
na03s02 TIMEBOOST_cell_20376 ( .a(TIMEBOOST_net_532), .b(g52631_da), .c(g52393_sb), .o(TIMEBOOST_net_5445) );
na02m02 TIMEBOOST_cell_32672 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__Q), .o(TIMEBOOST_net_10247) );
na02f02 TIMEBOOST_cell_32671 ( .a(FE_OFN1559_n_12042), .b(TIMEBOOST_net_10246), .o(TIMEBOOST_net_6527) );
in01s01 g62605_u0 ( .a(FE_OFN1223_n_6391), .o(g62605_sb) );
na02m04 TIMEBOOST_cell_3175 ( .a(n_2457), .b(TIMEBOOST_net_167), .o(n_2983) );
na03s02 TIMEBOOST_cell_37603 ( .a(n_1607), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__Q), .c(FE_OFN716_n_8176), .o(TIMEBOOST_net_11040) );
na02m02 TIMEBOOST_cell_3176 ( .a(n_2982), .b(n_2458), .o(TIMEBOOST_net_168) );
in01s01 g62606_u0 ( .a(FE_OFN1233_n_6391), .o(g62606_sb) );
na02s01 TIMEBOOST_cell_36459 ( .a(FE_RN_484_0), .b(FE_OFN596_n_9694), .o(TIMEBOOST_net_10468) );
na02f04 TIMEBOOST_cell_38797 ( .a(n_8552), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__Q), .o(TIMEBOOST_net_11637) );
in01s01 TIMEBOOST_cell_8847 ( .a(TIMEBOOST_net_983), .o(TIMEBOOST_net_984) );
in01s01 g62607_u0 ( .a(n_4098), .o(g62607_sb) );
na02f02 TIMEBOOST_cell_44002 ( .a(TIMEBOOST_net_14239), .b(FE_OFN1423_n_8567), .o(TIMEBOOST_net_12871) );
na02s01 g62607_u2 ( .a(n_4400), .b(n_4098), .o(g62607_db) );
na02f02 TIMEBOOST_cell_44003 ( .a(n_9028), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__Q), .o(TIMEBOOST_net_14240) );
in01s01 g62608_u0 ( .a(FE_OFN1294_n_4098), .o(g62608_sb) );
na03f04 TIMEBOOST_cell_39149 ( .a(n_16241), .b(n_14000), .c(n_13999), .o(TIMEBOOST_net_11813) );
na02m02 TIMEBOOST_cell_32670 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__Q), .o(TIMEBOOST_net_10246) );
na02f02 TIMEBOOST_cell_32669 ( .a(FE_OFN1559_n_12042), .b(TIMEBOOST_net_10245), .o(TIMEBOOST_net_6525) );
in01s01 g62609_u0 ( .a(FE_OFN1241_n_4092), .o(g62609_sb) );
na02s01 TIMEBOOST_cell_36605 ( .a(TIMEBOOST_net_3694), .b(FE_OFN1044_n_2037), .o(TIMEBOOST_net_10541) );
na02m02 TIMEBOOST_cell_32668 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__Q), .o(TIMEBOOST_net_10245) );
na02f02 TIMEBOOST_cell_32667 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_10244), .o(TIMEBOOST_net_6520) );
in01s01 g62610_u0 ( .a(FE_OFN1200_n_4090), .o(g62610_sb) );
na02s01 TIMEBOOST_cell_45677 ( .a(n_4219), .b(FE_RN_720_0), .o(TIMEBOOST_net_15077) );
na02m02 TIMEBOOST_cell_32666 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__Q), .o(TIMEBOOST_net_10244) );
na02f02 TIMEBOOST_cell_32665 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_10243), .o(TIMEBOOST_net_6519) );
in01s01 g62611_u0 ( .a(FE_OFN1222_n_6391), .o(g62611_sb) );
na02m02 TIMEBOOST_cell_3177 ( .a(TIMEBOOST_net_168), .b(n_2457), .o(n_2459) );
na03s02 TIMEBOOST_cell_37613 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__Q), .b(FE_OFN699_n_7845), .c(n_2194), .o(TIMEBOOST_net_11045) );
na02m01 TIMEBOOST_cell_3178 ( .a(n_1515), .b(wishbone_slave_unit_pcim_sm_rdy_in), .o(TIMEBOOST_net_169) );
in01s01 g62612_u0 ( .a(FE_OFN1315_n_6624), .o(g62612_sb) );
na02f02 TIMEBOOST_cell_44004 ( .a(TIMEBOOST_net_14240), .b(FE_OFN1405_n_8567), .o(TIMEBOOST_net_13000) );
na02f02 TIMEBOOST_cell_3787 ( .a(TIMEBOOST_net_473), .b(n_15435), .o(n_4188) );
na02m02 TIMEBOOST_cell_44343 ( .a(n_9535), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__Q), .o(TIMEBOOST_net_14410) );
in01s01 g62613_u0 ( .a(FE_OFN1197_n_4090), .o(g62613_sb) );
na03s02 TIMEBOOST_cell_33970 ( .a(n_8892), .b(FE_OFN1671_n_9477), .c(g58367_da), .o(n_9459) );
na02m02 TIMEBOOST_cell_32664 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__1__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__1__Q), .o(TIMEBOOST_net_10243) );
na02f02 TIMEBOOST_cell_45474 ( .a(TIMEBOOST_net_14975), .b(FE_OFN1349_n_8567), .o(TIMEBOOST_net_14096) );
in01s01 g62614_u0 ( .a(FE_OFN1233_n_6391), .o(g62614_sb) );
na02s01 TIMEBOOST_cell_36461 ( .a(pci_target_unit_fifos_pcir_data_in), .b(g65716_db), .o(TIMEBOOST_net_10469) );
na02f02 TIMEBOOST_cell_38987 ( .a(TIMEBOOST_net_10103), .b(FE_OFN2158_n_16439), .o(TIMEBOOST_net_11732) );
in01s01 TIMEBOOST_cell_8849 ( .a(TIMEBOOST_net_985), .o(TIMEBOOST_net_986) );
in01s01 g62615_u0 ( .a(FE_OFN1272_n_4096), .o(g62615_sb) );
na02f02 TIMEBOOST_cell_3179 ( .a(TIMEBOOST_net_169), .b(n_2245), .o(n_6965) );
na03s02 TIMEBOOST_cell_37615 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__Q), .b(FE_OFN2084_n_8407), .c(n_2045), .o(TIMEBOOST_net_11046) );
na03s02 TIMEBOOST_cell_34250 ( .a(TIMEBOOST_net_9796), .b(FE_OFN1171_n_5592), .c(g62139_sb), .o(n_5554) );
in01s01 g62616_u0 ( .a(FE_OFN1214_n_4151), .o(g62616_sb) );
na02m02 TIMEBOOST_cell_42247 ( .a(n_9585), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__Q), .o(TIMEBOOST_net_13362) );
na02f02 TIMEBOOST_cell_41294 ( .a(TIMEBOOST_net_12885), .b(g57075_sb), .o(n_11668) );
na02m02 TIMEBOOST_cell_45475 ( .a(n_2051), .b(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q), .o(TIMEBOOST_net_14976) );
in01s01 g62617_u0 ( .a(FE_OFN1200_n_4090), .o(g62617_sb) );
na03s02 TIMEBOOST_cell_36757 ( .a(g64108_da), .b(g64108_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__Q), .o(TIMEBOOST_net_10617) );
na02f02 TIMEBOOST_cell_41292 ( .a(TIMEBOOST_net_12884), .b(g57241_sb), .o(n_11517) );
na02f02 TIMEBOOST_cell_41258 ( .a(TIMEBOOST_net_12867), .b(g57131_sb), .o(n_10473) );
in01s01 g62618_u0 ( .a(FE_OFN1320_n_6436), .o(g62618_sb) );
na02m02 TIMEBOOST_cell_44005 ( .a(n_9098), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__Q), .o(TIMEBOOST_net_14241) );
na02s02 TIMEBOOST_cell_38370 ( .a(TIMEBOOST_net_11423), .b(g62827_sb), .o(n_5323) );
na02f02 TIMEBOOST_cell_37101 ( .a(FE_RN_197_0), .b(n_10918), .o(TIMEBOOST_net_10789) );
in01s01 g62619_u0 ( .a(n_6319), .o(g62619_sb) );
na02s01 TIMEBOOST_cell_36465 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(g65753_sb), .o(TIMEBOOST_net_10471) );
na02m02 TIMEBOOST_cell_43571 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q), .b(n_4373), .o(TIMEBOOST_net_14024) );
na02s02 TIMEBOOST_cell_44865 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__Q), .b(FE_OFN1643_n_4671), .o(TIMEBOOST_net_14671) );
in01s01 g62620_u0 ( .a(FE_OFN1276_n_4096), .o(g62620_sb) );
na02s01 TIMEBOOST_cell_3181 ( .a(TIMEBOOST_net_170), .b(g60688_sb), .o(n_3880) );
na03s02 TIMEBOOST_cell_37617 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__Q), .b(FE_OFN2084_n_8407), .c(n_1929), .o(TIMEBOOST_net_11047) );
na03s02 TIMEBOOST_cell_34251 ( .a(TIMEBOOST_net_9795), .b(FE_OFN1168_n_5592), .c(g62097_sb), .o(n_5607) );
in01s01 g62621_u0 ( .a(FE_OFN1294_n_4098), .o(g62621_sb) );
na03s02 TIMEBOOST_cell_36759 ( .a(g60676_da), .b(g60676_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__Q), .o(TIMEBOOST_net_10618) );
na02m02 TIMEBOOST_cell_32658 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__6__Q), .o(TIMEBOOST_net_10240) );
na02m02 TIMEBOOST_cell_41260 ( .a(TIMEBOOST_net_12868), .b(g57134_sb), .o(n_10469) );
in01s01 g62622_u0 ( .a(FE_OFN1315_n_6624), .o(g62622_sb) );
na02f02 TIMEBOOST_cell_44006 ( .a(TIMEBOOST_net_14241), .b(FE_OFN1396_n_8567), .o(TIMEBOOST_net_12863) );
na02s01 TIMEBOOST_cell_38372 ( .a(TIMEBOOST_net_11424), .b(g62721_sb), .o(n_5541) );
na02s01 TIMEBOOST_cell_40388 ( .a(TIMEBOOST_net_12432), .b(g64325_db), .o(n_3851) );
in01s01 g62623_u0 ( .a(FE_OFN1235_n_6391), .o(g62623_sb) );
na02s01 TIMEBOOST_cell_36373 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__Q), .b(g65865_sb), .o(TIMEBOOST_net_10425) );
na03s02 TIMEBOOST_cell_39361 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__Q), .b(FE_OFN707_n_8119), .c(n_1893), .o(TIMEBOOST_net_11919) );
in01s01 TIMEBOOST_cell_8851 ( .a(TIMEBOOST_net_987), .o(TIMEBOOST_net_988) );
in01s01 g62624_u0 ( .a(FE_OFN1218_n_6886), .o(g62624_sb) );
na02f02 TIMEBOOST_cell_42248 ( .a(TIMEBOOST_net_13362), .b(FE_OFN1408_n_8567), .o(TIMEBOOST_net_12320) );
na02s01 TIMEBOOST_cell_2889 ( .a(TIMEBOOST_net_24), .b(n_875), .o(n_876) );
na02s02 TIMEBOOST_cell_31410 ( .a(n_3792), .b(g65015_sb), .o(TIMEBOOST_net_9616) );
in01s01 g62625_u0 ( .a(FE_OFN1234_n_6391), .o(g62625_sb) );
na02s01 TIMEBOOST_cell_36437 ( .a(pci_target_unit_fifos_pciw_addr_data_in_123), .b(g64172_sb), .o(TIMEBOOST_net_10457) );
na02f04 TIMEBOOST_cell_38798 ( .a(TIMEBOOST_net_11637), .b(FE_OFN2185_n_8567), .o(TIMEBOOST_net_10692) );
in01s01 TIMEBOOST_cell_8853 ( .a(TIMEBOOST_net_989), .o(TIMEBOOST_net_990) );
in01s01 g62626_u0 ( .a(FE_OFN1232_n_6391), .o(g62626_sb) );
na02f02 TIMEBOOST_cell_39008 ( .a(TIMEBOOST_net_11742), .b(g52532_sb), .o(n_13687) );
na02f02 TIMEBOOST_cell_38814 ( .a(TIMEBOOST_net_11645), .b(n_10256), .o(TIMEBOOST_net_10695) );
in01s01 TIMEBOOST_cell_8855 ( .a(TIMEBOOST_net_991), .o(TIMEBOOST_net_992) );
in01s01 g62627_u0 ( .a(FE_OFN1236_n_6391), .o(g62627_sb) );
na02s01 TIMEBOOST_cell_3414 ( .a(g58112_sb), .b(g58112_db), .o(TIMEBOOST_net_287) );
na02f02 TIMEBOOST_cell_42200 ( .a(TIMEBOOST_net_13338), .b(FE_OFN1388_n_8567), .o(TIMEBOOST_net_12290) );
na02s01 TIMEBOOST_cell_15795 ( .a(TIMEBOOST_net_3154), .b(g67049_sb), .o(n_1470) );
in01s01 g62628_u0 ( .a(FE_OFN1283_n_4097), .o(g62628_sb) );
na02s01 TIMEBOOST_cell_3183 ( .a(TIMEBOOST_net_171), .b(g60688_sb), .o(n_3872) );
na02m02 TIMEBOOST_cell_42249 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__Q), .b(n_9554), .o(TIMEBOOST_net_13363) );
na02s02 TIMEBOOST_cell_45678 ( .a(TIMEBOOST_net_15077), .b(FE_OFN1250_n_4093), .o(TIMEBOOST_net_13302) );
in01s01 g62629_u0 ( .a(FE_OFN1213_n_4151), .o(g62629_sb) );
na02f02 TIMEBOOST_cell_38891 ( .a(TIMEBOOST_net_2805), .b(n_3037), .o(TIMEBOOST_net_11684) );
na02s01 TIMEBOOST_cell_17005 ( .a(TIMEBOOST_net_3759), .b(g65704_db), .o(n_1613) );
na02s02 TIMEBOOST_cell_43493 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__Q), .b(n_3606), .o(TIMEBOOST_net_13985) );
in01s01 g62630_u0 ( .a(n_6232), .o(g62630_sb) );
na02s01 TIMEBOOST_cell_36321 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__22__Q), .b(g65964_sb), .o(TIMEBOOST_net_10399) );
na02s02 TIMEBOOST_cell_45153 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__Q), .b(n_4325), .o(TIMEBOOST_net_14815) );
na02s02 TIMEBOOST_cell_42825 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__Q), .b(g58303_sb), .o(TIMEBOOST_net_13651) );
in01s01 g62631_u0 ( .a(FE_OFN1253_n_4143), .o(g62631_sb) );
na02f02 TIMEBOOST_cell_42250 ( .a(TIMEBOOST_net_13363), .b(FE_OFN1419_n_8567), .o(TIMEBOOST_net_12321) );
na02m02 TIMEBOOST_cell_32656 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q), .o(TIMEBOOST_net_10239) );
na02f02 TIMEBOOST_cell_41262 ( .a(TIMEBOOST_net_12869), .b(g57113_sb), .o(n_11633) );
in01s01 g62632_u0 ( .a(n_6287), .o(g62632_sb) );
na03s02 TIMEBOOST_cell_38059 ( .a(g64295_da), .b(g64295_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__Q), .o(TIMEBOOST_net_11268) );
na02s01 TIMEBOOST_cell_17126 ( .a(pci_target_unit_del_sync_addr_in_222), .b(parchk_pci_ad_reg_in_1223), .o(TIMEBOOST_net_3820) );
na02s01 TIMEBOOST_cell_31802 ( .a(configuration_wb_err_addr_544), .b(TIMEBOOST_net_974), .o(TIMEBOOST_net_9812) );
in01s01 g62633_u0 ( .a(FE_OFN1323_n_6436), .o(g62633_sb) );
na02m02 TIMEBOOST_cell_44007 ( .a(n_9415), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__Q), .o(TIMEBOOST_net_14242) );
na02s02 TIMEBOOST_cell_18541 ( .a(TIMEBOOST_net_4527), .b(g63176_sb), .o(n_4947) );
na02s01 TIMEBOOST_cell_40390 ( .a(TIMEBOOST_net_12433), .b(g65278_db), .o(n_4288) );
in01s01 g62634_u0 ( .a(FE_OFN1223_n_6391), .o(g62634_sb) );
na02s01 TIMEBOOST_cell_3185 ( .a(TIMEBOOST_net_172), .b(g60688_sb), .o(n_3524) );
na02s01 TIMEBOOST_cell_37455 ( .a(pci_target_unit_del_sync_addr_in_217), .b(parchk_pci_ad_reg_in_1218), .o(TIMEBOOST_net_10966) );
na02s01 TIMEBOOST_cell_42622 ( .a(TIMEBOOST_net_13549), .b(g64798_db), .o(n_3758) );
in01s01 g62635_u0 ( .a(FE_OFN1315_n_6624), .o(g62635_sb) );
na02s02 TIMEBOOST_cell_42962 ( .a(TIMEBOOST_net_13719), .b(g52634_da), .o(TIMEBOOST_net_13184) );
na02s01 TIMEBOOST_cell_38374 ( .a(TIMEBOOST_net_11425), .b(n_4528), .o(n_6135) );
na02s02 TIMEBOOST_cell_38678 ( .a(TIMEBOOST_net_11577), .b(g62478_sb), .o(n_6631) );
in01s02 g62636_u0 ( .a(FE_OFN1322_n_6436), .o(g62636_sb) );
na02f02 TIMEBOOST_cell_44008 ( .a(TIMEBOOST_net_14242), .b(FE_OFN1387_n_8567), .o(TIMEBOOST_net_12870) );
na02s01 TIMEBOOST_cell_18545 ( .a(TIMEBOOST_net_4529), .b(g63122_sb), .o(n_5012) );
na02s01 TIMEBOOST_cell_18055 ( .a(TIMEBOOST_net_4284), .b(g65367_db), .o(n_4251) );
in01s01 g62637_u0 ( .a(FE_OFN1289_n_4098), .o(g62637_sb) );
na02m02 TIMEBOOST_cell_42251 ( .a(n_9564), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__Q), .o(TIMEBOOST_net_13364) );
na02s02 TIMEBOOST_cell_45154 ( .a(TIMEBOOST_net_14815), .b(FE_OFN1207_n_6356), .o(TIMEBOOST_net_12025) );
in01s01 g62638_u0 ( .a(FE_OFN1248_n_4093), .o(g62638_sb) );
na02s01 TIMEBOOST_cell_3187 ( .a(TIMEBOOST_net_173), .b(g60688_sb), .o(n_3205) );
na02f02 g53867_u0 ( .a(n_13436), .b(n_2100), .o(n_13650) );
na02f02 TIMEBOOST_cell_44344 ( .a(TIMEBOOST_net_14410), .b(FE_OFN1400_n_8567), .o(TIMEBOOST_net_12692) );
in01s01 g62639_u0 ( .a(FE_OFN1293_n_4098), .o(g62639_sb) );
na02f02 TIMEBOOST_cell_44178 ( .a(TIMEBOOST_net_14327), .b(FE_OFN1368_n_8567), .o(TIMEBOOST_net_13398) );
na02s02 TIMEBOOST_cell_39898 ( .a(TIMEBOOST_net_12187), .b(g62646_sb), .o(n_6257) );
in01s01 g62640_u0 ( .a(FE_OFN1225_n_6391), .o(g62640_sb) );
na02s01 TIMEBOOST_cell_3189 ( .a(TIMEBOOST_net_174), .b(g60688_sb), .o(n_7217) );
na02s01 TIMEBOOST_cell_18295 ( .a(n_4753), .b(TIMEBOOST_net_4404), .o(n_7145) );
na02s01 TIMEBOOST_cell_31409 ( .a(TIMEBOOST_net_9615), .b(g65000_db), .o(n_3641) );
in01s01 g62641_u0 ( .a(FE_OFN1276_n_4096), .o(g62641_sb) );
na02s01 TIMEBOOST_cell_3191 ( .a(TIMEBOOST_net_175), .b(n_2420), .o(n_2491) );
na02s01 TIMEBOOST_cell_18289 ( .a(n_4768), .b(TIMEBOOST_net_4401), .o(n_7189) );
na02m02 TIMEBOOST_cell_44009 ( .a(n_9810), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__Q), .o(TIMEBOOST_net_14243) );
in01s01 g62642_u0 ( .a(FE_OFN1241_n_4092), .o(g62642_sb) );
na02m02 TIMEBOOST_cell_44179 ( .a(n_9407), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q), .o(TIMEBOOST_net_14328) );
na02s02 TIMEBOOST_cell_39900 ( .a(TIMEBOOST_net_12188), .b(g63155_sb), .o(n_5830) );
na02s01 TIMEBOOST_cell_2898 ( .a(n_519), .b(n_879), .o(TIMEBOOST_net_29) );
in01s01 g62643_u0 ( .a(FE_OFN1243_n_4092), .o(g62643_sb) );
na02f02 TIMEBOOST_cell_44180 ( .a(TIMEBOOST_net_14328), .b(FE_OFN1389_n_8567), .o(TIMEBOOST_net_12752) );
na02m02 TIMEBOOST_cell_32654 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__Q), .o(TIMEBOOST_net_10238) );
na02f02 TIMEBOOST_cell_41264 ( .a(TIMEBOOST_net_12870), .b(g57579_sb), .o(n_11173) );
in01s01 g62644_u0 ( .a(FE_OFN1233_n_6391), .o(g62644_sb) );
in01s01 TIMEBOOST_cell_45895 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_), .o(TIMEBOOST_net_15202) );
na02s02 TIMEBOOST_cell_39902 ( .a(TIMEBOOST_net_12189), .b(g62647_sb), .o(n_6254) );
in01s01 TIMEBOOST_cell_8857 ( .a(TIMEBOOST_net_993), .o(TIMEBOOST_net_994) );
in01s01 g62645_u0 ( .a(FE_OFN1284_n_4097), .o(g62645_sb) );
na02f02 TIMEBOOST_cell_44010 ( .a(TIMEBOOST_net_14243), .b(FE_OFN1388_n_8567), .o(TIMEBOOST_net_12869) );
na02s01 TIMEBOOST_cell_18291 ( .a(n_4770), .b(TIMEBOOST_net_4402), .o(n_7177) );
na02m02 TIMEBOOST_cell_3194 ( .a(n_1269), .b(n_3007), .o(TIMEBOOST_net_177) );
in01s01 g62646_u0 ( .a(FE_OFN1234_n_6391), .o(g62646_sb) );
na02s01 TIMEBOOST_cell_37975 ( .a(g61956_sb), .b(g61956_db), .o(TIMEBOOST_net_11226) );
na02s02 TIMEBOOST_cell_38626 ( .a(TIMEBOOST_net_11551), .b(g62670_sb), .o(n_6199) );
in01s01 TIMEBOOST_cell_8859 ( .a(TIMEBOOST_net_995), .o(TIMEBOOST_net_996) );
in01s01 g62647_u0 ( .a(n_6431), .o(g62647_sb) );
na02s01 TIMEBOOST_cell_37205 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(g65692_sb), .o(TIMEBOOST_net_10841) );
na02s01 TIMEBOOST_cell_17128 ( .a(pci_target_unit_del_sync_addr_in_224), .b(parchk_pci_ad_reg_in_1225), .o(TIMEBOOST_net_3821) );
na02f02 TIMEBOOST_cell_36926 ( .a(TIMEBOOST_net_10701), .b(g52608_sb), .o(n_10213) );
in01s01 g62648_u0 ( .a(FE_OFN1224_n_6391), .o(g62648_sb) );
na02m04 TIMEBOOST_cell_3195 ( .a(n_3013), .b(TIMEBOOST_net_177), .o(n_3359) );
na02s01 TIMEBOOST_cell_18305 ( .a(n_4772), .b(TIMEBOOST_net_4409), .o(n_7182) );
na03f04 TIMEBOOST_cell_22380 ( .a(n_14226), .b(n_14055), .c(n_13982), .o(TIMEBOOST_net_6447) );
in01s01 g62649_u0 ( .a(FE_OFN1223_n_6391), .o(g62649_sb) );
na02m02 TIMEBOOST_cell_3197 ( .a(TIMEBOOST_net_178), .b(n_2754), .o(n_3200) );
na02s01 TIMEBOOST_cell_18293 ( .a(n_4773), .b(TIMEBOOST_net_4403), .o(n_7161) );
na02s02 TIMEBOOST_cell_3198 ( .a(n_1436), .b(wishbone_slave_unit_pcim_if_del_burst_in), .o(TIMEBOOST_net_179) );
in01s01 g62650_u0 ( .a(FE_OFN1272_n_4096), .o(g62650_sb) );
na02m02 TIMEBOOST_cell_3199 ( .a(TIMEBOOST_net_179), .b(n_3313), .o(n_3436) );
na02s01 TIMEBOOST_cell_18303 ( .a(n_4774), .b(TIMEBOOST_net_4408), .o(n_7205) );
na02f02 TIMEBOOST_cell_43776 ( .a(TIMEBOOST_net_14126), .b(FE_OFN1368_n_8567), .o(TIMEBOOST_net_12943) );
in01s01 g62651_u0 ( .a(FE_OFN1200_n_4090), .o(g62651_sb) );
na02m02 TIMEBOOST_cell_44181 ( .a(n_9137), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__Q), .o(TIMEBOOST_net_14329) );
na02m02 TIMEBOOST_cell_32652 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q), .o(TIMEBOOST_net_10237) );
na02f02 TIMEBOOST_cell_41266 ( .a(TIMEBOOST_net_12871), .b(g57371_sb), .o(n_11379) );
in01s01 g62652_u0 ( .a(FE_OFN1242_n_4092), .o(g62652_sb) );
na02s01 TIMEBOOST_cell_36277 ( .a(TIMEBOOST_net_9281), .b(n_574), .o(TIMEBOOST_net_10377) );
na02m02 TIMEBOOST_cell_32650 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__Q), .o(TIMEBOOST_net_10236) );
na02f02 TIMEBOOST_cell_41268 ( .a(TIMEBOOST_net_12872), .b(g57142_sb), .o(n_10465) );
in01s01 g62653_u0 ( .a(FE_OFN1193_n_6935), .o(g62653_sb) );
na02m04 TIMEBOOST_cell_3201 ( .a(n_2993), .b(TIMEBOOST_net_180), .o(n_3353) );
na02s01 TIMEBOOST_cell_18307 ( .a(n_4775), .b(TIMEBOOST_net_4410), .o(n_7171) );
na02s01 TIMEBOOST_cell_3202 ( .a(n_2648), .b(n_8511), .o(TIMEBOOST_net_181) );
in01s01 g62654_u0 ( .a(n_6645), .o(g62654_sb) );
na02s01 TIMEBOOST_cell_36447 ( .a(pci_target_unit_fifos_pcir_data_in_172), .b(g65795_sb), .o(TIMEBOOST_net_10462) );
na02m02 TIMEBOOST_cell_44011 ( .a(n_9106), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__Q), .o(TIMEBOOST_net_14244) );
na02f02 TIMEBOOST_cell_41146 ( .a(TIMEBOOST_net_12811), .b(g57333_sb), .o(n_11417) );
in01s01 g62655_u0 ( .a(n_6232), .o(g62655_sb) );
na02s01 TIMEBOOST_cell_45064 ( .a(TIMEBOOST_net_14770), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_11193) );
na02s01 TIMEBOOST_cell_36491 ( .a(n_2526), .b(g66410_db), .o(TIMEBOOST_net_10484) );
na02s01 TIMEBOOST_cell_31408 ( .a(n_3749), .b(g65000_sb), .o(TIMEBOOST_net_9615) );
in01s01 g62656_u0 ( .a(FE_OFN1235_n_6391), .o(g62656_sb) );
na02f04 TIMEBOOST_cell_20682 ( .a(g75072_sb), .b(n_16070), .o(TIMEBOOST_net_5598) );
na02s02 TIMEBOOST_cell_38376 ( .a(TIMEBOOST_net_11426), .b(g62794_sb), .o(n_5399) );
na02s01 TIMEBOOST_cell_17004 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(g65704_sb), .o(TIMEBOOST_net_3759) );
in01s01 g62657_u0 ( .a(FE_OFN1247_n_4093), .o(g62657_sb) );
na02s02 TIMEBOOST_cell_36547 ( .a(n_4488), .b(g64826_sb), .o(TIMEBOOST_net_10512) );
na02m02 TIMEBOOST_cell_32648 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__Q), .o(TIMEBOOST_net_10235) );
na02f02 TIMEBOOST_cell_41270 ( .a(TIMEBOOST_net_12873), .b(g57493_sb), .o(n_11243) );
in01s01 g62658_u0 ( .a(FE_OFN1249_n_4093), .o(g62658_sb) );
na02s01 TIMEBOOST_cell_36549 ( .a(n_4452), .b(g64755_sb), .o(TIMEBOOST_net_10513) );
na02m02 TIMEBOOST_cell_32646 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q), .o(TIMEBOOST_net_10234) );
na02f02 TIMEBOOST_cell_41272 ( .a(TIMEBOOST_net_12874), .b(g57436_sb), .o(n_11300) );
in01s01 g62659_u0 ( .a(FE_OFN1212_n_4151), .o(g62659_sb) );
na02s01 TIMEBOOST_cell_36551 ( .a(n_4672), .b(g64748_sb), .o(TIMEBOOST_net_10514) );
na02f02 TIMEBOOST_cell_37055 ( .a(TIMEBOOST_net_10130), .b(n_13901), .o(TIMEBOOST_net_10766) );
na02f02 TIMEBOOST_cell_37054 ( .a(FE_OFN1593_n_13741), .b(TIMEBOOST_net_10765), .o(g53234_p) );
in01s02 g62660_u0 ( .a(FE_OFN1311_n_6624), .o(g62660_sb) );
na02m02 TIMEBOOST_cell_44012 ( .a(TIMEBOOST_net_14244), .b(FE_OFN1396_n_8567), .o(TIMEBOOST_net_12868) );
na02s02 TIMEBOOST_cell_38378 ( .a(TIMEBOOST_net_11427), .b(g62792_sb), .o(n_5404) );
in01s01 g62661_u0 ( .a(FE_OFN1283_n_4097), .o(g62661_sb) );
na02s01 TIMEBOOST_cell_36497 ( .a(pci_target_unit_del_sync_addr_in_233), .b(g66420_db), .o(TIMEBOOST_net_10487) );
na02m02 TIMEBOOST_cell_32644 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__Q), .o(TIMEBOOST_net_10233) );
na02f02 TIMEBOOST_cell_41274 ( .a(TIMEBOOST_net_12875), .b(g57592_sb), .o(n_10286) );
in01s01 g62662_u0 ( .a(FE_OFN1231_n_6391), .o(g62662_sb) );
na02m02 TIMEBOOST_cell_44013 ( .a(n_9721), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__Q), .o(TIMEBOOST_net_14245) );
na02s02 TIMEBOOST_cell_36555 ( .a(n_3764), .b(g64786_sb), .o(TIMEBOOST_net_10516) );
na02m02 TIMEBOOST_cell_37059 ( .a(g52476_da), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_10768) );
in01s02 g62663_u0 ( .a(FE_OFN1311_n_6624), .o(g62663_sb) );
na02f02 TIMEBOOST_cell_44014 ( .a(TIMEBOOST_net_14245), .b(FE_OFN1422_n_8567), .o(TIMEBOOST_net_12922) );
na02f04 TIMEBOOST_cell_3801 ( .a(TIMEBOOST_net_480), .b(n_7216), .o(n_7704) );
na02m02 TIMEBOOST_cell_41633 ( .a(n_9114), .b(wishbone_slave_unit_del_sync_addr_out_reg_5__Q), .o(TIMEBOOST_net_13055) );
in01s01 g62664_u0 ( .a(n_6287), .o(g62664_sb) );
na02s01 TIMEBOOST_cell_36333 ( .a(parchk_pci_ad_reg_in_1206), .b(g67040_db), .o(TIMEBOOST_net_10405) );
na02s01 TIMEBOOST_cell_3395 ( .a(TIMEBOOST_net_277), .b(FE_OFN1628_n_4438), .o(n_4433) );
na02s02 TIMEBOOST_cell_43431 ( .a(n_4901), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__Q), .o(TIMEBOOST_net_13954) );
in01s01 g62665_u0 ( .a(FE_OFN1269_n_4095), .o(g62665_sb) );
na02s01 TIMEBOOST_cell_36531 ( .a(TIMEBOOST_net_3397), .b(FE_OFN917_n_4725), .o(TIMEBOOST_net_10504) );
na02m02 TIMEBOOST_cell_32642 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__21__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__21__Q), .o(TIMEBOOST_net_10232) );
na02f02 TIMEBOOST_cell_41276 ( .a(TIMEBOOST_net_12876), .b(g57169_sb), .o(n_10455) );
in01s01 g62666_u0 ( .a(FE_OFN1314_n_6624), .o(g62666_sb) );
na02m02 TIMEBOOST_cell_44015 ( .a(n_9608), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__Q), .o(TIMEBOOST_net_14246) );
na02f02 TIMEBOOST_cell_3803 ( .a(TIMEBOOST_net_481), .b(n_16452), .o(n_7624) );
na02f02 TIMEBOOST_cell_45476 ( .a(TIMEBOOST_net_14976), .b(n_9144), .o(TIMEBOOST_net_14457) );
in01s01 g62667_u0 ( .a(FE_OFN1293_n_4098), .o(g62667_sb) );
na02s01 TIMEBOOST_cell_36557 ( .a(pci_target_unit_fifos_pciw_addr_data_in_143), .b(g64171_sb), .o(TIMEBOOST_net_10517) );
na03s02 TIMEBOOST_cell_36747 ( .a(g64093_da), .b(g64093_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__Q), .o(TIMEBOOST_net_10612) );
na02s01 g62000_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__Q), .b(FE_OFN2258_n_8060), .o(g62000_db) );
in01s01 g62668_u0 ( .a(FE_OFN1285_n_4097), .o(g62668_sb) );
na02s02 TIMEBOOST_cell_42022 ( .a(TIMEBOOST_net_13249), .b(g62357_sb), .o(n_6885) );
na02f02 TIMEBOOST_cell_44016 ( .a(TIMEBOOST_net_14246), .b(FE_OFN1411_n_8567), .o(TIMEBOOST_net_12903) );
na02m02 TIMEBOOST_cell_44017 ( .a(n_9497), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__Q), .o(TIMEBOOST_net_14247) );
in01s01 g62669_u0 ( .a(FE_OFN1202_n_4090), .o(g62669_sb) );
na02s01 TIMEBOOST_cell_3203 ( .a(TIMEBOOST_net_181), .b(n_3021), .o(n_3377) );
na02f02 TIMEBOOST_cell_37809 ( .a(TIMEBOOST_net_9677), .b(g54328_sb), .o(TIMEBOOST_net_11143) );
na02f02 TIMEBOOST_cell_44018 ( .a(TIMEBOOST_net_14247), .b(FE_OFN1374_n_8567), .o(TIMEBOOST_net_12841) );
in01s01 g62670_u0 ( .a(FE_OFN1247_n_4093), .o(g62670_sb) );
na02s01 TIMEBOOST_cell_17339 ( .a(TIMEBOOST_net_3926), .b(g58161_sb), .o(n_9627) );
na02f02 TIMEBOOST_cell_44390 ( .a(TIMEBOOST_net_14433), .b(FE_OFN1397_n_8567), .o(TIMEBOOST_net_12704) );
na02s02 TIMEBOOST_cell_43255 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q), .b(n_3629), .o(TIMEBOOST_net_13866) );
in01s01 g62671_u0 ( .a(FE_OFN1270_n_4095), .o(g62671_sb) );
na02s01 TIMEBOOST_cell_36561 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(g64160_sb), .o(TIMEBOOST_net_10519) );
na02s01 TIMEBOOST_cell_16816 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__Q), .b(g65315_sb), .o(TIMEBOOST_net_3665) );
na02m02 TIMEBOOST_cell_32640 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__Q), .o(TIMEBOOST_net_10231) );
in01s01 g62672_u0 ( .a(FE_OFN1261_n_4143), .o(g62672_sb) );
na02s01 TIMEBOOST_cell_36563 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__Q), .b(FE_OFN527_n_9899), .o(TIMEBOOST_net_10520) );
na02s02 TIMEBOOST_cell_43375 ( .a(n_351), .b(n_4909), .o(TIMEBOOST_net_13926) );
na02f02 TIMEBOOST_cell_41192 ( .a(TIMEBOOST_net_12834), .b(g57188_sb), .o(n_10449) );
in01s01 g62673_u0 ( .a(FE_OFN1312_n_6624), .o(g62673_sb) );
na02s01 TIMEBOOST_cell_45588 ( .a(TIMEBOOST_net_15032), .b(FE_OFN2254_n_9687), .o(TIMEBOOST_net_10928) );
na02f04 TIMEBOOST_cell_3805 ( .a(TIMEBOOST_net_482), .b(n_3202), .o(n_3491) );
na02f02 TIMEBOOST_cell_3806 ( .a(n_2754), .b(n_3192), .o(TIMEBOOST_net_483) );
in01s01 g62674_u0 ( .a(FE_OFN1249_n_4093), .o(g62674_sb) );
na02s01 TIMEBOOST_cell_36565 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__Q), .b(FE_OFN535_n_9823), .o(TIMEBOOST_net_10521) );
na02f02 TIMEBOOST_cell_21825 ( .a(TIMEBOOST_net_6169), .b(n_2870), .o(n_4172) );
na02m02 TIMEBOOST_cell_32526 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__Q), .o(TIMEBOOST_net_10174) );
in01s01 g62675_u0 ( .a(FE_OFN1202_n_4090), .o(g62675_sb) );
na02s04 TIMEBOOST_cell_3205 ( .a(n_1692), .b(TIMEBOOST_net_182), .o(n_2179) );
na03s02 TIMEBOOST_cell_37595 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__Q), .b(FE_OFN701_n_7845), .c(n_1605), .o(TIMEBOOST_net_11036) );
na02s02 TIMEBOOST_cell_31405 ( .a(TIMEBOOST_net_9613), .b(g65040_db), .o(n_4328) );
in01s01 g62676_u0 ( .a(FE_OFN365_n_4093), .o(g62676_sb) );
na02s01 TIMEBOOST_cell_36567 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q), .b(FE_OFN1631_n_9531), .o(TIMEBOOST_net_10522) );
na02s01 TIMEBOOST_cell_42937 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__Q), .b(FE_OFN584_n_9692), .o(TIMEBOOST_net_13707) );
na03s01 TIMEBOOST_cell_34283 ( .a(TIMEBOOST_net_9811), .b(FE_OFN1174_n_5592), .c(g62121_sb), .o(n_5575) );
in01s01 g62677_u0 ( .a(n_6554), .o(g62677_sb) );
na02s02 TIMEBOOST_cell_43643 ( .a(n_3548), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__Q), .o(TIMEBOOST_net_14060) );
na02m04 TIMEBOOST_cell_3397 ( .a(TIMEBOOST_net_278), .b(n_2691), .o(n_2915) );
na02m02 TIMEBOOST_cell_3398 ( .a(n_2316), .b(n_2308), .o(TIMEBOOST_net_279) );
in01s01 g62678_u0 ( .a(FE_OFN1268_n_4095), .o(g62678_sb) );
na02s01 TIMEBOOST_cell_36569 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__Q), .b(g65822_sb), .o(TIMEBOOST_net_10523) );
na03m02 TIMEBOOST_cell_45477 ( .a(TIMEBOOST_net_613), .b(g52403_sb), .c(g52403_db), .o(TIMEBOOST_net_14977) );
na02s02 TIMEBOOST_cell_41980 ( .a(TIMEBOOST_net_13228), .b(g62932_sb), .o(n_6017) );
in01s01 g62679_u0 ( .a(FE_OFN1230_n_6391), .o(g62679_sb) );
na02s01 TIMEBOOST_cell_36305 ( .a(parchk_pci_ad_reg_in_1232), .b(g67055_db), .o(TIMEBOOST_net_10391) );
na02s02 TIMEBOOST_cell_43592 ( .a(TIMEBOOST_net_14034), .b(FE_OFN1320_n_6436), .o(TIMEBOOST_net_12213) );
na03f02 TIMEBOOST_cell_3512 ( .a(n_4806), .b(n_2802), .c(n_2843), .o(TIMEBOOST_net_336) );
in01s01 g62680_u0 ( .a(FE_OFN1268_n_4095), .o(g62680_sb) );
na02s01 TIMEBOOST_cell_36603 ( .a(TIMEBOOST_net_3702), .b(FE_OFN1042_n_2037), .o(TIMEBOOST_net_10540) );
na02m02 TIMEBOOST_cell_32528 ( .a(n_271), .b(n_366), .o(TIMEBOOST_net_10175) );
in01s01 TIMEBOOST_cell_32829 ( .a(TIMEBOOST_net_10330), .o(TIMEBOOST_net_10329) );
in01s01 g62681_u0 ( .a(FE_OFN1268_n_4095), .o(g62681_sb) );
na02s01 TIMEBOOST_cell_36571 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__Q), .b(g64224_sb), .o(TIMEBOOST_net_10524) );
na02s02 TIMEBOOST_cell_43593 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__Q), .b(n_4519), .o(TIMEBOOST_net_14035) );
na02f02 TIMEBOOST_cell_41148 ( .a(TIMEBOOST_net_12812), .b(g57209_sb), .o(n_11547) );
in01s01 g62682_u0 ( .a(FE_OFN1208_n_6356), .o(g62682_sb) );
na02s01 TIMEBOOST_cell_36573 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__Q), .b(g65954_sb), .o(TIMEBOOST_net_10525) );
na02f02 TIMEBOOST_cell_32587 ( .a(n_12010), .b(TIMEBOOST_net_10204), .o(TIMEBOOST_net_6419) );
na03s02 TIMEBOOST_cell_34269 ( .a(TIMEBOOST_net_9810), .b(FE_OFN1171_n_5592), .c(g62137_sb), .o(n_5556) );
in01s01 g62683_u0 ( .a(FE_OFN1250_n_4093), .o(g62683_sb) );
na02m04 TIMEBOOST_cell_3207 ( .a(TIMEBOOST_net_183), .b(n_1694), .o(n_2175) );
na02s01 TIMEBOOST_cell_18285 ( .a(n_4779), .b(TIMEBOOST_net_4399), .o(n_7209) );
no02m01 TIMEBOOST_cell_3208 ( .a(wishbone_slave_unit_pcim_if_del_req_in), .b(wishbone_slave_unit_pci_initiator_if_err_recovery), .o(TIMEBOOST_net_184) );
in01s01 g62684_u0 ( .a(FE_OFN1264_n_4095), .o(g62684_sb) );
na02s02 TIMEBOOST_cell_36575 ( .a(g65230_sb), .b(pci_target_unit_del_sync_bc_in_201), .o(TIMEBOOST_net_10526) );
na02s01 TIMEBOOST_cell_30855 ( .a(TIMEBOOST_net_9338), .b(g65044_db), .o(n_3623) );
na02s01 TIMEBOOST_cell_15839 ( .a(TIMEBOOST_net_3176), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_385), .o(TIMEBOOST_net_73) );
in01s01 g62685_u0 ( .a(FE_OFN1269_n_4095), .o(g62685_sb) );
na02s01 TIMEBOOST_cell_36577 ( .a(wbu_latency_tim_val_in_248), .b(n_6986), .o(TIMEBOOST_net_10527) );
na02s01 TIMEBOOST_cell_15861 ( .a(TIMEBOOST_net_3187), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_395), .o(TIMEBOOST_net_77) );
na02m02 TIMEBOOST_cell_30797 ( .a(g58767_db), .b(TIMEBOOST_net_9309), .o(n_9865) );
oa12m02 g62686_u0 ( .a(n_2955), .b(n_2954), .c(wbu_addr_in_273), .o(n_3332) );
oa12m02 g62687_u0 ( .a(n_3148), .b(n_3147), .c(wbu_addr_in_276), .o(n_3465) );
in01s01 g62688_u0 ( .a(FE_OFN1231_n_6391), .o(g62688_sb) );
na02s02 TIMEBOOST_cell_43432 ( .a(TIMEBOOST_net_13954), .b(n_6431), .o(TIMEBOOST_net_12208) );
na02s01 TIMEBOOST_cell_36579 ( .a(TIMEBOOST_net_252), .b(g61870_sb), .o(TIMEBOOST_net_10528) );
na02f02 TIMEBOOST_cell_41278 ( .a(TIMEBOOST_net_12877), .b(g57295_sb), .o(n_11457) );
in01s01 g62689_u0 ( .a(FE_OFN1243_n_4092), .o(g62689_sb) );
na02s01 TIMEBOOST_cell_36533 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(g65754_sb), .o(TIMEBOOST_net_10505) );
na02m02 TIMEBOOST_cell_44391 ( .a(n_9526), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__Q), .o(TIMEBOOST_net_14434) );
na02s01 TIMEBOOST_cell_15875 ( .a(TIMEBOOST_net_3194), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_412), .o(TIMEBOOST_net_72) );
in01s01 g62690_u0 ( .a(FE_OFN1243_n_4092), .o(g62690_sb) );
no02m02 TIMEBOOST_cell_3209 ( .a(TIMEBOOST_net_184), .b(FE_OCPN1841_n_16089), .o(n_3160) );
na02s02 TIMEBOOST_cell_36581 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_64), .b(pci_target_unit_pcit_if_strd_addr_in_700), .o(TIMEBOOST_net_10529) );
na02s01 TIMEBOOST_cell_3210 ( .a(n_16151), .b(pci_target_unit_wishbone_master_first_wb_data_access), .o(TIMEBOOST_net_185) );
in01s01 g62691_u0 ( .a(FE_OFN1241_n_4092), .o(g62691_sb) );
na02s01 TIMEBOOST_cell_36529 ( .a(pci_target_unit_fifos_pcir_data_in_188), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__Q), .o(TIMEBOOST_net_10503) );
na02s01 TIMEBOOST_cell_2899 ( .a(TIMEBOOST_net_29), .b(n_1968), .o(n_1353) );
na02s08 TIMEBOOST_cell_2900 ( .a(conf_wb_err_addr_in_953), .b(conf_wb_err_addr_in_950), .o(TIMEBOOST_net_30) );
oa12s01 g62692_u0 ( .a(pci_target_unit_pcit_if_comp_flush_in), .b(FE_OFN781_n_2746), .c(n_15397), .o(n_4667) );
in01s01 g62693_u0 ( .a(FE_OFN1270_n_4095), .o(g62693_sb) );
na02s01 TIMEBOOST_cell_36499 ( .a(pci_target_unit_del_sync_addr_in_232), .b(g66422_db), .o(TIMEBOOST_net_10488) );
na03m02 TIMEBOOST_cell_33049 ( .a(TIMEBOOST_net_781), .b(n_4086), .c(n_15762), .o(n_4792) );
na03s04 TIMEBOOST_cell_33048 ( .a(FE_OFN1611_n_2122), .b(wishbone_slave_unit_pcim_sm_data_in_658), .c(FE_RN_580_0), .o(FE_RN_581_0) );
in01s01 g62695_u0 ( .a(n_15788), .o(n_4666) );
in01s01 g62697_u0 ( .a(FE_OFN1232_n_6391), .o(g62697_sb) );
na02s01 TIMEBOOST_cell_36329 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__Q), .b(g65810_sb), .o(TIMEBOOST_net_10403) );
na02f02 TIMEBOOST_cell_3513 ( .a(TIMEBOOST_net_336), .b(n_3236), .o(n_4808) );
na02s01 TIMEBOOST_cell_38380 ( .a(TIMEBOOST_net_11428), .b(g59380_sb), .o(n_7679) );
in01s01 g62698_u0 ( .a(FE_OFN1270_n_4095), .o(g62698_sb) );
na02s01 TIMEBOOST_cell_36493 ( .a(n_2507), .b(g66421_db), .o(TIMEBOOST_net_10485) );
na03s02 TIMEBOOST_cell_42003 ( .a(n_4343), .b(n_4344), .c(FE_OFN1270_n_4095), .o(TIMEBOOST_net_13240) );
na02s01 TIMEBOOST_cell_42004 ( .a(TIMEBOOST_net_13240), .b(g62671_sb), .o(n_6196) );
no02m02 g62699_u0 ( .a(n_2429), .b(conf_wb_err_addr_in_965), .o(g62699_p) );
ao12m02 g62699_u1 ( .a(g62699_p), .b(conf_wb_err_addr_in_965), .c(n_2429), .o(n_3154) );
oa12m02 g62700_u0 ( .a(n_3325), .b(n_3324), .c(wbm_adr_o_27_), .o(n_4160) );
in01s01 g62701_u0 ( .a(FE_OFN1234_n_6391), .o(g62701_sb) );
na02s01 TIMEBOOST_cell_36351 ( .a(pci_target_unit_del_sync_bc_in_203), .b(g66413_db), .o(TIMEBOOST_net_10414) );
na02s01 TIMEBOOST_cell_38382 ( .a(TIMEBOOST_net_11429), .b(g62730_sb), .o(n_5519) );
na02s02 TIMEBOOST_cell_37163 ( .a(n_808), .b(n_1009), .o(TIMEBOOST_net_10820) );
oa12s02 g62702_u0 ( .a(n_3446), .b(n_1098), .c(n_4662), .o(n_4664) );
oa12s01 g62703_u0 ( .a(n_3444), .b(n_1658), .c(n_4662), .o(n_4663) );
oa12s02 g62704_u0 ( .a(n_3445), .b(n_1688), .c(n_4662), .o(n_4661) );
oa12s02 g62705_u0 ( .a(n_3443), .b(n_2262), .c(n_4662), .o(n_4660) );
in01s01 g62706_u0 ( .a(FE_OFN1268_n_4095), .o(g62706_sb) );
na02s01 TIMEBOOST_cell_36495 ( .a(TIMEBOOST_net_1202), .b(FE_OFN989_n_574), .o(TIMEBOOST_net_10486) );
na03s01 TIMEBOOST_cell_34796 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__Q), .b(g62326_sb), .c(g62326_db), .o(n_6937) );
na02s01 TIMEBOOST_cell_16632 ( .a(pci_target_unit_fifos_pciw_addr_data_in_144), .b(g64118_sb), .o(TIMEBOOST_net_3573) );
in01s01 g62707_u0 ( .a(FE_OFN1250_n_4093), .o(g62707_sb) );
na02m01 TIMEBOOST_cell_3211 ( .a(TIMEBOOST_net_185), .b(n_4874), .o(n_3267) );
na02s01 TIMEBOOST_cell_18311 ( .a(n_4758), .b(TIMEBOOST_net_4412), .o(n_7149) );
na02s01 TIMEBOOST_cell_15874 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_99), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3194) );
oa12m01 g62708_u0 ( .a(n_2019), .b(n_2018), .c(pci_target_unit_wishbone_master_rty_counter_7_), .o(n_2451) );
oa12s02 g62709_u0 ( .a(n_2949), .b(n_2948), .c(wbm_adr_o_24_), .o(n_3331) );
in01s01 g62710_u0 ( .a(FE_OFN1244_n_4092), .o(g62710_sb) );
na02s01 TIMEBOOST_cell_17261 ( .a(TIMEBOOST_net_3887), .b(g58422_sb), .o(n_9425) );
na02s01 TIMEBOOST_cell_16633 ( .a(TIMEBOOST_net_3573), .b(g64118_db), .o(n_4042) );
na02s02 TIMEBOOST_cell_45190 ( .a(TIMEBOOST_net_14833), .b(FE_OFN1261_n_4143), .o(TIMEBOOST_net_12641) );
in01s01 g62711_u0 ( .a(FE_OFN1241_n_4092), .o(g62711_sb) );
na02s01 TIMEBOOST_cell_36583 ( .a(wbs_sel_i_3_), .b(g63587_db), .o(TIMEBOOST_net_10530) );
na02s02 TIMEBOOST_cell_39904 ( .a(TIMEBOOST_net_12190), .b(g62921_sb), .o(n_6039) );
in01s01 g62712_u0 ( .a(FE_OFN1206_n_6356), .o(g62712_sb) );
na02m02 TIMEBOOST_cell_44019 ( .a(n_9543), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__Q), .o(TIMEBOOST_net_14248) );
na02s02 TIMEBOOST_cell_39166 ( .a(TIMEBOOST_net_11821), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_9855) );
na02s01 TIMEBOOST_cell_3214 ( .a(g65733_db), .b(g61705_sb), .o(TIMEBOOST_net_187) );
in01s01 g62713_u0 ( .a(FE_OFN1246_n_4093), .o(g62713_sb) );
na02s01 TIMEBOOST_cell_36585 ( .a(wbs_sel_i_2_), .b(g63586_db), .o(TIMEBOOST_net_10531) );
na02s01 TIMEBOOST_cell_44866 ( .a(TIMEBOOST_net_14671), .b(g65399_sb), .o(TIMEBOOST_net_11870) );
in01s01 g62714_u0 ( .a(FE_OFN1288_n_4098), .o(g62714_sb) );
na02s01 TIMEBOOST_cell_36587 ( .a(wbs_sel_i_0_), .b(g63584_db), .o(TIMEBOOST_net_10532) );
na02f02 TIMEBOOST_cell_44697 ( .a(n_969), .b(n_14971), .o(TIMEBOOST_net_14587) );
na02m02 TIMEBOOST_cell_41634 ( .a(FE_OFN1439_n_9372), .b(TIMEBOOST_net_13055), .o(TIMEBOOST_net_11674) );
in01s01 g62715_u0 ( .a(FE_OFN1207_n_6356), .o(g62715_sb) );
na02s01 TIMEBOOST_cell_36589 ( .a(wbs_sel_i_1_), .b(g63585_db), .o(TIMEBOOST_net_10533) );
na03s02 TIMEBOOST_cell_2697 ( .a(n_4610), .b(g61840_sb), .c(g61840_db), .o(n_6971) );
na02f02 TIMEBOOST_cell_42516 ( .a(TIMEBOOST_net_13496), .b(g57144_sb), .o(n_10464) );
in01s01 g62716_u0 ( .a(n_4662), .o(g62716_sb) );
na03f02 TIMEBOOST_cell_34460 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_388), .b(g54197_sb), .c(TIMEBOOST_net_569), .o(n_13421) );
na02m02 TIMEBOOST_cell_38884 ( .a(TIMEBOOST_net_11680), .b(g58471_sb), .o(n_9374) );
na02s02 TIMEBOOST_cell_3313 ( .a(TIMEBOOST_net_236), .b(n_4470), .o(n_4376) );
ao12s02 g62717_u0 ( .a(n_3326), .b(conf_wb_err_addr_in_945), .c(FE_OFN1142_n_15261), .o(n_4158) );
ao12s02 g62718_u0 ( .a(n_3323), .b(conf_wb_err_addr_in_948), .c(FE_OFN1142_n_15261), .o(n_4157) );
in01s01 g62719_u0 ( .a(FE_OFN1192_n_6935), .o(g62719_sb) );
na02s02 TIMEBOOST_cell_31404 ( .a(n_4482), .b(g65040_sb), .o(TIMEBOOST_net_9613) );
na02s01 g62719_u2 ( .a(n_6136), .b(FE_OFN1192_n_6935), .o(g62719_db) );
na02s01 TIMEBOOST_cell_3216 ( .a(g65780_db), .b(g61705_sb), .o(TIMEBOOST_net_188) );
in01s01 g62720_u0 ( .a(FE_OFN881_g64577_p), .o(g62720_sb) );
na02f02 TIMEBOOST_cell_37056 ( .a(FE_OFN1593_n_13741), .b(TIMEBOOST_net_10766), .o(g53263_p) );
na02f02 TIMEBOOST_cell_36974 ( .a(TIMEBOOST_net_10725), .b(g58828_sb), .o(n_8611) );
na02m02 TIMEBOOST_cell_36808 ( .a(TIMEBOOST_net_10642), .b(n_4154), .o(n_13556) );
in01s01 g62721_u0 ( .a(FE_OFN1130_g64577_p), .o(g62721_sb) );
na02m02 TIMEBOOST_cell_32638 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__14__Q), .o(TIMEBOOST_net_10230) );
na02f02 TIMEBOOST_cell_39010 ( .a(TIMEBOOST_net_11743), .b(g52519_sb), .o(n_13740) );
na02f02 TIMEBOOST_cell_41280 ( .a(TIMEBOOST_net_12878), .b(g57267_sb), .o(n_11485) );
in01s01 g62722_u0 ( .a(FE_OFN2105_g64577_p), .o(g62722_sb) );
na02s01 TIMEBOOST_cell_18309 ( .a(n_4760), .b(TIMEBOOST_net_4411), .o(n_7159) );
na02s01 TIMEBOOST_cell_37441 ( .a(TIMEBOOST_net_3453), .b(g52647_sb), .o(TIMEBOOST_net_10959) );
na02m02 TIMEBOOST_cell_39478 ( .a(TIMEBOOST_net_1724), .b(TIMEBOOST_net_11977), .o(n_13666) );
in01s01 g62723_u0 ( .a(FE_OFN1132_g64577_p), .o(g62723_sb) );
na02m02 TIMEBOOST_cell_32636 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__Q), .o(TIMEBOOST_net_10229) );
na02s02 TIMEBOOST_cell_39339 ( .a(TIMEBOOST_net_9543), .b(FE_OFN948_n_2248), .o(TIMEBOOST_net_11908) );
na02f02 TIMEBOOST_cell_41282 ( .a(TIMEBOOST_net_12879), .b(g57251_sb), .o(n_11505) );
na02s02 TIMEBOOST_cell_39462 ( .a(TIMEBOOST_net_11969), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_4545) );
na02s01 g62724_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q), .b(FE_OFN1106_g64577_p), .o(g62724_db) );
na02s01 TIMEBOOST_cell_37604 ( .a(TIMEBOOST_net_11040), .b(g61802_sb), .o(n_8191) );
in01s01 g62725_u0 ( .a(FE_OFN2106_g64577_p), .o(g62725_sb) );
na02s01 TIMEBOOST_cell_18297 ( .a(n_4748), .b(TIMEBOOST_net_4405), .o(n_7139) );
no02s02 TIMEBOOST_cell_37168 ( .a(TIMEBOOST_net_10822), .b(g64630_BP), .o(g64630_p) );
na02s01 TIMEBOOST_cell_45589 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q), .b(g63568_sb), .o(TIMEBOOST_net_15033) );
in01s01 g62726_u0 ( .a(FE_OFN877_g64577_p), .o(g62726_sb) );
na02m02 TIMEBOOST_cell_32634 ( .a(n_384), .b(n_255), .o(TIMEBOOST_net_10228) );
in01s01 TIMEBOOST_cell_45918 ( .a(TIMEBOOST_net_15224), .o(TIMEBOOST_net_15225) );
na02f02 TIMEBOOST_cell_41284 ( .a(TIMEBOOST_net_12880), .b(g57145_sb), .o(n_11605) );
in01s01 g62727_u0 ( .a(FE_OFN1118_g64577_p), .o(g62727_sb) );
na02m02 TIMEBOOST_cell_32632 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__Q), .o(TIMEBOOST_net_10227) );
na02s02 TIMEBOOST_cell_39906 ( .a(TIMEBOOST_net_12191), .b(g63177_sb), .o(n_5794) );
na02m02 TIMEBOOST_cell_45478 ( .a(TIMEBOOST_net_14977), .b(n_4889), .o(n_14816) );
in01s01 g62728_u0 ( .a(FE_OFN1129_g64577_p), .o(g62728_sb) );
na03s02 TIMEBOOST_cell_37543 ( .a(TIMEBOOST_net_3808), .b(g65702_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__Q), .o(TIMEBOOST_net_11010) );
na02s02 TIMEBOOST_cell_38384 ( .a(TIMEBOOST_net_11430), .b(g63559_sb), .o(n_4115) );
na02f02 TIMEBOOST_cell_44298 ( .a(TIMEBOOST_net_14387), .b(FE_OFN1414_n_8567), .o(n_11592) );
in01s01 g62729_u0 ( .a(FE_OFN1106_g64577_p), .o(g62729_sb) );
na02s02 TIMEBOOST_cell_36786 ( .a(TIMEBOOST_net_10631), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_4601) );
na02s02 TIMEBOOST_cell_43625 ( .a(n_65), .b(n_3667), .o(TIMEBOOST_net_14051) );
na02s01 TIMEBOOST_cell_36788 ( .a(TIMEBOOST_net_10632), .b(g62851_sb), .o(n_5267) );
in01s01 g62730_u0 ( .a(FE_OFN1115_g64577_p), .o(g62730_sb) );
na02f02 TIMEBOOST_cell_41230 ( .a(TIMEBOOST_net_12853), .b(g57193_sb), .o(n_11560) );
na02s02 TIMEBOOST_cell_39908 ( .a(TIMEBOOST_net_12192), .b(g62409_sb), .o(n_6781) );
na02f02 TIMEBOOST_cell_41248 ( .a(TIMEBOOST_net_12862), .b(g57301_sb), .o(n_11449) );
in01s01 g62731_u0 ( .a(FE_OFN1120_g64577_p), .o(g62731_sb) );
na03f02 TIMEBOOST_cell_21820 ( .a(n_3054), .b(n_2924), .c(n_2868), .o(TIMEBOOST_net_6167) );
na02s01 TIMEBOOST_cell_37752 ( .a(TIMEBOOST_net_11114), .b(TIMEBOOST_net_288), .o(TIMEBOOST_net_10051) );
na02s02 TIMEBOOST_cell_37754 ( .a(TIMEBOOST_net_11115), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_10600) );
in01s01 g62732_u0 ( .a(FE_OFN1118_g64577_p), .o(g62732_sb) );
na02m02 TIMEBOOST_cell_32628 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__Q), .o(TIMEBOOST_net_10225) );
na02s02 TIMEBOOST_cell_39910 ( .a(TIMEBOOST_net_12193), .b(g62924_sb), .o(n_6033) );
na02f02 TIMEBOOST_cell_41250 ( .a(TIMEBOOST_net_12863), .b(g57168_sb), .o(n_10457) );
in01s01 g62733_u0 ( .a(FE_OFN1125_g64577_p), .o(g62733_sb) );
na02m02 TIMEBOOST_cell_32626 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__Q), .o(TIMEBOOST_net_10224) );
na02f02 TIMEBOOST_cell_44020 ( .a(TIMEBOOST_net_14248), .b(FE_OFN1404_n_8567), .o(TIMEBOOST_net_13374) );
na02f02 TIMEBOOST_cell_41252 ( .a(TIMEBOOST_net_12864), .b(g57409_sb), .o(n_11334) );
in01s01 g62734_u0 ( .a(FE_OFN881_g64577_p), .o(g62734_sb) );
na02s02 TIMEBOOST_cell_38386 ( .a(TIMEBOOST_net_11431), .b(g62728_sb), .o(n_5523) );
na02s01 g62734_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__Q), .b(FE_OFN881_g64577_p), .o(g62734_db) );
na02s01 TIMEBOOST_cell_39368 ( .a(TIMEBOOST_net_11922), .b(g65882_sb), .o(n_1864) );
in01s01 g62735_u0 ( .a(FE_OFN1137_g64577_p), .o(g62735_sb) );
na02m02 TIMEBOOST_cell_32624 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__Q), .o(TIMEBOOST_net_10223) );
na03s02 TIMEBOOST_cell_38349 ( .a(n_1293), .b(FE_OFN1117_g64577_p), .c(n_2247), .o(TIMEBOOST_net_11413) );
na02f02 TIMEBOOST_cell_41254 ( .a(TIMEBOOST_net_12865), .b(g57327_sb), .o(n_11423) );
in01s01 g62736_u0 ( .a(FE_OFN1132_g64577_p), .o(g62736_sb) );
na02f02 TIMEBOOST_cell_21821 ( .a(TIMEBOOST_net_6167), .b(n_2867), .o(n_4171) );
na03s02 TIMEBOOST_cell_38211 ( .a(TIMEBOOST_net_4007), .b(g64134_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__Q), .o(TIMEBOOST_net_11344) );
na02m02 TIMEBOOST_cell_32622 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__18__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__18__Q), .o(TIMEBOOST_net_10222) );
in01s01 g62737_u0 ( .a(FE_OFN1125_g64577_p), .o(g62737_sb) );
na02f02 TIMEBOOST_cell_43760 ( .a(TIMEBOOST_net_14118), .b(FE_OFN1412_n_8567), .o(TIMEBOOST_net_12947) );
na02s02 TIMEBOOST_cell_39912 ( .a(TIMEBOOST_net_12194), .b(g62625_sb), .o(n_6305) );
na02f02 TIMEBOOST_cell_22347 ( .a(TIMEBOOST_net_6430), .b(n_10054), .o(n_12146) );
in01s01 g62738_u0 ( .a(FE_OFN1097_g64577_p), .o(g62738_sb) );
na02s01 TIMEBOOST_cell_36467 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(g65787_sb), .o(TIMEBOOST_net_10472) );
na02s01 g62738_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__Q), .b(FE_OFN1097_g64577_p), .o(g62738_db) );
na02s01 TIMEBOOST_cell_36450 ( .a(TIMEBOOST_net_10463), .b(g58093_sb), .o(TIMEBOOST_net_9593) );
in01s01 g62739_u0 ( .a(FE_OFN1120_g64577_p), .o(g62739_sb) );
na03s02 TIMEBOOST_cell_37523 ( .a(TIMEBOOST_net_3788), .b(g65966_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__Q), .o(TIMEBOOST_net_11000) );
na02s02 TIMEBOOST_cell_10318 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_62), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_1726) );
na02s01 TIMEBOOST_cell_17399 ( .a(TIMEBOOST_net_3956), .b(g64259_db), .o(n_3914) );
in01s01 g62740_u0 ( .a(FE_OFN1112_g64577_p), .o(g62740_sb) );
na02s01 TIMEBOOST_cell_42705 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__Q), .b(g65910_sb), .o(TIMEBOOST_net_13591) );
na02s02 TIMEBOOST_cell_39914 ( .a(TIMEBOOST_net_12195), .b(g62441_sb), .o(n_6714) );
na02s01 TIMEBOOST_cell_42773 ( .a(FE_OFN213_n_9124), .b(g58174_sb), .o(TIMEBOOST_net_13625) );
in01s01 g62741_u0 ( .a(FE_OFN1116_g64577_p), .o(g62741_sb) );
na02s01 TIMEBOOST_cell_36334 ( .a(TIMEBOOST_net_10405), .b(g67040_sb), .o(n_1277) );
na02s01 TIMEBOOST_cell_39916 ( .a(TIMEBOOST_net_12196), .b(g62382_sb), .o(n_6837) );
na02s01 TIMEBOOST_cell_36336 ( .a(TIMEBOOST_net_10406), .b(g67040_sb), .o(n_1704) );
in01s01 g62742_u0 ( .a(FE_OFN2105_g64577_p), .o(g62742_sb) );
na03s02 TIMEBOOST_cell_37541 ( .a(TIMEBOOST_net_3790), .b(g65720_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__Q), .o(TIMEBOOST_net_11009) );
na02s02 TIMEBOOST_cell_37756 ( .a(TIMEBOOST_net_11116), .b(FE_OFN2022_n_4778), .o(TIMEBOOST_net_10606) );
na02f02 TIMEBOOST_cell_44609 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__Q), .b(n_9670), .o(TIMEBOOST_net_14543) );
in01s01 g62743_u0 ( .a(FE_OFN1119_g64577_p), .o(g62743_sb) );
na02s01 TIMEBOOST_cell_37521 ( .a(n_3755), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__Q), .o(TIMEBOOST_net_10999) );
na03s01 TIMEBOOST_cell_36803 ( .a(g64120_da), .b(g64120_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__Q), .o(TIMEBOOST_net_10640) );
na02s02 TIMEBOOST_cell_37758 ( .a(TIMEBOOST_net_11117), .b(FE_OFN2022_n_4778), .o(TIMEBOOST_net_10604) );
in01s01 g62744_u0 ( .a(FE_OFN1127_g64577_p), .o(g62744_sb) );
na02s01 TIMEBOOST_cell_36338 ( .a(TIMEBOOST_net_10407), .b(g67040_sb), .o(n_1502) );
na02s01 TIMEBOOST_cell_39331 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__12__Q), .b(g64229_sb), .o(TIMEBOOST_net_11904) );
na02m02 TIMEBOOST_cell_45479 ( .a(TIMEBOOST_net_4823), .b(g62068_sb), .o(TIMEBOOST_net_14978) );
in01s01 g62745_u0 ( .a(FE_OFN1118_g64577_p), .o(g62745_sb) );
na02s01 TIMEBOOST_cell_38388 ( .a(TIMEBOOST_net_11432), .b(g62787_sb), .o(n_5416) );
na02m02 TIMEBOOST_cell_38752 ( .a(TIMEBOOST_net_11614), .b(g53930_sb), .o(n_13515) );
na02s01 TIMEBOOST_cell_39356 ( .a(TIMEBOOST_net_11916), .b(g61871_sb), .o(n_8092) );
in01s01 g62746_u0 ( .a(FE_OFN1094_g64577_p), .o(g62746_sb) );
na02f02 TIMEBOOST_cell_42482 ( .a(TIMEBOOST_net_13479), .b(g57076_sb), .o(n_11667) );
na02s02 TIMEBOOST_cell_39918 ( .a(TIMEBOOST_net_12197), .b(g63042_sb), .o(n_5858) );
na02s02 TIMEBOOST_cell_39920 ( .a(TIMEBOOST_net_12198), .b(g62400_sb), .o(n_6799) );
in01s01 g62747_u0 ( .a(FE_OFN1139_g64577_p), .o(g62747_sb) );
na02m02 TIMEBOOST_cell_45480 ( .a(TIMEBOOST_net_14978), .b(TIMEBOOST_net_5527), .o(n_14811) );
na02s01 TIMEBOOST_cell_38390 ( .a(TIMEBOOST_net_11433), .b(g62793_sb), .o(n_5402) );
na02s01 TIMEBOOST_cell_30868 ( .a(pci_target_unit_pcit_if_strd_addr_in_686), .b(n_2598), .o(TIMEBOOST_net_9345) );
in01s01 g62748_u0 ( .a(FE_OFN1139_g64577_p), .o(g62748_sb) );
na02s01 TIMEBOOST_cell_36452 ( .a(TIMEBOOST_net_10464), .b(g64138_db), .o(n_4737) );
na02s02 TIMEBOOST_cell_39922 ( .a(TIMEBOOST_net_12199), .b(g62511_sb), .o(n_6556) );
na02f02 TIMEBOOST_cell_12667 ( .a(FE_OFN1586_n_13736), .b(TIMEBOOST_net_2900), .o(n_14430) );
in01s01 g62749_u0 ( .a(FE_OFN1125_g64577_p), .o(g62749_sb) );
na02m02 TIMEBOOST_cell_44021 ( .a(n_9859), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__Q), .o(TIMEBOOST_net_14249) );
na02s01 TIMEBOOST_cell_38392 ( .a(TIMEBOOST_net_11434), .b(g63139_sb), .o(n_4970) );
na02f02 TIMEBOOST_cell_44525 ( .a(n_9081), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__Q), .o(TIMEBOOST_net_14501) );
in01s01 g62750_u0 ( .a(FE_OFN1133_g64577_p), .o(g62750_sb) );
na02f02 TIMEBOOST_cell_44526 ( .a(TIMEBOOST_net_14501), .b(FE_OFN2167_n_8567), .o(TIMEBOOST_net_13457) );
na02s02 TIMEBOOST_cell_39924 ( .a(TIMEBOOST_net_12200), .b(g62938_sb), .o(n_6005) );
na02f02 TIMEBOOST_cell_44022 ( .a(TIMEBOOST_net_14249), .b(FE_OFN1415_n_8567), .o(TIMEBOOST_net_12840) );
in01s01 g62751_u0 ( .a(FE_OFN1124_g64577_p), .o(g62751_sb) );
na02m02 TIMEBOOST_cell_44023 ( .a(n_9619), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__Q), .o(TIMEBOOST_net_14250) );
na02s01 TIMEBOOST_cell_38754 ( .a(TIMEBOOST_net_11615), .b(g53919_sb), .o(n_13627) );
na02f02 TIMEBOOST_cell_12679 ( .a(TIMEBOOST_net_2906), .b(n_14035), .o(n_14252) );
in01s01 g62752_u0 ( .a(FE_OFN1120_g64577_p), .o(g62752_sb) );
na02s01 TIMEBOOST_cell_37519 ( .a(TIMEBOOST_net_9549), .b(FE_OFN1051_n_16657), .o(TIMEBOOST_net_10998) );
na02s01 TIMEBOOST_cell_38058 ( .a(TIMEBOOST_net_11267), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_4679) );
na02s02 TIMEBOOST_cell_37760 ( .a(TIMEBOOST_net_11118), .b(FE_OFN2022_n_4778), .o(TIMEBOOST_net_10603) );
in01s01 g62753_u0 ( .a(FE_OFN1119_g64577_p), .o(g62753_sb) );
na02s01 TIMEBOOST_cell_37517 ( .a(TIMEBOOST_net_9537), .b(FE_OFN1056_n_4727), .o(TIMEBOOST_net_10997) );
na02s02 TIMEBOOST_cell_38060 ( .a(TIMEBOOST_net_11268), .b(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_4573) );
na02s02 TIMEBOOST_cell_37762 ( .a(TIMEBOOST_net_11119), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_10593) );
in01s01 g62754_u0 ( .a(FE_OFN1265_n_4095), .o(g62754_sb) );
na02s01 TIMEBOOST_cell_36591 ( .a(wbs_adr_i_0_), .b(g63582_sb), .o(TIMEBOOST_net_10534) );
na02f02 TIMEBOOST_cell_39012 ( .a(TIMEBOOST_net_11744), .b(g52506_sb), .o(n_13724) );
na02f02 TIMEBOOST_cell_44024 ( .a(TIMEBOOST_net_14250), .b(FE_OFN1425_n_8567), .o(TIMEBOOST_net_12703) );
in01s01 g62755_u0 ( .a(FE_OFN1233_n_6391), .o(g62755_sb) );
na02s01 TIMEBOOST_cell_36327 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__Q), .b(g65861_sb), .o(TIMEBOOST_net_10402) );
na02m02 TIMEBOOST_cell_39157 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__Q), .b(n_13447), .o(TIMEBOOST_net_11817) );
na02f02 TIMEBOOST_cell_39014 ( .a(TIMEBOOST_net_11745), .b(g52534_sb), .o(n_13685) );
in01s01 g62756_u0 ( .a(FE_OFN1128_g64577_p), .o(g62756_sb) );
na03s01 TIMEBOOST_cell_33759 ( .a(FE_OFN215_n_9856), .b(g58045_sb), .c(g58045_db), .o(n_9745) );
na02s02 TIMEBOOST_cell_38394 ( .a(TIMEBOOST_net_11435), .b(g62785_sb), .o(n_5421) );
na02f02 TIMEBOOST_cell_44752 ( .a(TIMEBOOST_net_14614), .b(n_11973), .o(n_12507) );
in01s01 g62757_u0 ( .a(FE_OFN1092_g64577_p), .o(g62757_sb) );
na02s01 TIMEBOOST_cell_36870 ( .a(TIMEBOOST_net_10673), .b(g61796_db), .o(n_8205) );
na03s02 TIMEBOOST_cell_38239 ( .a(g64321_da), .b(g64321_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__Q), .o(TIMEBOOST_net_11358) );
na02s01 TIMEBOOST_cell_36872 ( .a(TIMEBOOST_net_10674), .b(g61779_db), .o(n_8248) );
in01s01 g62758_u0 ( .a(FE_OFN1320_n_6436), .o(g62758_sb) );
na02m02 TIMEBOOST_cell_44025 ( .a(n_9833), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__Q), .o(TIMEBOOST_net_14251) );
na02f04 TIMEBOOST_cell_3807 ( .a(TIMEBOOST_net_483), .b(n_3202), .o(n_3193) );
na02s02 TIMEBOOST_cell_45481 ( .a(n_13145), .b(pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_77), .o(TIMEBOOST_net_14979) );
in01s01 g62759_u0 ( .a(FE_OFN1116_g64577_p), .o(g62759_sb) );
na02s01 TIMEBOOST_cell_41788 ( .a(TIMEBOOST_net_13132), .b(g58267_db), .o(n_9037) );
na02f02 TIMEBOOST_cell_39016 ( .a(TIMEBOOST_net_11746), .b(g52504_sb), .o(n_13727) );
na03f06 TIMEBOOST_cell_45845 ( .a(n_11136), .b(n_11139), .c(n_11137), .o(TIMEBOOST_net_15161) );
in01s01 g62760_u0 ( .a(FE_OFN1252_n_4143), .o(g62760_sb) );
no03f04 TIMEBOOST_cell_36593 ( .a(n_2227), .b(n_1399), .c(FE_RN_150_0), .o(TIMEBOOST_net_10535) );
na03s02 TIMEBOOST_cell_2701 ( .a(n_4593), .b(g61961_sb), .c(g61961_db), .o(n_6951) );
na02s02 TIMEBOOST_cell_18847 ( .a(TIMEBOOST_net_4680), .b(g63135_sb), .o(n_4980) );
in01s01 g62761_u0 ( .a(FE_OFN1265_n_4095), .o(g62761_sb) );
na02s01 TIMEBOOST_cell_36595 ( .a(wbs_adr_i_1_), .b(g52466_sb), .o(TIMEBOOST_net_10536) );
na02s01 TIMEBOOST_cell_18901 ( .a(TIMEBOOST_net_4707), .b(g63123_sb), .o(n_5009) );
na02s01 TIMEBOOST_cell_18605 ( .a(TIMEBOOST_net_4559), .b(g62831_sb), .o(n_5313) );
in01s01 g62762_u0 ( .a(FE_OFN1121_g64577_p), .o(g62762_sb) );
na03f04 TIMEBOOST_cell_44753 ( .a(n_11841), .b(n_16404), .c(FE_RN_909_0), .o(TIMEBOOST_net_14615) );
na03s02 TIMEBOOST_cell_34254 ( .a(TIMEBOOST_net_9792), .b(FE_OFN1171_n_5592), .c(g62112_sb), .o(n_5585) );
na02s01 TIMEBOOST_cell_45679 ( .a(n_4365), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q), .o(TIMEBOOST_net_15078) );
in01s01 g62763_u0 ( .a(n_6554), .o(g62763_sb) );
na02s01 TIMEBOOST_cell_36353 ( .a(TIMEBOOST_net_3222), .b(n_8953), .o(TIMEBOOST_net_10415) );
na02f08 TIMEBOOST_cell_3399 ( .a(n_2777), .b(TIMEBOOST_net_279), .o(n_3278) );
na02f04 TIMEBOOST_cell_3400 ( .a(n_2380), .b(FE_RN_83_0), .o(TIMEBOOST_net_280) );
in01s01 g62764_u0 ( .a(FE_OFN1130_g64577_p), .o(g62764_sb) );
na02f02 TIMEBOOST_cell_42484 ( .a(TIMEBOOST_net_13480), .b(g57345_sb), .o(n_10390) );
na02f02 TIMEBOOST_cell_44182 ( .a(TIMEBOOST_net_14329), .b(FE_OFN1377_n_8567), .o(TIMEBOOST_net_13399) );
na02f04 TIMEBOOST_cell_45846 ( .a(TIMEBOOST_net_15161), .b(n_11140), .o(n_12554) );
in01s01 g62765_u0 ( .a(FE_OFN1132_g64577_p), .o(g62765_sb) );
na03f06 TIMEBOOST_cell_45847 ( .a(n_17016), .b(n_11157), .c(n_17017), .o(TIMEBOOST_net_15162) );
na02s01 TIMEBOOST_cell_38396 ( .a(TIMEBOOST_net_11436), .b(g63431_sb), .o(n_4934) );
na02f04 TIMEBOOST_cell_45848 ( .a(TIMEBOOST_net_15162), .b(n_11144), .o(n_12558) );
in01s01 g62766_u0 ( .a(FE_OFN1130_g64577_p), .o(g62766_sb) );
na03f06 TIMEBOOST_cell_45849 ( .a(n_11129), .b(n_11126), .c(n_16582), .o(TIMEBOOST_net_15163) );
na03s02 TIMEBOOST_cell_38245 ( .a(TIMEBOOST_net_3996), .b(g64107_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__Q), .o(TIMEBOOST_net_11361) );
na02f04 TIMEBOOST_cell_45850 ( .a(TIMEBOOST_net_15163), .b(n_16581), .o(n_12552) );
in01s01 g62767_u0 ( .a(FE_OFN1119_g64577_p), .o(g62767_sb) );
na03f06 TIMEBOOST_cell_45851 ( .a(n_11790), .b(n_11107), .c(n_11106), .o(TIMEBOOST_net_15164) );
na03s02 TIMEBOOST_cell_38247 ( .a(TIMEBOOST_net_3985), .b(g64090_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__Q), .o(TIMEBOOST_net_11362) );
na02f04 TIMEBOOST_cell_45852 ( .a(TIMEBOOST_net_15164), .b(n_11104), .o(n_12547) );
in01s01 g62768_u0 ( .a(FE_OFN1136_g64577_p), .o(g62768_sb) );
na02m02 TIMEBOOST_cell_42119 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__Q), .b(n_4388), .o(TIMEBOOST_net_13298) );
na03s02 TIMEBOOST_cell_38249 ( .a(TIMEBOOST_net_4013), .b(g64208_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__Q), .o(TIMEBOOST_net_11363) );
na02m02 TIMEBOOST_cell_44151 ( .a(n_9463), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__Q), .o(TIMEBOOST_net_14314) );
in01s01 g62769_u0 ( .a(FE_OFN1137_g64577_p), .o(g62769_sb) );
na02f02 TIMEBOOST_cell_44026 ( .a(TIMEBOOST_net_14251), .b(FE_OFN1401_n_8567), .o(TIMEBOOST_net_12760) );
na02s01 TIMEBOOST_cell_39168 ( .a(TIMEBOOST_net_11822), .b(g65835_sb), .o(n_2150) );
na02f04 TIMEBOOST_cell_44754 ( .a(TIMEBOOST_net_14615), .b(FE_RN_910_0), .o(n_16406) );
in01s01 g62770_u0 ( .a(FE_OFN1135_g64577_p), .o(g62770_sb) );
na03s02 TIMEBOOST_cell_43029 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__Q), .b(FE_OFN1120_g64577_p), .c(g62731_sb), .o(TIMEBOOST_net_13753) );
na02s01 TIMEBOOST_cell_38398 ( .a(TIMEBOOST_net_11437), .b(g63040_sb), .o(n_5170) );
na02m02 TIMEBOOST_cell_44027 ( .a(n_9472), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__Q), .o(TIMEBOOST_net_14252) );
in01s01 g62771_u0 ( .a(FE_OFN1131_g64577_p), .o(g62771_sb) );
na02m02 TIMEBOOST_cell_44527 ( .a(n_9452), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__Q), .o(TIMEBOOST_net_14502) );
na03s02 TIMEBOOST_cell_38251 ( .a(TIMEBOOST_net_3992), .b(g64127_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__Q), .o(TIMEBOOST_net_11364) );
na02f02 TIMEBOOST_cell_44028 ( .a(TIMEBOOST_net_14252), .b(FE_OFN1408_n_8567), .o(TIMEBOOST_net_12894) );
in01s01 g62772_u0 ( .a(FE_OFN1116_g64577_p), .o(g62772_sb) );
na02m02 TIMEBOOST_cell_44029 ( .a(n_9786), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__Q), .o(TIMEBOOST_net_14253) );
na02s01 TIMEBOOST_cell_39926 ( .a(TIMEBOOST_net_12201), .b(g62434_sb), .o(n_6729) );
na02s01 TIMEBOOST_cell_43433 ( .a(n_1916), .b(g61746_sb), .o(TIMEBOOST_net_13955) );
in01s01 g62773_u0 ( .a(FE_OFN881_g64577_p), .o(g62773_sb) );
na02s01 TIMEBOOST_cell_36874 ( .a(TIMEBOOST_net_10675), .b(g61767_db), .o(n_8277) );
na02f02 TIMEBOOST_cell_36976 ( .a(TIMEBOOST_net_10726), .b(g58802_sb), .o(n_8640) );
na02s01 TIMEBOOST_cell_36876 ( .a(TIMEBOOST_net_10676), .b(g58297_db), .o(n_9216) );
in01s01 g62774_u0 ( .a(FE_OFN1120_g64577_p), .o(g62774_sb) );
na03f02 TIMEBOOST_cell_21822 ( .a(n_3048), .b(n_2917), .c(n_2860), .o(TIMEBOOST_net_6168) );
na02f02 TIMEBOOST_cell_37115 ( .a(FE_OFN1605_n_13997), .b(TIMEBOOST_net_10183), .o(TIMEBOOST_net_10796) );
na02s01 TIMEBOOST_cell_39298 ( .a(TIMEBOOST_net_11887), .b(g65953_sb), .o(n_2167) );
in01s01 g62775_u0 ( .a(FE_OFN1136_g64577_p), .o(g62775_sb) );
na02s02 TIMEBOOST_cell_37986 ( .a(TIMEBOOST_net_11231), .b(n_4064), .o(n_5275) );
na03s02 TIMEBOOST_cell_38313 ( .a(n_3898), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__16__Q), .c(FE_OFN2104_g64577_p), .o(TIMEBOOST_net_11395) );
na02f02 TIMEBOOST_cell_44030 ( .a(TIMEBOOST_net_14253), .b(FE_OFN1411_n_8567), .o(TIMEBOOST_net_12848) );
in01s01 g62776_u0 ( .a(FE_OFN1112_g64577_p), .o(g62776_sb) );
na02m02 TIMEBOOST_cell_44031 ( .a(n_9011), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__Q), .o(TIMEBOOST_net_14254) );
na03s02 TIMEBOOST_cell_38315 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__Q), .b(FE_OFN1128_g64577_p), .c(n_3510), .o(TIMEBOOST_net_11396) );
na02s01 TIMEBOOST_cell_45590 ( .a(TIMEBOOST_net_15033), .b(g63568_db), .o(n_4594) );
in01s01 g62777_u0 ( .a(FE_OFN1106_g64577_p), .o(g62777_sb) );
na02s02 TIMEBOOST_cell_10530 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_10__Q), .b(FE_OFN2072_n_15978), .o(TIMEBOOST_net_1832) );
na02s01 g62777_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q), .b(FE_OFN1106_g64577_p), .o(g62777_db) );
na02s02 TIMEBOOST_cell_10531 ( .a(TIMEBOOST_net_1832), .b(FE_OFN1084_n_13221), .o(TIMEBOOST_net_570) );
in01s01 g62778_u0 ( .a(FE_OFN882_g64577_p), .o(g62778_sb) );
na02f02 TIMEBOOST_cell_44032 ( .a(TIMEBOOST_net_14254), .b(FE_OFN1405_n_8567), .o(TIMEBOOST_net_12902) );
na03s02 TIMEBOOST_cell_38317 ( .a(n_4012), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__Q), .c(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_11397) );
na02m02 TIMEBOOST_cell_44033 ( .a(n_9607), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__Q), .o(TIMEBOOST_net_14255) );
in01s01 g62779_u0 ( .a(FE_OFN1115_g64577_p), .o(g62779_sb) );
na02f02 TIMEBOOST_cell_44034 ( .a(TIMEBOOST_net_14255), .b(FE_OFN1407_n_8567), .o(TIMEBOOST_net_12906) );
na02s01 TIMEBOOST_cell_38400 ( .a(TIMEBOOST_net_11438), .b(g63069_sb), .o(n_5112) );
na02s01 TIMEBOOST_cell_43434 ( .a(TIMEBOOST_net_13955), .b(g61746_db), .o(n_8325) );
in01s01 g62780_u0 ( .a(FE_OFN1100_g64577_p), .o(g62780_sb) );
no02f04 TIMEBOOST_cell_36878 ( .a(TIMEBOOST_net_10677), .b(FE_RN_130_0), .o(TIMEBOOST_net_6402) );
na02s01 g62780_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__14__Q), .b(FE_OFN1100_g64577_p), .o(g62780_db) );
na02m02 TIMEBOOST_cell_36880 ( .a(TIMEBOOST_net_10678), .b(g59808_sb), .o(n_7615) );
in01s01 g62781_u0 ( .a(FE_OFN1123_g64577_p), .o(g62781_sb) );
na02s02 TIMEBOOST_cell_43435 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__Q), .b(n_4328), .o(TIMEBOOST_net_13956) );
na02s02 TIMEBOOST_cell_38680 ( .a(TIMEBOOST_net_11578), .b(g62632_sb), .o(n_6289) );
na02f02 TIMEBOOST_cell_44035 ( .a(n_9064), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__Q), .o(TIMEBOOST_net_14256) );
in01s01 g62782_u0 ( .a(FE_OFN1130_g64577_p), .o(g62782_sb) );
na02f02 TIMEBOOST_cell_44036 ( .a(TIMEBOOST_net_14256), .b(FE_OFN1416_n_8567), .o(TIMEBOOST_net_12973) );
na02s02 TIMEBOOST_cell_38682 ( .a(TIMEBOOST_net_11579), .b(g62421_sb), .o(n_6754) );
na02s02 TIMEBOOST_cell_43436 ( .a(TIMEBOOST_net_13956), .b(FE_OFN1234_n_6391), .o(TIMEBOOST_net_12639) );
in01s01 g62783_u0 ( .a(FE_OFN1097_g64577_p), .o(g62783_sb) );
na02s02 TIMEBOOST_cell_36882 ( .a(TIMEBOOST_net_10679), .b(g61858_db), .o(n_8123) );
na02s01 g62783_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__Q), .b(FE_OFN1097_g64577_p), .o(g62783_db) );
na02s02 TIMEBOOST_cell_36884 ( .a(TIMEBOOST_net_10680), .b(g61859_db), .o(n_8121) );
in01s01 g62784_u0 ( .a(FE_OFN1124_g64577_p), .o(g62784_sb) );
na02m02 TIMEBOOST_cell_44037 ( .a(n_9447), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__Q), .o(TIMEBOOST_net_14257) );
in01s01 TIMEBOOST_cell_45930 ( .a(TIMEBOOST_net_15236), .o(TIMEBOOST_net_15237) );
na02f02 TIMEBOOST_cell_44038 ( .a(TIMEBOOST_net_14257), .b(FE_OFN1374_n_8567), .o(TIMEBOOST_net_12905) );
in01s01 g62785_u0 ( .a(FE_OFN1119_g64577_p), .o(g62785_sb) );
na02s02 TIMEBOOST_cell_37515 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__Q), .b(g64339_sb), .o(TIMEBOOST_net_10996) );
na02s02 TIMEBOOST_cell_37764 ( .a(TIMEBOOST_net_11120), .b(FE_OFN2021_n_4778), .o(TIMEBOOST_net_10595) );
na02s01 TIMEBOOST_cell_37684 ( .a(TIMEBOOST_net_11080), .b(g61700_sb), .o(n_8428) );
in01s01 g62786_u0 ( .a(FE_OFN1132_g64577_p), .o(g62786_sb) );
na02f02 TIMEBOOST_cell_44528 ( .a(TIMEBOOST_net_14502), .b(FE_OFN2188_n_8567), .o(TIMEBOOST_net_13021) );
na03s02 TIMEBOOST_cell_38321 ( .a(n_3903), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__12__Q), .c(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_11399) );
na02m02 TIMEBOOST_cell_44039 ( .a(n_9551), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q), .o(TIMEBOOST_net_14258) );
in01s01 g62787_u0 ( .a(FE_OFN1124_g64577_p), .o(g62787_sb) );
na02f02 TIMEBOOST_cell_44040 ( .a(TIMEBOOST_net_14258), .b(FE_OFN1411_n_8567), .o(TIMEBOOST_net_12904) );
na02s01 TIMEBOOST_cell_38402 ( .a(TIMEBOOST_net_11439), .b(g63078_sb), .o(n_5096) );
na02f02 TIMEBOOST_cell_44041 ( .a(n_9067), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__Q), .o(TIMEBOOST_net_14259) );
in01s01 g62788_u0 ( .a(FE_OFN1121_g64577_p), .o(g62788_sb) );
na02f02 TIMEBOOST_cell_44042 ( .a(TIMEBOOST_net_14259), .b(FE_OFN1380_n_8567), .o(TIMEBOOST_net_13378) );
na03s02 TIMEBOOST_cell_38323 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__Q), .b(FE_OFN1136_g64577_p), .c(n_3917), .o(TIMEBOOST_net_11400) );
na02m02 TIMEBOOST_cell_44043 ( .a(n_9592), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__Q), .o(TIMEBOOST_net_14260) );
in01s01 g62789_u0 ( .a(FE_OFN1094_g64577_p), .o(g62789_sb) );
na02s02 TIMEBOOST_cell_39928 ( .a(TIMEBOOST_net_12202), .b(g62697_sb), .o(n_6160) );
na02s01 TIMEBOOST_cell_43394 ( .a(TIMEBOOST_net_13935), .b(n_6319), .o(TIMEBOOST_net_11569) );
in01s01 g62790_u0 ( .a(FE_OFN1123_g64577_p), .o(g62790_sb) );
na02f02 TIMEBOOST_cell_44044 ( .a(TIMEBOOST_net_14260), .b(FE_OFN1390_n_8567), .o(TIMEBOOST_net_12811) );
na02s02 TIMEBOOST_cell_42975 ( .a(g52624_da), .b(g52402_sb), .o(TIMEBOOST_net_13726) );
na02m02 TIMEBOOST_cell_44045 ( .a(n_9719), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__Q), .o(TIMEBOOST_net_14261) );
in01s01 g62791_u0 ( .a(FE_OFN877_g64577_p), .o(g62791_sb) );
na02s02 TIMEBOOST_cell_43395 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__Q), .b(n_4656), .o(TIMEBOOST_net_13936) );
na02s01 g62791_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__Q), .b(FE_OFN1100_g64577_p), .o(g62791_db) );
na02f02 TIMEBOOST_cell_44046 ( .a(TIMEBOOST_net_14261), .b(FE_OFN1384_n_8567), .o(TIMEBOOST_net_13022) );
in01s01 g62792_u0 ( .a(FE_OFN1112_g64577_p), .o(g62792_sb) );
na02s01 g64752_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__Q), .b(FE_OFN678_n_4460), .o(g64752_db) );
in01s01 TIMEBOOST_cell_45919 ( .a(wbm_dat_i_19_), .o(TIMEBOOST_net_15226) );
na02m02 TIMEBOOST_cell_44047 ( .a(n_9724), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__Q), .o(TIMEBOOST_net_14262) );
in01s01 g62793_u0 ( .a(FE_OFN1123_g64577_p), .o(g62793_sb) );
na02s01 TIMEBOOST_cell_39170 ( .a(TIMEBOOST_net_11823), .b(g65863_sb), .o(n_1572) );
na02s02 TIMEBOOST_cell_39930 ( .a(TIMEBOOST_net_12203), .b(g62563_sb), .o(n_6433) );
na02f02 TIMEBOOST_cell_44048 ( .a(TIMEBOOST_net_14262), .b(FE_OFN1387_n_8567), .o(TIMEBOOST_net_12940) );
in01s01 g62794_u0 ( .a(FE_OFN1112_g64577_p), .o(g62794_sb) );
na02s01 TIMEBOOST_cell_38404 ( .a(TIMEBOOST_net_11440), .b(g62823_sb), .o(n_5332) );
na02m02 TIMEBOOST_cell_44309 ( .a(n_9088), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__Q), .o(TIMEBOOST_net_14393) );
na02f02 TIMEBOOST_cell_12787 ( .a(n_14056), .b(TIMEBOOST_net_2960), .o(n_16250) );
in01s01 g62795_u0 ( .a(FE_OFN1130_g64577_p), .o(g62795_sb) );
na02s01 TIMEBOOST_cell_37826 ( .a(TIMEBOOST_net_11151), .b(FE_OFN561_n_9895), .o(TIMEBOOST_net_9688) );
na02s02 TIMEBOOST_cell_39932 ( .a(TIMEBOOST_net_12204), .b(g62701_sb), .o(n_6156) );
na02s02 TIMEBOOST_cell_19255 ( .a(TIMEBOOST_net_4884), .b(g60608_sb), .o(n_4846) );
in01s01 g62796_u0 ( .a(FE_OFN1136_g64577_p), .o(g62796_sb) );
na02f02 TIMEBOOST_cell_12623 ( .a(TIMEBOOST_net_2878), .b(n_13901), .o(TIMEBOOST_net_939) );
na02s02 TIMEBOOST_cell_39934 ( .a(TIMEBOOST_net_12205), .b(g62755_sb), .o(n_6127) );
na02s01 TIMEBOOST_cell_39420 ( .a(TIMEBOOST_net_11948), .b(FE_OFN1166_n_5615), .o(TIMEBOOST_net_11372) );
in01s01 g62797_u0 ( .a(FE_OFN1132_g64577_p), .o(g62797_sb) );
na02m02 TIMEBOOST_cell_44049 ( .a(n_9479), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q), .o(TIMEBOOST_net_14263) );
na02f02 TIMEBOOST_cell_38795 ( .a(n_2926), .b(n_2859), .o(TIMEBOOST_net_11636) );
na02f02 TIMEBOOST_cell_12621 ( .a(TIMEBOOST_net_2877), .b(n_13901), .o(TIMEBOOST_net_937) );
na03f03 TIMEBOOST_cell_21818 ( .a(n_5230), .b(n_2797), .c(n_2820), .o(TIMEBOOST_net_6166) );
na02s02 TIMEBOOST_cell_39394 ( .a(TIMEBOOST_net_11935), .b(FE_OFN270_n_9836), .o(n_9488) );
na02s01 TIMEBOOST_cell_37592 ( .a(TIMEBOOST_net_11034), .b(g61811_sb), .o(n_8171) );
in01s01 g62799_u0 ( .a(FE_OFN1100_g64577_p), .o(g62799_sb) );
na03f02 TIMEBOOST_cell_36215 ( .a(FE_OCP_RBN1973_n_12381), .b(TIMEBOOST_net_10303), .c(FE_OFN1755_n_12681), .o(n_15935) );
na02s01 g62799_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q), .b(FE_OFN1100_g64577_p), .o(g62799_db) );
na02s01 TIMEBOOST_cell_36838 ( .a(TIMEBOOST_net_10657), .b(FE_OFN1207_n_6356), .o(TIMEBOOST_net_5194) );
in01s01 g62800_u0 ( .a(FE_OFN1115_g64577_p), .o(g62800_sb) );
na02s01 TIMEBOOST_cell_37256 ( .a(TIMEBOOST_net_10866), .b(FE_OFN682_n_4460), .o(TIMEBOOST_net_9384) );
na02s02 TIMEBOOST_cell_42976 ( .a(TIMEBOOST_net_13726), .b(TIMEBOOST_net_462), .o(TIMEBOOST_net_5432) );
na02s01 TIMEBOOST_cell_43635 ( .a(n_1575), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__Q), .o(TIMEBOOST_net_14056) );
in01s01 g62801_u0 ( .a(FE_OFN2104_g64577_p), .o(g62801_sb) );
na02s01 TIMEBOOST_cell_37513 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__Q), .b(g64237_sb), .o(TIMEBOOST_net_10995) );
na02s01 TIMEBOOST_cell_37680 ( .a(TIMEBOOST_net_11078), .b(g61954_sb), .o(n_7917) );
na02s01 TIMEBOOST_cell_37682 ( .a(TIMEBOOST_net_11079), .b(g62022_sb), .o(n_7853) );
in01s01 g62802_u0 ( .a(FE_OFN2105_g64577_p), .o(g62802_sb) );
na02m02 TIMEBOOST_cell_32502 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__12__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__12__Q), .o(TIMEBOOST_net_10162) );
na02s01 TIMEBOOST_cell_37624 ( .a(TIMEBOOST_net_11050), .b(g61795_sb), .o(n_8208) );
na02s01 TIMEBOOST_cell_37626 ( .a(TIMEBOOST_net_11051), .b(g61770_sb), .o(n_8269) );
in01s01 g62803_u0 ( .a(FE_OFN1134_g64577_p), .o(g62803_sb) );
na02s01 TIMEBOOST_cell_16813 ( .a(TIMEBOOST_net_3663), .b(g65313_db), .o(n_3567) );
na02s01 g62803_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q), .b(FE_OFN1104_g64577_p), .o(g62803_db) );
na02f02 TIMEBOOST_cell_40946 ( .a(TIMEBOOST_net_12711), .b(g57470_sb), .o(n_10819) );
na02s02 TIMEBOOST_cell_17823 ( .a(TIMEBOOST_net_4168), .b(g62005_sb), .o(n_7885) );
na03s02 TIMEBOOST_cell_1551 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__Q), .b(g62468_sb), .c(g62468_db), .o(n_6657) );
na02s01 TIMEBOOST_cell_37628 ( .a(TIMEBOOST_net_11052), .b(g61789_sb), .o(n_8223) );
in01s01 g62805_u0 ( .a(FE_OFN1100_g64577_p), .o(g62805_sb) );
na02m04 TIMEBOOST_cell_36832 ( .a(g52400_sb), .b(TIMEBOOST_net_10654), .o(TIMEBOOST_net_9992) );
na02f02 TIMEBOOST_cell_44198 ( .a(TIMEBOOST_net_14337), .b(FE_OFN1404_n_8567), .o(TIMEBOOST_net_13401) );
na02m02 TIMEBOOST_cell_36810 ( .a(TIMEBOOST_net_10643), .b(n_3460), .o(n_13506) );
in01s01 g62806_u0 ( .a(FE_OFN1122_g64577_p), .o(g62806_sb) );
na02m02 TIMEBOOST_cell_32386 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_23__Q), .o(TIMEBOOST_net_10104) );
in01s01 TIMEBOOST_cell_45931 ( .a(wbm_dat_i_24_), .o(TIMEBOOST_net_15238) );
na02f02 TIMEBOOST_cell_40948 ( .a(TIMEBOOST_net_12712), .b(g57478_sb), .o(n_11259) );
in01s01 g62807_u0 ( .a(FE_OFN1100_g64577_p), .o(g62807_sb) );
na02s02 TIMEBOOST_cell_36812 ( .a(TIMEBOOST_net_10644), .b(g63036_db), .o(n_5176) );
na02s01 g62807_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__14__Q), .b(FE_OFN1100_g64577_p), .o(g62807_db) );
na02s02 TIMEBOOST_cell_36814 ( .a(TIMEBOOST_net_10645), .b(g62833_sb), .o(n_5308) );
in01s01 g62808_u0 ( .a(FE_OFN1106_g64577_p), .o(g62808_sb) );
na02f02 TIMEBOOST_cell_39018 ( .a(TIMEBOOST_net_11747), .b(g52529_sb), .o(n_13688) );
na02s01 g62808_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__13__Q), .b(FE_OFN1106_g64577_p), .o(g62808_db) );
na02f02 TIMEBOOST_cell_10535 ( .a(TIMEBOOST_net_1834), .b(g54155_da), .o(n_13444) );
in01s01 g62809_u0 ( .a(FE_OFN2105_g64577_p), .o(g62809_sb) );
na02s01 TIMEBOOST_cell_37511 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__Q), .b(g64232_sb), .o(TIMEBOOST_net_10994) );
na02s01 TIMEBOOST_cell_37630 ( .a(TIMEBOOST_net_11053), .b(g61784_sb), .o(n_8236) );
na02s02 TIMEBOOST_cell_37632 ( .a(TIMEBOOST_net_11054), .b(g61794_sb), .o(n_8210) );
in01s01 g62810_u0 ( .a(FE_OFN1129_g64577_p), .o(g62810_sb) );
na02s01 TIMEBOOST_cell_44886 ( .a(TIMEBOOST_net_14681), .b(n_4672), .o(TIMEBOOST_net_10977) );
na02s01 TIMEBOOST_cell_38406 ( .a(TIMEBOOST_net_11441), .b(g63556_sb), .o(n_4601) );
na02f02 TIMEBOOST_cell_37058 ( .a(FE_OCP_RBN1961_FE_OFN1591_n_13741), .b(TIMEBOOST_net_10767), .o(g53226_p) );
in01s01 g62811_u0 ( .a(FE_OFN1104_g64577_p), .o(g62811_sb) );
na02s01 TIMEBOOST_cell_36454 ( .a(TIMEBOOST_net_10465), .b(g65717_db), .o(n_1611) );
na02s01 g62811_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__Q), .b(FE_OFN1104_g64577_p), .o(g62811_db) );
na02s01 TIMEBOOST_cell_36456 ( .a(TIMEBOOST_net_10466), .b(g65212_db), .o(n_2676) );
in01s01 g62812_u0 ( .a(FE_OFN1112_g64577_p), .o(g62812_sb) );
na02m02 TIMEBOOST_cell_42566 ( .a(TIMEBOOST_net_13521), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_1__Q), .o(TIMEBOOST_net_10864) );
na02s01 TIMEBOOST_cell_38560 ( .a(TIMEBOOST_net_11518), .b(g62043_sb), .o(n_7769) );
na02m02 TIMEBOOST_cell_45482 ( .a(TIMEBOOST_net_14979), .b(FE_OFN1306_n_13124), .o(TIMEBOOST_net_14464) );
in01s01 g62813_u0 ( .a(FE_OFN1135_g64577_p), .o(g62813_sb) );
na02s01 TIMEBOOST_cell_44882 ( .a(TIMEBOOST_net_14679), .b(g65809_db), .o(n_1904) );
na02s02 TIMEBOOST_cell_39936 ( .a(TIMEBOOST_net_12206), .b(g62493_sb), .o(n_6598) );
na04f04 TIMEBOOST_cell_36232 ( .a(n_13055), .b(n_12792), .c(n_12906), .d(n_12907), .o(n_13138) );
in01s01 g62814_u0 ( .a(FE_OFN877_g64577_p), .o(g62814_sb) );
na04f04 TIMEBOOST_cell_36234 ( .a(n_13050), .b(n_12786), .c(n_12887), .d(n_12886), .o(n_13133) );
in01s01 TIMEBOOST_cell_45920 ( .a(TIMEBOOST_net_15226), .o(TIMEBOOST_net_15227) );
na02s01 TIMEBOOST_cell_17123 ( .a(TIMEBOOST_net_3818), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_1540) );
in01s01 g62815_u0 ( .a(FE_OFN882_g64577_p), .o(g62815_sb) );
no02f08 TIMEBOOST_cell_36258 ( .a(TIMEBOOST_net_10367), .b(n_16287), .o(TIMEBOOST_net_109) );
na02s01 TIMEBOOST_cell_17119 ( .a(TIMEBOOST_net_3816), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_1542) );
in01s01 g62816_u0 ( .a(FE_OFN1122_g64577_p), .o(g62816_sb) );
na02s01 TIMEBOOST_cell_17127 ( .a(TIMEBOOST_net_3820), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_1554) );
na02s01 TIMEBOOST_cell_39938 ( .a(TIMEBOOST_net_12207), .b(g62969_sb), .o(n_5944) );
na02s01 TIMEBOOST_cell_17129 ( .a(TIMEBOOST_net_3821), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_1539) );
in01s01 g62817_u0 ( .a(FE_OFN2105_g64577_p), .o(g62817_sb) );
na03s02 TIMEBOOST_cell_37545 ( .a(TIMEBOOST_net_3787), .b(g65965_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__Q), .o(TIMEBOOST_net_11011) );
na02s01 TIMEBOOST_cell_37634 ( .a(TIMEBOOST_net_11055), .b(g61774_sb), .o(n_8260) );
na02s01 TIMEBOOST_cell_37636 ( .a(TIMEBOOST_net_11056), .b(g61773_sb), .o(n_8262) );
in01s01 g62818_u0 ( .a(FE_OFN882_g64577_p), .o(g62818_sb) );
na02s01 TIMEBOOST_cell_17121 ( .a(TIMEBOOST_net_3817), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_1555) );
na03f02 TIMEBOOST_cell_21824 ( .a(n_3068), .b(n_2925), .c(n_2858), .o(TIMEBOOST_net_6169) );
na03f02 TIMEBOOST_cell_36200 ( .a(n_12357), .b(TIMEBOOST_net_10295), .c(n_11831), .o(n_12645) );
in01s01 g62819_u0 ( .a(FE_OFN2105_g64577_p), .o(g62819_sb) );
na03f02 TIMEBOOST_cell_36202 ( .a(n_12357), .b(TIMEBOOST_net_10293), .c(n_11831), .o(n_12728) );
na03s01 TIMEBOOST_cell_39449 ( .a(TIMEBOOST_net_3351), .b(g64085_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__Q), .o(TIMEBOOST_net_11963) );
na02s01 TIMEBOOST_cell_36340 ( .a(TIMEBOOST_net_10408), .b(g67040_sb), .o(n_1681) );
in01s01 g62820_u0 ( .a(FE_OFN1125_g64577_p), .o(g62820_sb) );
na02s01 TIMEBOOST_cell_36278 ( .a(TIMEBOOST_net_10377), .b(FE_OFN988_n_574), .o(n_1634) );
na02s02 TIMEBOOST_cell_39940 ( .a(TIMEBOOST_net_12208), .b(g62447_sb), .o(n_7385) );
na02s02 TIMEBOOST_cell_36260 ( .a(TIMEBOOST_net_10368), .b(n_2681), .o(TIMEBOOST_net_484) );
in01s01 g62821_u0 ( .a(FE_OFN1097_g64577_p), .o(g62821_sb) );
na02s02 TIMEBOOST_cell_36886 ( .a(TIMEBOOST_net_10681), .b(g61863_db), .o(n_8111) );
na02s01 g62821_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__Q), .b(FE_OFN1097_g64577_p), .o(g62821_db) );
na02f02 TIMEBOOST_cell_12643 ( .a(TIMEBOOST_net_2888), .b(n_14207), .o(n_14449) );
in01s01 g62822_u0 ( .a(FE_OFN1133_g64577_p), .o(g62822_sb) );
na02m02 TIMEBOOST_cell_36262 ( .a(wbu_addr_in_251), .b(TIMEBOOST_net_10369), .o(TIMEBOOST_net_3167) );
na02s01 TIMEBOOST_cell_44970 ( .a(TIMEBOOST_net_14723), .b(g58075_db), .o(n_9719) );
na03f02 TIMEBOOST_cell_36204 ( .a(n_12101), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__Q), .c(FE_OFN1757_n_12681), .o(n_12526) );
in01s01 g62823_u0 ( .a(FE_OFN1112_g64577_p), .o(g62823_sb) );
na03f02 TIMEBOOST_cell_36206 ( .a(n_12259), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__Q), .c(FE_OFN1577_n_12028), .o(n_12689) );
na02s02 TIMEBOOST_cell_39942 ( .a(TIMEBOOST_net_12209), .b(g62996_sb), .o(n_5890) );
na03f02 TIMEBOOST_cell_36208 ( .a(n_12058), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__Q), .c(FE_OFN1757_n_12681), .o(n_12481) );
in01s01 g62824_u0 ( .a(FE_OFN1116_g64577_p), .o(g62824_sb) );
na02m02 TIMEBOOST_cell_38886 ( .a(TIMEBOOST_net_11681), .b(g58485_sb), .o(n_9350) );
na02s02 TIMEBOOST_cell_45731 ( .a(n_3631), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__Q), .o(TIMEBOOST_net_15104) );
in01s01 g62825_u0 ( .a(FE_OFN1124_g64577_p), .o(g62825_sb) );
na02f02 TIMEBOOST_cell_18316 ( .a(n_2922), .b(n_3004), .o(TIMEBOOST_net_4415) );
na02f02 TIMEBOOST_cell_39172 ( .a(TIMEBOOST_net_11824), .b(FE_RN_333_0), .o(FE_RN_355_0) );
na02s01 g52468_u1 ( .a(wbs_adr_i_22_), .b(g52463_sb), .o(g52468_da) );
in01s01 g62826_u0 ( .a(FE_OFN2106_g64577_p), .o(g62826_sb) );
na02s01 TIMEBOOST_cell_37509 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__Q), .b(g64347_sb), .o(TIMEBOOST_net_10993) );
na02s01 TIMEBOOST_cell_37638 ( .a(TIMEBOOST_net_11057), .b(g61995_sb), .o(n_7905) );
na02s01 TIMEBOOST_cell_37640 ( .a(TIMEBOOST_net_11058), .b(g61993_sb), .o(n_7909) );
in01s01 g62827_u0 ( .a(FE_OFN1120_g64577_p), .o(g62827_sb) );
na03f03 TIMEBOOST_cell_45853 ( .a(n_11090), .b(n_11089), .c(n_10785), .o(TIMEBOOST_net_15165) );
na02s01 TIMEBOOST_cell_37642 ( .a(TIMEBOOST_net_11059), .b(g61886_sb), .o(n_8059) );
na02s01 TIMEBOOST_cell_37644 ( .a(TIMEBOOST_net_11060), .b(g61750_sb), .o(n_8316) );
in01s01 g62828_u0 ( .a(FE_OFN2106_g64577_p), .o(g62828_sb) );
na02s01 TIMEBOOST_cell_37507 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__Q), .b(g64265_sb), .o(TIMEBOOST_net_10992) );
na02s01 TIMEBOOST_cell_37646 ( .a(TIMEBOOST_net_11061), .b(g61910_sb), .o(n_8001) );
na02s01 TIMEBOOST_cell_37648 ( .a(TIMEBOOST_net_11062), .b(g61763_sb), .o(n_8285) );
in01s01 g62829_u0 ( .a(FE_OFN1124_g64577_p), .o(g62829_sb) );
na02s01 g52462_u1 ( .a(wbs_adr_i_16_), .b(g52462_sb), .o(g52462_da) );
na03s02 TIMEBOOST_cell_34799 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .b(g62719_sb), .c(g62719_db), .o(n_6138) );
na03f02 TIMEBOOST_cell_36196 ( .a(n_12068), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__Q), .c(n_11823), .o(n_12489) );
in01s01 g62830_u0 ( .a(FE_OFN1120_g64577_p), .o(g62830_sb) );
na02f02 TIMEBOOST_cell_44666 ( .a(TIMEBOOST_net_14571), .b(FE_OFN1417_n_8567), .o(TIMEBOOST_net_12785) );
na02s01 TIMEBOOST_cell_37650 ( .a(TIMEBOOST_net_11063), .b(g62069_sb), .o(n_7830) );
na02s02 TIMEBOOST_cell_36760 ( .a(TIMEBOOST_net_10618), .b(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_4494) );
in01s01 g62831_u0 ( .a(FE_OFN877_g64577_p), .o(g62831_sb) );
na03s01 TIMEBOOST_cell_33955 ( .a(n_1719), .b(g61903_sb), .c(g61903_db), .o(n_8017) );
na02s01 TIMEBOOST_cell_45065 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__Q), .b(FE_OFN543_n_9690), .o(TIMEBOOST_net_14771) );
na03s01 TIMEBOOST_cell_33956 ( .a(n_1879), .b(g61909_sb), .c(g61909_db), .o(n_8003) );
in01s01 g62832_u0 ( .a(FE_OFN1136_g64577_p), .o(g62832_sb) );
na03s01 TIMEBOOST_cell_33957 ( .a(n_1888), .b(g61893_sb), .c(g61893_db), .o(n_8041) );
na02s02 TIMEBOOST_cell_10902 ( .a(g54191_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_410), .o(TIMEBOOST_net_2018) );
na03s02 TIMEBOOST_cell_33958 ( .a(n_1844), .b(g61865_sb), .c(g61865_db), .o(n_8107) );
in01s01 g62833_u0 ( .a(FE_OFN1134_g64577_p), .o(g62833_sb) );
na02m02 TIMEBOOST_cell_43564 ( .a(TIMEBOOST_net_14020), .b(FE_OFN1313_n_6624), .o(TIMEBOOST_net_12240) );
na02s01 g62833_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__Q), .b(FE_OFN1104_g64577_p), .o(g62833_db) );
na02f02 TIMEBOOST_cell_44268 ( .a(TIMEBOOST_net_14372), .b(FE_OFN1423_n_8567), .o(TIMEBOOST_net_12832) );
in01s01 g62834_u0 ( .a(FE_OFN1118_g64577_p), .o(g62834_sb) );
na03s01 TIMEBOOST_cell_33961 ( .a(n_2160), .b(g62000_sb), .c(g62000_db), .o(n_7895) );
na02m02 TIMEBOOST_cell_21828 ( .a(g59126_db), .b(g59126_sb), .o(TIMEBOOST_net_6171) );
na03f02 TIMEBOOST_cell_36156 ( .a(FE_OFN2209_n_11027), .b(TIMEBOOST_net_10279), .c(FE_OFN1752_n_12086), .o(n_12745) );
in01s01 g62835_u0 ( .a(FE_OFN1106_g64577_p), .o(g62835_sb) );
na02s02 TIMEBOOST_cell_10536 ( .a(n_211), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_1835) );
na02s01 g62835_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN1106_g64577_p), .o(g62835_db) );
na02s02 TIMEBOOST_cell_37842 ( .a(TIMEBOOST_net_11159), .b(g58488_sb), .o(n_9345) );
in01s01 g62836_u0 ( .a(FE_OFN2105_g64577_p), .o(g62836_sb) );
na02s04 TIMEBOOST_cell_44755 ( .a(conf_wb_err_addr_in_969), .b(conf_wb_err_addr_in_970), .o(TIMEBOOST_net_14616) );
na02s01 TIMEBOOST_cell_37652 ( .a(TIMEBOOST_net_11064), .b(g61720_sb), .o(n_8384) );
na02s01 TIMEBOOST_cell_37654 ( .a(TIMEBOOST_net_11065), .b(g61946_sb), .o(n_7933) );
in01s01 g62837_u0 ( .a(FE_OFN1119_g64577_p), .o(g62837_sb) );
na02s02 TIMEBOOST_cell_42983 ( .a(TIMEBOOST_net_4302), .b(FE_OFN2212_n_8407), .o(TIMEBOOST_net_13730) );
na02s01 TIMEBOOST_cell_37656 ( .a(TIMEBOOST_net_11066), .b(g61727_sb), .o(n_8366) );
na02s02 TIMEBOOST_cell_37658 ( .a(TIMEBOOST_net_11067), .b(g62006_sb), .o(n_7883) );
in01s01 g62838_u0 ( .a(FE_OFN1122_g64577_p), .o(g62838_sb) );
na03f02 TIMEBOOST_cell_36158 ( .a(FE_OFN2209_n_11027), .b(TIMEBOOST_net_10277), .c(FE_OFN1752_n_12086), .o(n_12751) );
na03s02 TIMEBOOST_cell_38171 ( .a(TIMEBOOST_net_3355), .b(g64202_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__Q), .o(TIMEBOOST_net_11324) );
na03f02 TIMEBOOST_cell_36160 ( .a(FE_OFN2210_n_11027), .b(TIMEBOOST_net_10272), .c(FE_OFN1752_n_12086), .o(n_12618) );
in01s01 g62839_u0 ( .a(FE_OFN1135_g64577_p), .o(g62839_sb) );
na03f02 TIMEBOOST_cell_36162 ( .a(FE_OFN2210_n_11027), .b(TIMEBOOST_net_10264), .c(FE_OFN1753_n_12086), .o(n_12717) );
na04f02 TIMEBOOST_cell_34805 ( .a(g52395_db), .b(n_3317), .c(g52395_sb), .d(TIMEBOOST_net_593), .o(n_14826) );
na04f02 TIMEBOOST_cell_36164 ( .a(n_11793), .b(n_11149), .c(n_11148), .d(n_11152), .o(n_12556) );
in01s01 g62840_u0 ( .a(FE_OFN1135_g64577_p), .o(g62840_sb) );
na02s03 TIMEBOOST_cell_45763 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__Q), .b(n_13182), .o(TIMEBOOST_net_15120) );
na02m02 TIMEBOOST_cell_38981 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_4__Q), .o(TIMEBOOST_net_11729) );
na02s01 TIMEBOOST_cell_43437 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__Q), .b(n_3598), .o(TIMEBOOST_net_13957) );
in01s01 g62841_u0 ( .a(FE_OFN1115_g64577_p), .o(g62841_sb) );
na02m02 TIMEBOOST_cell_38718 ( .a(TIMEBOOST_net_11597), .b(g59806_sb), .o(n_7617) );
na02s01 TIMEBOOST_cell_19014 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q), .b(g58331_sb), .o(TIMEBOOST_net_4764) );
na02s01 TIMEBOOST_cell_37258 ( .a(TIMEBOOST_net_10867), .b(FE_OFN687_n_4417), .o(TIMEBOOST_net_9391) );
in01s01 g62842_u0 ( .a(FE_OFN2106_g64577_p), .o(g62842_sb) );
na02s02 TIMEBOOST_cell_37499 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__Q), .b(g58356_sb), .o(TIMEBOOST_net_10988) );
na02s01 TIMEBOOST_cell_37660 ( .a(TIMEBOOST_net_11068), .b(g61805_sb), .o(n_8184) );
na02s01 TIMEBOOST_cell_37209 ( .a(n_12179), .b(n_657), .o(TIMEBOOST_net_10843) );
in01s01 g62843_u0 ( .a(FE_OFN1104_g64577_p), .o(g62843_sb) );
na02f02 TIMEBOOST_cell_37070 ( .a(TIMEBOOST_net_10773), .b(FE_OFN1589_n_13736), .o(n_16238) );
na02s01 g62843_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__Q), .b(FE_OFN1104_g64577_p), .o(g62843_db) );
na02f02 TIMEBOOST_cell_37106 ( .a(TIMEBOOST_net_10791), .b(n_12561), .o(n_12823) );
in01s01 g62844_u0 ( .a(FE_OFN881_g64577_p), .o(g62844_sb) );
na02f02 TIMEBOOST_cell_36816 ( .a(TIMEBOOST_net_10646), .b(g54321_db), .o(n_13000) );
na02s01 g62844_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__Q), .b(FE_OFN881_g64577_p), .o(g62844_db) );
na02f02 TIMEBOOST_cell_37060 ( .a(g52614_db), .b(TIMEBOOST_net_10768), .o(TIMEBOOST_net_10194) );
in01s01 g62845_u0 ( .a(FE_OFN1135_g64577_p), .o(g62845_sb) );
na02s01 TIMEBOOST_cell_36342 ( .a(TIMEBOOST_net_10409), .b(g67051_sb), .o(n_1497) );
na02s02 TIMEBOOST_cell_10914 ( .a(g54179_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_399), .o(TIMEBOOST_net_2024) );
na02s01 TIMEBOOST_cell_41734 ( .a(TIMEBOOST_net_13105), .b(g57893_db), .o(n_9141) );
in01s01 g62846_u0 ( .a(FE_OFN1136_g64577_p), .o(g62846_sb) );
na02f02 TIMEBOOST_cell_12619 ( .a(TIMEBOOST_net_2876), .b(n_13901), .o(TIMEBOOST_net_938) );
na02s02 TIMEBOOST_cell_43055 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q), .b(n_4310), .o(TIMEBOOST_net_13766) );
na02s01 TIMEBOOST_cell_38408 ( .a(TIMEBOOST_net_11442), .b(g62786_sb), .o(n_5418) );
in01s01 g62847_u0 ( .a(FE_OFN1121_g64577_p), .o(g62847_sb) );
na02f02 TIMEBOOST_cell_41580 ( .a(TIMEBOOST_net_13028), .b(g57596_sb), .o(n_10797) );
na02s01 TIMEBOOST_cell_37418 ( .a(TIMEBOOST_net_10947), .b(FE_OFN1809_n_4454), .o(TIMEBOOST_net_10552) );
na02s01 TIMEBOOST_cell_31786 ( .a(parchk_pci_ad_out_in_1183), .b(configuration_wb_err_data_586), .o(TIMEBOOST_net_9804) );
in01s01 g62848_u0 ( .a(FE_OFN1106_g64577_p), .o(g62848_sb) );
na02s01 TIMEBOOST_cell_39362 ( .a(TIMEBOOST_net_11919), .b(g61882_sb), .o(n_8066) );
na02s01 g62848_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__13__Q), .b(FE_OFN1106_g64577_p), .o(g62848_db) );
na02f02 TIMEBOOST_cell_37090 ( .a(TIMEBOOST_net_10783), .b(FE_OFN1587_n_13736), .o(g53154_p) );
in01s01 g62849_u0 ( .a(FE_OFN877_g64577_p), .o(g62849_sb) );
na02s01 TIMEBOOST_cell_42850 ( .a(TIMEBOOST_net_13663), .b(FE_OFN720_n_8060), .o(TIMEBOOST_net_11248) );
na02m02 TIMEBOOST_cell_41607 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_6__Q), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_13042) );
na02s01 TIMEBOOST_cell_32030 ( .a(configuration_pci_err_addr_482), .b(wbm_adr_o_12_), .o(TIMEBOOST_net_9926) );
in01s01 g62850_u0 ( .a(FE_OFN1129_g64577_p), .o(g62850_sb) );
na02s02 TIMEBOOST_cell_32029 ( .a(TIMEBOOST_net_9925), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_4907) );
na02m02 TIMEBOOST_cell_10922 ( .a(g54030_sb), .b(n_12595), .o(TIMEBOOST_net_2028) );
na02m02 TIMEBOOST_cell_43719 ( .a(n_9523), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__Q), .o(TIMEBOOST_net_14098) );
in01s01 g62851_u0 ( .a(FE_OFN881_g64577_p), .o(g62851_sb) );
na02s01 TIMEBOOST_cell_36818 ( .a(TIMEBOOST_net_10647), .b(g61939_db), .o(n_7945) );
na02s01 TIMEBOOST_cell_19020 ( .a(wishbone_slave_unit_pcim_sm_data_in_652), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__Q), .o(TIMEBOOST_net_4767) );
na02s01 TIMEBOOST_cell_17531 ( .a(TIMEBOOST_net_4022), .b(g65920_sb), .o(n_1566) );
in01s01 g62852_u0 ( .a(FE_OFN1104_g64577_p), .o(g62852_sb) );
na02s02 TIMEBOOST_cell_36712 ( .a(TIMEBOOST_net_10594), .b(g63593_sb), .o(n_4775) );
na02s01 g62852_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__Q), .b(FE_OFN1104_g64577_p), .o(g62852_db) );
na02s02 TIMEBOOST_cell_36714 ( .a(TIMEBOOST_net_10595), .b(g63594_sb), .o(n_4774) );
in01s01 g62853_u0 ( .a(FE_OFN1120_g64577_p), .o(g62853_sb) );
na02f02 TIMEBOOST_cell_41150 ( .a(TIMEBOOST_net_12813), .b(g57220_sb), .o(n_11535) );
na02s02 TIMEBOOST_cell_37662 ( .a(TIMEBOOST_net_11069), .b(g61869_sb), .o(n_8097) );
na02s01 TIMEBOOST_cell_37664 ( .a(TIMEBOOST_net_11070), .b(g61905_sb), .o(n_8012) );
in01s01 g62854_u0 ( .a(FE_OFN1118_g64577_p), .o(g62854_sb) );
na02s01 TIMEBOOST_cell_18789 ( .a(TIMEBOOST_net_4651), .b(g62860_sb), .o(n_5246) );
na02s02 TIMEBOOST_cell_39396 ( .a(TIMEBOOST_net_11936), .b(g58377_sb), .o(n_9452) );
na02m02 TIMEBOOST_cell_36344 ( .a(TIMEBOOST_net_10410), .b(n_2256), .o(TIMEBOOST_net_131) );
in01s01 g62855_u0 ( .a(FE_OFN1112_g64577_p), .o(g62855_sb) );
na03f02 TIMEBOOST_cell_45483 ( .a(n_8548), .b(n_317), .c(FE_OFN1403_n_8567), .o(TIMEBOOST_net_14980) );
na02m02 TIMEBOOST_cell_39174 ( .a(g57795_da), .b(TIMEBOOST_net_11825), .o(TIMEBOOST_net_6243) );
na03s02 TIMEBOOST_cell_42063 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__Q), .b(n_3611), .c(FE_OFN1278_n_4097), .o(TIMEBOOST_net_13270) );
in01s01 g62856_u0 ( .a(FE_OFN1135_g64577_p), .o(g62856_sb) );
na03f02 TIMEBOOST_cell_32937 ( .a(n_2675), .b(n_1774), .c(n_16495), .o(n_3452) );
na02s02 TIMEBOOST_cell_38410 ( .a(TIMEBOOST_net_11443), .b(g62812_sb), .o(n_5354) );
na03f02 TIMEBOOST_cell_22350 ( .a(n_9311), .b(n_10176), .c(n_9312), .o(TIMEBOOST_net_6432) );
in01s01 g62857_u0 ( .a(FE_OFN1137_g64577_p), .o(g62857_sb) );
na02m02 TIMEBOOST_cell_44183 ( .a(n_9521), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__Q), .o(TIMEBOOST_net_14330) );
na02s02 TIMEBOOST_cell_44424 ( .a(TIMEBOOST_net_14450), .b(FE_OFN1306_n_13124), .o(TIMEBOOST_net_13417) );
na02s02 TIMEBOOST_cell_45194 ( .a(TIMEBOOST_net_14835), .b(FE_OFN1244_n_4092), .o(TIMEBOOST_net_12095) );
in01s01 g62858_u0 ( .a(FE_OFN1097_g64577_p), .o(g62858_sb) );
na02m02 TIMEBOOST_cell_36820 ( .a(TIMEBOOST_net_10648), .b(g54170_sb), .o(TIMEBOOST_net_9881) );
na02s01 g62858_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__Q), .b(FE_OFN1097_g64577_p), .o(g62858_db) );
na02s01 TIMEBOOST_cell_17521 ( .a(TIMEBOOST_net_4017), .b(g65856_sb), .o(n_1582) );
in01s01 g62859_u0 ( .a(FE_OFN1100_g64577_p), .o(g62859_sb) );
na02s01 TIMEBOOST_cell_36458 ( .a(TIMEBOOST_net_10467), .b(g58009_sb), .o(TIMEBOOST_net_9779) );
na02s01 g62859_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__14__Q), .b(FE_OFN1100_g64577_p), .o(g62859_db) );
na02s01 TIMEBOOST_cell_36460 ( .a(TIMEBOOST_net_10468), .b(g58206_sb), .o(TIMEBOOST_net_9774) );
in01s01 g62860_u0 ( .a(FE_OFN2104_g64577_p), .o(g62860_sb) );
na02s02 TIMEBOOST_cell_36762 ( .a(TIMEBOOST_net_10619), .b(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_4705) );
na02m02 TIMEBOOST_cell_44199 ( .a(n_1609), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .o(TIMEBOOST_net_14338) );
na02f02 TIMEBOOST_cell_12866 ( .a(FE_OFN1587_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__Q), .o(TIMEBOOST_net_3000) );
in01s01 g62861_u0 ( .a(FE_OFN2104_g64577_p), .o(g62861_sb) );
na02s01 TIMEBOOST_cell_37571 ( .a(parchk_pci_ad_reg_in_1235), .b(g65893_sb), .o(TIMEBOOST_net_11024) );
na02s01 TIMEBOOST_cell_37207 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(g65707_sb), .o(TIMEBOOST_net_10842) );
na02s01 TIMEBOOST_cell_37666 ( .a(TIMEBOOST_net_11071), .b(g61821_sb), .o(n_8147) );
in01s01 g62862_u0 ( .a(FE_OFN1136_g64577_p), .o(g62862_sb) );
na02f02 TIMEBOOST_cell_12868 ( .a(FE_OFN1586_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__Q), .o(TIMEBOOST_net_3001) );
na02s01 TIMEBOOST_cell_38412 ( .a(TIMEBOOST_net_11444), .b(g63554_sb), .o(n_4603) );
na02f02 TIMEBOOST_cell_44050 ( .a(TIMEBOOST_net_14263), .b(FE_OFN1421_n_8567), .o(TIMEBOOST_net_12941) );
in01s01 g62863_u0 ( .a(FE_OFN1131_g64577_p), .o(g62863_sb) );
na02s02 TIMEBOOST_cell_43438 ( .a(TIMEBOOST_net_13957), .b(FE_OFN1232_n_6391), .o(TIMEBOOST_net_12184) );
na02s01 TIMEBOOST_cell_39482 ( .a(TIMEBOOST_net_11979), .b(TIMEBOOST_net_9823), .o(n_7153) );
na02m02 TIMEBOOST_cell_44051 ( .a(n_9071), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q), .o(TIMEBOOST_net_14264) );
in01s01 g62864_u0 ( .a(FE_OFN1123_g64577_p), .o(g62864_sb) );
na03f02 TIMEBOOST_cell_35947 ( .a(TIMEBOOST_net_10100), .b(FE_OFN1472_g52675_p), .c(g52517_sb), .o(n_13798) );
na02s02 g62864_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__Q), .b(FE_OFN1115_g64577_p), .o(g62864_db) );
na02f04 TIMEBOOST_cell_39020 ( .a(TIMEBOOST_net_11748), .b(FE_OFN2243_g52675_p), .o(TIMEBOOST_net_10750) );
in01s01 g62865_u0 ( .a(FE_OFN882_g64577_p), .o(g62865_sb) );
na02f02 TIMEBOOST_cell_37108 ( .a(TIMEBOOST_net_10792), .b(n_12562), .o(n_12824) );
na02s02 TIMEBOOST_cell_18647 ( .a(TIMEBOOST_net_4580), .b(g63134_sb), .o(n_4982) );
na02s01 TIMEBOOST_cell_38642 ( .a(TIMEBOOST_net_11559), .b(g59109_sb), .o(n_8709) );
na02s01 TIMEBOOST_cell_30740 ( .a(pci_ad_i_15_), .b(parchk_pci_ad_reg_in_1219), .o(TIMEBOOST_net_9281) );
na02s01 TIMEBOOST_cell_30854 ( .a(n_3741), .b(g65044_sb), .o(TIMEBOOST_net_9338) );
ao22f02 g62868_u0 ( .a(n_4642), .b(n_16160), .c(n_1447), .d(pci_target_unit_wbm_sm_pci_tar_read_request), .o(n_17030) );
ao12f02 g62869_u0 ( .a(n_3321), .b(n_16000), .c(n_2833), .o(n_4155) );
ao12f02 g62870_u0 ( .a(n_4136), .b(FE_OFN1066_n_15808), .c(configuration_pci_err_data_504), .o(n_4803) );
ao12f02 g62871_u0 ( .a(n_4135), .b(FE_OFN1066_n_15808), .c(configuration_pci_err_data_506), .o(n_4802) );
oa12s02 g62872_u0 ( .a(n_3327), .b(conf_wb_err_addr_in_943), .c(FE_OFN1142_n_15261), .o(n_4154) );
no02s01 g62873_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_), .b(n_1419), .o(g62873_p) );
ao12s01 g62873_u1 ( .a(g62873_p), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_), .c(n_1419), .o(n_2274) );
no02s01 g62874_u0 ( .a(wbu_addr_in_254), .b(n_2013), .o(g62874_p) );
ao12s01 g62874_u1 ( .a(g62874_p), .b(wbu_addr_in_254), .c(n_2013), .o(n_2273) );
no02m02 g62875_u0 ( .a(n_2436), .b(conf_wb_err_addr_in_957), .o(g62875_p) );
ao12m02 g62875_u1 ( .a(g62875_p), .b(conf_wb_err_addr_in_957), .c(n_2436), .o(n_3153) );
no02s01 g62876_u0 ( .a(n_1463), .b(conf_wb_err_addr_in_946), .o(g62876_p) );
ao12s02 g62876_u1 ( .a(g62876_p), .b(conf_wb_err_addr_in_946), .c(n_1463), .o(n_2272) );
no02s01 g62877_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_3_), .b(n_1190), .o(g62877_p) );
ao12s01 g62877_u1 ( .a(g62877_p), .b(pci_target_unit_del_sync_comp_cycle_count_3_), .c(n_1190), .o(n_2024) );
oa12s01 g62878_u0 ( .a(n_3447), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_0_), .c(n_4662), .o(n_4659) );
no02s01 g62879_u0 ( .a(n_2012), .b(wbm_adr_o_5_), .o(g62879_p) );
ao12s01 g62879_u1 ( .a(g62879_p), .b(wbm_adr_o_5_), .c(n_2012), .o(n_2271) );
no02s01 g62880_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_3_), .b(n_1213), .o(g62880_p) );
ao12s01 g62880_u1 ( .a(g62880_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_3_), .c(n_1213), .o(n_2023) );
no02s02 g62881_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_3_), .b(n_1216), .o(g62881_p) );
ao12s01 g62881_u1 ( .a(g62881_p), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_3_), .c(n_1216), .o(n_2022) );
no02m01 g62882_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr), .b(FE_OFN1192_n_6935), .o(g62882_p) );
ao12m01 g62882_u1 ( .a(g62882_p), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .c(FE_OFN1192_n_6935), .o(n_6112) );
in01s01 g62883_u0 ( .a(FE_OFN1202_n_4090), .o(g62883_sb) );
na02s02 TIMEBOOST_cell_16368 ( .a(n_3744), .b(g65083_sb), .o(TIMEBOOST_net_3441) );
na03s02 TIMEBOOST_cell_37581 ( .a(n_2061), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__Q), .c(FE_OFN2081_n_8176), .o(TIMEBOOST_net_11029) );
na02s01 TIMEBOOST_cell_3218 ( .a(g65902_db), .b(g61705_sb), .o(TIMEBOOST_net_189) );
in01s01 g62884_u0 ( .a(FE_OFN1288_n_4098), .o(g62884_sb) );
na02s02 TIMEBOOST_cell_36597 ( .a(n_1117), .b(n_7835), .o(TIMEBOOST_net_10537) );
na02s02 TIMEBOOST_cell_31083 ( .a(TIMEBOOST_net_9452), .b(n_4479), .o(n_4330) );
na02f02 TIMEBOOST_cell_43720 ( .a(TIMEBOOST_net_14098), .b(FE_OFN1409_n_8567), .o(TIMEBOOST_net_12751) );
in01s01 g62885_u0 ( .a(FE_OFN1310_n_6624), .o(g62885_sb) );
na02f02 TIMEBOOST_cell_44052 ( .a(TIMEBOOST_net_14264), .b(FE_OFN1412_n_8567), .o(TIMEBOOST_net_12850) );
na02f04 TIMEBOOST_cell_3809 ( .a(TIMEBOOST_net_484), .b(n_2971), .o(n_3179) );
na02s02 TIMEBOOST_cell_17963 ( .a(TIMEBOOST_net_4238), .b(g65358_da), .o(n_4255) );
in01s01 g62886_u0 ( .a(FE_OFN1289_n_4098), .o(g62886_sb) );
na02s02 TIMEBOOST_cell_36599 ( .a(TIMEBOOST_net_775), .b(n_3395), .o(TIMEBOOST_net_10538) );
na02s01 TIMEBOOST_cell_30845 ( .a(TIMEBOOST_net_9333), .b(g64903_db), .o(n_3692) );
na02m02 TIMEBOOST_cell_44529 ( .a(n_9094), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__Q), .o(TIMEBOOST_net_14503) );
in01s01 g62887_u0 ( .a(FE_OFN1249_n_4093), .o(g62887_sb) );
na02s01 TIMEBOOST_cell_36601 ( .a(TIMEBOOST_net_3701), .b(FE_OFN1042_n_2037), .o(TIMEBOOST_net_10539) );
na02f02 TIMEBOOST_cell_44053 ( .a(n_9030), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__Q), .o(TIMEBOOST_net_14265) );
na02s02 TIMEBOOST_cell_30885 ( .a(TIMEBOOST_net_9353), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_3731) );
in01s01 g62888_u0 ( .a(FE_OFN1258_n_4143), .o(g62888_sb) );
na02s01 TIMEBOOST_cell_36607 ( .a(g58227_sb), .b(g58227_db), .o(TIMEBOOST_net_10542) );
na02f02 TIMEBOOST_cell_45484 ( .a(TIMEBOOST_net_14980), .b(g58608_sb), .o(n_8899) );
na02s02 TIMEBOOST_cell_30801 ( .a(TIMEBOOST_net_9311), .b(wbu_addr_in_263), .o(n_9124) );
in01s01 g62889_u0 ( .a(FE_OFN1253_n_4143), .o(g62889_sb) );
na02s01 TIMEBOOST_cell_36609 ( .a(pci_target_unit_del_sync_bc_in_203), .b(g65940_db), .o(TIMEBOOST_net_10543) );
na02s01 TIMEBOOST_cell_30853 ( .a(TIMEBOOST_net_9337), .b(g65026_sb), .o(n_3628) );
na02m02 TIMEBOOST_cell_30803 ( .a(TIMEBOOST_net_9312), .b(g58797_db), .o(n_9868) );
in01s01 g62890_u0 ( .a(FE_OFN1265_n_4095), .o(g62890_sb) );
na02s01 TIMEBOOST_cell_36611 ( .a(FE_OFN231_n_9839), .b(g58156_sb), .o(TIMEBOOST_net_10544) );
na02f02 TIMEBOOST_cell_43740 ( .a(TIMEBOOST_net_14108), .b(FE_OFN1374_n_8567), .o(TIMEBOOST_net_12768) );
na02s02 TIMEBOOST_cell_30883 ( .a(TIMEBOOST_net_9352), .b(FE_OFN784_n_2678), .o(TIMEBOOST_net_3732) );
in01s01 g62891_u0 ( .a(FE_OFN1272_n_4096), .o(g62891_sb) );
na02s01 TIMEBOOST_cell_42917 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__Q), .b(FE_OFN587_n_9692), .o(TIMEBOOST_net_13697) );
na02f02 TIMEBOOST_cell_45854 ( .a(TIMEBOOST_net_15165), .b(n_11088), .o(n_12543) );
na02s01 TIMEBOOST_cell_42640 ( .a(TIMEBOOST_net_13558), .b(g57973_db), .o(n_9115) );
in01s01 g62892_u0 ( .a(FE_OFN1219_n_6886), .o(g62892_sb) );
na02s01 TIMEBOOST_cell_36613 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__Q), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_10545) );
na02s02 TIMEBOOST_cell_30847 ( .a(TIMEBOOST_net_9334), .b(g64916_sb), .o(n_3687) );
na02s01 TIMEBOOST_cell_30859 ( .a(TIMEBOOST_net_9340), .b(FE_OFN223_n_9844), .o(n_9737) );
in01s01 g62893_u0 ( .a(FE_OFN1248_n_4093), .o(g62893_sb) );
na03f02 TIMEBOOST_cell_45485 ( .a(n_8550), .b(n_251), .c(FE_OFN2182_n_8567), .o(TIMEBOOST_net_14981) );
na03f04 TIMEBOOST_cell_45855 ( .a(n_10617), .b(n_10029), .c(n_10916), .o(TIMEBOOST_net_15166) );
na02m02 TIMEBOOST_cell_43721 ( .a(n_9066), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__Q), .o(TIMEBOOST_net_14099) );
in01s01 g62894_u0 ( .a(FE_OFN1202_n_4090), .o(g62894_sb) );
na02m04 TIMEBOOST_cell_3223 ( .a(n_2397), .b(TIMEBOOST_net_191), .o(n_2398) );
na02f02 TIMEBOOST_cell_37808 ( .a(TIMEBOOST_net_11142), .b(FE_OFN2128_n_16497), .o(n_12982) );
na02f02 TIMEBOOST_cell_45486 ( .a(TIMEBOOST_net_14981), .b(g58606_sb), .o(n_8955) );
in01s01 g62895_u0 ( .a(FE_OFN1260_n_4143), .o(g62895_sb) );
na02s01 TIMEBOOST_cell_36615 ( .a(g58225_sb), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_10546) );
na02s01 TIMEBOOST_cell_41762 ( .a(TIMEBOOST_net_13119), .b(TIMEBOOST_net_3575), .o(TIMEBOOST_net_5433) );
na02s01 TIMEBOOST_cell_39944 ( .a(TIMEBOOST_net_12210), .b(g62485_sb), .o(n_6617) );
in01s01 g62896_u0 ( .a(FE_OFN1284_n_4097), .o(g62896_sb) );
na02s01 TIMEBOOST_cell_36617 ( .a(pci_target_unit_del_sync_bc_in_202), .b(g65946_db), .o(TIMEBOOST_net_10547) );
na02s02 TIMEBOOST_cell_42006 ( .a(TIMEBOOST_net_13241), .b(g62525_sb), .o(n_6526) );
in01s01 g62897_u0 ( .a(FE_OFN1294_n_4098), .o(g62897_sb) );
na02s01 TIMEBOOST_cell_36537 ( .a(TIMEBOOST_net_9323), .b(FE_OFN951_n_2055), .o(TIMEBOOST_net_10507) );
na02s01 TIMEBOOST_cell_16820 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__Q), .b(g65323_sb), .o(TIMEBOOST_net_3667) );
na03s02 TIMEBOOST_cell_41809 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__Q), .b(g64306_da), .c(g64306_db), .o(TIMEBOOST_net_13143) );
in01s01 g62898_u0 ( .a(FE_OFN1310_n_6624), .o(g62898_sb) );
na02s02 TIMEBOOST_cell_43464 ( .a(TIMEBOOST_net_13970), .b(FE_OFN1233_n_6391), .o(TIMEBOOST_net_12169) );
na02s02 TIMEBOOST_cell_37559 ( .a(pci_target_unit_pcit_if_strd_addr_in_696), .b(g52625_sb), .o(TIMEBOOST_net_11018) );
na02s01 TIMEBOOST_cell_22304 ( .a(g52472_da), .b(FE_OFN1022_n_11877), .o(TIMEBOOST_net_6409) );
in01s01 g62899_u0 ( .a(FE_OFN1214_n_4151), .o(g62899_sb) );
na02s01 TIMEBOOST_cell_36619 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__Q), .b(FE_OFN515_n_9697), .o(TIMEBOOST_net_10548) );
na02f02 TIMEBOOST_cell_44234 ( .a(TIMEBOOST_net_14355), .b(FE_OFN1417_n_8567), .o(TIMEBOOST_net_12855) );
in01s01 g62900_u0 ( .a(FE_OFN1284_n_4097), .o(g62900_sb) );
na02s06 TIMEBOOST_cell_3225 ( .a(n_2562), .b(TIMEBOOST_net_192), .o(n_3388) );
na03s02 TIMEBOOST_cell_37583 ( .a(n_1927), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__Q), .c(FE_OFN714_n_8140), .o(TIMEBOOST_net_11030) );
na02m02 TIMEBOOST_cell_3226 ( .a(n_3503), .b(n_2308), .o(TIMEBOOST_net_193) );
in01s02 g62901_u0 ( .a(FE_OFN1322_n_6436), .o(g62901_sb) );
na02s02 TIMEBOOST_cell_43439 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__Q), .b(n_3536), .o(TIMEBOOST_net_13958) );
na03s02 TIMEBOOST_cell_34801 ( .a(n_3763), .b(g62366_sb), .c(g62366_db), .o(n_6869) );
na02s02 TIMEBOOST_cell_38414 ( .a(TIMEBOOST_net_11445), .b(g62796_sb), .o(n_5393) );
in01s02 g62902_u0 ( .a(FE_OFN1316_n_6624), .o(g62902_sb) );
na02f02 TIMEBOOST_cell_44054 ( .a(TIMEBOOST_net_14265), .b(FE_OFN1377_n_8567), .o(TIMEBOOST_net_12908) );
na02f02 TIMEBOOST_cell_3815 ( .a(TIMEBOOST_net_487), .b(g54139_da), .o(n_13362) );
na02s01 TIMEBOOST_cell_18439 ( .a(TIMEBOOST_net_4476), .b(g58369_db), .o(n_9012) );
in01s01 g62903_u0 ( .a(FE_OFN1264_n_4095), .o(g62903_sb) );
na02s01 TIMEBOOST_cell_36621 ( .a(FE_OFN1648_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__Q), .o(TIMEBOOST_net_10549) );
na03f02 TIMEBOOST_cell_45487 ( .a(n_8547), .b(n_393), .c(FE_OFN2185_n_8567), .o(TIMEBOOST_net_14982) );
na02f02 TIMEBOOST_cell_42486 ( .a(TIMEBOOST_net_13481), .b(g57157_sb), .o(n_11593) );
in01s01 g62904_u0 ( .a(FE_OFN1250_n_4093), .o(g62904_sb) );
na02f02 TIMEBOOST_cell_43722 ( .a(TIMEBOOST_net_14099), .b(FE_OFN1368_n_8567), .o(TIMEBOOST_net_12816) );
na02s01 TIMEBOOST_cell_44795 ( .a(FE_OFN219_n_9853), .b(g58046_sb), .o(TIMEBOOST_net_14636) );
na02s01 TIMEBOOST_cell_3228 ( .a(n_3783), .b(n_4671), .o(TIMEBOOST_net_194) );
in01s01 g62905_u0 ( .a(n_6287), .o(g62905_sb) );
na02f02 TIMEBOOST_cell_37127 ( .a(FE_RN_140_0), .b(n_10961), .o(TIMEBOOST_net_10802) );
na02f04 TIMEBOOST_cell_3401 ( .a(TIMEBOOST_net_280), .b(n_7092), .o(n_16325) );
na02f02 TIMEBOOST_cell_3402 ( .a(FE_RN_401_0), .b(FE_RN_403_0), .o(TIMEBOOST_net_281) );
in01s01 g62906_u0 ( .a(FE_OFN1315_n_6624), .o(g62906_sb) );
na02f02 TIMEBOOST_cell_44530 ( .a(TIMEBOOST_net_14503), .b(FE_OFN2180_n_8567), .o(TIMEBOOST_net_13458) );
na03m02 TIMEBOOST_cell_38919 ( .a(g52479_da), .b(FE_OFN1023_n_11877), .c(n_739), .o(TIMEBOOST_net_11698) );
na02s02 TIMEBOOST_cell_40392 ( .a(TIMEBOOST_net_12434), .b(g65366_db), .o(n_4252) );
in01s02 g62907_u0 ( .a(FE_OFN1248_n_4093), .o(g62907_sb) );
na02s01 TIMEBOOST_cell_3229 ( .a(TIMEBOOST_net_194), .b(g65371_da), .o(n_3531) );
na02f02 TIMEBOOST_cell_37810 ( .a(TIMEBOOST_net_11143), .b(FE_OFN2126_n_16497), .o(n_12988) );
na02s03 TIMEBOOST_cell_3230 ( .a(n_2680), .b(n_2681), .o(TIMEBOOST_net_195) );
in01s01 g62908_u0 ( .a(FE_OFN1258_n_4143), .o(g62908_sb) );
na02s01 TIMEBOOST_cell_36623 ( .a(g58050_sb), .b(g58050_db), .o(TIMEBOOST_net_10550) );
na02s02 TIMEBOOST_cell_43517 ( .a(n_3731), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__Q), .o(TIMEBOOST_net_13997) );
na02f02 TIMEBOOST_cell_44698 ( .a(TIMEBOOST_net_14587), .b(TIMEBOOST_net_6262), .o(n_9237) );
in01s01 g62909_u0 ( .a(FE_OFN1231_n_6391), .o(g62909_sb) );
na02m02 TIMEBOOST_cell_44055 ( .a(n_9113), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__Q), .o(TIMEBOOST_net_14266) );
na02s01 TIMEBOOST_cell_36625 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__Q), .b(FE_OFN207_n_9865), .o(TIMEBOOST_net_10551) );
na02s02 TIMEBOOST_cell_37812 ( .a(TIMEBOOST_net_11144), .b(g62018_sb), .o(n_7859) );
in01s01 g62910_u0 ( .a(FE_OFN1278_n_4097), .o(g62910_sb) );
na02m04 TIMEBOOST_cell_3231 ( .a(TIMEBOOST_net_195), .b(n_2461), .o(n_2991) );
na02s01 TIMEBOOST_cell_43030 ( .a(TIMEBOOST_net_13753), .b(n_4043), .o(n_5517) );
na02f02 TIMEBOOST_cell_22274 ( .a(n_9976), .b(n_10560), .o(TIMEBOOST_net_6394) );
in01s01 g62911_u0 ( .a(n_6287), .o(g62911_sb) );
na02f02 TIMEBOOST_cell_37135 ( .a(n_16253), .b(n_16248), .o(TIMEBOOST_net_10806) );
na02f02 TIMEBOOST_cell_3403 ( .a(TIMEBOOST_net_281), .b(FE_RN_402_0), .o(FE_RN_404_0) );
na02s01 TIMEBOOST_cell_16369 ( .a(TIMEBOOST_net_3441), .b(g65083_db), .o(n_3600) );
in01s01 g62912_u0 ( .a(FE_OFN1312_n_6624), .o(g62912_sb) );
na02f02 TIMEBOOST_cell_44056 ( .a(TIMEBOOST_net_14266), .b(FE_OFN1380_n_8567), .o(TIMEBOOST_net_12917) );
na02s01 TIMEBOOST_cell_39304 ( .a(TIMEBOOST_net_11890), .b(g65838_db), .o(n_1881) );
na02s01 TIMEBOOST_cell_40394 ( .a(TIMEBOOST_net_12435), .b(g61884_sb), .o(n_8062) );
in01s01 g62913_u0 ( .a(FE_OFN1212_n_4151), .o(g62913_sb) );
na02f02 TIMEBOOST_cell_36523 ( .a(n_4806), .b(n_3018), .o(TIMEBOOST_net_10500) );
na02s01 TIMEBOOST_cell_16811 ( .a(TIMEBOOST_net_3662), .b(g65334_db), .o(n_3552) );
in01s01 g62914_u0 ( .a(FE_OFN1276_n_4096), .o(g62914_sb) );
na02m04 TIMEBOOST_cell_3233 ( .a(TIMEBOOST_net_196), .b(n_2694), .o(n_3147) );
na03s02 TIMEBOOST_cell_37579 ( .a(n_2203), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__Q), .c(FE_OFN2081_n_8176), .o(TIMEBOOST_net_11028) );
na02s02 TIMEBOOST_cell_3234 ( .a(n_2427), .b(n_2431), .o(TIMEBOOST_net_197) );
in01s01 g62915_u0 ( .a(FE_OFN1204_n_4090), .o(g62915_sb) );
na02s02 TIMEBOOST_cell_36539 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__Q), .b(FE_OFN660_n_4392), .o(TIMEBOOST_net_10508) );
na02s01 TIMEBOOST_cell_42730 ( .a(TIMEBOOST_net_13603), .b(FE_OFN2256_n_8060), .o(TIMEBOOST_net_1755) );
na02s02 TIMEBOOST_cell_43138 ( .a(TIMEBOOST_net_13807), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_12119) );
in01s01 g62916_u0 ( .a(FE_OFN1193_n_6935), .o(g62916_sb) );
na02f02 TIMEBOOST_cell_3235 ( .a(n_2437), .b(TIMEBOOST_net_197), .o(n_2432) );
na02f02 TIMEBOOST_cell_45797 ( .a(n_9121), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__Q), .o(TIMEBOOST_net_15137) );
na02s01 TIMEBOOST_cell_3236 ( .a(n_3386), .b(FE_OFN197_n_2683), .o(TIMEBOOST_net_198) );
in01s01 g62917_u0 ( .a(FE_OFN1248_n_4093), .o(g62917_sb) );
na02s01 TIMEBOOST_cell_3237 ( .a(TIMEBOOST_net_198), .b(n_15762), .o(n_4533) );
na02f02 TIMEBOOST_cell_45798 ( .a(TIMEBOOST_net_15137), .b(FE_OFN1370_n_8567), .o(TIMEBOOST_net_14458) );
na02s01 TIMEBOOST_cell_3238 ( .a(g58042_sb), .b(g58054_db), .o(TIMEBOOST_net_199) );
in01s01 g62918_u0 ( .a(FE_OFN1248_n_4093), .o(g62918_sb) );
na02s01 TIMEBOOST_cell_3239 ( .a(TIMEBOOST_net_199), .b(FE_OFN229_n_9120), .o(n_9092) );
na02s02 TIMEBOOST_cell_39307 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__Q), .b(g58287_sb), .o(TIMEBOOST_net_11892) );
no02f02 TIMEBOOST_cell_22365 ( .a(TIMEBOOST_net_6439), .b(n_13564), .o(g53012_p) );
in01s01 g62919_u0 ( .a(n_6554), .o(g62919_sb) );
no03f02 TIMEBOOST_cell_37131 ( .a(FE_RN_843_0), .b(FE_RN_845_0), .c(FE_RN_844_0), .o(TIMEBOOST_net_10804) );
na02s01 g66422_u2 ( .a(parchk_pci_ad_reg_in_1233), .b(FE_OFN795_n_2520), .o(g66422_db) );
na02s01 TIMEBOOST_cell_3406 ( .a(FE_OFN211_n_9858), .b(g58110_sb), .o(TIMEBOOST_net_283) );
in01s01 g62920_u0 ( .a(FE_OFN1226_n_6391), .o(g62920_sb) );
na02f02 TIMEBOOST_cell_4069 ( .a(TIMEBOOST_net_614), .b(n_13828), .o(n_14087) );
na02s01 TIMEBOOST_cell_37573 ( .a(parchk_pci_ad_reg_in_1230), .b(g65893_sb), .o(TIMEBOOST_net_11025) );
na02s01 TIMEBOOST_cell_3242 ( .a(FE_OFN201_n_9230), .b(g58268_sb), .o(TIMEBOOST_net_201) );
in01s01 g62921_u0 ( .a(n_6232), .o(g62921_sb) );
na02s01 TIMEBOOST_cell_44883 ( .a(FE_OFN1678_n_4655), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__Q), .o(TIMEBOOST_net_14680) );
na02s01 TIMEBOOST_cell_3407 ( .a(TIMEBOOST_net_283), .b(g58110_db), .o(n_9684) );
na02s01 TIMEBOOST_cell_3408 ( .a(FE_OFN213_n_9124), .b(g58111_sb), .o(TIMEBOOST_net_284) );
in01s01 g62922_u0 ( .a(FE_OFN1244_n_4092), .o(g62922_sb) );
na02s02 TIMEBOOST_cell_42076 ( .a(TIMEBOOST_net_13276), .b(n_6287), .o(TIMEBOOST_net_11580) );
na02s01 TIMEBOOST_cell_42851 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__Q), .b(n_1868), .o(TIMEBOOST_net_13664) );
na02f02 TIMEBOOST_cell_36954 ( .a(TIMEBOOST_net_10715), .b(g58808_sb), .o(n_8633) );
in01s01 g62923_u0 ( .a(FE_OFN1272_n_4096), .o(g62923_sb) );
na02s01 TIMEBOOST_cell_3243 ( .a(TIMEBOOST_net_201), .b(g58268_db), .o(n_9219) );
na02s02 TIMEBOOST_cell_37561 ( .a(pci_target_unit_pcit_if_strd_addr_in_710), .b(g52639_sb), .o(TIMEBOOST_net_11019) );
na02s01 TIMEBOOST_cell_3244 ( .a(FE_OFN203_n_9228), .b(g58269_sb), .o(TIMEBOOST_net_202) );
in01s01 g62924_u0 ( .a(n_6645), .o(g62924_sb) );
na02s01 TIMEBOOST_cell_44884 ( .a(TIMEBOOST_net_14680), .b(n_4482), .o(TIMEBOOST_net_10981) );
na02s01 TIMEBOOST_cell_3409 ( .a(TIMEBOOST_net_284), .b(g58111_db), .o(n_9077) );
na02s01 TIMEBOOST_cell_9728 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__Q), .b(g65913_sb), .o(TIMEBOOST_net_1431) );
in01s01 g62925_u0 ( .a(FE_OFN1192_n_6935), .o(g62925_sb) );
na02s01 TIMEBOOST_cell_3245 ( .a(TIMEBOOST_net_202), .b(g58269_db), .o(n_9218) );
na02s01 g62925_u2 ( .a(n_4261), .b(FE_OFN1192_n_6935), .o(g62925_db) );
na02f02 TIMEBOOST_cell_45488 ( .a(TIMEBOOST_net_14982), .b(g58609_sb), .o(n_8898) );
in01s01 g62926_u0 ( .a(n_6232), .o(g62926_sb) );
in01s01 TIMEBOOST_cell_45941 ( .a(wbm_dat_i_29_), .o(TIMEBOOST_net_15248) );
na02s01 TIMEBOOST_cell_9729 ( .a(TIMEBOOST_net_1431), .b(g65913_db), .o(n_1853) );
na02s01 TIMEBOOST_cell_43499 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__Q), .b(n_3682), .o(TIMEBOOST_net_13988) );
in01s01 g62927_u0 ( .a(FE_OFN1244_n_4092), .o(g62927_sb) );
na02m02 TIMEBOOST_cell_43789 ( .a(n_9074), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__Q), .o(TIMEBOOST_net_14133) );
na02s01 TIMEBOOST_cell_42852 ( .a(TIMEBOOST_net_13664), .b(FE_OFN720_n_8060), .o(TIMEBOOST_net_11245) );
na02f02 TIMEBOOST_cell_36956 ( .a(TIMEBOOST_net_10716), .b(g58821_sb), .o(n_8620) );
in01s01 g62928_u0 ( .a(FE_OFN1202_n_4090), .o(g62928_sb) );
na02s01 TIMEBOOST_cell_40853 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__Q), .b(n_13106), .o(TIMEBOOST_net_12665) );
na02f02 TIMEBOOST_cell_44722 ( .a(TIMEBOOST_net_14599), .b(FE_OFN1600_n_13995), .o(n_14493) );
na02s02 TIMEBOOST_cell_40688 ( .a(TIMEBOOST_net_12582), .b(g62665_sb), .o(n_6208) );
in01s01 g62929_u0 ( .a(FE_OFN1248_n_4093), .o(g62929_sb) );
na02s01 TIMEBOOST_cell_3249 ( .a(TIMEBOOST_net_204), .b(n_4473), .o(n_4485) );
na03s02 TIMEBOOST_cell_37537 ( .a(TIMEBOOST_net_3804), .b(g65909_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__Q), .o(TIMEBOOST_net_11007) );
na02s01 TIMEBOOST_cell_40839 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__Q), .b(n_13164), .o(TIMEBOOST_net_12658) );
in01s01 g62930_u0 ( .a(FE_OFN1264_n_4095), .o(g62930_sb) );
na02s01 TIMEBOOST_cell_39187 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__Q), .b(g65851_sb), .o(TIMEBOOST_net_11832) );
na02s02 TIMEBOOST_cell_42853 ( .a(n_1571), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__Q), .o(TIMEBOOST_net_13665) );
na02f02 TIMEBOOST_cell_36958 ( .a(TIMEBOOST_net_10717), .b(g58834_sb), .o(n_8603) );
in01s01 g62931_u0 ( .a(FE_OFN1235_n_6391), .o(g62931_sb) );
na02s01 TIMEBOOST_cell_42587 ( .a(g58026_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__Q), .o(TIMEBOOST_net_13532) );
na02s01 TIMEBOOST_cell_18581 ( .a(TIMEBOOST_net_4547), .b(g63112_sb), .o(n_5031) );
na02f02 TIMEBOOST_cell_41664 ( .a(TIMEBOOST_net_13070), .b(FE_OFN2158_n_16439), .o(TIMEBOOST_net_11738) );
in01s01 g62932_u0 ( .a(FE_OFN1283_n_4097), .o(g62932_sb) );
na02f02 TIMEBOOST_cell_43790 ( .a(TIMEBOOST_net_14133), .b(FE_OFN1413_n_8567), .o(TIMEBOOST_net_12982) );
na02s02 TIMEBOOST_cell_42854 ( .a(TIMEBOOST_net_13665), .b(FE_OFN2212_n_8407), .o(TIMEBOOST_net_11244) );
na02f02 TIMEBOOST_cell_36960 ( .a(TIMEBOOST_net_10718), .b(g58827_sb), .o(n_8613) );
in01s01 g62933_u0 ( .a(FE_OFN1276_n_4096), .o(g62933_sb) );
na02s02 TIMEBOOST_cell_40832 ( .a(TIMEBOOST_net_12654), .b(FE_OFN1331_n_13547), .o(TIMEBOOST_net_11603) );
na02s02 TIMEBOOST_cell_37563 ( .a(pci_target_unit_pcit_if_strd_addr_in_709), .b(g52638_sb), .o(TIMEBOOST_net_11020) );
na02s01 TIMEBOOST_cell_41736 ( .a(TIMEBOOST_net_13106), .b(g65272_da), .o(n_4292) );
in01s01 g62934_u0 ( .a(FE_OFN1275_n_4096), .o(g62934_sb) );
na02s02 TIMEBOOST_cell_3253 ( .a(TIMEBOOST_net_206), .b(n_2329), .o(n_8448) );
na02s01 TIMEBOOST_cell_37565 ( .a(g65893_sb), .b(parchk_pci_ad_reg_in_1226), .o(TIMEBOOST_net_11021) );
na03f02 TIMEBOOST_cell_36050 ( .a(FE_OCP_RBN1962_FE_OFN1591_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__Q), .c(n_13888), .o(n_14268) );
in01s01 g62935_u0 ( .a(FE_OFN1276_n_4096), .o(g62935_sb) );
na02s02 TIMEBOOST_cell_45708 ( .a(TIMEBOOST_net_15092), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_12582) );
na02f04 TIMEBOOST_cell_38800 ( .a(TIMEBOOST_net_11638), .b(FE_OFN2185_n_8567), .o(TIMEBOOST_net_10691) );
na02m02 TIMEBOOST_cell_3256 ( .a(n_16474), .b(n_7114), .o(TIMEBOOST_net_208) );
in01s01 g62936_u0 ( .a(FE_OFN1234_n_6391), .o(g62936_sb) );
na02s01 TIMEBOOST_cell_36307 ( .a(parchk_pci_ad_reg_in_1207), .b(g67073_db), .o(TIMEBOOST_net_10392) );
na02m02 TIMEBOOST_cell_3521 ( .a(TIMEBOOST_net_340), .b(n_3413), .o(n_4894) );
na02s02 TIMEBOOST_cell_3522 ( .a(n_3391), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_341) );
in01s01 g62937_u0 ( .a(FE_OFN1194_n_6935), .o(g62937_sb) );
na02m02 TIMEBOOST_cell_44057 ( .a(n_9584), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__Q), .o(TIMEBOOST_net_14267) );
na03s02 TIMEBOOST_cell_37535 ( .a(TIMEBOOST_net_3789), .b(g65969_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__Q), .o(TIMEBOOST_net_11006) );
na02f06 TIMEBOOST_cell_3258 ( .a(FE_RN_528_0), .b(FE_RN_527_0), .o(TIMEBOOST_net_209) );
in01s01 g62938_u0 ( .a(FE_OFN1236_n_6391), .o(g62938_sb) );
na02s01 TIMEBOOST_cell_42588 ( .a(TIMEBOOST_net_13532), .b(g58026_db), .o(TIMEBOOST_net_12427) );
na03s02 TIMEBOOST_cell_37567 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__Q), .b(FE_OFN1803_n_9690), .c(FE_OFN243_n_9116), .o(TIMEBOOST_net_11022) );
na02s01 TIMEBOOST_cell_42855 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__Q), .b(n_2178), .o(TIMEBOOST_net_13666) );
in01s01 g62939_u0 ( .a(n_6431), .o(g62939_sb) );
na02f02 TIMEBOOST_cell_12552 ( .a(g75418_da), .b(g75418_db), .o(TIMEBOOST_net_2843) );
na02m02 TIMEBOOST_cell_38834 ( .a(TIMEBOOST_net_11655), .b(g58840_sb), .o(n_8674) );
na02s02 TIMEBOOST_cell_40549 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_), .b(n_1678), .o(TIMEBOOST_net_12513) );
in01s01 g62940_u0 ( .a(FE_OFN1289_n_4098), .o(g62940_sb) );
na02s02 TIMEBOOST_cell_43500 ( .a(TIMEBOOST_net_13988), .b(FE_OFN1234_n_6391), .o(TIMEBOOST_net_12194) );
na02f02 TIMEBOOST_cell_36962 ( .a(TIMEBOOST_net_10719), .b(g58806_sb), .o(n_8635) );
na02f02 TIMEBOOST_cell_42829 ( .a(TIMEBOOST_net_9664), .b(g54326_sb), .o(TIMEBOOST_net_13653) );
in01s01 g62941_u0 ( .a(FE_OFN1233_n_6391), .o(g62941_sb) );
na02f02 TIMEBOOST_cell_44610 ( .a(TIMEBOOST_net_14543), .b(FE_OFN2190_n_8567), .o(TIMEBOOST_net_12995) );
na02f02 TIMEBOOST_cell_36928 ( .a(TIMEBOOST_net_10702), .b(g52611_sb), .o(n_10190) );
na04s02 TIMEBOOST_cell_34238 ( .a(g64349_da), .b(g64349_db), .c(g63117_sb), .d(g63117_db), .o(n_7117) );
in01s01 g62942_u0 ( .a(FE_OFN1222_n_6391), .o(g62942_sb) );
na02f06 TIMEBOOST_cell_3259 ( .a(TIMEBOOST_net_209), .b(FE_RN_529_0), .o(FE_OFN1060_n_16720) );
na02s02 TIMEBOOST_cell_43376 ( .a(TIMEBOOST_net_13926), .b(n_6431), .o(TIMEBOOST_net_12157) );
na02s01 TIMEBOOST_cell_3260 ( .a(n_3764), .b(n_4671), .o(TIMEBOOST_net_210) );
in01s01 g62943_u0 ( .a(FE_OFN1283_n_4097), .o(g62943_sb) );
no02s02 TIMEBOOST_cell_44769 ( .a(n_564), .b(n_2263), .o(TIMEBOOST_net_14623) );
na02s01 TIMEBOOST_cell_36347 ( .a(parchk_pci_ad_reg_in_1220), .b(g67071_db), .o(TIMEBOOST_net_10412) );
na02s01 TIMEBOOST_cell_36346 ( .a(TIMEBOOST_net_10411), .b(g66399_sb), .o(n_2543) );
in01s01 g62944_u0 ( .a(FE_OFN1264_n_4095), .o(g62944_sb) );
na02m02 TIMEBOOST_cell_43791 ( .a(n_9773), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__Q), .o(TIMEBOOST_net_14134) );
na02s02 TIMEBOOST_cell_42826 ( .a(TIMEBOOST_net_13651), .b(g58303_db), .o(n_9027) );
na02f02 TIMEBOOST_cell_36930 ( .a(TIMEBOOST_net_10703), .b(FE_OFN2200_n_10256), .o(n_10277) );
in01s01 g62945_u0 ( .a(FE_OFN1234_n_6391), .o(g62945_sb) );
na02f02 TIMEBOOST_cell_44058 ( .a(TIMEBOOST_net_14267), .b(FE_OFN1385_n_8567), .o(TIMEBOOST_net_13379) );
na02s02 TIMEBOOST_cell_43440 ( .a(TIMEBOOST_net_13958), .b(FE_OFN1230_n_6391), .o(TIMEBOOST_net_12632) );
na02s01 TIMEBOOST_cell_39262 ( .a(TIMEBOOST_net_11869), .b(g64150_db), .o(n_4015) );
in01s01 g62946_u0 ( .a(FE_OFN1243_n_4092), .o(g62946_sb) );
na02f02 TIMEBOOST_cell_43792 ( .a(TIMEBOOST_net_14134), .b(FE_OFN1388_n_8567), .o(TIMEBOOST_net_12898) );
na02s01 TIMEBOOST_cell_32186 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__Q), .b(n_13176), .o(TIMEBOOST_net_10004) );
na02s01 TIMEBOOST_cell_39214 ( .a(TIMEBOOST_net_11845), .b(n_1653), .o(TIMEBOOST_net_11474) );
in01s01 g62947_u0 ( .a(FE_OFN1315_n_6624), .o(g62947_sb) );
na02m02 TIMEBOOST_cell_44059 ( .a(n_9583), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__Q), .o(TIMEBOOST_net_14268) );
na02m02 TIMEBOOST_cell_10551 ( .a(TIMEBOOST_net_1842), .b(FE_OFN1085_n_13221), .o(TIMEBOOST_net_569) );
na02s02 TIMEBOOST_cell_10553 ( .a(TIMEBOOST_net_1843), .b(FE_OFN1083_n_13221), .o(TIMEBOOST_net_878) );
in01s01 g62948_u0 ( .a(FE_OFN1312_n_6624), .o(g62948_sb) );
na02f02 TIMEBOOST_cell_44060 ( .a(TIMEBOOST_net_14268), .b(FE_OFN1384_n_8567), .o(TIMEBOOST_net_12830) );
na02s02 TIMEBOOST_cell_18519 ( .a(TIMEBOOST_net_4516), .b(g62824_sb), .o(n_5330) );
na02f02 TIMEBOOST_cell_22586 ( .a(n_14384), .b(n_14087), .o(TIMEBOOST_net_6550) );
in01s01 g62949_u0 ( .a(FE_OFN1293_n_4098), .o(g62949_sb) );
na02s01 TIMEBOOST_cell_39189 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__22__Q), .b(n_8176), .o(TIMEBOOST_net_11833) );
na02s01 TIMEBOOST_cell_32184 ( .a(configuration_sync_command_bit2), .b(wbu_wb_init_complete_in), .o(TIMEBOOST_net_10003) );
na02m02 TIMEBOOST_cell_32183 ( .a(n_3482), .b(TIMEBOOST_net_10002), .o(n_14810) );
in01s01 g62950_u0 ( .a(FE_OFN1243_n_4092), .o(g62950_sb) );
na02f02 TIMEBOOST_cell_43793 ( .a(TIMEBOOST_net_10047), .b(g57143_sb), .o(TIMEBOOST_net_14135) );
na03s02 TIMEBOOST_cell_37859 ( .a(FE_OFN262_n_9851), .b(FE_OFN1690_n_9528), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__Q), .o(TIMEBOOST_net_11168) );
no02m04 TIMEBOOST_cell_32181 ( .a(FE_OFN1706_n_4868), .b(TIMEBOOST_net_10001), .o(TIMEBOOST_net_5288) );
in01s01 g62951_u0 ( .a(FE_OFN1272_n_4096), .o(g62951_sb) );
na02s01 TIMEBOOST_cell_3261 ( .a(TIMEBOOST_net_210), .b(g65325_da), .o(n_3558) );
na02s01 TIMEBOOST_cell_44796 ( .a(TIMEBOOST_net_14636), .b(g58046_db), .o(n_9744) );
na02s01 TIMEBOOST_cell_3262 ( .a(n_3780), .b(n_4677), .o(TIMEBOOST_net_211) );
in01s01 g62952_u0 ( .a(FE_OFN1260_n_4143), .o(g62952_sb) );
na02f02 TIMEBOOST_cell_43794 ( .a(TIMEBOOST_net_14135), .b(FE_OFN1415_n_8567), .o(n_11606) );
no02m04 TIMEBOOST_cell_32180 ( .a(n_13784), .b(FE_RN_396_0), .o(TIMEBOOST_net_10001) );
na02s01 TIMEBOOST_cell_37421 ( .a(wbu_latency_tim_val_in_243), .b(n_6986), .o(TIMEBOOST_net_10949) );
in01s01 g62953_u0 ( .a(FE_OFN2063_n_6391), .o(g62953_sb) );
na02s01 TIMEBOOST_cell_36357 ( .a(pci_target_unit_del_sync_addr_in_213), .b(g66414_db), .o(TIMEBOOST_net_10417) );
na02m02 TIMEBOOST_cell_44345 ( .a(n_9087), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__Q), .o(TIMEBOOST_net_14411) );
na02m02 TIMEBOOST_cell_39176 ( .a(g53892_db), .b(TIMEBOOST_net_11826), .o(TIMEBOOST_net_10573) );
in01s01 g62954_u0 ( .a(FE_OFN1295_n_4098), .o(g62954_sb) );
na02m02 TIMEBOOST_cell_43795 ( .a(n_9009), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__Q), .o(TIMEBOOST_net_14136) );
na02s01 TIMEBOOST_cell_37420 ( .a(TIMEBOOST_net_10948), .b(g60671_sb), .o(TIMEBOOST_net_857) );
na02s01 TIMEBOOST_cell_36717 ( .a(g61962_sb), .b(g61962_db), .o(TIMEBOOST_net_10597) );
in01s01 g62955_u0 ( .a(FE_OFN1312_n_6624), .o(g62955_sb) );
na02m02 TIMEBOOST_cell_44061 ( .a(n_9651), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__Q), .o(TIMEBOOST_net_14269) );
na02s01 TIMEBOOST_cell_38416 ( .a(TIMEBOOST_net_11446), .b(g63397_sb), .o(n_4130) );
na02s02 TIMEBOOST_cell_39946 ( .a(TIMEBOOST_net_12211), .b(g62454_sb), .o(n_6689) );
in01s01 g62956_u0 ( .a(FE_OFN1313_n_6624), .o(g62956_sb) );
na02f02 TIMEBOOST_cell_44062 ( .a(TIMEBOOST_net_14269), .b(FE_OFN1405_n_8567), .o(TIMEBOOST_net_12829) );
na02s01 TIMEBOOST_cell_39419 ( .a(conf_wb_err_addr_in_950), .b(configuration_wb_err_addr_541), .o(TIMEBOOST_net_11948) );
na02s01 TIMEBOOST_cell_40396 ( .a(TIMEBOOST_net_12436), .b(g61872_sb), .o(n_8089) );
in01s01 g62957_u0 ( .a(FE_OFN1250_n_4093), .o(g62957_sb) );
na02s01 TIMEBOOST_cell_3263 ( .a(TIMEBOOST_net_211), .b(g65411_da), .o(n_3515) );
na03s02 TIMEBOOST_cell_37539 ( .a(TIMEBOOST_net_3791), .b(g65732_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__Q), .o(TIMEBOOST_net_11008) );
na02s01 TIMEBOOST_cell_39219 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__Q), .b(n_8232), .o(TIMEBOOST_net_11848) );
in01s01 g62958_u0 ( .a(FE_OFN1294_n_4098), .o(g62958_sb) );
na02f02 TIMEBOOST_cell_38899 ( .a(n_4708), .b(wbu_addr_in_275), .o(TIMEBOOST_net_11688) );
na02s02 TIMEBOOST_cell_36716 ( .a(TIMEBOOST_net_10596), .b(g63595_sb), .o(n_4773) );
na02s01 TIMEBOOST_cell_36719 ( .a(g61885_sb), .b(g61989_db), .o(TIMEBOOST_net_10598) );
in01s01 g62959_u0 ( .a(FE_OFN1294_n_4098), .o(g62959_sb) );
no03f02 TIMEBOOST_cell_37137 ( .a(FE_RN_831_0), .b(FE_RN_832_0), .c(FE_RN_833_0), .o(TIMEBOOST_net_10807) );
na02s02 TIMEBOOST_cell_36718 ( .a(TIMEBOOST_net_10597), .b(g63601_sb), .o(TIMEBOOST_net_9825) );
na02s01 TIMEBOOST_cell_36721 ( .a(g61880_sb), .b(g61983_db), .o(TIMEBOOST_net_10599) );
in01s01 g62960_u0 ( .a(FE_OFN1323_n_6436), .o(g62960_sb) );
na02m02 TIMEBOOST_cell_44063 ( .a(n_9042), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__Q), .o(TIMEBOOST_net_14270) );
na02s02 TIMEBOOST_cell_10545 ( .a(TIMEBOOST_net_1839), .b(FE_OFN1085_n_13221), .o(TIMEBOOST_net_563) );
na02s01 TIMEBOOST_cell_10245 ( .a(TIMEBOOST_net_1689), .b(g64136_sb), .o(n_4026) );
in01s01 g62961_u0 ( .a(FE_OFN1312_n_6624), .o(g62961_sb) );
na02s02 TIMEBOOST_cell_37962 ( .a(TIMEBOOST_net_11219), .b(g58240_sb), .o(n_9551) );
na02f02 TIMEBOOST_cell_43738 ( .a(TIMEBOOST_net_14107), .b(FE_OFN1423_n_8567), .o(TIMEBOOST_net_12698) );
na02s02 TIMEBOOST_cell_19287 ( .a(TIMEBOOST_net_4900), .b(g60647_sb), .o(n_5679) );
in01s01 g62962_u0 ( .a(FE_OFN1293_n_4098), .o(g62962_sb) );
na02s01 TIMEBOOST_cell_38418 ( .a(TIMEBOOST_net_11447), .b(g62836_sb), .o(n_5300) );
na02s02 TIMEBOOST_cell_36720 ( .a(TIMEBOOST_net_10598), .b(g63618_sb), .o(TIMEBOOST_net_9824) );
na02f02 TIMEBOOST_cell_44064 ( .a(TIMEBOOST_net_14270), .b(FE_OFN1401_n_8567), .o(TIMEBOOST_net_12764) );
in01s01 g62963_u0 ( .a(FE_OFN1223_n_6391), .o(g62963_sb) );
na02s02 TIMEBOOST_cell_39264 ( .a(TIMEBOOST_net_11870), .b(n_4476), .o(n_4238) );
na03s02 TIMEBOOST_cell_37533 ( .a(TIMEBOOST_net_3802), .b(g65773_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__Q), .o(TIMEBOOST_net_11005) );
na02s01 TIMEBOOST_cell_37988 ( .a(TIMEBOOST_net_11232), .b(g61812_sb), .o(n_7887) );
in01s01 g62964_u0 ( .a(n_6287), .o(g62964_sb) );
no03f06 TIMEBOOST_cell_36297 ( .a(FE_RN_686_0), .b(n_2864), .c(n_436), .o(TIMEBOOST_net_10387) );
na02s01 TIMEBOOST_cell_40524 ( .a(TIMEBOOST_net_12500), .b(FE_OFN1300_n_5763), .o(TIMEBOOST_net_11515) );
na02s01 TIMEBOOST_cell_3416 ( .a(FE_OFN221_n_9846), .b(g58118_sb), .o(TIMEBOOST_net_288) );
in01s01 g62965_u0 ( .a(FE_OFN1270_n_4095), .o(g62965_sb) );
na02s01 TIMEBOOST_cell_36501 ( .a(pci_target_unit_del_sync_addr_in_227), .b(g66424_db), .o(TIMEBOOST_net_10489) );
na02f02 TIMEBOOST_cell_38806 ( .a(TIMEBOOST_net_11641), .b(FE_OFN2187_n_8567), .o(n_11634) );
na02f04 TIMEBOOST_cell_32169 ( .a(n_16322), .b(TIMEBOOST_net_9995), .o(TIMEBOOST_net_6374) );
in01s01 g62966_u0 ( .a(FE_OFN1226_n_6391), .o(g62966_sb) );
na02f02 TIMEBOOST_cell_3267 ( .a(TIMEBOOST_net_213), .b(FE_RN_356_0), .o(n_5747) );
na02s01 TIMEBOOST_cell_36631 ( .a(TIMEBOOST_net_269), .b(g61797_sb), .o(TIMEBOOST_net_10554) );
na02s01 TIMEBOOST_cell_31401 ( .a(TIMEBOOST_net_9611), .b(n_4450), .o(n_4339) );
in01s01 g62967_u0 ( .a(FE_OFN1323_n_6436), .o(g62967_sb) );
na02m02 TIMEBOOST_cell_44065 ( .a(n_9065), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__Q), .o(TIMEBOOST_net_14271) );
na03s02 TIMEBOOST_cell_39491 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__Q), .b(FE_OFN1128_g64577_p), .c(n_4524), .o(TIMEBOOST_net_11984) );
na02s02 TIMEBOOST_cell_38420 ( .a(TIMEBOOST_net_11448), .b(g63105_sb), .o(n_5044) );
in01s02 g62968_u0 ( .a(FE_OFN1317_n_6624), .o(g62968_sb) );
na02f02 TIMEBOOST_cell_44066 ( .a(TIMEBOOST_net_14271), .b(FE_OFN1401_n_8567), .o(TIMEBOOST_net_12765) );
na02s02 TIMEBOOST_cell_10557 ( .a(TIMEBOOST_net_1845), .b(g52879_sb), .o(TIMEBOOST_net_889) );
na02s01 TIMEBOOST_cell_43096 ( .a(TIMEBOOST_net_13786), .b(FE_OFN1225_n_6391), .o(TIMEBOOST_net_12058) );
in01s01 g62969_u0 ( .a(n_6287), .o(g62969_sb) );
na02s01 TIMEBOOST_cell_36303 ( .a(parchk_pci_ad_reg_in_1224), .b(g67041_db), .o(TIMEBOOST_net_10390) );
na02f02 TIMEBOOST_cell_37034 ( .a(TIMEBOOST_net_10755), .b(FE_OFN1774_n_13800), .o(g74872_p) );
na02s01 TIMEBOOST_cell_3418 ( .a(FE_OFN231_n_9839), .b(g58124_sb), .o(TIMEBOOST_net_289) );
in01s01 g62970_u0 ( .a(FE_OFN1257_n_4143), .o(g62970_sb) );
na02s01 TIMEBOOST_cell_36553 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__Q), .b(g58391_sb), .o(TIMEBOOST_net_10515) );
na02m04 TIMEBOOST_cell_32168 ( .a(n_440), .b(n_46), .o(TIMEBOOST_net_9995) );
na02s01 TIMEBOOST_cell_32028 ( .a(configuration_pci_err_data_529), .b(wbm_dat_o_28_), .o(TIMEBOOST_net_9925) );
in01s01 g62971_u0 ( .a(FE_OFN1234_n_6391), .o(g62971_sb) );
na02m02 TIMEBOOST_cell_44067 ( .a(n_9036), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q), .o(TIMEBOOST_net_14272) );
na02s02 TIMEBOOST_cell_42679 ( .a(n_3777), .b(g65094_sb), .o(TIMEBOOST_net_13578) );
na02m02 TIMEBOOST_cell_32500 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__Q), .o(TIMEBOOST_net_10161) );
in01s01 g62972_u0 ( .a(FE_OFN1218_n_6886), .o(g62972_sb) );
na02s01 TIMEBOOST_cell_36633 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(g63547_sb), .o(TIMEBOOST_net_10555) );
na02s02 TIMEBOOST_cell_32027 ( .a(TIMEBOOST_net_9924), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_4906) );
na02s01 TIMEBOOST_cell_32026 ( .a(configuration_pci_err_data_526), .b(wbm_dat_o_25_), .o(TIMEBOOST_net_9924) );
in01s01 g62973_u0 ( .a(n_6232), .o(g62973_sb) );
na02s02 TIMEBOOST_cell_43441 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__Q), .b(n_3513), .o(TIMEBOOST_net_13959) );
na02s02 TIMEBOOST_cell_3419 ( .a(TIMEBOOST_net_289), .b(g58124_db), .o(n_9669) );
na02s01 TIMEBOOST_cell_3420 ( .a(FE_OFN233_n_9876), .b(g58125_sb), .o(TIMEBOOST_net_290) );
in01s01 g62974_u0 ( .a(FE_OFN1213_n_4151), .o(g62974_sb) );
na02s01 TIMEBOOST_cell_36635 ( .a(wbs_we_i), .b(g63588_sb), .o(TIMEBOOST_net_10556) );
na02f02 TIMEBOOST_cell_44700 ( .a(TIMEBOOST_net_14588), .b(g54472_sb), .o(n_13618) );
in01s01 g62975_u0 ( .a(FE_OFN1230_n_6391), .o(g62975_sb) );
na02s02 TIMEBOOST_cell_43256 ( .a(TIMEBOOST_net_13866), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_12044) );
na02s04 TIMEBOOST_cell_44756 ( .a(TIMEBOOST_net_14616), .b(n_1409), .o(TIMEBOOST_net_10817) );
na03s02 TIMEBOOST_cell_38041 ( .a(g65376_da), .b(g65376_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__Q), .o(TIMEBOOST_net_11259) );
in01s01 g62976_u0 ( .a(FE_OFN1285_n_4097), .o(g62976_sb) );
na02f02 TIMEBOOST_cell_36637 ( .a(n_3115), .b(configuration_icr_bit2_0), .o(TIMEBOOST_net_10557) );
na02s02 TIMEBOOST_cell_44835 ( .a(FE_OFN640_n_4669), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__Q), .o(TIMEBOOST_net_14656) );
na02s01 TIMEBOOST_cell_37912 ( .a(TIMEBOOST_net_11194), .b(g58140_sb), .o(n_9655) );
in01s01 g62977_u0 ( .a(FE_OFN1236_n_6391), .o(g62977_sb) );
na02f02 TIMEBOOST_cell_44068 ( .a(TIMEBOOST_net_14272), .b(FE_OFN1391_n_8567), .o(TIMEBOOST_net_12755) );
na03f02 TIMEBOOST_cell_45489 ( .a(n_8553), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__Q), .c(FE_OFN2184_n_8567), .o(TIMEBOOST_net_14983) );
na02f02 TIMEBOOST_cell_44214 ( .a(TIMEBOOST_net_14345), .b(FE_OFN1380_n_8567), .o(TIMEBOOST_net_12886) );
in01s01 g62978_u0 ( .a(n_6232), .o(g62978_sb) );
na02s01 g65679_u3 ( .a(g65679_da), .b(g65679_db), .o(n_1956) );
na02s01 TIMEBOOST_cell_3421 ( .a(TIMEBOOST_net_290), .b(g58125_db), .o(n_9668) );
na02f02 TIMEBOOST_cell_44392 ( .a(TIMEBOOST_net_14434), .b(FE_OFN1414_n_8567), .o(TIMEBOOST_net_12725) );
in01s01 g62979_u0 ( .a(n_6319), .o(g62979_sb) );
na02s02 TIMEBOOST_cell_43442 ( .a(TIMEBOOST_net_13959), .b(FE_OFN1234_n_6391), .o(TIMEBOOST_net_12181) );
na02s01 TIMEBOOST_cell_3423 ( .a(TIMEBOOST_net_291), .b(FE_OFN254_n_9825), .o(n_9659) );
na02s01 TIMEBOOST_cell_44852 ( .a(TIMEBOOST_net_14664), .b(g64762_db), .o(n_4491) );
in01s01 g62980_u0 ( .a(FE_OFN1231_n_6391), .o(g62980_sb) );
na02s01 TIMEBOOST_cell_39430 ( .a(TIMEBOOST_net_11953), .b(g61999_sb), .o(n_7897) );
na02s01 TIMEBOOST_cell_36639 ( .a(pci_target_unit_pcit_if_strd_addr_in_712), .b(g52641_sb), .o(TIMEBOOST_net_10558) );
na02s01 TIMEBOOST_cell_15799 ( .a(TIMEBOOST_net_3156), .b(g67049_sb), .o(n_1429) );
in01s01 g62981_u0 ( .a(FE_OFN1236_n_6391), .o(g62981_sb) );
na02m02 TIMEBOOST_cell_44069 ( .a(n_9790), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__Q), .o(TIMEBOOST_net_14273) );
na02m02 TIMEBOOST_cell_44531 ( .a(n_9405), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__8__Q), .o(TIMEBOOST_net_14504) );
na02f02 TIMEBOOST_cell_45490 ( .a(TIMEBOOST_net_14983), .b(g58595_sb), .o(n_8957) );
in01s01 g62982_u0 ( .a(FE_OFN1231_n_6391), .o(g62982_sb) );
na02f02 TIMEBOOST_cell_44070 ( .a(TIMEBOOST_net_14273), .b(FE_OFN1400_n_8567), .o(TIMEBOOST_net_12713) );
na02s01 TIMEBOOST_cell_36525 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__Q), .b(FE_OFN1795_n_9904), .o(TIMEBOOST_net_10501) );
na02s01 TIMEBOOST_cell_44855 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__Q), .b(FE_OFN580_n_9531), .o(TIMEBOOST_net_14666) );
in01s02 g62983_u0 ( .a(FE_OFN1311_n_6624), .o(g62983_sb) );
na02f02 TIMEBOOST_cell_44532 ( .a(TIMEBOOST_net_14504), .b(FE_OFN1427_n_8567), .o(TIMEBOOST_net_13498) );
na02s01 TIMEBOOST_cell_38422 ( .a(TIMEBOOST_net_11449), .b(g63436_sb), .o(n_4623) );
na02s01 TIMEBOOST_cell_38562 ( .a(TIMEBOOST_net_11519), .b(g62036_sb), .o(n_7780) );
in01s01 g62984_u0 ( .a(FE_OFN1219_n_6886), .o(g62984_sb) );
na02s01 TIMEBOOST_cell_36397 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(g65745_sb), .o(TIMEBOOST_net_10437) );
na02s02 TIMEBOOST_cell_38070 ( .a(TIMEBOOST_net_11273), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_4687) );
na02s01 TIMEBOOST_cell_31914 ( .a(FE_OFN203_n_9228), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q), .o(TIMEBOOST_net_9868) );
in01s01 g62985_u0 ( .a(FE_OFN1230_n_6391), .o(g62985_sb) );
na02m02 TIMEBOOST_cell_44071 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q), .b(n_9214), .o(TIMEBOOST_net_14274) );
na02s02 TIMEBOOST_cell_3539 ( .a(TIMEBOOST_net_349), .b(FE_OFN258_n_9862), .o(n_9722) );
na02s01 TIMEBOOST_cell_3540 ( .a(n_2313), .b(n_2314), .o(TIMEBOOST_net_350) );
in01s01 g62986_u0 ( .a(FE_OFN1207_n_6356), .o(g62986_sb) );
na02m02 TIMEBOOST_cell_44335 ( .a(n_9596), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q), .o(TIMEBOOST_net_14406) );
in01s01 TIMEBOOST_cell_45909 ( .a(wbm_dat_i_14_), .o(TIMEBOOST_net_15216) );
na02s02 TIMEBOOST_cell_37914 ( .a(TIMEBOOST_net_11195), .b(g58001_sb), .o(n_9791) );
in01s01 g62987_u0 ( .a(FE_OFN1230_n_6391), .o(g62987_sb) );
na03s02 TIMEBOOST_cell_5438 ( .a(n_3747), .b(g65076_sb), .c(g65076_db), .o(n_3603) );
na02m02 TIMEBOOST_cell_3541 ( .a(n_7039), .b(TIMEBOOST_net_350), .o(n_7711) );
na02m02 TIMEBOOST_cell_3542 ( .a(n_2756), .b(n_1229), .o(TIMEBOOST_net_351) );
in01s01 g62988_u0 ( .a(FE_OFN1314_n_6624), .o(g62988_sb) );
na03s02 TIMEBOOST_cell_5430 ( .a(n_3764), .b(g64939_sb), .c(g64939_db), .o(n_3675) );
na02f02 TIMEBOOST_cell_3837 ( .a(TIMEBOOST_net_498), .b(g54157_da), .o(n_13442) );
na02f02 TIMEBOOST_cell_18261 ( .a(TIMEBOOST_net_4387), .b(FE_OCPN1909_n_16497), .o(TIMEBOOST_net_2037) );
in01s01 g62989_u0 ( .a(FE_OFN1295_n_4098), .o(g62989_sb) );
na02s01 TIMEBOOST_cell_36469 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(g65714_sb), .o(TIMEBOOST_net_10473) );
na02s02 TIMEBOOST_cell_44836 ( .a(TIMEBOOST_net_14656), .b(n_4447), .o(TIMEBOOST_net_10910) );
na02s02 TIMEBOOST_cell_37916 ( .a(TIMEBOOST_net_11196), .b(g58027_sb), .o(n_9761) );
in01s01 g62990_u0 ( .a(n_6319), .o(g62990_sb) );
in01s01 TIMEBOOST_cell_45932 ( .a(TIMEBOOST_net_15238), .o(TIMEBOOST_net_15239) );
na02s01 TIMEBOOST_cell_40736 ( .a(TIMEBOOST_net_12606), .b(g62965_sb), .o(n_5952) );
na02s01 TIMEBOOST_cell_3426 ( .a(FE_OFN247_n_9112), .b(g57942_sb), .o(TIMEBOOST_net_293) );
in01s01 g62991_u0 ( .a(FE_OFN1276_n_4096), .o(g62991_sb) );
na02m02 TIMEBOOST_cell_3269 ( .a(n_2485), .b(TIMEBOOST_net_214), .o(n_3195) );
na03s02 TIMEBOOST_cell_37531 ( .a(TIMEBOOST_net_3806), .b(g64145_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__Q), .o(TIMEBOOST_net_11004) );
na02s01 TIMEBOOST_cell_39948 ( .a(TIMEBOOST_net_12212), .b(g62369_sb), .o(n_6865) );
in01s01 g62992_u0 ( .a(n_6319), .o(g62992_sb) );
na02m02 TIMEBOOST_cell_44533 ( .a(n_9714), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q), .o(TIMEBOOST_net_14505) );
na02s01 TIMEBOOST_cell_3427 ( .a(TIMEBOOST_net_293), .b(g57942_db), .o(n_9128) );
na02m02 TIMEBOOST_cell_17495 ( .a(FE_OFN2127_n_16497), .b(TIMEBOOST_net_4004), .o(TIMEBOOST_net_466) );
in01s01 g62993_u0 ( .a(FE_OFN1272_n_4096), .o(g62993_sb) );
na02s01 TIMEBOOST_cell_18611 ( .a(TIMEBOOST_net_4562), .b(g62850_sb), .o(n_5269) );
na03s02 TIMEBOOST_cell_37529 ( .a(TIMEBOOST_net_3803), .b(g65807_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__Q), .o(TIMEBOOST_net_11003) );
na02s01 TIMEBOOST_cell_3272 ( .a(n_3783), .b(n_4677), .o(TIMEBOOST_net_216) );
in01s01 g62994_u0 ( .a(FE_OFN1225_n_6391), .o(g62994_sb) );
na02s01 TIMEBOOST_cell_3273 ( .a(TIMEBOOST_net_216), .b(g65291_da), .o(n_4163) );
na02f02 TIMEBOOST_cell_44728 ( .a(TIMEBOOST_net_14602), .b(FE_OFN1577_n_12028), .o(TIMEBOOST_net_678) );
na02s01 TIMEBOOST_cell_42641 ( .a(FE_OFN209_n_9126), .b(g58172_sb), .o(TIMEBOOST_net_13559) );
in01s01 g62995_u0 ( .a(FE_OFN1193_n_6935), .o(g62995_sb) );
na02s01 TIMEBOOST_cell_3275 ( .a(TIMEBOOST_net_217), .b(g64355_sb), .o(n_3823) );
na02s02 TIMEBOOST_cell_43078 ( .a(TIMEBOOST_net_13777), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_11548) );
na02s02 TIMEBOOST_cell_43320 ( .a(TIMEBOOST_net_13898), .b(g63174_sb), .o(n_5796) );
in01s01 g62996_u0 ( .a(n_6319), .o(g62996_sb) );
na03s02 TIMEBOOST_cell_5411 ( .a(n_3764), .b(g64856_sb), .c(g64856_db), .o(n_3720) );
na02s02 TIMEBOOST_cell_3429 ( .a(TIMEBOOST_net_294), .b(g57968_sb), .o(n_9113) );
na02s01 TIMEBOOST_cell_3430 ( .a(FE_OFN239_n_9832), .b(g58129_sb), .o(TIMEBOOST_net_295) );
in01s01 g62997_u0 ( .a(FE_OFN1225_n_6391), .o(g62997_sb) );
na02s01 TIMEBOOST_cell_3277 ( .a(TIMEBOOST_net_218), .b(n_4488), .o(n_4296) );
na02s02 TIMEBOOST_cell_37981 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_395), .b(g54175_sb), .o(TIMEBOOST_net_11229) );
na03f02 TIMEBOOST_cell_36001 ( .a(TIMEBOOST_net_10109), .b(n_13617), .c(g54484_sb), .o(n_13616) );
in01s01 g62998_u0 ( .a(FE_OFN1320_n_6436), .o(g62998_sb) );
na02s02 TIMEBOOST_cell_45597 ( .a(TIMEBOOST_net_9359), .b(FE_OFN789_n_2678), .o(TIMEBOOST_net_15037) );
na02s02 TIMEBOOST_cell_42856 ( .a(TIMEBOOST_net_13666), .b(FE_OFN2212_n_8407), .o(TIMEBOOST_net_11144) );
na02s01 TIMEBOOST_cell_38564 ( .a(TIMEBOOST_net_11520), .b(g62057_sb), .o(n_7752) );
in01s01 g62999_u0 ( .a(FE_OFN1200_n_4090), .o(g62999_sb) );
na02s01 TIMEBOOST_cell_36471 ( .a(pci_target_unit_fifos_pcir_data_in_174), .b(g65770_sb), .o(TIMEBOOST_net_10474) );
na02f02 TIMEBOOST_cell_41244 ( .a(TIMEBOOST_net_12860), .b(g57085_sb), .o(n_11657) );
na02f02 TIMEBOOST_cell_42328 ( .a(TIMEBOOST_net_13402), .b(g57155_sb), .o(n_11595) );
na02f02 g62_u0 ( .a(FE_OCPN1888_FE_OFN473_n_16992), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__Q), .o(n_15533) );
in01s01 g63000_u0 ( .a(FE_OFN1230_n_6391), .o(g63000_sb) );
na02s01 TIMEBOOST_cell_40822 ( .a(TIMEBOOST_net_12649), .b(g63181_sb), .o(n_5788) );
na02m04 TIMEBOOST_cell_3543 ( .a(n_2761), .b(TIMEBOOST_net_351), .o(n_3197) );
na02s01 TIMEBOOST_cell_38424 ( .a(TIMEBOOST_net_11450), .b(g63552_sb), .o(n_4605) );
in01s01 g63001_u0 ( .a(FE_OFN1214_n_4151), .o(g63001_sb) );
na02s01 TIMEBOOST_cell_36393 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__Q), .b(g65891_sb), .o(TIMEBOOST_net_10435) );
na02s02 TIMEBOOST_cell_44867 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__Q), .b(FE_OFN1642_n_4671), .o(TIMEBOOST_net_14672) );
na02s01 TIMEBOOST_cell_37574 ( .a(TIMEBOOST_net_11025), .b(g65928_db), .o(n_2583) );
in01s01 g63002_u0 ( .a(FE_OFN1272_n_4096), .o(g63002_sb) );
na02s01 TIMEBOOST_cell_3279 ( .a(TIMEBOOST_net_219), .b(n_4479), .o(n_4284) );
na03s02 TIMEBOOST_cell_37527 ( .a(TIMEBOOST_net_3807), .b(g65693_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__Q), .o(TIMEBOOST_net_11002) );
na02s02 TIMEBOOST_cell_43460 ( .a(TIMEBOOST_net_13968), .b(FE_OFN1230_n_6391), .o(TIMEBOOST_net_12165) );
in01s02 g63003_u0 ( .a(n_6645), .o(g63003_sb) );
na02s02 TIMEBOOST_cell_40824 ( .a(TIMEBOOST_net_12650), .b(g63173_sb), .o(n_5798) );
na02s01 TIMEBOOST_cell_3431 ( .a(TIMEBOOST_net_295), .b(g58129_db), .o(n_9665) );
na02s01 TIMEBOOST_cell_3432 ( .a(FE_OFN241_n_9830), .b(g58130_sb), .o(TIMEBOOST_net_296) );
in01s02 g63004_u0 ( .a(FE_OFN1317_n_6624), .o(g63004_sb) );
na02f02 TIMEBOOST_cell_44072 ( .a(TIMEBOOST_net_14274), .b(FE_OFN1373_n_8567), .o(TIMEBOOST_net_12711) );
na02s02 TIMEBOOST_cell_10563 ( .a(TIMEBOOST_net_1848), .b(g59097_sb), .o(TIMEBOOST_net_891) );
na02s01 TIMEBOOST_cell_38566 ( .a(TIMEBOOST_net_11521), .b(g62037_sb), .o(n_7779) );
in01s01 g63005_u0 ( .a(FE_OFN1234_n_6391), .o(g63005_sb) );
na02s02 TIMEBOOST_cell_40826 ( .a(TIMEBOOST_net_12651), .b(g62929_sb), .o(n_6023) );
na02s02 TIMEBOOST_cell_3545 ( .a(TIMEBOOST_net_352), .b(FE_OFN264_n_9849), .o(n_9886) );
na02s01 TIMEBOOST_cell_42567 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__Q), .b(FE_OFN602_n_9687), .o(TIMEBOOST_net_13522) );
in01s01 g63006_u0 ( .a(FE_OFN1196_n_4090), .o(g63006_sb) );
na02s01 TIMEBOOST_cell_36395 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(g65699_sb), .o(TIMEBOOST_net_10436) );
na03s01 TIMEBOOST_cell_6613 ( .a(n_1894), .b(g61879_sb), .c(g61879_db), .o(n_8071) );
in01s01 g63007_u0 ( .a(FE_OFN1258_n_4143), .o(g63007_sb) );
na02s01 TIMEBOOST_cell_36535 ( .a(TIMEBOOST_net_9324), .b(FE_OFN953_n_2055), .o(TIMEBOOST_net_10506) );
in01s01 TIMEBOOST_cell_45910 ( .a(TIMEBOOST_net_15216), .o(TIMEBOOST_net_15217) );
na02f02 TIMEBOOST_cell_42330 ( .a(TIMEBOOST_net_13403), .b(g57550_sb), .o(n_11194) );
in01s02 g63008_u0 ( .a(FE_OFN1311_n_6624), .o(g63008_sb) );
na03s02 TIMEBOOST_cell_5400 ( .a(n_3780), .b(g64752_sb), .c(g64752_db), .o(n_3791) );
in01s01 TIMEBOOST_cell_45911 ( .a(wbm_dat_i_15_), .o(TIMEBOOST_net_15218) );
na02s01 TIMEBOOST_cell_38568 ( .a(TIMEBOOST_net_11522), .b(g62052_sb), .o(n_7757) );
in01s01 g63009_u0 ( .a(FE_OFN1235_n_6391), .o(g63009_sb) );
na02f02 TIMEBOOST_cell_12594 ( .a(n_2740), .b(FE_OFN2198_n_10256), .o(TIMEBOOST_net_2864) );
na02f02 TIMEBOOST_cell_21603 ( .a(TIMEBOOST_net_6058), .b(g57404_sb), .o(n_11337) );
in01s01 TIMEBOOST_cell_32846 ( .a(TIMEBOOST_net_10347), .o(wbs_dat_i_6_) );
in01s01 g63010_u0 ( .a(FE_OFN1134_g64577_p), .o(g63010_sb) );
na02s02 TIMEBOOST_cell_45096 ( .a(TIMEBOOST_net_14786), .b(n_13825), .o(TIMEBOOST_net_12470) );
na02s01 TIMEBOOST_cell_17198 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__Q), .b(g65365_sb), .o(TIMEBOOST_net_3856) );
na02s02 TIMEBOOST_cell_36764 ( .a(TIMEBOOST_net_10620), .b(FE_OFN2106_g64577_p), .o(TIMEBOOST_net_4694) );
in01s01 g63011_u0 ( .a(FE_OFN1207_n_6356), .o(g63011_sb) );
na03s02 TIMEBOOST_cell_6554 ( .a(n_4476), .b(g64972_sb), .c(g64972_db), .o(n_4371) );
na02s01 TIMEBOOST_cell_42008 ( .a(TIMEBOOST_net_13242), .b(g62963_sb), .o(n_5956) );
na02m02 TIMEBOOST_cell_42263 ( .a(n_9822), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__Q), .o(TIMEBOOST_net_13370) );
in01s01 g63012_u0 ( .a(FE_OFN1121_g64577_p), .o(g63012_sb) );
na04f02 TIMEBOOST_cell_36166 ( .a(n_10782), .b(n_11066), .c(n_11067), .d(n_11065), .o(n_12537) );
no02m02 TIMEBOOST_cell_10944 ( .a(n_13784), .b(FE_RN_370_0), .o(TIMEBOOST_net_2039) );
na02s04 TIMEBOOST_cell_45492 ( .a(TIMEBOOST_net_14984), .b(g54368_sb), .o(n_13075) );
in01s01 g63013_u0 ( .a(FE_OFN1104_g64577_p), .o(g63013_sb) );
na02f02 TIMEBOOST_cell_36942 ( .a(TIMEBOOST_net_10709), .b(TIMEBOOST_net_2864), .o(TIMEBOOST_net_10083) );
na02s01 g63013_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__Q), .b(FE_OFN1104_g64577_p), .o(g63013_db) );
na02m02 TIMEBOOST_cell_36822 ( .a(TIMEBOOST_net_10649), .b(g54168_sb), .o(TIMEBOOST_net_9880) );
in01s01 g63014_u0 ( .a(FE_OFN2105_g64577_p), .o(g63014_sb) );
na03s02 TIMEBOOST_cell_37525 ( .a(TIMEBOOST_net_3798), .b(g65967_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__Q), .o(TIMEBOOST_net_11001) );
na02s01 TIMEBOOST_cell_37668 ( .a(TIMEBOOST_net_11072), .b(g61814_sb), .o(n_8163) );
na02s01 TIMEBOOST_cell_37670 ( .a(TIMEBOOST_net_11073), .b(g62002_sb), .o(n_7891) );
in01s01 g63015_u0 ( .a(FE_OFN1122_g64577_p), .o(g63015_sb) );
na02s01 TIMEBOOST_cell_37575 ( .a(parchk_pci_ad_reg_in_1231), .b(g65893_sb), .o(TIMEBOOST_net_11026) );
na02s01 TIMEBOOST_cell_37672 ( .a(TIMEBOOST_net_11074), .b(g61729_sb), .o(n_8362) );
na02s01 TIMEBOOST_cell_37674 ( .a(TIMEBOOST_net_11075), .b(g61883_sb), .o(n_8064) );
in01s01 g63016_u0 ( .a(FE_OFN1100_g64577_p), .o(g63016_sb) );
na02s01 TIMEBOOST_cell_36602 ( .a(TIMEBOOST_net_10539), .b(g65841_sb), .o(n_1879) );
na02s01 g63016_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__Q), .b(FE_OFN1100_g64577_p), .o(g63016_db) );
na02s01 TIMEBOOST_cell_19723 ( .a(TIMEBOOST_net_5118), .b(g62653_sb), .o(n_6238) );
in01s01 g63017_u0 ( .a(FE_OFN1134_g64577_p), .o(g63017_sb) );
na02f02 TIMEBOOST_cell_12885 ( .a(TIMEBOOST_net_3009), .b(n_10792), .o(TIMEBOOST_net_960) );
na02f02 TIMEBOOST_cell_38995 ( .a(TIMEBOOST_net_10105), .b(FE_OFN2158_n_16439), .o(TIMEBOOST_net_11736) );
na02f02 TIMEBOOST_cell_18315 ( .a(TIMEBOOST_net_4414), .b(g54150_da), .o(n_13450) );
in01s01 g63018_u0 ( .a(FE_OFN2104_g64577_p), .o(g63018_sb) );
na03s06 TIMEBOOST_cell_44757 ( .a(conf_wb_err_addr_in_970), .b(conf_wb_err_addr_in_971), .c(n_1441), .o(TIMEBOOST_net_14617) );
na02s01 TIMEBOOST_cell_19955 ( .a(TIMEBOOST_net_5234), .b(g62536_sb), .o(n_6498) );
no02m01 TIMEBOOST_cell_18228 ( .a(TIMEBOOST_net_788), .b(n_15645), .o(TIMEBOOST_net_4371) );
in01s01 g63019_u0 ( .a(FE_OFN2105_g64577_p), .o(g63019_sb) );
na02s02 TIMEBOOST_cell_39950 ( .a(TIMEBOOST_net_12213), .b(g62618_sb), .o(n_7374) );
na02f02 TIMEBOOST_cell_39001 ( .a(TIMEBOOST_net_10104), .b(FE_OFN2158_n_16439), .o(TIMEBOOST_net_11739) );
na02s02 TIMEBOOST_cell_38426 ( .a(TIMEBOOST_net_11451), .b(g63571_sb), .o(n_4111) );
in01s01 g63020_u0 ( .a(FE_OFN1100_g64577_p), .o(g63020_sb) );
na02s02 TIMEBOOST_cell_36766 ( .a(TIMEBOOST_net_10621), .b(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_4502) );
na02s01 g63020_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__Q), .b(FE_OFN1100_g64577_p), .o(g63020_db) );
na02s02 TIMEBOOST_cell_38428 ( .a(TIMEBOOST_net_11452), .b(g63099_sb), .o(n_5056) );
in01s01 g63021_u0 ( .a(FE_OFN1116_g64577_p), .o(g63021_sb) );
no02m02 TIMEBOOST_cell_10950 ( .a(FE_RN_541_0), .b(n_13784), .o(TIMEBOOST_net_2042) );
na03s02 TIMEBOOST_cell_33962 ( .a(n_2054), .b(g62025_sb), .c(g62025_db), .o(n_7847) );
in01s01 g63022_u0 ( .a(FE_OFN882_g64577_p), .o(g63022_sb) );
na02s02 TIMEBOOST_cell_43074 ( .a(TIMEBOOST_net_13775), .b(FE_OFN1197_n_4090), .o(TIMEBOOST_net_12030) );
na02s02 TIMEBOOST_cell_43472 ( .a(TIMEBOOST_net_13974), .b(FE_OFN1234_n_6391), .o(TIMEBOOST_net_12150) );
na02f02 TIMEBOOST_cell_12899 ( .a(FE_OCP_RBN1985_FE_OFN1591_n_13741), .b(TIMEBOOST_net_3016), .o(g53158_p) );
in01s01 g63023_u0 ( .a(FE_OFN882_g64577_p), .o(g63023_sb) );
na02f02 TIMEBOOST_cell_12901 ( .a(FE_OCP_RBN1985_FE_OFN1591_n_13741), .b(TIMEBOOST_net_3017), .o(g74859_p) );
na02s02 TIMEBOOST_cell_44425 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_0__Q), .o(TIMEBOOST_net_14451) );
na02f02 TIMEBOOST_cell_12903 ( .a(FE_OCP_RBN1984_FE_OFN1591_n_13741), .b(TIMEBOOST_net_3018), .o(g53230_p) );
in01s01 g63024_u0 ( .a(FE_OFN1122_g64577_p), .o(g63024_sb) );
na02s01 TIMEBOOST_cell_37936 ( .a(TIMEBOOST_net_11206), .b(g58360_sb), .o(n_9463) );
na02m02 TIMEBOOST_cell_44629 ( .a(n_9733), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q), .o(TIMEBOOST_net_14553) );
na02f02 TIMEBOOST_cell_12905 ( .a(FE_OCP_RBN1985_FE_OFN1591_n_13741), .b(TIMEBOOST_net_3019), .o(g53251_p) );
na02m02 TIMEBOOST_cell_38714 ( .a(TIMEBOOST_net_11595), .b(g62408_sb), .o(n_6783) );
na02s01 g63025_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__21__Q), .b(FE_OFN1106_g64577_p), .o(g63025_db) );
na02s02 TIMEBOOST_cell_38430 ( .a(TIMEBOOST_net_11453), .b(g63092_sb), .o(n_5068) );
in01s01 g63026_u0 ( .a(FE_OFN1122_g64577_p), .o(g63026_sb) );
na02s02 TIMEBOOST_cell_37557 ( .a(pci_target_unit_pcit_if_strd_addr_in_707), .b(g52636_sb), .o(TIMEBOOST_net_11017) );
na02s01 TIMEBOOST_cell_37606 ( .a(TIMEBOOST_net_11041), .b(g61712_sb), .o(n_8402) );
na03s02 TIMEBOOST_cell_1582 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__Q), .b(g62575_sb), .c(g62575_db), .o(n_6402) );
in01s01 g63027_u0 ( .a(FE_OFN877_g64577_p), .o(g63027_sb) );
na03s01 TIMEBOOST_cell_33964 ( .a(n_1936), .b(g61766_sb), .c(g61766_db), .o(n_8279) );
na02s01 g63027_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__Q), .b(FE_OFN1100_g64577_p), .o(g63027_db) );
no02f02 TIMEBOOST_cell_12909 ( .a(TIMEBOOST_net_3021), .b(FE_RN_816_0), .o(n_14438) );
in01s01 g63028_u0 ( .a(FE_OFN1123_g64577_p), .o(g63028_sb) );
na02s02 TIMEBOOST_cell_16800 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__Q), .b(g65393_sb), .o(TIMEBOOST_net_3657) );
na02s02 TIMEBOOST_cell_45155 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__Q), .b(n_4282), .o(TIMEBOOST_net_14816) );
na02s01 TIMEBOOST_cell_16803 ( .a(TIMEBOOST_net_3658), .b(g65025_db), .o(n_3629) );
in01s01 g63029_u0 ( .a(n_6645), .o(g63029_sb) );
na02s02 TIMEBOOST_cell_43443 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__Q), .b(n_4393), .o(TIMEBOOST_net_13960) );
na02s01 TIMEBOOST_cell_3433 ( .a(TIMEBOOST_net_296), .b(g58130_db), .o(n_9663) );
na02s01 TIMEBOOST_cell_3434 ( .a(FE_OFN247_n_9112), .b(g58064_db), .o(TIMEBOOST_net_297) );
in01s01 g63030_u0 ( .a(FE_OFN1118_g64577_p), .o(g63030_sb) );
na03s02 TIMEBOOST_cell_34256 ( .a(TIMEBOOST_net_9819), .b(FE_OFN1169_n_5592), .c(g62109_sb), .o(n_5589) );
na02f02 TIMEBOOST_cell_44713 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__Q), .b(FE_OFN1746_n_12004), .o(TIMEBOOST_net_14595) );
in01s01 g63031_u0 ( .a(FE_OFN1123_g64577_p), .o(g63031_sb) );
na02s02 TIMEBOOST_cell_39952 ( .a(TIMEBOOST_net_12214), .b(g62898_sb), .o(n_6081) );
na02s02 g63031_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__Q), .b(FE_OFN1123_g64577_p), .o(g63031_db) );
in01s01 g63032_u0 ( .a(FE_OFN1131_g64577_p), .o(g63032_sb) );
na02s01 TIMEBOOST_cell_16642 ( .a(pci_target_unit_fifos_pciw_addr_data_in_147), .b(g64161_sb), .o(TIMEBOOST_net_3578) );
na02m02 TIMEBOOST_cell_10962 ( .a(n_1161), .b(n_1162), .o(TIMEBOOST_net_2048) );
na02m02 TIMEBOOST_cell_39954 ( .a(TIMEBOOST_net_12215), .b(g62967_sb), .o(n_5948) );
in01s01 g63033_u0 ( .a(FE_OFN1121_g64577_p), .o(g63033_sb) );
na02s02 TIMEBOOST_cell_39956 ( .a(TIMEBOOST_net_12216), .b(g62663_sb), .o(n_6213) );
na03s02 TIMEBOOST_cell_34257 ( .a(TIMEBOOST_net_9818), .b(FE_OFN1174_n_5592), .c(g62108_sb), .o(n_5591) );
na02f02 TIMEBOOST_cell_44152 ( .a(TIMEBOOST_net_14314), .b(FE_OFN1419_n_8567), .o(TIMEBOOST_net_12846) );
in01s01 g63034_u0 ( .a(FE_OFN1116_g64577_p), .o(g63034_sb) );
no02f04 TIMEBOOST_cell_12917 ( .a(FE_RN_807_0), .b(TIMEBOOST_net_3025), .o(n_14273) );
na02f02 TIMEBOOST_cell_18206 ( .a(FE_OFN1069_n_15729), .b(configuration_wb_err_data_582), .o(TIMEBOOST_net_4360) );
na02f04 TIMEBOOST_cell_37110 ( .a(TIMEBOOST_net_10793), .b(n_12573), .o(n_12835) );
in01s01 g63035_u0 ( .a(FE_OFN1127_g64577_p), .o(g63035_sb) );
no02f02 TIMEBOOST_cell_12921 ( .a(TIMEBOOST_net_3027), .b(n_7823), .o(g53078_p) );
na02f02 TIMEBOOST_cell_44184 ( .a(TIMEBOOST_net_14330), .b(FE_OFN1390_n_8567), .o(TIMEBOOST_net_12750) );
na02f02 TIMEBOOST_cell_44073 ( .a(n_9032), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__Q), .o(TIMEBOOST_net_14275) );
in01s01 g63036_u0 ( .a(FE_OFN1120_g64577_p), .o(g63036_sb) );
na02s01 TIMEBOOST_cell_38432 ( .a(TIMEBOOST_net_11454), .b(g61894_sb), .o(n_7967) );
na02s02 g63036_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__Q), .b(FE_OFN1129_g64577_p), .o(g63036_db) );
na02f02 TIMEBOOST_cell_44074 ( .a(TIMEBOOST_net_14275), .b(FE_OFN1381_n_8567), .o(TIMEBOOST_net_13380) );
in01s01 g63037_u0 ( .a(FE_OFN1121_g64577_p), .o(g63037_sb) );
na02s01 TIMEBOOST_cell_38434 ( .a(TIMEBOOST_net_11455), .b(g61925_sb), .o(n_7973) );
na02s01 TIMEBOOST_cell_37608 ( .a(TIMEBOOST_net_11042), .b(g61723_sb), .o(n_8376) );
na02s01 TIMEBOOST_cell_38436 ( .a(TIMEBOOST_net_11456), .b(g61932_sb), .o(n_7959) );
in01s01 g63038_u0 ( .a(FE_OFN1122_g64577_p), .o(g63038_sb) );
na04f02 TIMEBOOST_cell_36170 ( .a(n_11061), .b(n_11777), .c(n_11060), .d(n_11062), .o(n_12535) );
na02s01 TIMEBOOST_cell_18212 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_408), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_4363) );
na03f02 TIMEBOOST_cell_36172 ( .a(n_14128), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__Q), .c(FE_OFN1601_n_13995), .o(n_14451) );
in01s01 g63039_u0 ( .a(FE_OFN1097_g64577_p), .o(g63039_sb) );
na02f02 TIMEBOOST_cell_42955 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_400), .b(g54134_sb), .o(TIMEBOOST_net_13716) );
na02s01 g63039_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__Q), .b(FE_OFN1097_g64577_p), .o(g63039_db) );
na02s01 TIMEBOOST_cell_38438 ( .a(TIMEBOOST_net_11457), .b(g61934_sb), .o(n_7955) );
in01s01 g63040_u0 ( .a(FE_OFN1133_g64577_p), .o(g63040_sb) );
na02f02 TIMEBOOST_cell_44638 ( .a(TIMEBOOST_net_14557), .b(FE_OFN2174_n_8567), .o(TIMEBOOST_net_13484) );
na02s01 TIMEBOOST_cell_18214 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_390), .b(FE_OFN2070_n_15978), .o(TIMEBOOST_net_4364) );
na02s02 TIMEBOOST_cell_38440 ( .a(TIMEBOOST_net_11458), .b(FE_OFN1801_n_9690), .o(TIMEBOOST_net_4725) );
in01s01 g63041_u0 ( .a(FE_OFN1133_g64577_p), .o(g63041_sb) );
no02f06 TIMEBOOST_cell_12943 ( .a(TIMEBOOST_net_3038), .b(n_13340), .o(n_13907) );
na02s02 TIMEBOOST_cell_37964 ( .a(TIMEBOOST_net_11220), .b(g61892_sb), .o(n_8044) );
na02s01 TIMEBOOST_cell_39178 ( .a(TIMEBOOST_net_11827), .b(g58079_sb), .o(TIMEBOOST_net_356) );
in01s01 g63042_u0 ( .a(FE_OFN2064_n_6391), .o(g63042_sb) );
na02m02 TIMEBOOST_cell_44075 ( .a(n_9516), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__Q), .o(TIMEBOOST_net_14276) );
na02f02 TIMEBOOST_cell_44076 ( .a(TIMEBOOST_net_14276), .b(FE_OFN1424_n_8567), .o(TIMEBOOST_net_13381) );
na02s02 TIMEBOOST_cell_43475 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__Q), .b(n_3574), .o(TIMEBOOST_net_13976) );
in01s01 g63043_u0 ( .a(FE_OFN1119_g64577_p), .o(g63043_sb) );
na02s01 TIMEBOOST_cell_37483 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__Q), .b(g65887_sb), .o(TIMEBOOST_net_10980) );
na02s01 TIMEBOOST_cell_37610 ( .a(TIMEBOOST_net_11043), .b(g61927_sb), .o(n_7969) );
na02f04 TIMEBOOST_cell_11683 ( .a(TIMEBOOST_net_2408), .b(n_8566), .o(n_8819) );
in01s01 g63044_u0 ( .a(FE_OFN1128_g64577_p), .o(g63044_sb) );
na02s02 TIMEBOOST_cell_9048 ( .a(FE_OFN2055_n_8831), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_22__Q), .o(TIMEBOOST_net_1091) );
na02s02 TIMEBOOST_cell_38594 ( .a(TIMEBOOST_net_11535), .b(n_2234), .o(n_4859) );
na02s02 TIMEBOOST_cell_38442 ( .a(TIMEBOOST_net_11459), .b(FE_OFN569_n_9528), .o(TIMEBOOST_net_4722) );
in01s01 g63045_u0 ( .a(FE_OFN1097_g64577_p), .o(g63045_sb) );
na02s02 TIMEBOOST_cell_37766 ( .a(TIMEBOOST_net_11121), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_10596) );
na02f02 TIMEBOOST_cell_39151 ( .a(n_12313), .b(TIMEBOOST_net_10189), .o(TIMEBOOST_net_11814) );
na02s02 TIMEBOOST_cell_37768 ( .a(TIMEBOOST_net_11122), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_10594) );
in01s01 g63046_u0 ( .a(FE_OFN1123_g64577_p), .o(g63046_sb) );
na03s02 TIMEBOOST_cell_6314 ( .a(FE_OFN254_n_9825), .b(g58168_db), .c(g58140_sb), .o(n_9623) );
na02m02 TIMEBOOST_cell_10980 ( .a(wbm_adr_o_26_), .b(FE_OFN1700_n_5751), .o(TIMEBOOST_net_2057) );
na02f02 TIMEBOOST_cell_12789 ( .a(TIMEBOOST_net_2961), .b(n_14140), .o(n_14461) );
in01s01 g63047_u0 ( .a(FE_OFN881_g64577_p), .o(g63047_sb) );
na02m02 TIMEBOOST_cell_38888 ( .a(TIMEBOOST_net_11682), .b(g58837_sb), .o(n_8677) );
na02s01 g63047_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__Q), .b(FE_OFN881_g64577_p), .o(g63047_db) );
na02s02 TIMEBOOST_cell_36768 ( .a(TIMEBOOST_net_10622), .b(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_4627) );
in01s01 g63048_u0 ( .a(FE_OFN1094_g64577_p), .o(g63048_sb) );
na02f02 TIMEBOOST_cell_22570 ( .a(FE_OFN1739_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__Q), .o(TIMEBOOST_net_6542) );
na02s01 TIMEBOOST_cell_15833 ( .a(TIMEBOOST_net_3173), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_405), .o(TIMEBOOST_net_67) );
na03s02 TIMEBOOST_cell_33810 ( .a(FE_OFN215_n_9856), .b(g58234_sb), .c(g58234_db), .o(n_9557) );
in01s01 g63049_u0 ( .a(FE_OFN1129_g64577_p), .o(g63049_sb) );
na02s01 TIMEBOOST_cell_38444 ( .a(TIMEBOOST_net_11460), .b(g61931_sb), .o(n_7961) );
na02s01 TIMEBOOST_cell_19034 ( .a(wishbone_slave_unit_pcim_sm_data_in_662), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__Q), .o(TIMEBOOST_net_4774) );
na02s01 TIMEBOOST_cell_16804 ( .a(n_3770), .b(g64970_sb), .o(TIMEBOOST_net_3659) );
in01s01 g63050_u0 ( .a(FE_OFN1112_g64577_p), .o(g63050_sb) );
na03s02 TIMEBOOST_cell_43321 ( .a(n_3716), .b(FE_OFN1278_n_4097), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__15__Q), .o(TIMEBOOST_net_13899) );
na02f02 TIMEBOOST_cell_39093 ( .a(FE_OCP_RBN1999_n_13971), .b(TIMEBOOST_net_10228), .o(TIMEBOOST_net_11785) );
na02s01 TIMEBOOST_cell_41735 ( .a(n_4498), .b(n_4677), .o(TIMEBOOST_net_13106) );
in01s01 g63051_u0 ( .a(FE_OFN1134_g64577_p), .o(g63051_sb) );
na02s01 TIMEBOOST_cell_16810 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__Q), .b(g65334_sb), .o(TIMEBOOST_net_3662) );
na02s01 g63051_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__Q), .b(FE_OFN882_g64577_p), .o(g63051_db) );
na02s02 TIMEBOOST_cell_43559 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__Q), .b(n_4336), .o(TIMEBOOST_net_14018) );
in01s01 g63052_u0 ( .a(FE_OFN881_g64577_p), .o(g63052_sb) );
na02s02 TIMEBOOST_cell_39300 ( .a(TIMEBOOST_net_11888), .b(g65683_sb), .o(n_2039) );
na02s01 g63052_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__Q), .b(FE_OFN1104_g64577_p), .o(g63052_db) );
na02f02 TIMEBOOST_cell_37125 ( .a(n_13997), .b(TIMEBOOST_net_6241), .o(TIMEBOOST_net_10801) );
in01s01 g63053_u0 ( .a(FE_OFN1135_g64577_p), .o(g63053_sb) );
na02s01 TIMEBOOST_cell_38446 ( .a(TIMEBOOST_net_11461), .b(FE_OFN1651_n_9428), .o(TIMEBOOST_net_2032) );
na03s02 TIMEBOOST_cell_38043 ( .a(g64290_da), .b(g64290_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__Q), .o(TIMEBOOST_net_11260) );
na02s01 TIMEBOOST_cell_43257 ( .a(n_3675), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__Q), .o(TIMEBOOST_net_13867) );
in01s01 g63054_u0 ( .a(FE_OFN1128_g64577_p), .o(g63054_sb) );
na02f02 TIMEBOOST_cell_43810 ( .a(TIMEBOOST_net_14143), .b(FE_OFN1398_n_8567), .o(TIMEBOOST_net_12958) );
no02m04 TIMEBOOST_cell_19038 ( .a(FE_RN_710_0), .b(n_13784), .o(TIMEBOOST_net_4776) );
na02s01 g65962_u3 ( .a(g65962_da), .b(g65962_db), .o(n_2160) );
in01s01 g63055_u0 ( .a(FE_OFN1115_g64577_p), .o(g63055_sb) );
na02f02 TIMEBOOST_cell_44534 ( .a(TIMEBOOST_net_14505), .b(FE_OFN2177_n_8567), .o(TIMEBOOST_net_13495) );
na02m02 TIMEBOOST_cell_38941 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_16__Q), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__Q), .o(TIMEBOOST_net_11709) );
na02s02 TIMEBOOST_cell_43390 ( .a(TIMEBOOST_net_13933), .b(n_6232), .o(TIMEBOOST_net_12156) );
in01s01 g63056_u0 ( .a(FE_OFN1104_g64577_p), .o(g63056_sb) );
na02s01 TIMEBOOST_cell_36824 ( .a(TIMEBOOST_net_10650), .b(g54173_sb), .o(TIMEBOOST_net_9879) );
na02s01 g63056_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__Q), .b(FE_OFN1104_g64577_p), .o(g63056_db) );
na02f10 TIMEBOOST_cell_36241 ( .a(conf_wb_err_bc_in_846), .b(g67048_sb), .o(TIMEBOOST_net_10359) );
na02s02 TIMEBOOST_cell_36790 ( .a(TIMEBOOST_net_10633), .b(FE_OFN1126_g64577_p), .o(TIMEBOOST_net_4668) );
no02f02 TIMEBOOST_cell_39180 ( .a(TIMEBOOST_net_11828), .b(FE_RN_619_0), .o(TIMEBOOST_net_323) );
na02f02 TIMEBOOST_cell_37036 ( .a(TIMEBOOST_net_10756), .b(FE_OFN1774_n_13800), .o(g74879_p) );
in01s01 g63058_u0 ( .a(FE_OFN1104_g64577_p), .o(g63058_sb) );
na02f02 TIMEBOOST_cell_37038 ( .a(TIMEBOOST_net_10757), .b(FE_OFN1774_n_13800), .o(g74886_p) );
na02f02 TIMEBOOST_cell_44408 ( .a(TIMEBOOST_net_14442), .b(FE_OFN1389_n_8567), .o(TIMEBOOST_net_12818) );
na02f02 TIMEBOOST_cell_37040 ( .a(TIMEBOOST_net_10758), .b(FE_OFN1774_n_13800), .o(g53175_p) );
in01s01 g63059_u0 ( .a(FE_OFN882_g64577_p), .o(g63059_sb) );
na02m02 TIMEBOOST_cell_44077 ( .a(n_9469), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__Q), .o(TIMEBOOST_net_14277) );
na02s02 TIMEBOOST_cell_39266 ( .a(TIMEBOOST_net_11871), .b(n_4442), .o(n_4233) );
na02s02 TIMEBOOST_cell_43391 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__Q), .b(n_1959), .o(TIMEBOOST_net_13934) );
in01s01 g63060_u0 ( .a(FE_OFN877_g64577_p), .o(g63060_sb) );
na02s02 TIMEBOOST_cell_43392 ( .a(TIMEBOOST_net_13934), .b(n_6554), .o(TIMEBOOST_net_12152) );
na02s01 g63060_u2 ( .a(FE_OFN1100_g64577_p), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__Q), .o(g63060_db) );
na02f04 TIMEBOOST_cell_39022 ( .a(TIMEBOOST_net_11749), .b(FE_OFN2241_g52675_p), .o(TIMEBOOST_net_10751) );
in01s01 g63061_u0 ( .a(FE_OFN1140_g64577_p), .o(g63061_sb) );
na02f02 TIMEBOOST_cell_44078 ( .a(TIMEBOOST_net_14277), .b(FE_OFN1406_n_8567), .o(TIMEBOOST_net_12839) );
na02m02 TIMEBOOST_cell_39958 ( .a(TIMEBOOST_net_12217), .b(g62345_sb), .o(n_6910) );
na02m02 TIMEBOOST_cell_44551 ( .a(n_9777), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__Q), .o(TIMEBOOST_net_14514) );
in01s01 g63062_u0 ( .a(FE_OFN1122_g64577_p), .o(g63062_sb) );
na02f02 TIMEBOOST_cell_44552 ( .a(TIMEBOOST_net_14514), .b(FE_OFN2182_n_8567), .o(TIMEBOOST_net_13465) );
na02m02 TIMEBOOST_cell_45799 ( .a(n_9436), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__Q), .o(TIMEBOOST_net_15138) );
na02s02 TIMEBOOST_cell_42760 ( .a(TIMEBOOST_net_13618), .b(g64176_da), .o(TIMEBOOST_net_11349) );
in01s01 g63063_u0 ( .a(FE_OFN1122_g64577_p), .o(g63063_sb) );
na02m02 TIMEBOOST_cell_44553 ( .a(n_9814), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__Q), .o(TIMEBOOST_net_14515) );
na02s01 g63063_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__Q), .b(FE_OFN1106_g64577_p), .o(g63063_db) );
na02s02 TIMEBOOST_cell_42761 ( .a(g58127_sb), .b(g58127_db), .o(TIMEBOOST_net_13619) );
in01s01 g63064_u0 ( .a(FE_OFN1135_g64577_p), .o(g63064_sb) );
na02f02 TIMEBOOST_cell_38448 ( .a(TIMEBOOST_net_11462), .b(FE_OCP_RBN2223_n_15347), .o(n_15377) );
na02m02 TIMEBOOST_cell_32546 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__Q), .o(TIMEBOOST_net_10184) );
na02s02 TIMEBOOST_cell_42762 ( .a(TIMEBOOST_net_13619), .b(FE_OFN235_n_9834), .o(n_9666) );
in01s01 g63065_u0 ( .a(FE_OFN1140_g64577_p), .o(g63065_sb) );
na02s02 TIMEBOOST_cell_38450 ( .a(TIMEBOOST_net_11463), .b(g54190_sb), .o(n_13490) );
na02s01 TIMEBOOST_cell_39233 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(g65682_sb), .o(TIMEBOOST_net_11855) );
na02f02 TIMEBOOST_cell_44554 ( .a(TIMEBOOST_net_14515), .b(FE_OFN2182_n_8567), .o(TIMEBOOST_net_13466) );
in01s01 g63066_u0 ( .a(FE_OFN2105_g64577_p), .o(g63066_sb) );
na02m02 TIMEBOOST_cell_43811 ( .a(n_9019), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__Q), .o(TIMEBOOST_net_14144) );
na02s01 TIMEBOOST_cell_39235 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(g65728_sb), .o(TIMEBOOST_net_11856) );
na02s01 TIMEBOOST_cell_42764 ( .a(TIMEBOOST_net_13620), .b(g63545_da), .o(TIMEBOOST_net_11319) );
in01s01 g63067_u0 ( .a(FE_OFN877_g64577_p), .o(g63067_sb) );
na02s01 TIMEBOOST_cell_43393 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__Q), .b(n_4474), .o(TIMEBOOST_net_13935) );
na02s02 TIMEBOOST_cell_39960 ( .a(TIMEBOOST_net_12218), .b(g62504_sb), .o(n_6572) );
na02m02 TIMEBOOST_cell_44555 ( .a(n_9473), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__Q), .o(TIMEBOOST_net_14516) );
in01s01 g63068_u0 ( .a(FE_OFN1123_g64577_p), .o(g63068_sb) );
na03f08 TIMEBOOST_cell_2089 ( .a(FE_RN_302_0), .b(n_16977), .c(n_15458), .o(n_16131) );
na02s01 TIMEBOOST_cell_39237 ( .a(n_4444), .b(g64931_sb), .o(TIMEBOOST_net_11857) );
na02s01 TIMEBOOST_cell_16799 ( .a(TIMEBOOST_net_3656), .b(g65056_db), .o(n_3615) );
in01s01 g63069_u0 ( .a(FE_OFN1137_g64577_p), .o(g63069_sb) );
na03f02 TIMEBOOST_cell_36078 ( .a(n_11972), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__Q), .c(FE_OFN1749_n_12004), .o(n_12684) );
na02s02 TIMEBOOST_cell_45787 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__Q), .b(n_4449), .o(TIMEBOOST_net_15132) );
na02m04 TIMEBOOST_cell_45494 ( .a(TIMEBOOST_net_14985), .b(g54369_sb), .o(n_13074) );
in01s01 g63070_u0 ( .a(FE_OFN882_g64577_p), .o(g63070_sb) );
na03f02 TIMEBOOST_cell_35990 ( .a(TIMEBOOST_net_10120), .b(n_13617), .c(g54491_sb), .o(n_13603) );
na02f02 TIMEBOOST_cell_41152 ( .a(TIMEBOOST_net_12814), .b(g57512_sb), .o(n_10319) );
na03f02 TIMEBOOST_cell_35992 ( .a(TIMEBOOST_net_10118), .b(n_13617), .c(g54471_sb), .o(n_13619) );
in01s01 g63071_u0 ( .a(FE_OFN1131_g64577_p), .o(g63071_sb) );
na02s01 TIMEBOOST_cell_9762 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__Q), .b(g65908_sb), .o(TIMEBOOST_net_1448) );
na02s01 TIMEBOOST_cell_39241 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__Q), .b(g58314_sb), .o(TIMEBOOST_net_11859) );
na03f02 TIMEBOOST_cell_35994 ( .a(TIMEBOOST_net_10116), .b(n_13617), .c(g54493_sb), .o(n_13599) );
in01s01 g63072_u0 ( .a(FE_OFN1121_g64577_p), .o(g63072_sb) );
na02s01 TIMEBOOST_cell_42866 ( .a(TIMEBOOST_net_13671), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_11212) );
na02m02 TIMEBOOST_cell_32544 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q), .o(TIMEBOOST_net_10183) );
na02f02 TIMEBOOST_cell_41861 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_388), .b(g54153_sb), .o(TIMEBOOST_net_13169) );
in01s01 g63073_u0 ( .a(FE_OFN1116_g64577_p), .o(g63073_sb) );
na02f02 TIMEBOOST_cell_13035 ( .a(FE_OFN1577_n_12028), .b(TIMEBOOST_net_3084), .o(n_12752) );
na02f02 TIMEBOOST_cell_41154 ( .a(TIMEBOOST_net_12815), .b(g57279_sb), .o(n_10413) );
na02f02 TIMEBOOST_cell_13037 ( .a(FE_OFN1577_n_12028), .b(TIMEBOOST_net_3085), .o(n_12686) );
in01s01 g63074_u0 ( .a(FE_OFN1136_g64577_p), .o(g63074_sb) );
na02s01 TIMEBOOST_cell_39243 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q), .b(g58425_sb), .o(TIMEBOOST_net_11860) );
na02s01 TIMEBOOST_cell_19050 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__Q), .b(g65432_sb), .o(TIMEBOOST_net_4782) );
in01s01 g63075_u0 ( .a(FE_OFN1129_g64577_p), .o(g63075_sb) );
na02s01 TIMEBOOST_cell_42798 ( .a(TIMEBOOST_net_13637), .b(g64091_db), .o(n_4064) );
na02s01 TIMEBOOST_cell_39245 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__Q), .b(g58338_sb), .o(TIMEBOOST_net_11861) );
na02s02 TIMEBOOST_cell_42799 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__Q), .b(g58398_sb), .o(TIMEBOOST_net_13638) );
in01s01 g63076_u0 ( .a(FE_OFN1130_g64577_p), .o(g63076_sb) );
na02s02 TIMEBOOST_cell_42800 ( .a(TIMEBOOST_net_13638), .b(g58398_db), .o(n_9436) );
na02m02 TIMEBOOST_cell_32542 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__Q), .o(TIMEBOOST_net_10182) );
na02s01 TIMEBOOST_cell_42801 ( .a(TIMEBOOST_net_9566), .b(FE_OFN1801_n_9690), .o(TIMEBOOST_net_13639) );
in01s01 g63077_u0 ( .a(FE_OFN1097_g64577_p), .o(g63077_sb) );
na02f02 TIMEBOOST_cell_37042 ( .a(TIMEBOOST_net_10759), .b(FE_OFN1596_n_13741), .o(g53238_p) );
na02s01 g63077_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q), .b(FE_OFN1095_g64577_p), .o(g63077_db) );
na02f02 TIMEBOOST_cell_37044 ( .a(TIMEBOOST_net_10760), .b(FE_OFN1768_n_14054), .o(g53242_p) );
in01s01 g63078_u0 ( .a(FE_OFN1133_g64577_p), .o(g63078_sb) );
na02f02 TIMEBOOST_cell_44556 ( .a(TIMEBOOST_net_14516), .b(FE_OFN2178_n_8567), .o(TIMEBOOST_net_13467) );
na02f02 TIMEBOOST_cell_32541 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_10181), .o(TIMEBOOST_net_6341) );
na02s02 TIMEBOOST_cell_42802 ( .a(TIMEBOOST_net_13639), .b(g58263_sb), .o(n_9038) );
in01s01 g63079_u0 ( .a(FE_OFN1132_g64577_p), .o(g63079_sb) );
na02m02 TIMEBOOST_cell_42803 ( .a(g52483_da), .b(FE_OFN8_n_11877), .o(TIMEBOOST_net_13640) );
na02m02 TIMEBOOST_cell_32540 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__Q), .o(TIMEBOOST_net_10181) );
na02f02 TIMEBOOST_cell_13059 ( .a(n_11920), .b(TIMEBOOST_net_3096), .o(n_12639) );
in01s01 g63080_u0 ( .a(FE_OFN1119_g64577_p), .o(g63080_sb) );
na02s04 TIMEBOOST_cell_45809 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_9__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_774), .o(TIMEBOOST_net_15143) );
na02m02 TIMEBOOST_cell_11685 ( .a(n_8529), .b(TIMEBOOST_net_2409), .o(n_8531) );
na02s02 TIMEBOOST_cell_37940 ( .a(TIMEBOOST_net_11208), .b(g58386_sb), .o(n_9445) );
in01s01 g63081_u0 ( .a(FE_OFN2106_g64577_p), .o(g63081_sb) );
na02s01 TIMEBOOST_cell_37487 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__Q), .b(n_4452), .o(TIMEBOOST_net_10982) );
na02s02 TIMEBOOST_cell_38452 ( .a(TIMEBOOST_net_11464), .b(g54193_sb), .o(n_13424) );
na02s02 TIMEBOOST_cell_37918 ( .a(TIMEBOOST_net_11197), .b(g58171_sb), .o(n_9619) );
in01s01 g63082_u0 ( .a(FE_OFN1133_g64577_p), .o(g63082_sb) );
na02m02 TIMEBOOST_cell_42804 ( .a(TIMEBOOST_net_13640), .b(n_2226), .o(TIMEBOOST_net_11687) );
na02f02 TIMEBOOST_cell_41156 ( .a(TIMEBOOST_net_12816), .b(g57298_sb), .o(n_10408) );
na02s01 TIMEBOOST_cell_42805 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__13__Q), .b(g64283_sb), .o(TIMEBOOST_net_13641) );
in01s01 g63083_u0 ( .a(FE_OFN1120_g64577_p), .o(g63083_sb) );
na02s01 TIMEBOOST_cell_37489 ( .a(TIMEBOOST_net_9504), .b(FE_OFN1043_n_2037), .o(TIMEBOOST_net_10983) );
na02s01 TIMEBOOST_cell_36348 ( .a(TIMEBOOST_net_10412), .b(g67051_sb), .o(n_1499) );
na02s01 TIMEBOOST_cell_37612 ( .a(TIMEBOOST_net_11044), .b(g61818_sb), .o(n_8154) );
in01s01 g63084_u0 ( .a(FE_OFN1123_g64577_p), .o(g63084_sb) );
na02f02 TIMEBOOST_cell_13065 ( .a(TIMEBOOST_net_3099), .b(n_11978), .o(n_12692) );
na02s01 TIMEBOOST_cell_18966 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q), .b(g58339_sb), .o(TIMEBOOST_net_4740) );
na02s01 TIMEBOOST_cell_42806 ( .a(TIMEBOOST_net_13641), .b(g64283_db), .o(n_3890) );
in01s01 g63085_u0 ( .a(FE_OFN881_g64577_p), .o(g63085_sb) );
na02f02 TIMEBOOST_cell_36994 ( .a(TIMEBOOST_net_10735), .b(g58810_sb), .o(n_8631) );
na02f02 TIMEBOOST_cell_36978 ( .a(TIMEBOOST_net_10727), .b(g58804_sb), .o(n_8637) );
na02f02 TIMEBOOST_cell_36996 ( .a(TIMEBOOST_net_10736), .b(g58818_sb), .o(n_8623) );
in01s01 g63086_u0 ( .a(FE_OFN1094_g64577_p), .o(g63086_sb) );
na02f02 TIMEBOOST_cell_22571 ( .a(n_11890), .b(TIMEBOOST_net_6542), .o(n_12607) );
na02s01 g63086_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q), .b(FE_OFN1094_g64577_p), .o(g63086_db) );
na03s02 TIMEBOOST_cell_33811 ( .a(FE_OFN215_n_9856), .b(g58204_sb), .c(g58204_db), .o(n_9583) );
in01s01 g63087_u0 ( .a(FE_OFN1123_g64577_p), .o(g63087_sb) );
na02s01 TIMEBOOST_cell_42807 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__Q), .b(g65303_sb), .o(TIMEBOOST_net_13642) );
na03s02 TIMEBOOST_cell_34270 ( .a(TIMEBOOST_net_9809), .b(FE_OFN1174_n_5592), .c(g62105_sb), .o(n_5595) );
na02s01 TIMEBOOST_cell_42808 ( .a(TIMEBOOST_net_13642), .b(g65303_db), .o(n_4276) );
in01s01 g63088_u0 ( .a(FE_OFN1137_g64577_p), .o(g63088_sb) );
na03s02 TIMEBOOST_cell_42809 ( .a(g61868_sb), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__Q), .c(FE_OFN704_n_8069), .o(TIMEBOOST_net_13643) );
na03s02 TIMEBOOST_cell_34271 ( .a(TIMEBOOST_net_9808), .b(FE_OFN1169_n_5592), .c(g62081_sb), .o(n_5628) );
na02s01 TIMEBOOST_cell_42810 ( .a(TIMEBOOST_net_13643), .b(n_1900), .o(n_8100) );
in01s01 g63089_u0 ( .a(FE_OFN1104_g64577_p), .o(g63089_sb) );
na02f02 TIMEBOOST_cell_36998 ( .a(TIMEBOOST_net_10737), .b(g58829_sb), .o(n_8609) );
na02f02 TIMEBOOST_cell_44409 ( .a(TIMEBOOST_net_10048), .b(g57322_sb), .o(TIMEBOOST_net_14443) );
na02f02 TIMEBOOST_cell_36980 ( .a(TIMEBOOST_net_10728), .b(g58801_sb), .o(n_8641) );
in01s01 g63090_u0 ( .a(FE_OFN1131_g64577_p), .o(g63090_sb) );
na02m02 TIMEBOOST_cell_41649 ( .a(wishbone_slave_unit_del_sync_bc_out_reg_1__Q), .b(n_1721), .o(TIMEBOOST_net_13063) );
na03s02 TIMEBOOST_cell_38237 ( .a(g64219_da), .b(g64219_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__Q), .o(TIMEBOOST_net_11357) );
in01s01 g63091_u0 ( .a(FE_OFN1104_g64577_p), .o(g63091_sb) );
na02s02 TIMEBOOST_cell_39444 ( .a(TIMEBOOST_net_11960), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_4499) );
na02s01 g63091_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__Q), .b(FE_OFN1104_g64577_p), .o(g63091_db) );
na02s01 TIMEBOOST_cell_37257 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__Q), .b(n_3739), .o(TIMEBOOST_net_10867) );
in01s01 g63092_u0 ( .a(FE_OFN2106_g64577_p), .o(g63092_sb) );
na02f02 TIMEBOOST_cell_41158 ( .a(TIMEBOOST_net_12817), .b(g57507_sb), .o(n_10325) );
na02s01 TIMEBOOST_cell_37614 ( .a(TIMEBOOST_net_11045), .b(g61731_sb), .o(n_8358) );
na02s01 TIMEBOOST_cell_37616 ( .a(TIMEBOOST_net_11046), .b(g61780_sb), .o(n_8246) );
in01s01 g63093_u0 ( .a(FE_OFN1119_g64577_p), .o(g63093_sb) );
na02s01 TIMEBOOST_cell_37491 ( .a(TIMEBOOST_net_9506), .b(FE_OFN1043_n_2037), .o(TIMEBOOST_net_10984) );
na02s01 TIMEBOOST_cell_37454 ( .a(TIMEBOOST_net_10965), .b(FE_OFN775_n_15366), .o(TIMEBOOST_net_10565) );
na02m02 TIMEBOOST_cell_38890 ( .a(TIMEBOOST_net_11683), .b(g58458_sb), .o(n_8989) );
in01s01 g63094_u0 ( .a(FE_OFN1200_n_4090), .o(g63094_sb) );
na02s01 TIMEBOOST_cell_36405 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__Q), .b(FE_OFN600_n_9687), .o(TIMEBOOST_net_10441) );
na03s01 TIMEBOOST_cell_34005 ( .a(conf_wb_err_addr_in_959), .b(g62119_sb), .c(g62119_db), .o(n_5577) );
na02s02 TIMEBOOST_cell_41770 ( .a(TIMEBOOST_net_13123), .b(g58285_db), .o(n_9033) );
in01s01 g63095_u0 ( .a(FE_OFN1106_g64577_p), .o(g63095_sb) );
na02s01 TIMEBOOST_cell_37259 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__Q), .b(n_3749), .o(TIMEBOOST_net_10868) );
na02s01 g63095_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__13__Q), .b(FE_OFN1106_g64577_p), .o(g63095_db) );
na02s02 TIMEBOOST_cell_39446 ( .a(TIMEBOOST_net_11961), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_4517) );
in01s01 g63096_u0 ( .a(FE_OFN881_g64577_p), .o(g63096_sb) );
na02s01 TIMEBOOST_cell_39464 ( .a(TIMEBOOST_net_11970), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_4609) );
na02m02 TIMEBOOST_cell_42201 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__Q), .b(n_9631), .o(TIMEBOOST_net_13339) );
na02s02 TIMEBOOST_cell_37215 ( .a(wishbone_slave_unit_pcim_if_del_we_in), .b(FE_OCPN1832_n_16949), .o(TIMEBOOST_net_10846) );
in01s01 g63097_u0 ( .a(FE_OFN1134_g64577_p), .o(g63097_sb) );
na03f02 TIMEBOOST_cell_35892 ( .a(TIMEBOOST_net_6209), .b(FE_OCPN1903_FE_OFN1061_n_16720), .c(FE_RN_411_0), .o(FE_RN_415_0) );
na02s02 TIMEBOOST_cell_38454 ( .a(TIMEBOOST_net_11465), .b(g54192_sb), .o(n_13425) );
no02f02 TIMEBOOST_cell_13083 ( .a(n_12220), .b(TIMEBOOST_net_3108), .o(n_12647) );
in01s01 g63098_u0 ( .a(FE_OFN1135_g64577_p), .o(g63098_sb) );
na03f02 TIMEBOOST_cell_35996 ( .a(TIMEBOOST_net_10114), .b(n_13617), .c(g54495_sb), .o(n_13595) );
na02m02 TIMEBOOST_cell_39159 ( .a(wbu_addr_in_270), .b(g58789_sb), .o(TIMEBOOST_net_11818) );
na03f02 TIMEBOOST_cell_35998 ( .a(TIMEBOOST_net_10112), .b(n_13617), .c(g54486_sb), .o(n_13613) );
in01s01 g63099_u0 ( .a(FE_OFN2106_g64577_p), .o(g63099_sb) );
na02s01 TIMEBOOST_cell_37493 ( .a(TIMEBOOST_net_9507), .b(FE_OFN1044_n_2037), .o(TIMEBOOST_net_10985) );
na02s01 TIMEBOOST_cell_42881 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q), .b(FE_OFN579_n_9531), .o(TIMEBOOST_net_13679) );
na02s01 TIMEBOOST_cell_42882 ( .a(TIMEBOOST_net_13679), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_11157) );
in01s01 g63100_u0 ( .a(FE_OFN877_g64577_p), .o(g63100_sb) );
na02f02 TIMEBOOST_cell_41650 ( .a(FE_OFN1437_n_9372), .b(TIMEBOOST_net_13063), .o(TIMEBOOST_net_11682) );
na02s02 TIMEBOOST_cell_43603 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__Q), .b(n_4338), .o(TIMEBOOST_net_14040) );
na02s01 TIMEBOOST_cell_41832 ( .a(g63614_da), .b(TIMEBOOST_net_13154), .o(n_7147) );
in01s01 g63101_u0 ( .a(FE_OFN1139_g64577_p), .o(g63101_sb) );
na02f04 TIMEBOOST_cell_45862 ( .a(TIMEBOOST_net_15169), .b(n_11913), .o(n_12810) );
na02s01 g63101_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__Q), .b(FE_OFN1107_g64577_p), .o(g63101_db) );
na02s01 TIMEBOOST_cell_41834 ( .a(g63611_da), .b(TIMEBOOST_net_13155), .o(n_7193) );
in01s01 g63102_u0 ( .a(FE_OFN1123_g64577_p), .o(g63102_sb) );
in01s01 TIMEBOOST_cell_45863 ( .a(TIMEBOOST_net_15170), .o(pci_target_unit_del_sync_sync_req_comp_pending) );
na02m02 TIMEBOOST_cell_32524 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__Q), .o(TIMEBOOST_net_10173) );
na02s04 TIMEBOOST_cell_45496 ( .a(TIMEBOOST_net_14986), .b(g54355_sb), .o(n_13125) );
in01s01 g63103_u0 ( .a(FE_OFN2104_g64577_p), .o(g63103_sb) );
na02s01 TIMEBOOST_cell_41836 ( .a(g63602_da), .b(TIMEBOOST_net_13156), .o(n_7185) );
na02s01 TIMEBOOST_cell_42568 ( .a(TIMEBOOST_net_13522), .b(g58126_sb), .o(TIMEBOOST_net_11198) );
na02f02 TIMEBOOST_cell_13103 ( .a(TIMEBOOST_net_3118), .b(n_12352), .o(n_12635) );
in01s01 g63104_u0 ( .a(FE_OFN1140_g64577_p), .o(g63104_sb) );
na02m02 TIMEBOOST_cell_41837 ( .a(FE_OFN1150_n_13249), .b(TIMEBOOST_net_9629), .o(TIMEBOOST_net_13157) );
na02s01 TIMEBOOST_cell_42569 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__Q), .b(FE_OFN602_n_9687), .o(TIMEBOOST_net_13523) );
in01s01 g63105_u0 ( .a(FE_OFN2105_g64577_p), .o(g63105_sb) );
na02s01 TIMEBOOST_cell_18169 ( .a(TIMEBOOST_net_4341), .b(g61915_sb), .o(n_7991) );
na02s01 TIMEBOOST_cell_42883 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__Q), .b(FE_OFN1651_n_9428), .o(TIMEBOOST_net_13680) );
na02s01 TIMEBOOST_cell_42884 ( .a(TIMEBOOST_net_13680), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_11159) );
in01s01 g63106_u0 ( .a(FE_OFN877_g64577_p), .o(g63106_sb) );
na02s04 TIMEBOOST_cell_45498 ( .a(TIMEBOOST_net_14987), .b(g54356_sb), .o(n_13086) );
na02s02 TIMEBOOST_cell_43119 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__31__Q), .b(n_4478), .o(TIMEBOOST_net_13798) );
na02m02 TIMEBOOST_cell_42827 ( .a(n_2710), .b(n_2301), .o(TIMEBOOST_net_13652) );
in01s01 g63107_u0 ( .a(FE_OFN1115_g64577_p), .o(g63107_sb) );
na02s02 TIMEBOOST_cell_43474 ( .a(TIMEBOOST_net_13975), .b(FE_OFN2064_n_6391), .o(TIMEBOOST_net_12195) );
na02s01 TIMEBOOST_cell_42570 ( .a(TIMEBOOST_net_13523), .b(g58117_sb), .o(TIMEBOOST_net_11938) );
in01s01 TIMEBOOST_cell_45880 ( .a(TIMEBOOST_net_15186), .o(TIMEBOOST_net_15187) );
in01s01 g63108_u0 ( .a(FE_OFN1242_n_4092), .o(g63108_sb) );
na02s01 TIMEBOOST_cell_36407 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__Q), .b(g65847_sb), .o(TIMEBOOST_net_10442) );
na02f02 TIMEBOOST_cell_41030 ( .a(TIMEBOOST_net_12753), .b(g57473_sb), .o(n_11261) );
in01s01 g63109_u0 ( .a(FE_OFN1118_g64577_p), .o(g63109_sb) );
na03s02 TIMEBOOST_cell_35912 ( .a(n_4609), .b(g61841_sb), .c(g61841_db), .o(n_6969) );
na02s01 TIMEBOOST_cell_42571 ( .a(FE_OFN205_n_9140), .b(g58270_sb), .o(TIMEBOOST_net_13524) );
na03f02 TIMEBOOST_cell_35914 ( .a(wbu_addr_in_274), .b(g52609_sb), .c(TIMEBOOST_net_10082), .o(n_11862) );
in01s01 g63110_u0 ( .a(FE_OFN1134_g64577_p), .o(g63110_sb) );
na03f02 TIMEBOOST_cell_35916 ( .a(wbu_addr_in_256), .b(g52620_sb), .c(TIMEBOOST_net_10084), .o(n_11850) );
na02s01 TIMEBOOST_cell_42572 ( .a(TIMEBOOST_net_13524), .b(g58270_db), .o(n_9036) );
na02f02 TIMEBOOST_cell_13123 ( .a(n_12049), .b(TIMEBOOST_net_3128), .o(n_12762) );
in01s01 g63111_u0 ( .a(FE_OFN1131_g64577_p), .o(g63111_sb) );
na02s02 TIMEBOOST_cell_45721 ( .a(n_4303), .b(n_26), .o(TIMEBOOST_net_15099) );
na02s01 TIMEBOOST_cell_42573 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__Q), .b(FE_OFN603_n_9687), .o(TIMEBOOST_net_13525) );
na02m04 TIMEBOOST_cell_45500 ( .a(TIMEBOOST_net_14988), .b(g54351_sb), .o(n_13090) );
in01s01 g63112_u0 ( .a(FE_OFN1121_g64577_p), .o(g63112_sb) );
na02f02 TIMEBOOST_cell_13129 ( .a(n_11838), .b(TIMEBOOST_net_3131), .o(n_17035) );
na02s01 TIMEBOOST_cell_42574 ( .a(TIMEBOOST_net_13525), .b(g58123_sb), .o(TIMEBOOST_net_11933) );
na03f06 TIMEBOOST_cell_35920 ( .a(g75178_db), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_), .c(FE_OCP_RBN2232_n_16273), .o(n_16550) );
in01s01 g63113_u0 ( .a(FE_OFN1137_g64577_p), .o(g63113_sb) );
no03f02 TIMEBOOST_cell_35922 ( .a(n_4649), .b(n_12595), .c(n_4877), .o(g59347_p) );
no02s02 TIMEBOOST_cell_42575 ( .a(TIMEBOOST_net_107), .b(n_1696), .o(TIMEBOOST_net_13526) );
na03s01 TIMEBOOST_cell_35924 ( .a(n_3226), .b(g60692_sb), .c(g60692_db), .o(n_7575) );
in01s01 g63114_u0 ( .a(FE_OFN1130_g64577_p), .o(g63114_sb) );
na02s01 TIMEBOOST_cell_42833 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__18__Q), .b(g65351_sb), .o(TIMEBOOST_net_13655) );
na02f02 TIMEBOOST_cell_41160 ( .a(TIMEBOOST_net_12818), .b(g57320_sb), .o(n_11431) );
na03s02 TIMEBOOST_cell_45715 ( .a(n_4276), .b(FE_OFN1248_n_4093), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__Q), .o(TIMEBOOST_net_15096) );
in01s01 g63115_u0 ( .a(FE_OFN1137_g64577_p), .o(g63115_sb) );
na02s01 TIMEBOOST_cell_37495 ( .a(TIMEBOOST_net_9509), .b(FE_OFN1044_n_2037), .o(TIMEBOOST_net_10986) );
na02s02 TIMEBOOST_cell_45716 ( .a(TIMEBOOST_net_15096), .b(g62907_sb), .o(n_6063) );
in01s01 g63116_u0 ( .a(FE_OFN1130_g64577_p), .o(g63116_sb) );
na02m02 TIMEBOOST_cell_44611 ( .a(n_9223), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__Q), .o(TIMEBOOST_net_14544) );
na02s01 TIMEBOOST_cell_37445 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__Q), .b(g58430_sb), .o(TIMEBOOST_net_10961) );
na02f02 TIMEBOOST_cell_44612 ( .a(TIMEBOOST_net_14544), .b(FE_OFN1427_n_8567), .o(TIMEBOOST_net_13017) );
in01s01 g63117_u0 ( .a(FE_OFN1095_g64577_p), .o(g63117_sb) );
na03s02 TIMEBOOST_cell_37183 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_26__Q), .b(FE_OFN2055_n_8831), .c(g58785_sb), .o(TIMEBOOST_net_10830) );
na02s01 g63117_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__Q), .b(FE_OFN1095_g64577_p), .o(g63117_db) );
na02s02 TIMEBOOST_cell_19157 ( .a(TIMEBOOST_net_4835), .b(g52876_sb), .o(TIMEBOOST_net_2310) );
in01s01 g63118_u0 ( .a(FE_OFN1136_g64577_p), .o(g63118_sb) );
na02s04 TIMEBOOST_cell_45502 ( .a(TIMEBOOST_net_14989), .b(g54352_sb), .o(n_13089) );
na02s01 TIMEBOOST_cell_37461 ( .a(pci_target_unit_del_sync_addr_in_213), .b(parchk_pci_ad_reg_in_1214), .o(TIMEBOOST_net_10969) );
in01s01 g63119_u0 ( .a(FE_OFN1132_g64577_p), .o(g63119_sb) );
na02m02 TIMEBOOST_cell_44613 ( .a(n_9501), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__Q), .o(TIMEBOOST_net_14545) );
na02f02 TIMEBOOST_cell_44714 ( .a(TIMEBOOST_net_14595), .b(n_11924), .o(n_12646) );
na02f02 TIMEBOOST_cell_44614 ( .a(TIMEBOOST_net_14545), .b(FE_OFN2188_n_8567), .o(TIMEBOOST_net_13012) );
in01s01 g63120_u0 ( .a(FE_OFN1119_g64577_p), .o(g63120_sb) );
na02f02 TIMEBOOST_cell_44715 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__Q), .b(FE_OFN1747_n_12004), .o(TIMEBOOST_net_14596) );
na02s01 TIMEBOOST_cell_42885 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__Q), .b(FE_OFN523_n_9428), .o(TIMEBOOST_net_13681) );
na02s01 TIMEBOOST_cell_42886 ( .a(TIMEBOOST_net_13681), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_11203) );
in01s01 g63121_u0 ( .a(FE_OFN1125_g64577_p), .o(g63121_sb) );
na02m02 TIMEBOOST_cell_44615 ( .a(n_9712), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__Q), .o(TIMEBOOST_net_14546) );
na02s01 TIMEBOOST_cell_37497 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__Q), .b(n_3774), .o(TIMEBOOST_net_10987) );
na02s01 TIMEBOOST_cell_42768 ( .a(TIMEBOOST_net_13622), .b(g65408_da), .o(TIMEBOOST_net_5439) );
in01s01 g63122_u0 ( .a(FE_OFN1112_g64577_p), .o(g63122_sb) );
na02s01 TIMEBOOST_cell_43079 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__Q), .b(n_4224), .o(TIMEBOOST_net_13778) );
na02f02 TIMEBOOST_cell_44729 ( .a(n_12283), .b(n_12002), .o(TIMEBOOST_net_14603) );
na02s04 TIMEBOOST_cell_45812 ( .a(TIMEBOOST_net_15144), .b(FE_OFN2136_n_13124), .o(TIMEBOOST_net_14986) );
in01s01 g63123_u0 ( .a(FE_OFN1131_g64577_p), .o(g63123_sb) );
na02s01 TIMEBOOST_cell_43258 ( .a(TIMEBOOST_net_13867), .b(FE_OFN1224_n_6391), .o(TIMEBOOST_net_12528) );
na02f02 TIMEBOOST_cell_44730 ( .a(TIMEBOOST_net_14603), .b(n_15936), .o(TIMEBOOST_net_679) );
na02s01 TIMEBOOST_cell_42680 ( .a(TIMEBOOST_net_13578), .b(g65094_db), .o(n_3596) );
in01s01 g63124_u0 ( .a(FE_OFN1106_g64577_p), .o(g63124_sb) );
na02s02 TIMEBOOST_cell_38305 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__Q), .b(g58357_sb), .o(TIMEBOOST_net_11391) );
na02s01 g63124_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__13__Q), .b(FE_OFN1106_g64577_p), .o(g63124_db) );
na02f04 TIMEBOOST_cell_39024 ( .a(TIMEBOOST_net_11750), .b(FE_OFN2243_g52675_p), .o(TIMEBOOST_net_10746) );
in01s01 g63125_u0 ( .a(FE_OFN1134_g64577_p), .o(g63125_sb) );
na02s02 TIMEBOOST_cell_44435 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_792), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_27__Q), .o(TIMEBOOST_net_14456) );
na02m04 TIMEBOOST_cell_45815 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_786), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_21__Q), .o(TIMEBOOST_net_15146) );
na02s04 TIMEBOOST_cell_45504 ( .a(TIMEBOOST_net_14990), .b(g54348_sb), .o(n_13094) );
in01s01 g63126_u0 ( .a(FE_OFN1106_g64577_p), .o(g63126_sb) );
na02f02 TIMEBOOST_cell_36982 ( .a(TIMEBOOST_net_10729), .b(g58813_sb), .o(n_8628) );
na02s01 g63126_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__16__Q), .b(FE_OFN1106_g64577_p), .o(g63126_db) );
na02f02 TIMEBOOST_cell_36984 ( .a(TIMEBOOST_net_10730), .b(g58812_sb), .o(n_8629) );
na02s02 TIMEBOOST_cell_10538 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_13__Q), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_1836) );
na02s01 g63127_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__Q), .b(FE_OFN1107_g64577_p), .o(g63127_db) );
na02s02 TIMEBOOST_cell_10539 ( .a(TIMEBOOST_net_1836), .b(FE_OFN1085_n_13221), .o(TIMEBOOST_net_557) );
in01s01 g63128_u0 ( .a(FE_OFN1115_g64577_p), .o(g63128_sb) );
na02s08 TIMEBOOST_cell_3025 ( .a(TIMEBOOST_net_92), .b(n_1715), .o(n_2218) );
na02m04 TIMEBOOST_cell_45816 ( .a(TIMEBOOST_net_15146), .b(FE_OFN2134_n_13124), .o(TIMEBOOST_net_14988) );
na02f02 TIMEBOOST_cell_36986 ( .a(TIMEBOOST_net_10731), .b(g58826_sb), .o(n_8615) );
na02s01 TIMEBOOST_cell_37475 ( .a(TIMEBOOST_net_9512), .b(FE_OFN1043_n_2037), .o(TIMEBOOST_net_10976) );
na02f02 TIMEBOOST_cell_36988 ( .a(TIMEBOOST_net_10732), .b(g58836_sb), .o(n_8601) );
in01s01 g63130_u0 ( .a(FE_OFN877_g64577_p), .o(g63130_sb) );
na02m02 TIMEBOOST_cell_43723 ( .a(n_9768), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__Q), .o(TIMEBOOST_net_14100) );
na02s01 TIMEBOOST_cell_37479 ( .a(TIMEBOOST_net_9510), .b(FE_OFN1043_n_2037), .o(TIMEBOOST_net_10978) );
na02f02 TIMEBOOST_cell_22169 ( .a(TIMEBOOST_net_6341), .b(FE_OFN1600_n_13995), .o(FE_RN_890_0) );
in01s01 g63131_u0 ( .a(FE_OFN1115_g64577_p), .o(g63131_sb) );
na02f02 TIMEBOOST_cell_41488 ( .a(TIMEBOOST_net_12982), .b(g57266_sb), .o(n_10418) );
na02s01 TIMEBOOST_cell_42887 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__Q), .b(FE_OFN533_n_9823), .o(TIMEBOOST_net_13682) );
na04m02 TIMEBOOST_cell_34766 ( .a(TIMEBOOST_net_4826), .b(g59801_sb), .c(g52451_sb), .d(g52451_db), .o(n_14840) );
in01s01 g63132_u0 ( .a(FE_OFN1118_g64577_p), .o(g63132_sb) );
na03s01 TIMEBOOST_cell_13185 ( .a(pci_target_unit_fifos_pcir_whole_waddr_94), .b(pci_target_unit_fifos_pcir_flush_in), .c(g57780_sb), .o(TIMEBOOST_net_620) );
na02m04 TIMEBOOST_cell_45810 ( .a(TIMEBOOST_net_15143), .b(FE_OFN2135_n_13124), .o(TIMEBOOST_net_14985) );
na02m04 TIMEBOOST_cell_45506 ( .a(TIMEBOOST_net_14991), .b(g54350_sb), .o(n_13091) );
in01s01 g63133_u0 ( .a(FE_OFN1131_g64577_p), .o(g63133_sb) );
na02f02 TIMEBOOST_cell_43724 ( .a(TIMEBOOST_net_14100), .b(FE_OFN1392_n_8567), .o(TIMEBOOST_net_12948) );
na02s01 TIMEBOOST_cell_18197 ( .a(TIMEBOOST_net_4355), .b(g61916_sb), .o(n_7989) );
na02m04 TIMEBOOST_cell_45825 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_783), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_18__Q), .o(TIMEBOOST_net_15151) );
in01s01 g63134_u0 ( .a(FE_OFN1137_g64577_p), .o(g63134_sb) );
in01s01 TIMEBOOST_cell_45876 ( .a(TIMEBOOST_net_15182), .o(TIMEBOOST_net_15183) );
na02s02 TIMEBOOST_cell_37447 ( .a(FE_OFN245_n_9114), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__Q), .o(TIMEBOOST_net_10962) );
na02f02 TIMEBOOST_cell_41204 ( .a(TIMEBOOST_net_12840), .b(g57073_sb), .o(n_11669) );
in01s01 g63135_u0 ( .a(FE_OFN1137_g64577_p), .o(g63135_sb) );
na02f02 TIMEBOOST_cell_44642 ( .a(TIMEBOOST_net_14559), .b(FE_OFN2175_n_8567), .o(TIMEBOOST_net_12334) );
na02s01 TIMEBOOST_cell_37449 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q), .b(FE_OFN217_n_9889), .o(TIMEBOOST_net_10963) );
na02m02 TIMEBOOST_cell_41509 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__Q), .b(n_9811), .o(TIMEBOOST_net_12993) );
in01s01 g63136_u0 ( .a(FE_OFN2105_g64577_p), .o(g63136_sb) );
na02s02 TIMEBOOST_cell_10559 ( .a(TIMEBOOST_net_1846), .b(g52881_sb), .o(TIMEBOOST_net_887) );
na02s01 TIMEBOOST_cell_42888 ( .a(TIMEBOOST_net_13682), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_11202) );
na02s01 TIMEBOOST_cell_42889 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__Q), .b(FE_OFN563_n_9895), .o(TIMEBOOST_net_13683) );
in01s01 g63137_u0 ( .a(FE_OFN1120_g64577_p), .o(g63137_sb) );
na02s02 TIMEBOOST_cell_10555 ( .a(TIMEBOOST_net_1844), .b(g52880_sb), .o(TIMEBOOST_net_888) );
na02s01 TIMEBOOST_cell_37594 ( .a(TIMEBOOST_net_11035), .b(g61730_sb), .o(n_8360) );
na02s02 TIMEBOOST_cell_36770 ( .a(TIMEBOOST_net_10623), .b(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_4580) );
in01s01 g63138_u0 ( .a(FE_OFN881_g64577_p), .o(g63138_sb) );
na02f02 TIMEBOOST_cell_36990 ( .a(TIMEBOOST_net_10733), .b(g58814_sb), .o(n_8627) );
na02s01 TIMEBOOST_cell_37453 ( .a(pci_target_unit_del_sync_addr_in_227), .b(parchk_pci_ad_reg_in_1228), .o(TIMEBOOST_net_10965) );
na02f02 TIMEBOOST_cell_37046 ( .a(TIMEBOOST_net_10761), .b(FE_OFN1769_n_14054), .o(g53239_p) );
in01s01 g63139_u0 ( .a(FE_OFN1125_g64577_p), .o(g63139_sb) );
na02s01 TIMEBOOST_cell_43135 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__Q), .b(n_3699), .o(TIMEBOOST_net_13806) );
na02s01 TIMEBOOST_cell_37385 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__Q), .b(n_3770), .o(TIMEBOOST_net_10931) );
na02s02 TIMEBOOST_cell_43097 ( .a(n_4357), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q), .o(TIMEBOOST_net_13787) );
in01s01 g63140_u0 ( .a(FE_OFN1129_g64577_p), .o(g63140_sb) );
na02s01 TIMEBOOST_cell_42623 ( .a(n_3783), .b(g64799_sb), .o(TIMEBOOST_net_13550) );
na02s01 TIMEBOOST_cell_37373 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__Q), .b(g58431_sb), .o(TIMEBOOST_net_10925) );
in01s01 g63141_u0 ( .a(FE_OFN881_g64577_p), .o(g63141_sb) );
na02s01 TIMEBOOST_cell_36792 ( .a(TIMEBOOST_net_10634), .b(FE_OFN1139_g64577_p), .o(TIMEBOOST_net_4398) );
na02s02 TIMEBOOST_cell_43259 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__Q), .b(n_1960), .o(TIMEBOOST_net_13868) );
na02s02 TIMEBOOST_cell_36794 ( .a(TIMEBOOST_net_10635), .b(n_3931), .o(n_4993) );
in01s01 g63142_u0 ( .a(FE_OFN1121_g64577_p), .o(g63142_sb) );
na02m02 TIMEBOOST_cell_44645 ( .a(n_9881), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__Q), .o(TIMEBOOST_net_14561) );
na02m02 TIMEBOOST_cell_32498 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__Q), .o(TIMEBOOST_net_10160) );
na02f02 TIMEBOOST_cell_45036 ( .a(TIMEBOOST_net_14756), .b(g54133_sb), .o(n_13466) );
in01s01 g63143_u0 ( .a(FE_OFN1129_g64577_p), .o(g63143_sb) );
na02f04 TIMEBOOST_cell_45508 ( .a(TIMEBOOST_net_14992), .b(g54345_sb), .o(n_12968) );
na02s01 TIMEBOOST_cell_37375 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__Q), .b(g58429_sb), .o(TIMEBOOST_net_10926) );
na02s02 TIMEBOOST_cell_30877 ( .a(TIMEBOOST_net_9349), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_3733) );
in01s01 g63144_u0 ( .a(FE_OFN1236_n_6391), .o(g63144_sb) );
na02m02 TIMEBOOST_cell_44079 ( .a(n_9458), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__Q), .o(TIMEBOOST_net_14278) );
na02f02 TIMEBOOST_cell_44080 ( .a(TIMEBOOST_net_14278), .b(FE_OFN1400_n_8567), .o(TIMEBOOST_net_12748) );
na02s01 TIMEBOOST_cell_44890 ( .a(TIMEBOOST_net_14683), .b(g65766_db), .o(n_1646) );
in01s01 g63145_u0 ( .a(FE_OFN1202_n_4090), .o(g63145_sb) );
na02s02 TIMEBOOST_cell_3281 ( .a(TIMEBOOST_net_220), .b(n_2424), .o(n_2490) );
na03s01 TIMEBOOST_cell_37377 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__25__Q), .b(FE_OFN666_n_4495), .c(n_3785), .o(TIMEBOOST_net_10927) );
na02s02 TIMEBOOST_cell_40833 ( .a(n_16763), .b(n_2328), .o(TIMEBOOST_net_12655) );
in01s01 g63146_u0 ( .a(FE_OFN1197_n_4090), .o(g63146_sb) );
na02s01 TIMEBOOST_cell_36409 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__Q), .b(FE_OFN600_n_9687), .o(TIMEBOOST_net_10443) );
na02s02 TIMEBOOST_cell_44971 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__Q), .b(FE_OFN252_n_9868), .o(TIMEBOOST_net_14724) );
na03f02 TIMEBOOST_cell_36000 ( .a(TIMEBOOST_net_10110), .b(n_13617), .c(g54488_sb), .o(n_13609) );
in01s01 g63147_u0 ( .a(FE_OFN1214_n_4151), .o(g63147_sb) );
na02s01 TIMEBOOST_cell_36411 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(g65718_sb), .o(TIMEBOOST_net_10444) );
na02f02 TIMEBOOST_cell_38786 ( .a(TIMEBOOST_net_11631), .b(g57300_db), .o(n_11451) );
na02s02 TIMEBOOST_cell_32164 ( .a(wbm_adr_o_21_), .b(FE_OFN1699_n_5751), .o(TIMEBOOST_net_9993) );
in01s01 g63148_u0 ( .a(FE_OFN1270_n_4095), .o(g63148_sb) );
no03f02 TIMEBOOST_cell_36413 ( .a(FE_RN_659_0), .b(FE_RN_665_0), .c(FE_RN_653_0), .o(TIMEBOOST_net_10445) );
na02s02 TIMEBOOST_cell_38756 ( .a(TIMEBOOST_net_11616), .b(g53928_sb), .o(n_13517) );
na02s02 TIMEBOOST_cell_41783 ( .a(g65093_sb), .b(g65093_db), .o(TIMEBOOST_net_13130) );
in01s01 g63149_u0 ( .a(FE_OFN1203_n_4090), .o(g63149_sb) );
na02s01 TIMEBOOST_cell_36415 ( .a(n_3030), .b(g67051_sb), .o(TIMEBOOST_net_10446) );
na03f02 TIMEBOOST_cell_36097 ( .a(FE_OCP_RBN1979_n_10273), .b(TIMEBOOST_net_10206), .c(FE_OFN1554_n_12104), .o(n_12760) );
na02f02 TIMEBOOST_cell_42332 ( .a(TIMEBOOST_net_13404), .b(g57090_sb), .o(n_11651) );
in01s01 g63150_u0 ( .a(FE_OFN1216_n_4151), .o(g63150_sb) );
na02s01 TIMEBOOST_cell_36417 ( .a(n_8511), .b(g65997_db), .o(TIMEBOOST_net_10447) );
na02s01 TIMEBOOST_cell_45066 ( .a(TIMEBOOST_net_14771), .b(FE_OFN270_n_9836), .o(TIMEBOOST_net_11179) );
in01s01 g63151_u0 ( .a(FE_OFN1276_n_4096), .o(g63151_sb) );
na02s01 TIMEBOOST_cell_3283 ( .a(TIMEBOOST_net_221), .b(n_4476), .o(n_4486) );
na02s01 TIMEBOOST_cell_37401 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__Q), .b(g58454_sb), .o(TIMEBOOST_net_10939) );
na02m02 TIMEBOOST_cell_40834 ( .a(TIMEBOOST_net_12655), .b(FE_OFN1330_n_13547), .o(TIMEBOOST_net_11604) );
in01s01 g63152_u0 ( .a(FE_OFN2104_g64577_p), .o(g63152_sb) );
na02s02 TIMEBOOST_cell_39297 ( .a(TIMEBOOST_net_3508), .b(FE_OFN1797_n_2299), .o(TIMEBOOST_net_11887) );
na02s01 TIMEBOOST_cell_42890 ( .a(TIMEBOOST_net_13683), .b(FE_OFN262_n_9851), .o(TIMEBOOST_net_11187) );
na02s01 TIMEBOOST_cell_42891 ( .a(FE_OFN258_n_9862), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__Q), .o(TIMEBOOST_net_13684) );
in01s01 g63153_u0 ( .a(FE_OFN1215_n_4151), .o(g63153_sb) );
na02s01 TIMEBOOST_cell_36419 ( .a(n_15302), .b(g65996_db), .o(TIMEBOOST_net_10448) );
na02s01 TIMEBOOST_cell_41810 ( .a(TIMEBOOST_net_13143), .b(FE_OFN1104_g64577_p), .o(TIMEBOOST_net_4311) );
na02s01 TIMEBOOST_cell_16796 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__Q), .b(g65343_sb), .o(TIMEBOOST_net_3655) );
in01s01 g63154_u0 ( .a(FE_OFN1192_n_6935), .o(g63154_sb) );
na02s01 TIMEBOOST_cell_3285 ( .a(TIMEBOOST_net_222), .b(n_4470), .o(n_4484) );
na02s01 g63154_u2 ( .a(n_3568), .b(FE_OFN1192_n_6935), .o(g63154_db) );
na02s01 TIMEBOOST_cell_42756 ( .a(TIMEBOOST_net_13616), .b(g57951_db), .o(n_9125) );
in01s01 g63155_u0 ( .a(FE_OFN1233_n_6391), .o(g63155_sb) );
na02s02 TIMEBOOST_cell_43444 ( .a(TIMEBOOST_net_13960), .b(FE_OFN1235_n_6391), .o(TIMEBOOST_net_12161) );
na02s02 TIMEBOOST_cell_3553 ( .a(TIMEBOOST_net_356), .b(FE_OFN264_n_9849), .o(n_9715) );
na02f02 TIMEBOOST_cell_32565 ( .a(n_12313), .b(TIMEBOOST_net_10193), .o(TIMEBOOST_net_6567) );
in01s01 g63156_u0 ( .a(FE_OFN1272_n_4096), .o(g63156_sb) );
na02s01 TIMEBOOST_cell_3287 ( .a(TIMEBOOST_net_223), .b(n_4482), .o(n_4483) );
na02s01 TIMEBOOST_cell_37395 ( .a(g64907_db), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__22__Q), .o(TIMEBOOST_net_10936) );
na02m02 TIMEBOOST_cell_32480 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__Q), .o(TIMEBOOST_net_10151) );
in01s01 g63157_u0 ( .a(FE_OFN1288_n_4098), .o(g63157_sb) );
na02s01 TIMEBOOST_cell_36421 ( .a(n_2648), .b(g65994_db), .o(TIMEBOOST_net_10449) );
na03s02 TIMEBOOST_cell_33039 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__17__Q), .b(FE_OFN671_n_4505), .c(g64750_sb), .o(TIMEBOOST_net_308) );
na02s02 TIMEBOOST_cell_42984 ( .a(TIMEBOOST_net_13730), .b(g61733_sb), .o(n_8353) );
in01s01 g63158_u0 ( .a(FE_OFN1243_n_4092), .o(g63158_sb) );
na02s01 TIMEBOOST_cell_36423 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__Q), .b(n_4417), .o(TIMEBOOST_net_10450) );
na02f02 TIMEBOOST_cell_42334 ( .a(TIMEBOOST_net_13405), .b(g57440_sb), .o(n_10351) );
na02s01 TIMEBOOST_cell_44837 ( .a(g65902_da), .b(g61953_db), .o(TIMEBOOST_net_14657) );
in01s02 g63159_u0 ( .a(FE_OFN1316_n_6624), .o(g63159_sb) );
na03s02 TIMEBOOST_cell_38143 ( .a(TIMEBOOST_net_4243), .b(g64209_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__Q), .o(TIMEBOOST_net_11310) );
na02s01 TIMEBOOST_cell_18505 ( .a(TIMEBOOST_net_4509), .b(g62806_sb), .o(n_5368) );
na02f02 TIMEBOOST_cell_38892 ( .a(TIMEBOOST_net_11684), .b(n_4641), .o(n_5728) );
in01s01 g63160_u0 ( .a(FE_OFN1313_n_6624), .o(g63160_sb) );
na02m02 TIMEBOOST_cell_44081 ( .a(n_9520), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__Q), .o(TIMEBOOST_net_14279) );
na02s02 TIMEBOOST_cell_43260 ( .a(TIMEBOOST_net_13868), .b(FE_OFN1264_n_4095), .o(TIMEBOOST_net_12054) );
na02s01 TIMEBOOST_cell_39182 ( .a(TIMEBOOST_net_11829), .b(g64315_db), .o(n_4515) );
in01s02 g63161_u0 ( .a(FE_OFN1317_n_6624), .o(g63161_sb) );
na03f02 TIMEBOOST_cell_39171 ( .a(FE_RN_313_0), .b(FE_RN_323_0), .c(FE_RN_354_0), .o(TIMEBOOST_net_11824) );
na02s01 TIMEBOOST_cell_38456 ( .a(TIMEBOOST_net_11466), .b(g58409_db), .o(n_9431) );
na02s01 TIMEBOOST_cell_18641 ( .a(TIMEBOOST_net_4577), .b(g63128_sb), .o(n_4996) );
in01s01 g63162_u0 ( .a(FE_OFN1242_n_4092), .o(g63162_sb) );
na02s01 TIMEBOOST_cell_36425 ( .a(g64896_sb), .b(g64896_db), .o(TIMEBOOST_net_10451) );
na02s02 TIMEBOOST_cell_37828 ( .a(TIMEBOOST_net_11152), .b(g58116_sb), .o(n_9677) );
na02s01 TIMEBOOST_cell_44838 ( .a(TIMEBOOST_net_14657), .b(TIMEBOOST_net_189), .o(n_7919) );
in01s01 g63163_u0 ( .a(FE_OFN1279_n_4097), .o(g63163_sb) );
na02f06 TIMEBOOST_cell_36427 ( .a(FE_RN_883_0), .b(FE_RN_836_0), .o(TIMEBOOST_net_10452) );
na02s02 TIMEBOOST_cell_37876 ( .a(TIMEBOOST_net_11176), .b(g57939_sb), .o(n_9871) );
na02s01 TIMEBOOST_cell_37423 ( .a(wbu_latency_tim_val_in), .b(n_6986), .o(TIMEBOOST_net_10950) );
in01s01 g63164_u0 ( .a(FE_OFN1225_n_6391), .o(g63164_sb) );
na02s02 TIMEBOOST_cell_3289 ( .a(TIMEBOOST_net_224), .b(n_4645), .o(n_4478) );
na02s01 TIMEBOOST_cell_37405 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__Q), .b(g58336_sb), .o(TIMEBOOST_net_10941) );
na02s02 TIMEBOOST_cell_40838 ( .a(TIMEBOOST_net_12657), .b(FE_OFN1331_n_13547), .o(TIMEBOOST_net_11606) );
in01s01 g63165_u0 ( .a(FE_OFN881_g64577_p), .o(g63165_sb) );
na02s02 TIMEBOOST_cell_19159 ( .a(TIMEBOOST_net_4836), .b(g52878_sb), .o(TIMEBOOST_net_2301) );
na02s01 TIMEBOOST_cell_39247 ( .a(pci_target_unit_fifos_pciw_addr_data_in_125), .b(g64153_sb), .o(TIMEBOOST_net_11862) );
na02s02 TIMEBOOST_cell_19161 ( .a(TIMEBOOST_net_4837), .b(g52877_sb), .o(TIMEBOOST_net_2309) );
in01s01 g63166_u0 ( .a(FE_OFN1295_n_4098), .o(g63166_sb) );
na03s02 TIMEBOOST_cell_36429 ( .a(n_1037), .b(n_1208), .c(n_1189), .o(TIMEBOOST_net_10453) );
na02s01 TIMEBOOST_cell_37422 ( .a(TIMEBOOST_net_10949), .b(g60674_sb), .o(TIMEBOOST_net_856) );
na02s01 TIMEBOOST_cell_37425 ( .a(wbu_latency_tim_val_in_247), .b(n_6986), .o(TIMEBOOST_net_10951) );
in01s01 g63167_u0 ( .a(FE_OFN1276_n_4096), .o(g63167_sb) );
na02s01 TIMEBOOST_cell_3291 ( .a(TIMEBOOST_net_225), .b(n_4442), .o(n_4468) );
na02s01 TIMEBOOST_cell_37407 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__Q), .b(g58451_sb), .o(TIMEBOOST_net_10942) );
na03f02 TIMEBOOST_cell_36096 ( .a(FE_RN_146_0), .b(n_10912), .c(n_12571), .o(n_12833) );
in01s01 g63168_u0 ( .a(FE_OFN1242_n_4092), .o(g63168_sb) );
na02s01 TIMEBOOST_cell_36431 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(g65713_sb), .o(TIMEBOOST_net_10454) );
na02s01 TIMEBOOST_cell_37424 ( .a(TIMEBOOST_net_10950), .b(g60690_sb), .o(TIMEBOOST_net_855) );
na02s01 TIMEBOOST_cell_37427 ( .a(wbu_latency_tim_val_in_245), .b(n_6986), .o(TIMEBOOST_net_10952) );
in01s01 g63169_u0 ( .a(FE_OFN1132_g64577_p), .o(g63169_sb) );
na02s01 TIMEBOOST_cell_30878 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__Q), .b(pci_target_unit_fifos_pcir_data_in_188), .o(TIMEBOOST_net_9350) );
na02s01 TIMEBOOST_cell_37409 ( .a(pci_target_unit_fifos_pcir_data_in_175), .b(g65788_sb), .o(TIMEBOOST_net_10943) );
na02m02 TIMEBOOST_cell_43725 ( .a(n_9704), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__Q), .o(TIMEBOOST_net_14101) );
in01s01 g63170_u0 ( .a(FE_OFN1118_g64577_p), .o(g63170_sb) );
na02m04 TIMEBOOST_cell_45510 ( .a(TIMEBOOST_net_14993), .b(g54347_sb), .o(n_13095) );
na02f02 TIMEBOOST_cell_22204 ( .a(FE_OCPN1877_n_13903), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q), .o(TIMEBOOST_net_6359) );
in01s01 g63171_u0 ( .a(FE_OFN1225_n_6391), .o(g63171_sb) );
na02s01 TIMEBOOST_cell_43261 ( .a(n_1718), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__Q), .o(TIMEBOOST_net_13869) );
na02f02 TIMEBOOST_cell_39113 ( .a(TIMEBOOST_net_10180), .b(FE_OCPN2219_n_13997), .o(TIMEBOOST_net_11795) );
na02s01 TIMEBOOST_cell_15866 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_89), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3190) );
in01s01 g63172_u0 ( .a(FE_OFN1112_g64577_p), .o(g63172_sb) );
na02m02 TIMEBOOST_cell_44279 ( .a(n_9013), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__Q), .o(TIMEBOOST_net_14378) );
na02s02 TIMEBOOST_cell_37411 ( .a(pci_target_unit_del_sync_bc_in_203), .b(g65211_sb), .o(TIMEBOOST_net_10944) );
in01s01 g63173_u0 ( .a(FE_OFN1194_n_6935), .o(g63173_sb) );
na02s01 TIMEBOOST_cell_15867 ( .a(TIMEBOOST_net_3190), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_402), .o(TIMEBOOST_net_62) );
na02f02 TIMEBOOST_cell_44716 ( .a(TIMEBOOST_net_14596), .b(n_11893), .o(n_12612) );
na02s01 TIMEBOOST_cell_3296 ( .a(FE_OFN611_n_4501), .b(g64981_db), .o(TIMEBOOST_net_228) );
in01s01 g63174_u0 ( .a(FE_OFN1206_n_6356), .o(g63174_sb) );
na02s01 TIMEBOOST_cell_3297 ( .a(TIMEBOOST_net_228), .b(n_4488), .o(n_4364) );
na02s02 TIMEBOOST_cell_37413 ( .a(g65225_sb), .b(pci_target_unit_del_sync_bc_in_202), .o(TIMEBOOST_net_10945) );
na02m02 TIMEBOOST_cell_38459 ( .a(g54187_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_406), .o(TIMEBOOST_net_11468) );
in01s01 g63175_u0 ( .a(FE_OFN1136_g64577_p), .o(g63175_sb) );
na02f02 TIMEBOOST_cell_43726 ( .a(TIMEBOOST_net_14101), .b(FE_OFN1399_n_8567), .o(TIMEBOOST_net_12697) );
na02s01 TIMEBOOST_cell_37415 ( .a(TIMEBOOST_net_9350), .b(FE_OFN956_n_1699), .o(TIMEBOOST_net_10946) );
na02s01 TIMEBOOST_cell_45698 ( .a(TIMEBOOST_net_15087), .b(FE_OFN1222_n_6391), .o(TIMEBOOST_net_13254) );
in01s01 g63176_u0 ( .a(FE_OFN1116_g64577_p), .o(g63176_sb) );
na02s02 TIMEBOOST_cell_39962 ( .a(TIMEBOOST_net_12219), .b(g62351_sb), .o(n_6898) );
na02s01 TIMEBOOST_cell_37383 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__Q), .b(n_3785), .o(TIMEBOOST_net_10930) );
na02m02 TIMEBOOST_cell_44223 ( .a(n_9867), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__Q), .o(TIMEBOOST_net_14350) );
in01s01 g63177_u0 ( .a(FE_OFN1230_n_6391), .o(g63177_sb) );
in01s01 TIMEBOOST_cell_45933 ( .a(wbm_dat_i_25_), .o(TIMEBOOST_net_15240) );
na02f02 TIMEBOOST_cell_44082 ( .a(TIMEBOOST_net_14279), .b(FE_OFN1411_n_8567), .o(TIMEBOOST_net_12749) );
na02m02 TIMEBOOST_cell_32564 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__Q), .o(TIMEBOOST_net_10193) );
in01s01 g63178_u0 ( .a(FE_OFN1310_n_6624), .o(g63178_sb) );
na02f02 TIMEBOOST_cell_12786 ( .a(n_13903), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q), .o(TIMEBOOST_net_2960) );
na03s02 TIMEBOOST_cell_38069 ( .a(TIMEBOOST_net_3711), .b(g64289_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q), .o(TIMEBOOST_net_11273) );
na02s02 TIMEBOOST_cell_22295 ( .a(n_10157), .b(TIMEBOOST_net_6404), .o(n_11855) );
in01s01 g63179_u0 ( .a(FE_OFN1095_g64577_p), .o(g63179_sb) );
na02s02 TIMEBOOST_cell_36796 ( .a(TIMEBOOST_net_10636), .b(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_4626) );
na02s01 g63179_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__Q), .b(FE_OFN1095_g64577_p), .o(g63179_db) );
na02s02 TIMEBOOST_cell_36798 ( .a(TIMEBOOST_net_10637), .b(FE_OFN1126_g64577_p), .o(TIMEBOOST_net_4495) );
in01s01 g63180_u0 ( .a(FE_OFN1215_n_4151), .o(g63180_sb) );
na02s01 TIMEBOOST_cell_36433 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(g65782_sb), .o(TIMEBOOST_net_10455) );
na02s01 TIMEBOOST_cell_37426 ( .a(TIMEBOOST_net_10951), .b(g60672_sb), .o(TIMEBOOST_net_864) );
na02f02 TIMEBOOST_cell_41112 ( .a(TIMEBOOST_net_12794), .b(g57095_sb), .o(n_10843) );
in01s01 g63181_u0 ( .a(FE_OFN1272_n_4096), .o(g63181_sb) );
na02s02 TIMEBOOST_cell_43026 ( .a(TIMEBOOST_net_13751), .b(g62864_db), .o(n_5237) );
na02s01 TIMEBOOST_cell_37387 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__Q), .b(n_3777), .o(TIMEBOOST_net_10932) );
na02s02 TIMEBOOST_cell_38458 ( .a(TIMEBOOST_net_11467), .b(g58340_db), .o(n_9480) );
in01s01 g63182_u0 ( .a(FE_OFN1130_g64577_p), .o(g63182_sb) );
na02s01 TIMEBOOST_cell_43262 ( .a(TIMEBOOST_net_13869), .b(FE_OFN1225_n_6391), .o(TIMEBOOST_net_12536) );
na02s01 TIMEBOOST_cell_37417 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__Q), .b(n_3749), .o(TIMEBOOST_net_10947) );
na02s01 TIMEBOOST_cell_4280 ( .a(configuration_sync_command_bit2), .b(wbu_wb_init_complete_in), .o(TIMEBOOST_net_720) );
in01s01 g63183_u0 ( .a(FE_OFN1194_n_6935), .o(g63183_sb) );
na02s01 TIMEBOOST_cell_3301 ( .a(TIMEBOOST_net_230), .b(n_4498), .o(n_4338) );
na02s01 TIMEBOOST_cell_37389 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__Q), .b(n_3777), .o(TIMEBOOST_net_10933) );
na02s06 TIMEBOOST_cell_3302 ( .a(n_3222), .b(n_4743), .o(TIMEBOOST_net_231) );
in01s01 g63184_u0 ( .a(FE_OFN1212_n_4151), .o(g63184_sb) );
na02s01 TIMEBOOST_cell_36435 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(g65760_sb), .o(TIMEBOOST_net_10456) );
na02f02 TIMEBOOST_cell_44725 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__Q), .b(n_13873), .o(TIMEBOOST_net_14601) );
na02s01 TIMEBOOST_cell_37428 ( .a(TIMEBOOST_net_10952), .b(g59226_sb), .o(TIMEBOOST_net_851) );
in01s01 g63185_u0 ( .a(FE_OFN1203_n_4090), .o(g63185_sb) );
na02s01 TIMEBOOST_cell_36441 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(g63537_sb), .o(TIMEBOOST_net_10459) );
na02s01 TIMEBOOST_cell_36463 ( .a(pci_target_unit_fifos_pcir_data_in_172), .b(g65784_sb), .o(TIMEBOOST_net_10470) );
na02s01 TIMEBOOST_cell_36462 ( .a(TIMEBOOST_net_10469), .b(g65761_sb), .o(n_1943) );
in01s01 g63186_u0 ( .a(n_6431), .o(g63186_sb) );
na03s02 TIMEBOOST_cell_38141 ( .a(TIMEBOOST_net_4003), .b(g64223_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__Q), .o(TIMEBOOST_net_11309) );
na02s01 TIMEBOOST_cell_3435 ( .a(TIMEBOOST_net_297), .b(g58051_sb), .o(n_9088) );
na02f02 TIMEBOOST_cell_44636 ( .a(TIMEBOOST_net_14556), .b(FE_OFN2169_n_8567), .o(TIMEBOOST_net_13483) );
in01s01 g63187_u0 ( .a(FE_OFN1285_n_4097), .o(g63187_sb) );
na02s01 TIMEBOOST_cell_36443 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(g64199_sb), .o(TIMEBOOST_net_10460) );
na02f02 TIMEBOOST_cell_44727 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__20__Q), .b(TIMEBOOST_net_6570), .o(TIMEBOOST_net_14602) );
na02m02 TIMEBOOST_cell_43727 ( .a(n_9878), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q), .o(TIMEBOOST_net_14102) );
in01s01 g63188_u0 ( .a(FE_OFN1130_g64577_p), .o(g63188_sb) );
na02s01 TIMEBOOST_cell_4281 ( .a(TIMEBOOST_net_720), .b(n_709), .o(TIMEBOOST_net_485) );
na02f02 g53813_u0 ( .a(n_13466), .b(n_2114), .o(n_13672) );
na02s01 TIMEBOOST_cell_40738 ( .a(TIMEBOOST_net_12607), .b(g62471_sb), .o(n_6649) );
in01s01 g63189_u0 ( .a(FE_OFN1269_n_4095), .o(g63189_sb) );
na02s02 TIMEBOOST_cell_19083 ( .a(TIMEBOOST_net_4798), .b(g58361_db), .o(n_9462) );
na02m04 TIMEBOOST_cell_45512 ( .a(TIMEBOOST_net_14994), .b(g54344_sb), .o(n_13097) );
na02s02 TIMEBOOST_cell_42010 ( .a(TIMEBOOST_net_13243), .b(g62650_sb), .o(n_6246) );
in01s01 g63190_u0 ( .a(FE_OFN1212_n_4151), .o(g63190_sb) );
no02m02 TIMEBOOST_cell_36365 ( .a(n_2430), .b(TIMEBOOST_net_116), .o(TIMEBOOST_net_10421) );
na02f02 TIMEBOOST_cell_41620 ( .a(FE_OFN1440_n_9372), .b(TIMEBOOST_net_13048), .o(TIMEBOOST_net_11663) );
na02s01 TIMEBOOST_cell_42731 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__Q), .b(n_1578), .o(TIMEBOOST_net_13604) );
in01s01 g63191_u0 ( .a(FE_OFN1121_g64577_p), .o(g63191_sb) );
na02m02 g53820_u0 ( .a(n_13460), .b(n_2116), .o(n_13667) );
na02s02 TIMEBOOST_cell_43120 ( .a(TIMEBOOST_net_13798), .b(FE_OFN1212_n_4151), .o(TIMEBOOST_net_12100) );
in01s01 g63192_u0 ( .a(FE_OFN1202_n_4090), .o(g63192_sb) );
na02m02 TIMEBOOST_cell_3303 ( .a(TIMEBOOST_net_231), .b(n_2447), .o(n_8521) );
na02s02 TIMEBOOST_cell_43644 ( .a(TIMEBOOST_net_14060), .b(FE_OFN1316_n_6624), .o(TIMEBOOST_net_12227) );
na02s01 TIMEBOOST_cell_43322 ( .a(TIMEBOOST_net_13899), .b(g62526_sb), .o(n_6523) );
in01s01 g63193_u0 ( .a(FE_OFN1142_n_15261), .o(g63193_sb) );
na02s02 TIMEBOOST_cell_37686 ( .a(TIMEBOOST_net_11081), .b(g61944_sb), .o(n_7937) );
na02f02 TIMEBOOST_cell_44701 ( .a(TIMEBOOST_net_10098), .b(FE_OFN1472_g52675_p), .o(TIMEBOOST_net_14589) );
na02f04 TIMEBOOST_cell_45856 ( .a(TIMEBOOST_net_15166), .b(n_12440), .o(n_12773) );
in01s01 g63194_u0 ( .a(n_5546), .o(g63194_sb) );
na02s01 TIMEBOOST_cell_37253 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__Q), .b(wishbone_slave_unit_fifos_wbr_control_in), .o(TIMEBOOST_net_10865) );
na02s01 TIMEBOOST_cell_16041 ( .a(TIMEBOOST_net_3277), .b(n_2499), .o(n_2500) );
in01m01 g63195_u0 ( .a(FE_OFN1142_n_15261), .o(g63195_sb) );
na02s01 TIMEBOOST_cell_39184 ( .a(TIMEBOOST_net_11830), .b(g65904_db), .o(n_2177) );
na02s02 g63195_u2 ( .a(FE_OFN1142_n_15261), .b(conf_wb_err_addr_in_944), .o(g63195_db) );
na02s01 TIMEBOOST_cell_18465 ( .a(TIMEBOOST_net_4489), .b(g63102_sb), .o(n_5050) );
in01s01 g63196_u0 ( .a(FE_OFN1143_n_15261), .o(g63196_sb) );
na03s02 TIMEBOOST_cell_38223 ( .a(TIMEBOOST_net_3999), .b(g64098_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__Q), .o(TIMEBOOST_net_11350) );
na02s02 g63196_u2 ( .a(conf_wb_err_addr_in_949), .b(FE_OFN1144_n_15261), .o(g63196_db) );
na02m02 TIMEBOOST_cell_38836 ( .a(TIMEBOOST_net_11656), .b(g58480_sb), .o(n_9355) );
in01s01 g63197_u0 ( .a(FE_OFN1192_n_6935), .o(g63197_sb) );
na02s02 TIMEBOOST_cell_3305 ( .a(TIMEBOOST_net_232), .b(n_4488), .o(n_4489) );
na02s01 g63197_u2 ( .a(n_5769), .b(FE_OFN1192_n_6935), .o(g63197_db) );
na03s02 TIMEBOOST_cell_34478 ( .a(wbm_adr_o_19_), .b(FE_OFN1699_n_5751), .c(g61856_sb), .o(TIMEBOOST_net_593) );
in01s01 g63198_u0 ( .a(FE_OFN1192_n_6935), .o(g63198_sb) );
na02s01 TIMEBOOST_cell_31241 ( .a(TIMEBOOST_net_9531), .b(g64952_db), .o(n_4378) );
na02s01 g63198_u2 ( .a(n_1199), .b(FE_OFN1192_n_6935), .o(g63198_db) );
na02s01 TIMEBOOST_cell_31240 ( .a(n_4479), .b(g64952_sb), .o(TIMEBOOST_net_9531) );
in01s01 g63199_u0 ( .a(FE_OFN1192_n_6935), .o(g63199_sb) );
na02s01 TIMEBOOST_cell_31239 ( .a(TIMEBOOST_net_9530), .b(g64950_db), .o(n_3666) );
na02s01 g63199_u2 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .b(FE_OFN1192_n_6935), .o(g63199_db) );
na02s02 TIMEBOOST_cell_15908 ( .a(wbs_we_i), .b(n_1347), .o(TIMEBOOST_net_3211) );
no02m02 g63200_u0 ( .a(wbm_adr_o_16_), .b(n_2442), .o(g63200_p) );
ao12m02 g63200_u1 ( .a(g63200_p), .b(wbm_adr_o_16_), .c(n_2442), .o(n_3152) );
no02s02 g63201_u0 ( .a(wbu_addr_in_265), .b(n_2438), .o(g63201_p) );
ao12m02 g63201_u1 ( .a(g63201_p), .b(wbu_addr_in_265), .c(n_2438), .o(n_3151) );
in01m01 g63202_u0 ( .a(FE_OFN1697_n_5751), .o(g63202_sb) );
na02s01 TIMEBOOST_cell_37241 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__23__Q), .b(n_3741), .o(TIMEBOOST_net_10859) );
na02s01 TIMEBOOST_cell_19022 ( .a(wishbone_slave_unit_pcim_sm_data_in_648), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__Q), .o(TIMEBOOST_net_4768) );
na02s01 TIMEBOOST_cell_37260 ( .a(TIMEBOOST_net_10868), .b(FE_OFN687_n_4417), .o(TIMEBOOST_net_9390) );
in01m01 g63203_u0 ( .a(FE_OFN1697_n_5751), .o(g63203_sb) );
na02s01 TIMEBOOST_cell_37261 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__Q), .b(n_3761), .o(TIMEBOOST_net_10869) );
na02s01 TIMEBOOST_cell_19024 ( .a(wishbone_slave_unit_pcim_sm_data_in_644), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__Q), .o(TIMEBOOST_net_4769) );
na02s01 TIMEBOOST_cell_37262 ( .a(TIMEBOOST_net_10869), .b(FE_OFN686_n_4417), .o(TIMEBOOST_net_9388) );
in01m01 g63204_u0 ( .a(FE_OFN1700_n_5751), .o(g63204_sb) );
no02s01 TIMEBOOST_cell_42576 ( .a(TIMEBOOST_net_13526), .b(n_1635), .o(TIMEBOOST_net_3369) );
na02s02 TIMEBOOST_cell_11480 ( .a(n_2693), .b(FE_OFN1700_n_5751), .o(TIMEBOOST_net_2307) );
na02s02 TIMEBOOST_cell_19243 ( .a(TIMEBOOST_net_4878), .b(g60652_sb), .o(n_5672) );
no02s01 g63206_u0 ( .a(n_416), .b(n_1659), .o(g63206_p) );
ao12s02 g63206_u1 ( .a(g63206_p), .b(n_416), .c(n_1659), .o(n_2014) );
no02s01 g63207_u0 ( .a(pci_target_unit_fifos_pciw_inTransactionCount_0_), .b(n_5546), .o(g63207_p) );
ao12s01 g63207_u1 ( .a(g63207_p), .b(pci_target_unit_fifos_pciw_inTransactionCount_0_), .c(n_5546), .o(n_4797) );
no02s01 g63208_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_10_), .b(n_2473), .o(g63208_p) );
ao12s01 g63208_u1 ( .a(g63208_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_10_), .c(n_2473), .o(n_2965) );
no02s01 g63209_u0 ( .a(n_207), .b(n_2477), .o(g63209_p) );
ao12s01 g63209_u1 ( .a(g63209_p), .b(n_207), .c(n_2477), .o(n_2964) );
in01s01 g63213_u0 ( .a(FE_OFN191_n_1193), .o(n_2284) );
ao22s06 g63214_u0 ( .a(pci_irdy_i), .b(n_961), .c(parchk_pci_irdy_en_in), .d(out_bckp_irdy_out), .o(n_1193) );
no02f02 g63215_u0 ( .a(n_2254), .b(n_2249), .o(g63215_p) );
ao12f02 g63215_u1 ( .a(g63215_p), .b(n_2254), .c(n_2249), .o(n_2963) );
no02f03 g63216_u0 ( .a(n_2253), .b(n_2251), .o(g63216_p) );
ao12f04 g63216_u1 ( .a(g63216_p), .b(n_2253), .c(n_2251), .o(n_2962) );
no02f02 g63217_u0 ( .a(n_2252), .b(n_2255), .o(g63217_p) );
ao12f04 g63217_u1 ( .a(g63217_p), .b(n_2252), .c(n_2255), .o(n_2961) );
na02s01 g63226_u0 ( .a(n_4795), .b(n_1684), .o(n_4796) );
no02s01 g63227_u0 ( .a(n_2959), .b(n_2412), .o(n_2960) );
in01s01 g63228_u0 ( .a(n_3157), .o(n_2958) );
no02m01 g63229_u0 ( .a(n_15390), .b(n_705), .o(TIMEBOOST_net_10322) );
in01f06 g63230_u0 ( .a(n_4149), .o(n_5592) );
in01f03 g63245_u0 ( .a(n_4149), .o(n_5633) );
no02f04 g63250_u0 ( .a(n_3120), .b(FE_OCPN1838_n_1238), .o(n_4149) );
na02m02 g63251_u0 ( .a(n_3271), .b(n_4743), .o(n_8450) );
na02f06 g63252_u0 ( .a(n_2013), .b(wbu_addr_in_254), .o(g63252_p) );
in01f04 g63252_u1 ( .a(g63252_p), .o(n_2487) );
na02m04 g63253_u0 ( .a(n_2012), .b(wbm_adr_o_5_), .o(g63253_p) );
in01m04 g63253_u1 ( .a(g63253_p), .o(n_2485) );
na02m08 g63254_u0 ( .a(n_1669), .b(conf_wb_err_addr_in_946), .o(n_2035) );
na02s06 g63255_u0 ( .a(FE_OFN2245_n_4792), .b(n_2950), .o(n_4793) );
na02f08 g63256_u0 ( .a(n_2897), .b(n_4743), .o(g63256_p) );
in01f10 g63256_u1 ( .a(g63256_p), .o(n_16916) );
na02f02 TIMEBOOST_cell_44717 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__Q), .b(FE_OFN1747_n_12004), .o(TIMEBOOST_net_14597) );
na03s02 TIMEBOOST_cell_33373 ( .a(n_4465), .b(g64940_sb), .c(g64940_db), .o(n_4382) );
na02s03 g63259_u0 ( .a(n_1438), .b(pci_target_unit_del_sync_comp_cycle_count_3_), .o(g63259_p) );
in01s02 g63259_u1 ( .a(g63259_p), .o(n_1692) );
no02s03 g63261_u0 ( .a(n_1226), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_3_), .o(n_1714) );
na02m02 g63263_u0 ( .a(n_1476), .b(wishbone_slave_unit_del_sync_comp_cycle_count_3_), .o(g63263_p) );
in01m02 g63263_u1 ( .a(g63263_p), .o(n_1694) );
na02m01 g63264_u0 ( .a(n_4939), .b(FE_OFN1192_n_6935), .o(n_7136) );
in01f02 g63265_u0 ( .a(n_2956), .o(n_2957) );
no02f04 g63266_u0 ( .a(n_15390), .b(n_2215), .o(n_2956) );
no02m01 g63267_u0 ( .a(n_15390), .b(n_3267), .o(n_4177) );
na02f02 g63268_u0 ( .a(n_5230), .b(n_3406), .o(g63268_p) );
in01f02 g63268_u1 ( .a(g63268_p), .o(n_4654) );
na02f02 g63269_u0 ( .a(n_3117), .b(n_3245), .o(n_4146) );
na02s01 g63270_u0 ( .a(n_4662), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_3_), .o(n_3455) );
no02m06 g63271_u0 ( .a(n_15390), .b(n_2966), .o(g63271_p) );
in01f02 g63271_u1 ( .a(g63271_p), .o(n_3342) );
no02s06 g63272_u0 ( .a(n_8440), .b(n_3388), .o(n_7809) );
na02f02 TIMEBOOST_cell_41534 ( .a(TIMEBOOST_net_13005), .b(g57283_sb), .o(n_11472) );
no02f04 g63275_u0 ( .a(n_3090), .b(n_8440), .o(n_7803) );
na02s01 g63276_u0 ( .a(n_8440), .b(configuration_interrupt_line_39), .o(n_7565) );
na02s01 g63277_u0 ( .a(n_8440), .b(configuration_interrupt_line_40), .o(n_7564) );
na02s01 g63278_u0 ( .a(n_8440), .b(configuration_interrupt_line_41), .o(n_7562) );
na02s01 TIMEBOOST_cell_37180 ( .a(TIMEBOOST_net_10828), .b(g56934_sb), .o(TIMEBOOST_net_6388) );
in01f06 g63280_u0 ( .a(n_4685), .o(n_7398) );
in01f06 g63284_u0 ( .a(n_15919), .o(n_4685) );
na02f02 g63287_u0 ( .a(n_3109), .b(n_3247), .o(n_4144) );
na02s01 g63288_u0 ( .a(n_8440), .b(configuration_interrupt_line_43), .o(n_7561) );
na02f02 g63289_u0 ( .a(n_3409), .b(n_16160), .o(n_7321) );
na03f02 g63290_u0 ( .a(n_2852), .b(n_3285), .c(n_3057), .o(n_4649) );
na02f02 g63291_u0 ( .a(n_2920), .b(n_3116), .o(g63291_p) );
in01f02 g63291_u1 ( .a(g63291_p), .o(n_3454) );
na02f04 g63292_u0 ( .a(n_2013), .b(n_964), .o(g63292_p) );
in01f04 g63292_u1 ( .a(g63292_p), .o(n_2680) );
no02s02 g63293_u0 ( .a(n_8440), .b(n_4720), .o(g63293_p) );
in01s02 g63293_u1 ( .a(g63293_p), .o(n_8446) );
na02s01 g63294_u0 ( .a(n_8440), .b(wbu_cache_line_size_in_208), .o(n_7560) );
na02s01 TIMEBOOST_cell_42064 ( .a(TIMEBOOST_net_13270), .b(g62350_sb), .o(n_6900) );
na02m02 g63297_u0 ( .a(n_2954), .b(wbu_addr_in_273), .o(n_2955) );
na02m02 g63298_u0 ( .a(n_3147), .b(wbu_addr_in_276), .o(n_3148) );
na03s02 TIMEBOOST_cell_36781 ( .a(g64356_da), .b(g64356_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__Q), .o(TIMEBOOST_net_10629) );
no02f04 TIMEBOOST_cell_30834 ( .a(n_1403), .b(n_1397), .o(TIMEBOOST_net_9328) );
no02s10 g63301_u0 ( .a(n_3278), .b(n_8440), .o(n_7466) );
na02s01 TIMEBOOST_cell_45015 ( .a(n_15), .b(g65304_sb), .o(TIMEBOOST_net_14746) );
na02m02 TIMEBOOST_cell_30750 ( .a(n_976), .b(g66457_sb), .o(TIMEBOOST_net_9286) );
na02s02 TIMEBOOST_cell_42728 ( .a(TIMEBOOST_net_13602), .b(n_8892), .o(TIMEBOOST_net_10979) );
na02m02 TIMEBOOST_cell_38460 ( .a(TIMEBOOST_net_11468), .b(TIMEBOOST_net_563), .o(n_13428) );
in01s02 g63307_u1 ( .a(g63307_p), .o(n_3450) );
na02s02 g63309_u0 ( .a(n_8440), .b(wbu_cache_line_size_in_207), .o(n_7559) );
na02s03 g63310_u0 ( .a(n_853), .b(n_5546), .o(n_5545) );
in01s01 g63313_u0 ( .a(n_3448), .o(n_3449) );
no02f08 g63314_u0 ( .a(n_16280), .b(n_3319), .o(n_3448) );
na02m04 g63315_u0 ( .a(FE_OFN1143_n_15261), .b(n_4535), .o(g63315_p) );
in01m06 g63315_u1 ( .a(g63315_p), .o(n_13825) );
na02s02 g63316_u0 ( .a(FE_OFN1142_n_15261), .b(conf_wb_err_addr_in_943), .o(n_3327) );
in01m02 g63318_u0 ( .a(n_2011), .o(n_2458) );
na02f02 TIMEBOOST_cell_42262 ( .a(TIMEBOOST_net_13369), .b(FE_OFN1421_n_8567), .o(TIMEBOOST_net_12323) );
no02s01 g63320_u0 ( .a(n_1424), .b(FE_OFN778_n_4152), .o(n_2953) );
no02s01 g63321_u0 ( .a(FE_OCPN1841_n_16089), .b(n_8498), .o(n_2725) );
no02s02 g63322_u0 ( .a(n_2423), .b(FE_OFN778_n_4152), .o(n_2952) );
no02s02 g63323_u0 ( .a(n_1673), .b(FE_OFN1143_n_15261), .o(n_3326) );
ao12s01 g63324_u0 ( .a(n_4536), .b(n_2370), .c(n_4718), .o(n_4936) );
no02f04 g63338_u0 ( .a(n_15054), .b(n_2354), .o(g63338_p) );
in01f04 g63338_u1 ( .a(g63338_p), .o(n_5763) );
na02s01 g63339_u0 ( .a(n_8440), .b(wbu_cache_line_size_in_209), .o(n_7558) );
na02s02 g63340_u0 ( .a(n_2280), .b(FE_OFN199_n_3298), .o(g63340_p) );
in01s01 g63340_u1 ( .a(g63340_p), .o(n_4142) );
na02m02 g63341_u0 ( .a(n_3324), .b(wbm_adr_o_27_), .o(n_3325) );
na02s01 g63342_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_0_), .b(n_4662), .o(n_3447) );
na02s02 g63343_u0 ( .a(n_4662), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_1_), .o(n_3446) );
na02s01 g63344_u0 ( .a(n_4662), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_5_), .o(n_3445) );
na02s02 TIMEBOOST_cell_38591 ( .a(TIMEBOOST_net_9944), .b(FE_OFN1179_n_3476), .o(TIMEBOOST_net_11534) );
na02f02 g63348_u0 ( .a(n_2012), .b(n_1116), .o(g63348_p) );
in01f02 g63348_u1 ( .a(g63348_p), .o(n_2738) );
na02f08 g63349_u0 ( .a(n_2950), .b(n_1435), .o(n_2951) );
na02m01 g63350_u0 ( .a(n_2018), .b(pci_target_unit_wishbone_master_rty_counter_7_), .o(n_2019) );
no02m02 g63351_u0 ( .a(FE_OFN1142_n_15261), .b(n_2395), .o(n_3323) );
na02s01 g63352_u0 ( .a(n_8440), .b(wbu_cache_line_size_in_211), .o(n_7557) );
na02s01 g63353_u0 ( .a(n_4662), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_2_), .o(n_3444) );
na02s01 g63354_u0 ( .a(n_3020), .b(parity_checker_check_for_serr_on_second), .o(n_7396) );
na02s02 g63355_u0 ( .a(n_2948), .b(wbm_adr_o_24_), .o(n_2949) );
na02s01 g63356_u0 ( .a(n_4662), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_6_), .o(n_3443) );
in01s01 g63358_u0 ( .a(n_7795), .o(n_7785) );
no02m08 g63359_u0 ( .a(n_8440), .b(n_3261), .o(n_7795) );
na02s02 TIMEBOOST_cell_39964 ( .a(TIMEBOOST_net_12220), .b(g62622_sb), .o(n_6313) );
na02s01 g63361_u0 ( .a(wishbone_slave_unit_del_sync_comp_rty_exp_clr), .b(wishbone_slave_unit_del_sync_comp_rty_exp_reg), .o(g63361_p) );
in01s01 g63361_u1 ( .a(g63361_p), .o(n_4140) );
na02f02 g63362_u0 ( .a(n_15733), .b(n_5230), .o(g63362_p) );
in01f02 g63362_u1 ( .a(g63362_p), .o(n_4641) );
na02s01 TIMEBOOST_cell_39434 ( .a(TIMEBOOST_net_11955), .b(g62007_sb), .o(n_7881) );
no02m02 g63364_u0 ( .a(n_8440), .b(FE_OFN2100_n_3281), .o(g63364_p) );
in01m02 g63364_u1 ( .a(g63364_p), .o(n_8444) );
na02m02 TIMEBOOST_cell_41635 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_30__Q), .b(FE_OFN239_n_9832), .o(TIMEBOOST_net_13056) );
na02f02 g63373_u0 ( .a(n_2921), .b(n_2625), .o(n_3321) );
ao12f02 g63374_u0 ( .a(n_3111), .b(configuration_wb_err_addr_560), .c(n_15444), .o(n_3440) );
ao12f02 g63375_u0 ( .a(n_3114), .b(configuration_wb_err_addr_562), .c(n_15444), .o(n_3438) );
na02s01 TIMEBOOST_cell_37264 ( .a(TIMEBOOST_net_10870), .b(FE_OFN686_n_4417), .o(TIMEBOOST_net_9387) );
na02s02 g63377_u0 ( .a(n_3417), .b(n_4637), .o(n_4638) );
in01s01 g63378_u0 ( .a(FE_OFN1117_g64577_p), .o(g63378_sb) );
na03f02 TIMEBOOST_cell_22254 ( .a(n_16984), .b(n_16985), .c(n_9997), .o(TIMEBOOST_net_6384) );
na02s01 g63378_u2 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_1_), .b(FE_OFN1092_g64577_p), .o(g63378_db) );
na02f02 TIMEBOOST_cell_22255 ( .a(TIMEBOOST_net_6384), .b(n_10584), .o(n_12139) );
in01m02 g63379_u0 ( .a(n_4137), .o(n_4636) );
ao12m02 g63380_u0 ( .a(n_4131), .b(FE_OFN1117_g64577_p), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_), .o(n_4137) );
na02f02 g63381_u0 ( .a(n_3297), .b(n_2624), .o(n_4136) );
na03s02 TIMEBOOST_cell_5954 ( .a(n_4476), .b(g64860_sb), .c(g64860_db), .o(n_4430) );
na02f02 g63383_u0 ( .a(n_3294), .b(n_2620), .o(n_4135) );
no02f02 g63385_u0 ( .a(n_2432), .b(n_1372), .o(n_2947) );
in01s01 g63386_u0 ( .a(n_3436), .o(n_3437) );
na02m02 TIMEBOOST_cell_44083 ( .a(n_9590), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__Q), .o(TIMEBOOST_net_14280) );
na03s01 TIMEBOOST_cell_33511 ( .a(n_1579), .b(g61949_sb), .c(g61949_db), .o(n_7927) );
ao12f01 g63390_u0 ( .a(n_2443), .b(n_3260), .c(conf_wb_err_bc_in), .o(n_4635) );
in01s01 g63392_u0 ( .a(FE_OFN1117_g64577_p), .o(g63392_sb) );
na03f02 TIMEBOOST_cell_22256 ( .a(n_9280), .b(n_10081), .c(n_9283), .o(TIMEBOOST_net_6385) );
na02m04 TIMEBOOST_cell_39025 ( .a(wbs_wbb3_2_wbb2_dat_o_i_125), .b(wbs_dat_o_26_), .o(TIMEBOOST_net_11751) );
na02f02 TIMEBOOST_cell_22257 ( .a(TIMEBOOST_net_6385), .b(n_10084), .o(n_11846) );
na02m02 TIMEBOOST_cell_41636 ( .a(TIMEBOOST_net_13056), .b(FE_OFN1439_n_9372), .o(TIMEBOOST_net_11657) );
in01s02 g63394_u0 ( .a(n_4132), .o(n_4634) );
ao12m02 g63395_u0 ( .a(n_4131), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .c(FE_OFN1117_g64577_p), .o(n_4132) );
in01s01 g63397_u0 ( .a(FE_OFN1117_g64577_p), .o(g63397_sb) );
na02s02 TIMEBOOST_cell_30881 ( .a(TIMEBOOST_net_9351), .b(FE_OFN784_n_2678), .o(TIMEBOOST_net_3729) );
na03s02 TIMEBOOST_cell_34272 ( .a(TIMEBOOST_net_9807), .b(FE_OFN1165_n_5615), .c(g62110_sb), .o(n_5588) );
na02s01 TIMEBOOST_cell_30882 ( .a(pci_target_unit_pcit_if_strd_addr_in_716), .b(pci_target_unit_del_sync_addr_in_234), .o(TIMEBOOST_net_9352) );
oa12s01 g63398_u0 ( .a(n_16330), .b(n_653), .c(FE_OFN2093_n_2301), .o(n_2946) );
na02f02 TIMEBOOST_cell_37814 ( .a(TIMEBOOST_net_11145), .b(TIMEBOOST_net_1760), .o(n_12983) );
in01m01 g63400_u0 ( .a(n_3160), .o(n_2943) );
na02s01 TIMEBOOST_cell_30906 ( .a(pci_target_unit_pcit_if_strd_addr_in_693), .b(n_2507), .o(TIMEBOOST_net_9364) );
no02m02 g63402_u0 ( .a(n_1382), .b(n_2434), .o(n_2942) );
ao12f02 g63403_u0 ( .a(n_3112), .b(configuration_wb_err_addr_559), .c(n_15444), .o(n_17049) );
oa12f02 g63404_u0 ( .a(n_2701), .b(n_3304), .c(n_1998), .o(n_3432) );
ao12f02 g63406_u0 ( .a(n_3110), .b(configuration_wb_err_addr_561), .c(n_15444), .o(n_17040) );
no02m04 g63407_u0 ( .a(n_2930), .b(n_880), .o(n_3318) );
no02s02 g63409_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_13_), .b(n_1990), .o(g63409_p) );
ao12s02 g63409_u1 ( .a(g63409_p), .b(pci_target_unit_del_sync_comp_cycle_count_13_), .c(n_1990), .o(n_2721) );
ao12s02 g63410_u0 ( .a(n_3384), .b(n_4783), .c(configuration_interrupt_line_40), .o(n_4785) );
ao12s02 g63411_u0 ( .a(n_3381), .b(n_4783), .c(configuration_interrupt_line_39), .o(n_4784) );
ao12s02 g63412_u0 ( .a(n_3389), .b(n_4783), .c(configuration_interrupt_line_41), .o(n_4782) );
ao12s02 g63413_u0 ( .a(n_3387), .b(n_4783), .c(configuration_interrupt_line_43), .o(n_4781) );
oa12s02 g63414_u0 ( .a(n_2935), .b(n_2934), .c(wbm_adr_o_19_), .o(n_3317) );
oa12m02 g63415_u0 ( .a(n_2717), .b(n_2716), .c(wbu_addr_in_268), .o(n_3140) );
oa12m02 g63416_u0 ( .a(n_2715), .b(n_2714), .c(wbu_addr_in_269), .o(n_3139) );
ao12s02 g63417_u0 ( .a(n_3276), .b(n_4630), .c(wbu_cache_line_size_in_209), .o(n_4633) );
oa12m02 g63418_u0 ( .a(n_2713), .b(n_2712), .c(wbu_addr_in_272), .o(n_3138) );
oa12s02 g63419_u0 ( .a(n_3419), .b(n_1752), .c(FE_OFN1117_g64577_p), .o(n_4632) );
oa12s02 g63420_u0 ( .a(n_2707), .b(n_2706), .c(wbm_adr_o_20_), .o(n_3137) );
ao12s02 g63421_u0 ( .a(n_3274), .b(n_4630), .c(wbu_cache_line_size_in_208), .o(n_4631) );
no02m02 g63422_u0 ( .a(n_2398), .b(conf_wb_err_addr_in_964), .o(g63422_p) );
ao12m02 g63422_u1 ( .a(g63422_p), .b(conf_wb_err_addr_in_964), .c(n_2398), .o(n_3136) );
no02m02 g63423_u0 ( .a(n_2230), .b(conf_wb_err_addr_in_961), .o(g63423_p) );
ao12m02 g63423_u1 ( .a(g63423_p), .b(conf_wb_err_addr_in_961), .c(n_2230), .o(n_2941) );
no02f02 g63424_u0 ( .a(conf_wb_err_addr_in_960), .b(n_2266), .o(g63424_p) );
ao12f02 g63424_u1 ( .a(g63424_p), .b(conf_wb_err_addr_in_960), .c(n_2266), .o(n_2940) );
ao12s02 g63425_u0 ( .a(n_3279), .b(n_4630), .c(wbu_cache_line_size_in_207), .o(n_4629) );
no02s01 g63426_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_6_), .b(n_2009), .o(g63426_p) );
ao12s01 g63426_u1 ( .a(g63426_p), .b(pci_target_unit_del_sync_comp_cycle_count_6_), .c(n_2009), .o(n_2010) );
ao12s02 g63427_u0 ( .a(n_3266), .b(n_4630), .c(wbu_cache_line_size_in_211), .o(n_4628) );
no02s02 g63428_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q), .b(n_1994), .o(g63428_p) );
ao12s02 g63428_u1 ( .a(g63428_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q), .c(n_1994), .o(n_2731) );
no02s01 g63429_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_6_), .b(n_2007), .o(g63429_p) );
ao12s01 g63429_u1 ( .a(g63429_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_6_), .c(n_2007), .o(n_2008) );
na03s02 TIMEBOOST_cell_42765 ( .a(g58100_sb), .b(g58100_db), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__Q), .o(TIMEBOOST_net_13621) );
in01s01 g63431_u0 ( .a(FE_OFN1126_g64577_p), .o(g63431_sb) );
in01s01 TIMEBOOST_cell_32845 ( .a(TIMEBOOST_net_10346), .o(TIMEBOOST_net_10345) );
na02s01 TIMEBOOST_cell_37263 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__Q), .b(n_3747), .o(TIMEBOOST_net_10870) );
na02s06 TIMEBOOST_cell_44758 ( .a(TIMEBOOST_net_14617), .b(n_1442), .o(n_1443) );
in01s01 g63432_u0 ( .a(FE_OFN1133_g64577_p), .o(g63432_sb) );
na02s01 TIMEBOOST_cell_42589 ( .a(FE_OFN205_n_9140), .b(g57902_sb), .o(TIMEBOOST_net_13533) );
na02s02 TIMEBOOST_cell_37221 ( .a(n_276), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_0_), .o(TIMEBOOST_net_10849) );
na02s02 TIMEBOOST_cell_43271 ( .a(n_3778), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__Q), .o(TIMEBOOST_net_13874) );
in01s01 g63433_u0 ( .a(FE_OFN1126_g64577_p), .o(g63433_sb) );
na02m02 TIMEBOOST_cell_41595 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_20__Q), .b(FE_OFN221_n_9846), .o(TIMEBOOST_net_13036) );
na02s01 TIMEBOOST_cell_37223 ( .a(parchk_pci_ad_reg_in_1224), .b(pci_target_unit_del_sync_addr_in_223), .o(TIMEBOOST_net_10850) );
na02s01 TIMEBOOST_cell_45680 ( .a(TIMEBOOST_net_15078), .b(FE_OFN1194_n_6935), .o(TIMEBOOST_net_13256) );
in01s01 g63434_u0 ( .a(FE_OFN1126_g64577_p), .o(g63434_sb) );
na03s02 TIMEBOOST_cell_34244 ( .a(TIMEBOOST_net_9802), .b(FE_OFN1170_n_5592), .c(g62138_sb), .o(n_5555) );
na02s01 TIMEBOOST_cell_37225 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__Q), .b(n_4671), .o(TIMEBOOST_net_10851) );
na02s02 TIMEBOOST_cell_42750 ( .a(TIMEBOOST_net_13613), .b(g58175_db), .o(n_9615) );
in01s01 g63435_u0 ( .a(FE_OFN1125_g64577_p), .o(g63435_sb) );
na02s02 TIMEBOOST_cell_42951 ( .a(TIMEBOOST_net_9637), .b(FE_OFN1671_n_9477), .o(TIMEBOOST_net_13714) );
na02s01 g63435_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__Q), .b(FE_OFN1125_g64577_p), .o(g63435_db) );
na02f02 TIMEBOOST_cell_41536 ( .a(TIMEBOOST_net_13006), .b(g57563_sb), .o(n_11188) );
in01s01 g63436_u0 ( .a(FE_OFN1124_g64577_p), .o(g63436_sb) );
na02s02 TIMEBOOST_cell_45681 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__Q), .b(n_4309), .o(TIMEBOOST_net_15079) );
na02m02 TIMEBOOST_cell_39375 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_781), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_16__Q), .o(TIMEBOOST_net_11926) );
na02f02 TIMEBOOST_cell_41538 ( .a(TIMEBOOST_net_13007), .b(g57259_sb), .o(n_11495) );
in01s01 g63437_u0 ( .a(FE_OFN1128_g64577_p), .o(g63437_sb) );
na02m02 TIMEBOOST_cell_44393 ( .a(n_9514), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__Q), .o(TIMEBOOST_net_14435) );
na02s01 TIMEBOOST_cell_39377 ( .a(g58211_db), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q), .o(TIMEBOOST_net_11927) );
na03s02 TIMEBOOST_cell_41991 ( .a(n_3586), .b(FE_OFN1248_n_4093), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__Q), .o(TIMEBOOST_net_13234) );
in01s01 g63438_u0 ( .a(FE_OFN1125_g64577_p), .o(g63438_sb) );
na02s02 TIMEBOOST_cell_43263 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__Q), .b(n_3779), .o(TIMEBOOST_net_13870) );
na02s02 TIMEBOOST_cell_39379 ( .a(n_3269), .b(TIMEBOOST_net_603), .o(TIMEBOOST_net_11928) );
na02s01 TIMEBOOST_cell_41992 ( .a(TIMEBOOST_net_13234), .b(g62893_sb), .o(n_6091) );
in01s04 g63458_u0 ( .a(n_7350), .o(n_8272) );
in01s04 g63463_u0 ( .a(n_7350), .o(n_7845) );
in01m08 g63466_u0 ( .a(n_7350), .o(n_8069) );
in01s08 g63479_u0 ( .a(n_7350), .o(n_8119) );
in01s06 g63488_u0 ( .a(n_7350), .o(n_8232) );
in01s06 g63511_u0 ( .a(n_7350), .o(n_8140) );
in01s06 g63516_u0 ( .a(n_7350), .o(n_8176) );
in01s04 g63517_u0 ( .a(n_7350), .o(n_8060) );
in01s08 g63519_u0 ( .a(n_7350), .o(n_8407) );
in01m10 g63523_u0 ( .a(n_7102), .o(n_7350) );
ao22m08 g63524_u0 ( .a(n_1036), .b(pci_target_unit_fifos_pcir_wenable_in), .c(n_659), .d(pci_target_unit_fifos_pcir_wenable_in), .o(n_7102) );
no02s02 g63525_u0 ( .a(wbm_adr_o_23_), .b(n_2414), .o(g63525_p) );
ao12m02 g63525_u1 ( .a(g63525_p), .b(wbm_adr_o_23_), .c(n_2414), .o(n_3135) );
ao12f02 g63528_u0 ( .a(n_3301), .b(n_16543), .c(configuration_wb_err_cs_bit9), .o(n_4125) );
ao12f02 g63529_u0 ( .a(n_3407), .b(FE_OFN1066_n_15808), .c(configuration_pci_err_data_503), .o(n_4619) );
in01m01 g63530_u0 ( .a(n_15262), .o(g63530_sb) );
na02s01 TIMEBOOST_cell_9076 ( .a(pci_target_unit_fifos_pciw_cbe_in_153), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__Q), .o(TIMEBOOST_net_1105) );
na02f01 g63530_u2 ( .a(n_15262), .b(n_16763), .o(g63530_db) );
na02s01 TIMEBOOST_cell_9077 ( .a(TIMEBOOST_net_1105), .b(n_4725), .o(TIMEBOOST_net_217) );
ao12f02 g63531_u0 ( .a(n_3302), .b(FE_OCPN1845_n_16427), .c(n_3592), .o(n_4123) );
ao12f02 g63532_u0 ( .a(n_4088), .b(FE_OFN1695_n_3368), .c(wbu_cache_line_size_in_210), .o(n_4780) );
in01m01 g63533_u0 ( .a(FE_OFN1148_n_13249), .o(g63533_sb) );
na02s02 TIMEBOOST_cell_43594 ( .a(TIMEBOOST_net_14035), .b(FE_OFN1315_n_6624), .o(TIMEBOOST_net_12251) );
na02s02 TIMEBOOST_cell_39966 ( .a(TIMEBOOST_net_12221), .b(g62571_sb), .o(n_6413) );
na02f02 TIMEBOOST_cell_36932 ( .a(TIMEBOOST_net_10704), .b(g52599_sb), .o(n_10274) );
ao12f02 g63534_u0 ( .a(n_3306), .b(n_16791), .c(pciu_bar0_in_361), .o(n_4119) );
in01s01 g63537_u0 ( .a(FE_OFN904_n_4736), .o(g63537_sb) );
na02s01 TIMEBOOST_cell_17432 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__15__Q), .b(g64233_sb), .o(TIMEBOOST_net_3973) );
na02s01 g63537_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__Q), .b(FE_OFN904_n_4736), .o(g63537_db) );
na02s01 TIMEBOOST_cell_17433 ( .a(TIMEBOOST_net_3973), .b(g64233_db), .o(n_3939) );
in01s01 g63538_u0 ( .a(FE_OFN1074_n_4740), .o(g63538_sb) );
na03s02 TIMEBOOST_cell_38197 ( .a(TIMEBOOST_net_3704), .b(g64317_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__Q), .o(TIMEBOOST_net_11337) );
na02s01 g63538_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__Q), .b(FE_OFN1074_n_4740), .o(g63538_db) );
na02s02 TIMEBOOST_cell_38462 ( .a(TIMEBOOST_net_11469), .b(g58266_db), .o(n_9532) );
no02s01 g63539_u0 ( .a(wbm_adr_o_12_), .b(n_2441), .o(g63539_p) );
ao12s02 g63539_u1 ( .a(g63539_p), .b(wbm_adr_o_12_), .c(n_2441), .o(n_2720) );
oa12s01 g63540_u0 ( .a(n_3420), .b(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_), .c(FE_OFN1117_g64577_p), .o(n_4616) );
oa12s02 g63541_u0 ( .a(n_3416), .b(n_3415), .c(FE_OFN1117_g64577_p), .o(n_4614) );
no02s01 g63542_u0 ( .a(wbu_addr_in_261), .b(n_2437), .o(g63542_p) );
ao12m01 g63542_u1 ( .a(g63542_p), .b(wbu_addr_in_261), .c(n_2437), .o(n_2719) );
in01s01 g63543_u0 ( .a(FE_OFN1013_n_4734), .o(g63543_sb) );
na02s01 g63543_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(g63543_sb), .o(g63543_da) );
na02s01 g63543_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__Q), .b(FE_OFN1013_n_4734), .o(g63543_db) );
na02s01 TIMEBOOST_cell_39253 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__Q), .b(g58383_sb), .o(TIMEBOOST_net_11865) );
in01s01 g63544_u0 ( .a(FE_OFN1074_n_4740), .o(g63544_sb) );
na03s02 TIMEBOOST_cell_41973 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__Q), .b(n_3656), .c(FE_OFN1219_n_6886), .o(TIMEBOOST_net_13225) );
na02s01 g63544_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__Q), .b(FE_OFN1074_n_4740), .o(g63544_db) );
na02s02 TIMEBOOST_cell_38464 ( .a(TIMEBOOST_net_11470), .b(TIMEBOOST_net_568), .o(n_13423) );
in01s01 g63545_u0 ( .a(FE_OFN1013_n_4734), .o(g63545_sb) );
na02s01 g63545_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(g63545_sb), .o(g63545_da) );
na02s01 g63545_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__Q), .b(FE_OFN1013_n_4734), .o(g63545_db) );
na02m02 TIMEBOOST_cell_38939 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_31__Q), .o(TIMEBOOST_net_11708) );
no02m01 g63546_u0 ( .a(n_2931), .b(wbm_adr_o_15_), .o(g63546_p) );
ao12s02 g63546_u1 ( .a(g63546_p), .b(wbm_adr_o_15_), .c(n_2931), .o(n_3134) );
in01s01 g63547_u0 ( .a(FE_OFN1046_n_16657), .o(g63547_sb) );
na02s02 TIMEBOOST_cell_37770 ( .a(TIMEBOOST_net_11123), .b(FE_OFN2021_n_4778), .o(TIMEBOOST_net_10602) );
na02s01 g63547_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__Q), .b(FE_OFN1046_n_16657), .o(g63547_db) );
na02s02 TIMEBOOST_cell_38684 ( .a(TIMEBOOST_net_11580), .b(g62368_sb), .o(n_6867) );
in01s01 g63548_u0 ( .a(FE_OFN904_n_4736), .o(g63548_sb) );
na02s01 TIMEBOOST_cell_43483 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__Q), .b(n_3677), .o(TIMEBOOST_net_13980) );
na02s01 g63548_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__Q), .b(FE_OFN904_n_4736), .o(g63548_db) );
na02s01 TIMEBOOST_cell_42941 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__Q), .b(FE_OFN562_n_9895), .o(TIMEBOOST_net_13709) );
in01s01 g63549_u0 ( .a(FE_OFN1046_n_16657), .o(g63549_sb) );
na02s02 TIMEBOOST_cell_41763 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__Q), .b(g58372_sb), .o(TIMEBOOST_net_13120) );
na02s01 g63549_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__Q), .b(FE_OFN1046_n_16657), .o(g63549_db) );
na02s02 TIMEBOOST_cell_38466 ( .a(TIMEBOOST_net_11471), .b(g58437_db), .o(TIMEBOOST_net_10055) );
in01s01 g63550_u0 ( .a(FE_OFN1125_g64577_p), .o(g63550_sb) );
na02f02 TIMEBOOST_cell_22275 ( .a(TIMEBOOST_net_6394), .b(FE_RN_233_0), .o(n_12133) );
na02s01 TIMEBOOST_cell_44787 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__Q), .b(FE_OFN575_n_9902), .o(TIMEBOOST_net_14632) );
na02f02 TIMEBOOST_cell_44346 ( .a(TIMEBOOST_net_14411), .b(FE_OFN1397_n_8567), .o(TIMEBOOST_net_12735) );
in01s01 g63551_u0 ( .a(FE_OFN1128_g64577_p), .o(g63551_sb) );
na04f10 TIMEBOOST_cell_13291 ( .a(FE_RN_510_0), .b(FE_RN_508_0), .c(FE_RN_512_0), .d(FE_RN_514_0), .o(n_16560) );
na02s01 TIMEBOOST_cell_44788 ( .a(TIMEBOOST_net_14632), .b(g58093_sb), .o(TIMEBOOST_net_12447) );
na02f02 TIMEBOOST_cell_41572 ( .a(TIMEBOOST_net_13024), .b(g57039_sb), .o(n_10513) );
in01s01 g63552_u0 ( .a(FE_OFN1133_g64577_p), .o(g63552_sb) );
na02f02 TIMEBOOST_cell_22241 ( .a(TIMEBOOST_net_6377), .b(n_9968), .o(n_12132) );
na02s01 TIMEBOOST_cell_37227 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__Q), .b(n_3755), .o(TIMEBOOST_net_10852) );
na02s01 TIMEBOOST_cell_30931 ( .a(TIMEBOOST_net_9376), .b(g65671_sb), .o(n_2379) );
in01s01 g63553_u0 ( .a(FE_OFN1128_g64577_p), .o(g63553_sb) );
na02s02 TIMEBOOST_cell_45709 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__Q), .b(n_1849), .o(TIMEBOOST_net_15093) );
na02s01 TIMEBOOST_cell_39385 ( .a(g64164_da), .b(g64164_db), .o(TIMEBOOST_net_11931) );
na02m04 TIMEBOOST_cell_45514 ( .a(TIMEBOOST_net_14995), .b(g54341_sb), .o(n_12974) );
in01s01 g63554_u0 ( .a(FE_OFN1133_g64577_p), .o(g63554_sb) );
na02f02 TIMEBOOST_cell_44084 ( .a(TIMEBOOST_net_14280), .b(FE_OFN1420_n_8567), .o(TIMEBOOST_net_12833) );
na02s01 TIMEBOOST_cell_37229 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__Q), .b(n_3780), .o(TIMEBOOST_net_10853) );
na02s02 TIMEBOOST_cell_42111 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__Q), .b(n_3630), .o(TIMEBOOST_net_13294) );
in01s01 g63555_u0 ( .a(FE_OFN1126_g64577_p), .o(g63555_sb) );
na02s01 TIMEBOOST_cell_37231 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__Q), .b(FE_OFN577_n_9902), .o(TIMEBOOST_net_10854) );
na02s01 TIMEBOOST_cell_22276 ( .a(g52473_da), .b(FE_OFN1022_n_11877), .o(TIMEBOOST_net_6395) );
in01s01 g63556_u0 ( .a(FE_OFN1125_g64577_p), .o(g63556_sb) );
na02m02 TIMEBOOST_cell_44347 ( .a(n_9527), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__Q), .o(TIMEBOOST_net_14412) );
na02s01 TIMEBOOST_cell_37233 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__31__Q), .b(FE_OFN606_n_9904), .o(TIMEBOOST_net_10855) );
na02s01 TIMEBOOST_cell_22288 ( .a(g52456_da), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_6401) );
in01s01 g63557_u0 ( .a(FE_OFN1126_g64577_p), .o(g63557_sb) );
na02f02 TIMEBOOST_cell_22323 ( .a(TIMEBOOST_net_6418), .b(FE_OFN1748_n_12004), .o(n_12605) );
na02s01 TIMEBOOST_cell_37235 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(g65792_sb), .o(TIMEBOOST_net_10856) );
na02m02 TIMEBOOST_cell_44085 ( .a(n_9465), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__Q), .o(TIMEBOOST_net_14281) );
ao12f02 g63558_u0 ( .a(n_3125), .b(n_15808), .c(configuration_pci_err_data), .o(n_3428) );
in01s01 g63559_u0 ( .a(FE_OFN1117_g64577_p), .o(g63559_sb) );
na02s02 TIMEBOOST_cell_43067 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__Q), .b(n_3768), .o(TIMEBOOST_net_13772) );
na02s01 g63559_u2 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_), .b(FE_OFN1092_g64577_p), .o(g63559_db) );
na02s01 TIMEBOOST_cell_30856 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(g65889_sb), .o(TIMEBOOST_net_9339) );
in01s01 g63560_u0 ( .a(FE_OFN1092_g64577_p), .o(g63560_sb) );
na03s02 TIMEBOOST_cell_38387 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__Q), .b(FE_OFN1124_g64577_p), .c(n_4030), .o(TIMEBOOST_net_11432) );
na02s01 g63560_u2 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_), .b(FE_OFN1092_g64577_p), .o(g63560_db) );
na02f01 TIMEBOOST_cell_38468 ( .a(TIMEBOOST_net_11472), .b(n_13814), .o(n_14073) );
in01s01 g63561_u0 ( .a(FE_OFN1092_g64577_p), .o(g63561_sb) );
na02s02 TIMEBOOST_cell_38470 ( .a(TIMEBOOST_net_11473), .b(FE_OFN1699_n_5751), .o(TIMEBOOST_net_4823) );
na02s01 g63561_u2 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_0_), .b(FE_OFN1092_g64577_p), .o(g63561_db) );
na02s01 TIMEBOOST_cell_18497 ( .a(TIMEBOOST_net_4505), .b(g63555_sb), .o(n_4922) );
in01s01 g63562_u0 ( .a(FE_OFN1092_g64577_p), .o(g63562_sb) );
na02s02 TIMEBOOST_cell_38686 ( .a(TIMEBOOST_net_11581), .b(g62664_sb), .o(n_6211) );
na02s01 g63562_u2 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_2_), .b(FE_OFN1092_g64577_p), .o(g63562_db) );
na02s02 TIMEBOOST_cell_18499 ( .a(TIMEBOOST_net_4506), .b(g62784_sb), .o(n_5424) );
in01s01 g63563_u0 ( .a(FE_OFN1058_n_4727), .o(g63563_sb) );
na02s01 g63563_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__Q), .b(g63563_sb), .o(g63563_da) );
na02s01 g63563_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(FE_OFN1058_n_4727), .o(g63563_db) );
na02s02 TIMEBOOST_cell_38463 ( .a(g54195_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_414), .o(TIMEBOOST_net_11470) );
in01s01 g63564_u0 ( .a(FE_OFN1057_n_4727), .o(g63564_sb) );
na02m02 TIMEBOOST_cell_44185 ( .a(n_9680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__Q), .o(TIMEBOOST_net_14331) );
na02s01 g63564_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(FE_OFN1057_n_4727), .o(g63564_db) );
na02f04 TIMEBOOST_cell_39026 ( .a(TIMEBOOST_net_11751), .b(FE_OFN2242_g52675_p), .o(TIMEBOOST_net_10749) );
in01s01 g63565_u0 ( .a(FE_OFN918_n_4725), .o(g63565_sb) );
na02s01 g63565_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__Q), .b(g63565_sb), .o(g63565_da) );
na02s01 g63565_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(FE_OFN918_n_4725), .o(g63565_db) );
na02s01 TIMEBOOST_cell_17278 ( .a(n_3752), .b(FE_OFN651_n_4508), .o(TIMEBOOST_net_3896) );
in01s01 g63566_u0 ( .a(FE_OFN1031_n_4732), .o(g63566_sb) );
na02s01 g63566_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__Q), .b(g63566_sb), .o(g63566_da) );
na02s01 g63566_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(FE_OFN1031_n_4732), .o(g63566_db) );
na02f02 TIMEBOOST_cell_39107 ( .a(TIMEBOOST_net_10165), .b(FE_OFN1606_n_13997), .o(TIMEBOOST_net_11792) );
in01s01 g63567_u0 ( .a(FE_OFN929_n_4730), .o(g63567_sb) );
na02s01 TIMEBOOST_cell_16904 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__Q), .b(g64346_sb), .o(TIMEBOOST_net_3709) );
na02s01 g63567_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(FE_OFN929_n_4730), .o(g63567_db) );
na02s01 TIMEBOOST_cell_45097 ( .a(n_2206), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__Q), .o(TIMEBOOST_net_14787) );
in01s01 g63568_u0 ( .a(FE_OFN929_n_4730), .o(g63568_sb) );
na02s02 TIMEBOOST_cell_45156 ( .a(TIMEBOOST_net_14816), .b(FE_OFN1264_n_4095), .o(TIMEBOOST_net_12026) );
na02s01 g63568_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(FE_OFN929_n_4730), .o(g63568_db) );
na02s01 TIMEBOOST_cell_16905 ( .a(TIMEBOOST_net_3709), .b(g64346_db), .o(n_3831) );
in01s01 g63569_u0 ( .a(FE_OFN1031_n_4732), .o(g63569_sb) );
na02s01 TIMEBOOST_cell_45043 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__Q), .b(n_1722), .o(TIMEBOOST_net_14760) );
na02s01 g63569_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(FE_OFN1031_n_4732), .o(g63569_db) );
na03s01 TIMEBOOST_cell_38169 ( .a(g64188_da), .b(g64188_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__Q), .o(TIMEBOOST_net_11323) );
in01s01 g63570_u0 ( .a(FE_OFN918_n_4725), .o(g63570_sb) );
na02s01 g63570_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__Q), .b(g63570_sb), .o(g63570_da) );
na02s01 g63570_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(FE_OFN918_n_4725), .o(g63570_db) );
na02s01 TIMEBOOST_cell_40445 ( .a(parchk_pci_ad_out_in_1185), .b(configuration_wb_err_data_588), .o(TIMEBOOST_net_12461) );
in01s01 g63571_u0 ( .a(FE_OFN1117_g64577_p), .o(g63571_sb) );
na02s01 TIMEBOOST_cell_36629 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(g64116_sb), .o(TIMEBOOST_net_10553) );
na02s01 g63571_u2 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_), .b(FE_OFN1092_g64577_p), .o(g63571_db) );
na02s01 TIMEBOOST_cell_42577 ( .a(TIMEBOOST_net_1104), .b(n_4725), .o(TIMEBOOST_net_13527) );
in01s01 g63572_u0 ( .a(FE_OFN1092_g64577_p), .o(g63572_sb) );
na02m02 TIMEBOOST_cell_10540 ( .a(FE_OFN2072_n_15978), .b(wishbone_slave_unit_del_sync_addr_out_reg_16__Q), .o(TIMEBOOST_net_1837) );
na02s01 g63572_u2 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_2_), .b(FE_OFN1092_g64577_p), .o(g63572_db) );
na03s02 TIMEBOOST_cell_34258 ( .a(TIMEBOOST_net_9817), .b(FE_OFN1168_n_5592), .c(g62093_sb), .o(n_5612) );
in01s01 g63573_u0 ( .a(FE_OFN1092_g64577_p), .o(g63573_sb) );
na03s02 TIMEBOOST_cell_38193 ( .a(TIMEBOOST_net_3955), .b(g64251_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__Q), .o(TIMEBOOST_net_11335) );
na02s01 g63573_u2 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_1_), .b(FE_OFN1092_g64577_p), .o(g63573_db) );
na02f02 TIMEBOOST_cell_38894 ( .a(TIMEBOOST_net_11685), .b(FE_OFN2200_n_10256), .o(TIMEBOOST_net_10706) );
in01s01 g63574_u0 ( .a(FE_OFN1092_g64577_p), .o(g63574_sb) );
na02s01 TIMEBOOST_cell_38614 ( .a(TIMEBOOST_net_11545), .b(g62420_sb), .o(n_6757) );
na02s01 g63574_u2 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_), .b(FE_OFN1092_g64577_p), .o(g63574_db) );
na02s02 TIMEBOOST_cell_18503 ( .a(TIMEBOOST_net_4508), .b(g62800_sb), .o(n_5383) );
ao22s01 g63575_u0 ( .a(n_1180), .b(n_1999), .c(n_3250), .d(pci_target_unit_wishbone_master_read_count_reg_2__Q), .o(n_3316) );
in01s01 g63576_u0 ( .a(FE_OFN1698_n_5751), .o(g63576_sb) );
na02s01 TIMEBOOST_cell_37237 ( .a(pci_target_unit_fifos_pcir_data_in_187), .b(g65806_sb), .o(TIMEBOOST_net_10857) );
na02s01 TIMEBOOST_cell_19026 ( .a(wishbone_slave_unit_pcim_sm_data_in_649), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__Q), .o(TIMEBOOST_net_4770) );
na02s01 TIMEBOOST_cell_37266 ( .a(TIMEBOOST_net_10871), .b(FE_OFN1625_n_4438), .o(TIMEBOOST_net_9408) );
in01m01 g63577_u0 ( .a(FE_OFN1700_n_5751), .o(g63577_sb) );
na02s01 TIMEBOOST_cell_42706 ( .a(TIMEBOOST_net_13591), .b(g65910_db), .o(n_1854) );
na02s02 TIMEBOOST_cell_38596 ( .a(TIMEBOOST_net_11536), .b(g60669_sb), .o(n_5649) );
na02s03 TIMEBOOST_cell_37182 ( .a(TIMEBOOST_net_10829), .b(wbu_addr_in_262), .o(n_9858) );
no02m02 g63578_u0 ( .a(wbu_addr_in_264), .b(n_3132), .o(g63578_p) );
ao12m02 g63578_u1 ( .a(g63578_p), .b(wbu_addr_in_264), .c(n_3132), .o(n_3133) );
no02m01 g63579_u0 ( .a(n_2722), .b(conf_wb_err_addr_in_953), .o(g63579_p) );
ao12s02 g63579_u1 ( .a(g63579_p), .b(conf_wb_err_addr_in_953), .c(n_2722), .o(n_2744) );
no02m01 g63580_u0 ( .a(n_3130), .b(conf_wb_err_addr_in_956), .o(g63580_p) );
ao12m02 g63580_u1 ( .a(g63580_p), .b(conf_wb_err_addr_in_956), .c(n_3130), .o(n_3131) );
no02m02 g63581_u0 ( .a(FE_OFN1698_n_5751), .b(wbm_adr_o_2_), .o(g63581_p) );
ao12m02 g63581_u1 ( .a(g63581_p), .b(wbm_adr_o_2_), .c(FE_OFN1698_n_5751), .o(n_3425) );
in01s01 g63582_u0 ( .a(FE_OFN1021_n_11877), .o(g63582_sb) );
na02s01 TIMEBOOST_cell_17252 ( .a(n_4444), .b(FE_OFN1644_n_4671), .o(TIMEBOOST_net_3883) );
na02s01 g63582_u2 ( .a(wbu_addr_in), .b(FE_OFN1021_n_11877), .o(g63582_db) );
na02s02 TIMEBOOST_cell_17253 ( .a(TIMEBOOST_net_3883), .b(g65320_da), .o(n_4270) );
na02f02 TIMEBOOST_cell_42336 ( .a(TIMEBOOST_net_13406), .b(g57438_sb), .o(n_10355) );
na02s01 TIMEBOOST_cell_17834 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__Q), .b(g65815_sb), .o(TIMEBOOST_net_4174) );
na02s01 TIMEBOOST_cell_36604 ( .a(TIMEBOOST_net_10540), .b(g65899_sb), .o(n_1719) );
in01s01 g63584_u0 ( .a(FE_OFN1025_n_11877), .o(g63584_sb) );
na02m02 TIMEBOOST_cell_39968 ( .a(TIMEBOOST_net_12222), .b(g62901_sb), .o(n_6075) );
na02s01 g63584_u2 ( .a(wbu_sel_in), .b(FE_OFN1025_n_11877), .o(g63584_db) );
na02f02 TIMEBOOST_cell_44086 ( .a(TIMEBOOST_net_14281), .b(FE_OFN1383_n_8567), .o(TIMEBOOST_net_12822) );
na02s01 TIMEBOOST_cell_39255 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__Q), .b(g58444_sb), .o(TIMEBOOST_net_11866) );
na02s01 g63585_u2 ( .a(wbu_sel_in_312), .b(FE_OFN1025_n_11877), .o(g63585_db) );
na02s01 TIMEBOOST_cell_39268 ( .a(TIMEBOOST_net_11872), .b(g64166_db), .o(n_3999) );
in01s01 g63586_u0 ( .a(FE_OFN1025_n_11877), .o(g63586_sb) );
na02s01 TIMEBOOST_cell_39269 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__Q), .b(n_8176), .o(TIMEBOOST_net_11873) );
na02s01 g63586_u2 ( .a(wbu_sel_in_313), .b(FE_OFN1025_n_11877), .o(g63586_db) );
na02s01 TIMEBOOST_cell_39270 ( .a(TIMEBOOST_net_11873), .b(n_1603), .o(TIMEBOOST_net_11563) );
na02f04 TIMEBOOST_cell_45516 ( .a(TIMEBOOST_net_14996), .b(g54342_sb), .o(n_12972) );
na02s01 g63587_u2 ( .a(wbu_sel_in_314), .b(FE_OFN1025_n_11877), .o(g63587_db) );
na02m02 TIMEBOOST_cell_44087 ( .a(n_9464), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__Q), .o(TIMEBOOST_net_14282) );
in01s01 g63588_u0 ( .a(FE_OFN9_n_11877), .o(g63588_sb) );
na02f02 TIMEBOOST_cell_44088 ( .a(TIMEBOOST_net_14282), .b(FE_OFN1414_n_8567), .o(TIMEBOOST_net_12795) );
na02s01 g63588_u2 ( .a(n_16945), .b(FE_OFN9_n_11877), .o(g63588_db) );
na02m02 TIMEBOOST_cell_44089 ( .a(n_9492), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__Q), .o(TIMEBOOST_net_14283) );
in01s01 g63589_u0 ( .a(FE_OFN2_n_4778), .o(g63589_sb) );
na02s01 TIMEBOOST_cell_36606 ( .a(TIMEBOOST_net_10541), .b(g65828_sb), .o(n_1888) );
na02f06 TIMEBOOST_cell_37000 ( .a(TIMEBOOST_net_10738), .b(FE_OCP_RBN2016_n_16970), .o(n_13807) );
na02s01 TIMEBOOST_cell_36608 ( .a(TIMEBOOST_net_10542), .b(FE_OFN252_n_9868), .o(n_9562) );
in01s01 g63590_u0 ( .a(FE_OFN989_n_574), .o(g63590_sb) );
na02f02 TIMEBOOST_cell_43728 ( .a(TIMEBOOST_net_14102), .b(FE_OFN1383_n_8567), .o(TIMEBOOST_net_12695) );
na02m02 TIMEBOOST_cell_44535 ( .a(n_9613), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__Q), .o(TIMEBOOST_net_14506) );
na02s02 TIMEBOOST_cell_43264 ( .a(TIMEBOOST_net_13870), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_11539) );
in01s02 g63591_u0 ( .a(FE_OFN2021_n_4778), .o(g63591_sb) );
na02s01 g63591_u1 ( .a(wbs_dat_i_27_), .b(g63591_sb), .o(g63591_da) );
na02s02 TIMEBOOST_cell_39970 ( .a(TIMEBOOST_net_12223), .b(g62518_sb), .o(n_6541) );
na02s01 TIMEBOOST_cell_36464 ( .a(TIMEBOOST_net_10470), .b(g65784_db), .o(n_2006) );
in01s01 g63592_u0 ( .a(FE_OFN2_n_4778), .o(g63592_sb) );
na02s01 TIMEBOOST_cell_36610 ( .a(TIMEBOOST_net_10543), .b(g65940_sb), .o(n_2579) );
na02s01 g63592_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__Q), .b(FE_OFN2_n_4778), .o(g63592_db) );
na02s02 TIMEBOOST_cell_36612 ( .a(TIMEBOOST_net_10544), .b(g58156_db), .o(n_9635) );
in01s01 g63593_u0 ( .a(FE_OFN2_n_4778), .o(g63593_sb) );
na02s01 TIMEBOOST_cell_36614 ( .a(TIMEBOOST_net_10545), .b(FE_OFN552_n_9864), .o(TIMEBOOST_net_294) );
na02f04 TIMEBOOST_cell_37002 ( .a(TIMEBOOST_net_10739), .b(g52503_sb), .o(n_13823) );
na02s01 TIMEBOOST_cell_36616 ( .a(TIMEBOOST_net_10546), .b(g58225_db), .o(n_9048) );
in01s01 g63594_u0 ( .a(FE_OFN2021_n_4778), .o(g63594_sb) );
na02s01 TIMEBOOST_cell_36618 ( .a(TIMEBOOST_net_10547), .b(g65940_sb), .o(n_2575) );
na02f04 TIMEBOOST_cell_37004 ( .a(TIMEBOOST_net_10740), .b(g52505_sb), .o(n_13822) );
na02s01 TIMEBOOST_cell_36620 ( .a(TIMEBOOST_net_10548), .b(FE_OFN239_n_9832), .o(TIMEBOOST_net_3926) );
in01s01 g63595_u0 ( .a(FE_OFN2_n_4778), .o(g63595_sb) );
na02s01 TIMEBOOST_cell_36622 ( .a(TIMEBOOST_net_10549), .b(FE_OFN211_n_9858), .o(TIMEBOOST_net_3887) );
na02f04 TIMEBOOST_cell_37006 ( .a(TIMEBOOST_net_10741), .b(g52507_sb), .o(n_13719) );
na02s01 TIMEBOOST_cell_36624 ( .a(TIMEBOOST_net_10550), .b(FE_OFN221_n_9846), .o(n_9738) );
in01s01 g63596_u0 ( .a(FE_OFN2_n_4778), .o(g63596_sb) );
na02s01 TIMEBOOST_cell_36626 ( .a(TIMEBOOST_net_10551), .b(FE_OFN1635_n_9531), .o(TIMEBOOST_net_4032) );
na02f04 TIMEBOOST_cell_37008 ( .a(TIMEBOOST_net_10742), .b(g52508_sb), .o(n_13717) );
na02s01 TIMEBOOST_cell_36628 ( .a(TIMEBOOST_net_10552), .b(g64835_sb), .o(n_3729) );
in01s01 g63597_u0 ( .a(FE_OFN1079_n_4778), .o(g63597_sb) );
na02s01 g63597_u1 ( .a(wbs_dat_i_23_), .b(g63597_sb), .o(g63597_da) );
na02s02 TIMEBOOST_cell_39972 ( .a(TIMEBOOST_net_12224), .b(g62395_sb), .o(n_7390) );
na02s01 TIMEBOOST_cell_39186 ( .a(TIMEBOOST_net_11831), .b(g65934_db), .o(n_2170) );
in01s01 g63598_u0 ( .a(FE_OFN2022_n_4778), .o(g63598_sb) );
na02s01 TIMEBOOST_cell_39432 ( .a(TIMEBOOST_net_11954), .b(g62003_sb), .o(n_7889) );
na02f04 TIMEBOOST_cell_37010 ( .a(TIMEBOOST_net_10743), .b(g52510_sb), .o(n_13816) );
na02f02 TIMEBOOST_cell_38896 ( .a(TIMEBOOST_net_11686), .b(FE_OFN2198_n_10256), .o(TIMEBOOST_net_10082) );
in01s01 g63599_u0 ( .a(FE_OFN1079_n_4778), .o(g63599_sb) );
na02s01 g63599_u1 ( .a(wbs_dat_i_12_), .b(g63599_sb), .o(g63599_da) );
na02s01 g63599_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__Q), .b(FE_OFN1079_n_4778), .o(g63599_db) );
na02s01 TIMEBOOST_cell_38472 ( .a(TIMEBOOST_net_11474), .b(g61918_sb), .o(n_7953) );
in01s01 g63600_u0 ( .a(FE_OFN2021_n_4778), .o(g63600_sb) );
na02s02 TIMEBOOST_cell_38758 ( .a(TIMEBOOST_net_11617), .b(g53921_sb), .o(n_13523) );
na02f04 TIMEBOOST_cell_37012 ( .a(TIMEBOOST_net_10744), .b(g52511_sb), .o(n_13712) );
na02s02 TIMEBOOST_cell_38760 ( .a(TIMEBOOST_net_11618), .b(g53904_sb), .o(n_13537) );
in01s01 g63601_u0 ( .a(FE_OFN2022_n_4778), .o(g63601_sb) );
na02s01 TIMEBOOST_cell_39188 ( .a(TIMEBOOST_net_11832), .b(g65851_db), .o(n_2184) );
na02s01 g63601_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__Q), .b(FE_OFN1079_n_4778), .o(g63601_db) );
na02s02 TIMEBOOST_cell_38762 ( .a(TIMEBOOST_net_11619), .b(g53922_sb), .o(n_13522) );
in01s01 g63602_u0 ( .a(FE_OFN1079_n_4778), .o(g63602_sb) );
na02s01 g63602_u1 ( .a(wbs_dat_i_21_), .b(g63602_sb), .o(g63602_da) );
na02s01 g63602_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__Q), .b(FE_OFN1079_n_4778), .o(g63602_db) );
na03s01 TIMEBOOST_cell_963 ( .a(n_3994), .b(g62791_sb), .c(g62791_db), .o(n_5406) );
in01s01 g63603_u0 ( .a(FE_OFN1079_n_4778), .o(g63603_sb) );
na02s01 g63603_u1 ( .a(wbs_dat_i_28_), .b(g63603_sb), .o(g63603_da) );
na02s01 g63603_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__Q), .b(FE_OFN1079_n_4778), .o(g63603_db) );
na02s02 TIMEBOOST_cell_10861 ( .a(TIMEBOOST_net_1997), .b(g63172_sb), .o(n_4951) );
in01s02 g63604_u0 ( .a(FE_OFN2021_n_4778), .o(g63604_sb) );
na02s01 g63604_u1 ( .a(wbs_dat_i_30_), .b(g63604_sb), .o(g63604_da) );
na02f02 TIMEBOOST_cell_10342 ( .a(g54317_db), .b(n_12595), .o(TIMEBOOST_net_1738) );
na02s01 TIMEBOOST_cell_36466 ( .a(TIMEBOOST_net_10471), .b(g65753_db), .o(n_1922) );
in01s01 g63605_u0 ( .a(FE_OFN1079_n_4778), .o(g63605_sb) );
na02s01 g63605_u1 ( .a(wbs_dat_i_31_), .b(g63605_sb), .o(g63605_da) );
na02s01 g63605_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__Q), .b(FE_OFN1079_n_4778), .o(g63605_db) );
na02s02 TIMEBOOST_cell_18909 ( .a(TIMEBOOST_net_4711), .b(g62853_sb), .o(n_5263) );
in01s02 g63606_u0 ( .a(FE_OFN2_n_4778), .o(g63606_sb) );
na02s01 g63606_u1 ( .a(wbs_dat_i_3_), .b(g63606_sb), .o(g63606_da) );
na02s01 TIMEBOOST_cell_18284 ( .a(g61880_sb), .b(g61880_db), .o(TIMEBOOST_net_4399) );
na02s01 TIMEBOOST_cell_38062 ( .a(TIMEBOOST_net_11269), .b(FE_OFN1129_g64577_p), .o(TIMEBOOST_net_4685) );
in01s01 g63607_u0 ( .a(FE_OFN1079_n_4778), .o(g63607_sb) );
na02s01 g63607_u1 ( .a(wbs_dat_i_15_), .b(g63607_sb), .o(g63607_da) );
na02s01 g63607_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__Q), .b(FE_OFN1079_n_4778), .o(g63607_db) );
na02s01 TIMEBOOST_cell_38474 ( .a(TIMEBOOST_net_11475), .b(g61732_sb), .o(n_7947) );
in01s01 g63608_u0 ( .a(FE_OFN2022_n_4778), .o(g63608_sb) );
na02s01 TIMEBOOST_cell_38764 ( .a(TIMEBOOST_net_11620), .b(g53899_sb), .o(n_13546) );
na02f04 TIMEBOOST_cell_37014 ( .a(TIMEBOOST_net_10745), .b(g52512_sb), .o(n_13815) );
na02s02 TIMEBOOST_cell_38766 ( .a(TIMEBOOST_net_11621), .b(g53914_sb), .o(n_13470) );
in01s02 g63609_u0 ( .a(FE_OFN2_n_4778), .o(g63609_sb) );
na02s01 g63609_u1 ( .a(wbs_dat_i_7_), .b(g63609_sb), .o(g63609_da) );
na02f02 TIMEBOOST_cell_10346 ( .a(n_13763), .b(FE_OFN2251_n_2101), .o(TIMEBOOST_net_1740) );
na02f04 TIMEBOOST_cell_20683 ( .a(TIMEBOOST_net_5598), .b(g75072_db), .o(n_16441) );
in01s01 g63610_u0 ( .a(FE_OFN2021_n_4778), .o(g63610_sb) );
na02f02 TIMEBOOST_cell_38898 ( .a(TIMEBOOST_net_11687), .b(FE_OFN2198_n_10256), .o(TIMEBOOST_net_10084) );
na02f04 TIMEBOOST_cell_37016 ( .a(TIMEBOOST_net_10746), .b(g52513_sb), .o(n_13812) );
na02s01 TIMEBOOST_cell_39448 ( .a(TIMEBOOST_net_11962), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_4663) );
in01s01 g63611_u0 ( .a(FE_OFN1079_n_4778), .o(g63611_sb) );
na02s01 g63611_u1 ( .a(wbs_dat_i_11_), .b(g63611_sb), .o(g63611_da) );
na02s01 g63611_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__Q), .b(FE_OFN1079_n_4778), .o(g63611_db) );
na02s01 TIMEBOOST_cell_18591 ( .a(TIMEBOOST_net_4552), .b(g63038_sb), .o(n_5172) );
in01s01 g63612_u0 ( .a(FE_OFN1079_n_4778), .o(g63612_sb) );
na02s01 g63612_u1 ( .a(wbs_dat_i_17_), .b(g63612_sb), .o(g63612_da) );
na02s01 TIMEBOOST_cell_39271 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__12__Q), .b(g64270_sb), .o(TIMEBOOST_net_11874) );
na02s01 TIMEBOOST_cell_37156 ( .a(TIMEBOOST_net_10816), .b(pci_target_unit_del_sync_comp_rty_exp_reg), .o(TIMEBOOST_net_3181) );
in01s01 g63613_u0 ( .a(FE_OFN1079_n_4778), .o(g63613_sb) );
na02s01 g63613_u1 ( .a(wbs_dat_i_14_), .b(g63613_sb), .o(g63613_da) );
na02s01 g63613_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__Q), .b(FE_OFN1079_n_4778), .o(g63613_db) );
na02s01 TIMEBOOST_cell_18921 ( .a(TIMEBOOST_net_4717), .b(g63090_sb), .o(n_5074) );
in01s01 g63614_u0 ( .a(FE_OFN1079_n_4778), .o(g63614_sb) );
na02s01 g63614_u1 ( .a(wbs_dat_i_0_), .b(g63614_sb), .o(g63614_da) );
na02s01 g63614_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__Q), .b(FE_OFN1079_n_4778), .o(g63614_db) );
na02s01 TIMEBOOST_cell_18925 ( .a(TIMEBOOST_net_4719), .b(g63053_sb), .o(n_5143) );
in01s01 g63615_u0 ( .a(FE_OFN2022_n_4778), .o(g63615_sb) );
na02s01 TIMEBOOST_cell_36630 ( .a(TIMEBOOST_net_10553), .b(g64116_db), .o(n_4044) );
na02f04 TIMEBOOST_cell_37018 ( .a(TIMEBOOST_net_10747), .b(g52514_sb), .o(n_13809) );
na02s01 TIMEBOOST_cell_36632 ( .a(TIMEBOOST_net_10554), .b(g61797_db), .o(n_8203) );
in01s01 g63616_u0 ( .a(FE_OFN2_n_4778), .o(g63616_sb) );
na02s01 TIMEBOOST_cell_36634 ( .a(TIMEBOOST_net_10555), .b(g63547_db), .o(n_4610) );
na02s01 g63616_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__Q), .b(FE_OFN1079_n_4778), .o(g63616_db) );
na02s01 TIMEBOOST_cell_36636 ( .a(TIMEBOOST_net_10556), .b(g63588_db), .o(n_4100) );
in01s02 g63617_u0 ( .a(FE_OFN2021_n_4778), .o(g63617_sb) );
na02s01 g63617_u1 ( .a(wbs_dat_i_19_), .b(g63617_sb), .o(g63617_da) );
na02s02 TIMEBOOST_cell_38469 ( .a(wbm_adr_o_12_), .b(n_2720), .o(TIMEBOOST_net_11473) );
na02s01 TIMEBOOST_cell_36350 ( .a(TIMEBOOST_net_10413), .b(g67051_sb), .o(n_1452) );
in01s01 g63618_u0 ( .a(FE_OFN2022_n_4778), .o(g63618_sb) );
na02f02 TIMEBOOST_cell_36638 ( .a(TIMEBOOST_net_10557), .b(n_15436), .o(TIMEBOOST_net_473) );
na02s01 g63618_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__Q), .b(FE_OFN1079_n_4778), .o(g63618_db) );
na02s01 TIMEBOOST_cell_36468 ( .a(TIMEBOOST_net_10472), .b(g65787_db), .o(n_1908) );
in01s01 g63619_u0 ( .a(FE_OFN1079_n_4778), .o(g63619_sb) );
na02s01 g63619_u1 ( .a(wbs_dat_i_8_), .b(g63619_sb), .o(g63619_da) );
na02s01 g63619_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__Q), .b(FE_OFN1079_n_4778), .o(g63619_db) );
na02f02 TIMEBOOST_cell_10881 ( .a(TIMEBOOST_net_2007), .b(n_15406), .o(n_13124) );
in01s01 g63620_u0 ( .a(FE_OFN2022_n_4778), .o(g63620_sb) );
na02f02 TIMEBOOST_cell_45800 ( .a(TIMEBOOST_net_15138), .b(FE_OFN2167_n_8567), .o(TIMEBOOST_net_14581) );
na02f04 TIMEBOOST_cell_37020 ( .a(TIMEBOOST_net_10748), .b(g52518_sb), .o(n_13705) );
na02s01 TIMEBOOST_cell_36470 ( .a(TIMEBOOST_net_10473), .b(g65714_db), .o(TIMEBOOST_net_246) );
in01s02 g63621_u0 ( .a(FE_OFN2021_n_4778), .o(g63621_sb) );
na02s01 g63621_u1 ( .a(wbs_dat_i_29_), .b(g63621_sb), .o(g63621_da) );
na02s02 TIMEBOOST_cell_45682 ( .a(TIMEBOOST_net_15079), .b(FE_OFN1218_n_6886), .o(TIMEBOOST_net_12570) );
na02s01 TIMEBOOST_cell_36352 ( .a(TIMEBOOST_net_10414), .b(FE_OFN2094_n_2520), .o(n_2521) );
in01f20 g63667_u0 ( .a(pciu_cache_lsize_not_zero_in), .o(n_3319) );
na02s02 g63682_u0 ( .a(n_3809), .b(n_1472), .o(n_4746) );
in01m02 g63695_u0 ( .a(FE_OFN1155_n_3464), .o(n_4098) );
in01m02 g63708_u0 ( .a(FE_OFN1154_n_3464), .o(n_4097) );
in01m02 g63721_u0 ( .a(FE_OFN1155_n_3464), .o(n_4096) );
in01m02 g63734_u0 ( .a(FE_OFN1154_n_3464), .o(n_4095) );
in01m02 g63747_u0 ( .a(FE_OFN1155_n_3464), .o(n_4143) );
in01m02 g63773_u0 ( .a(FE_OFN1154_n_3464), .o(n_4093) );
in01m02 g63786_u0 ( .a(FE_OFN1155_n_3464), .o(n_4092) );
in01m04 g63799_u0 ( .a(FE_OFN1155_n_3464), .o(n_6391) );
in01s02 g63803_u0 ( .a(FE_OFN1154_n_3464), .o(n_6886) );
in01m02 g63834_u0 ( .a(FE_OFN1154_n_3464), .o(n_4151) );
in01s02 g63838_u0 ( .a(FE_OFN1154_n_3464), .o(n_6356) );
in01m01 g63847_u0 ( .a(FE_OFN1155_n_3464), .o(n_4090) );
in01s06 g63853_u0 ( .a(n_4658), .o(n_6431) );
in01f06 g63860_u0 ( .a(n_4658), .o(n_6436) );
in01s06 g63861_u0 ( .a(n_4658), .o(n_6554) );
in01s06 g63862_u0 ( .a(n_4658), .o(n_6319) );
in01s06 g63864_u0 ( .a(n_4658), .o(n_6287) );
in01s06 g63868_u0 ( .a(n_4658), .o(n_6645) );
in01s06 g63870_u0 ( .a(n_4658), .o(n_6232) );
in01m20 g63881_u0 ( .a(n_4658), .o(n_6624) );
in01f20 g63888_u0 ( .a(FE_OFN1192_n_6935), .o(n_4658) );
in01f08 g63889_u0 ( .a(FE_OFN1155_n_3464), .o(n_6935) );
na02f06 g63890_u0 ( .a(n_3314), .b(n_3313), .o(n_3464) );
no02s02 g63891_u0 ( .a(n_868), .b(FE_OFN1117_g64577_p), .o(g63891_p) );
in01s02 g63891_u1 ( .a(g63891_p), .o(n_4637) );
na02s01 g63892_u0 ( .a(n_646), .b(n_1825), .o(g63892_p) );
in01s01 g63892_u1 ( .a(g63892_p), .o(n_2445) );
no02s01 g63894_u0 ( .a(n_963), .b(FE_OFN778_n_4152), .o(n_2938) );
na02f02 g63895_u0 ( .a(n_3053), .b(n_4806), .o(g63895_p) );
in01f02 g63895_u1 ( .a(g63895_p), .o(n_3424) );
in01m01 g63896_u0 ( .a(n_2950), .o(n_14389) );
no02f08 g63897_u0 ( .a(n_1964), .b(n_2443), .o(n_2950) );
na02s01 g63899_u0 ( .a(FE_OFN1024_n_11877), .b(n_16818), .o(n_3423) );
in01f01 g63900_u0 ( .a(n_3421), .o(n_3422) );
na02m02 g63902_u0 ( .a(n_2441), .b(n_2433), .o(g63902_p) );
in01f02 g63902_u1 ( .a(g63902_p), .o(n_2442) );
na02f02 g63905_u0 ( .a(n_2727), .b(FE_OFN1619_n_1787), .o(n_2728) );
na02f02 g63907_u0 ( .a(n_2814), .b(n_2813), .o(n_3306) );
no02s02 g63908_u0 ( .a(n_1701), .b(FE_OFN778_n_4152), .o(n_2937) );
na02s01 g63909_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_), .b(FE_OFN1117_g64577_p), .o(n_3420) );
na02f02 g63910_u0 ( .a(n_3235), .b(n_2847), .o(n_4088) );
na02s02 g63911_u0 ( .a(n_2716), .b(wbu_addr_in_268), .o(n_2717) );
na02s02 g63912_u0 ( .a(n_2714), .b(wbu_addr_in_269), .o(n_2715) );
na02s02 TIMEBOOST_cell_45221 ( .a(n_4252), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__Q), .o(TIMEBOOST_net_14849) );
no02s01 g63914_u0 ( .a(n_4533), .b(wishbone_slave_unit_pci_initiator_sm_decode_count_0_), .o(n_4537) );
na02m02 g63915_u0 ( .a(n_2712), .b(wbu_addr_in_272), .o(n_2713) );
na02f04 g63916_u0 ( .a(n_2727), .b(wishbone_slave_unit_pci_initiator_if_current_byte_address), .o(g63916_p) );
in01f02 g63916_u1 ( .a(g63916_p), .o(n_2711) );
na02s02 TIMEBOOST_cell_42112 ( .a(TIMEBOOST_net_13294), .b(FE_OFN1317_n_6624), .o(TIMEBOOST_net_11598) );
na02s02 g63919_u0 ( .a(FE_OFN1117_g64577_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_), .o(n_3419) );
na02s01 g63920_u0 ( .a(FE_OFN1092_g64577_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_0_), .o(n_3417) );
na02s02 g63921_u0 ( .a(n_3415), .b(FE_OFN1117_g64577_p), .o(n_3416) );
na02s02 g63922_u0 ( .a(n_2437), .b(n_2431), .o(g63922_p) );
in01s02 g63922_u1 ( .a(g63922_p), .o(n_2438) );
na02s01 TIMEBOOST_cell_37267 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__Q), .b(n_3792), .o(TIMEBOOST_net_10872) );
in01s01 g63924_u0 ( .a(n_4535), .o(n_4536) );
no02m01 g63925_u0 ( .a(wishbone_slave_unit_pcim_sm_rdy_in), .b(FE_OFN999_n_15978), .o(g63925_p) );
in01s02 g63925_u1 ( .a(g63925_p), .o(n_4535) );
no02m02 g63926_u0 ( .a(FE_OFN967_n_2233), .b(n_3080), .o(n_3413) );
no02s06 g63927_u0 ( .a(FE_OFN1117_g64577_p), .b(pci_target_unit_fifos_pciw_control_in), .o(n_5546) );
no02s02 g63929_u0 ( .a(n_2231), .b(n_2232), .o(n_2710) );
na02m04 g63930_u0 ( .a(n_2722), .b(n_2435), .o(n_2436) );
na02s02 g63933_u0 ( .a(n_2934), .b(wbm_adr_o_19_), .o(n_2935) );
no02s01 g63934_u0 ( .a(n_1204), .b(n_4533), .o(n_4534) );
no02m02 g63935_u0 ( .a(n_2402), .b(n_2401), .o(g63935_p) );
in01s02 g63935_u1 ( .a(g63935_p), .o(n_2933) );
no02m02 g63936_u0 ( .a(n_2400), .b(n_2876), .o(n_3305) );
no02f04 g63938_u0 ( .a(n_2214), .b(FE_OCP_RBN2239_g74749_p), .o(n_4642) );
na02f02 g63939_u0 ( .a(pci_target_unit_wishbone_master_burst_chopped), .b(FE_OCP_RBN2237_g74749_p), .o(g63939_p) );
in01f02 g63939_u1 ( .a(g63939_p), .o(n_3410) );
na02f03 g63940_u0 ( .a(n_3304), .b(n_16159), .o(n_4674) );
no02f02 g63941_u0 ( .a(n_1998), .b(FE_OCP_RBN2239_g74749_p), .o(n_3409) );
no02s01 g63942_u0 ( .a(FE_OFN778_n_4152), .b(pci_target_unit_del_sync_comp_cycle_count_0_), .o(n_2932) );
na02s02 TIMEBOOST_cell_39974 ( .a(TIMEBOOST_net_12225), .b(g62885_sb), .o(n_6107) );
na02s01 TIMEBOOST_cell_42600 ( .a(TIMEBOOST_net_13538), .b(g65684_db), .o(n_1954) );
in01m02 g63943_u3 ( .a(g63943_p), .o(n_2264) );
no02f06 g63944_u0 ( .a(n_3047), .b(n_1192), .o(n_3408) );
na02s02 TIMEBOOST_cell_43608 ( .a(TIMEBOOST_net_14042), .b(FE_OFN1316_n_6624), .o(TIMEBOOST_net_12224) );
na02f02 TIMEBOOST_cell_41608 ( .a(FE_OFN1440_n_9372), .b(TIMEBOOST_net_13042), .o(TIMEBOOST_net_11653) );
na02m08 g63947_u0 ( .a(n_2218), .b(n_6986), .o(n_4662) );
no02s02 g63948_u0 ( .a(n_1484), .b(n_2009), .o(n_2477) );
na02s04 TIMEBOOST_cell_45518 ( .a(TIMEBOOST_net_14997), .b(g54339_sb), .o(n_12978) );
no02s02 g63950_u0 ( .a(n_1485), .b(n_2007), .o(n_2473) );
na02s02 g63951_u0 ( .a(n_2706), .b(wbm_adr_o_20_), .o(n_2707) );
na02s01 TIMEBOOST_cell_15858 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_81), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3186) );
na02f02 g63954_u0 ( .a(n_5230), .b(n_3077), .o(n_3407) );
na02m02 TIMEBOOST_cell_22424 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__Q), .o(TIMEBOOST_net_6469) );
ao12f02 g63957_u0 ( .a(n_3071), .b(FE_OCPN1845_n_16427), .c(n_3404), .o(n_3406) );
na02f02 g63958_u0 ( .a(n_2840), .b(n_2621), .o(n_3302) );
na02f02 g63959_u0 ( .a(FE_OFN1944_n_15813), .b(n_2984), .o(n_3301) );
na02s01 TIMEBOOST_cell_43012 ( .a(TIMEBOOST_net_13744), .b(n_4008), .o(n_5446) );
ao12f02 g63963_u0 ( .a(n_3042), .b(FE_OCPN1845_n_16427), .c(n_3078), .o(n_3403) );
na02s01 TIMEBOOST_cell_21939 ( .a(TIMEBOOST_net_6226), .b(g63048_sb), .o(n_5156) );
ao12s01 g63965_u0 ( .a(pci_target_unit_del_sync_req_comp_pending_sample), .b(n_3795), .c(g66433_sb), .o(n_4532) );
na02m02 TIMEBOOST_cell_44243 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__Q), .b(n_9130), .o(TIMEBOOST_net_14360) );
na02m02 TIMEBOOST_cell_38688 ( .a(TIMEBOOST_net_11582), .b(n_7618), .o(TIMEBOOST_net_10678) );
oa12s01 g63969_u0 ( .a(n_4084), .b(n_3386), .c(FE_OFN2121_n_2687), .o(n_4085) );
na02s02 TIMEBOOST_cell_43563 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__Q), .b(n_4232), .o(TIMEBOOST_net_14020) );
ao22f02 g63976_u0 ( .a(n_1013), .b(n_1626), .c(n_2430), .d(wishbone_slave_unit_pci_initiator_if_current_byte_address_36), .o(n_2959) );
na02s02 TIMEBOOST_cell_39498 ( .a(TIMEBOOST_net_11987), .b(g63081_sb), .o(n_5090) );
ao12f02 g63980_u0 ( .a(n_3084), .b(n_3372), .c(wbu_pref_en_in_137), .o(n_3399) );
ao12s04 g63981_u0 ( .a(FE_OFN1125_g64577_p), .b(n_980), .c(n_813), .o(n_4131) );
ao12f02 g63982_u0 ( .a(n_3119), .b(n_4718), .c(n_2344), .o(n_3120) );
na02f02 TIMEBOOST_cell_42202 ( .a(TIMEBOOST_net_13339), .b(FE_OFN1419_n_8567), .o(TIMEBOOST_net_12291) );
oa12s01 g63985_u0 ( .a(n_1488), .b(n_4904), .c(FE_OFN672_n_4505), .o(n_4918) );
oa12s01 g63986_u0 ( .a(n_2138), .b(n_4904), .c(FE_OFN665_n_4495), .o(n_4917) );
oa12s01 g63987_u0 ( .a(n_4510), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_14__583), .c(FE_OFN1640_n_4671), .o(n_4915) );
oa12s01 g63988_u0 ( .a(n_1642), .b(n_4904), .c(FE_OFN634_n_4454), .o(n_4914) );
no02s02 g63989_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_6_), .b(n_1417), .o(g63989_p) );
ao12s02 g63989_u1 ( .a(g63989_p), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_6_), .c(n_1417), .o(n_2262) );
oa12s01 g63990_u0 ( .a(n_1559), .b(n_4904), .c(FE_OFN614_n_4501), .o(n_4913) );
oa12s01 g63991_u0 ( .a(n_1555), .b(n_4904), .c(FE_OFN622_n_4409), .o(n_4912) );
oa12s02 g63992_u0 ( .a(n_1546), .b(n_4904), .c(FE_OFN659_n_4392), .o(n_4911) );
oa12s01 g63993_u0 ( .a(n_4513), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_11__466), .c(n_4677), .o(n_4909) );
ao22f02 g63_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__Q), .b(n_15568), .c(n_15566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__Q), .o(n_15529) );
in01m10 g64011_u0 ( .a(n_4743), .o(n_8440) );
oa12s01 g64016_u0 ( .a(n_1553), .b(n_4904), .c(FE_OFN648_n_4497), .o(n_4908) );
oa12s01 g64017_u0 ( .a(n_4511), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_7__310), .c(FE_OFN1678_n_4655), .o(n_4907) );
oa12s01 g64018_u0 ( .a(n_2131), .b(n_4904), .c(n_4417), .o(n_4906) );
oa12s02 g64019_u0 ( .a(n_1547), .b(n_4904), .c(FE_OFN1623_n_4438), .o(n_4905) );
oa12s01 g64020_u0 ( .a(n_4509), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_15__622), .c(FE_OFN651_n_4508), .o(n_4903) );
oa12s01 g64021_u0 ( .a(n_4514), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__544), .c(n_4669), .o(n_4902) );
no02s01 g64022_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_5_), .b(n_1015), .o(g64022_p) );
ao12s02 g64022_u1 ( .a(g64022_p), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_5_), .c(n_1015), .o(n_1688) );
oa12s01 g64023_u0 ( .a(n_1537), .b(n_4904), .c(FE_OFN682_n_4460), .o(n_4901) );
oa12s01 g64024_u0 ( .a(n_1377), .b(n_4904), .c(FE_OFN1660_n_4490), .o(n_4900) );
na04f04 TIMEBOOST_cell_36227 ( .a(n_13060), .b(n_12917), .c(n_12918), .d(n_12797), .o(n_13140) );
ao22m02 g64027_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_486), .c(configuration_wb_err_addr_548), .d(n_15445), .o(n_2927) );
ao22f02 g64028_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_492), .c(n_16791), .d(pciu_bar0_in_370), .o(n_2926) );
ao22f02 g64029_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_487), .c(n_16791), .d(pciu_bar0_in_365), .o(n_2925) );
ao22f02 g64030_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_488), .c(n_16791), .d(pciu_bar0_in_366), .o(n_2924) );
ao22f02 g64031_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_473), .c(configuration_interrupt_line_39), .d(n_3295), .o(n_3297) );
ao22f01 g64033_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_471), .c(configuration_interrupt_line_37), .d(n_3295), .o(n_3296) );
ao22m01 g64034_u0 ( .a(n_3115), .b(configuration_icr_bit_2961), .c(configuration_wb_err_addr_533), .d(n_15444), .o(n_3117) );
ao22f02 g64035_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_493), .c(configuration_wb_err_addr_555), .d(n_15445), .o(n_2922) );
ao22f02 g64036_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_495), .c(n_3252), .d(configuration_pci_err_cs_bit_464), .o(n_2921) );
in01f01 g64038_u0 ( .a(n_15645), .o(n_4795) );
ao22f02 g64041_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_501), .c(n_3252), .d(configuration_pci_err_cs_bit_470), .o(n_2920) );
ao22f02 g64042_u0 ( .a(n_3115), .b(pci_resi_conf_soft_res_in), .c(configuration_wb_err_addr_563), .d(n_15444), .o(n_3116) );
ao22f02 g64043_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_505), .c(FE_OFN1006_n_16288), .d(configuration_pci_err_addr_474), .o(n_2919) );
ao22m02 g64044_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_508), .c(FE_OFN1006_n_16288), .d(configuration_pci_err_addr_477), .o(n_2918) );
na02f02 TIMEBOOST_cell_42152 ( .a(TIMEBOOST_net_13314), .b(g57044_sb), .o(n_11690) );
na02s02 TIMEBOOST_cell_39976 ( .a(TIMEBOOST_net_12226), .b(g62433_sb), .o(n_6731) );
na02m04 TIMEBOOST_cell_45826 ( .a(TIMEBOOST_net_15151), .b(FE_OFN2134_n_13124), .o(TIMEBOOST_net_14993) );
ao22f02 g64048_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_475), .c(configuration_interrupt_line_41), .d(n_3295), .o(n_3294) );
ao22f02 g64049_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_491), .c(n_16791), .d(pciu_bar0_in_369), .o(n_2917) );
ao22f02 g64050_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_476), .c(configuration_interrupt_line_42), .d(n_3295), .o(n_3393) );
in01f02 g64051_u0 ( .a(n_2916), .o(n_3114) );
ao22f02 g64052_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_500), .c(n_3252), .d(configuration_pci_err_cs_bit_469), .o(n_2916) );
na03s02 TIMEBOOST_cell_5971 ( .a(n_4645), .b(g64974_sb), .c(g64974_db), .o(n_4369) );
na02s01 TIMEBOOST_cell_41692 ( .a(TIMEBOOST_net_13084), .b(wishbone_slave_unit_pci_initiator_sm_transfer), .o(TIMEBOOST_net_1098) );
ao22f02 g64055_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_490), .c(n_16791), .d(pciu_bar0_in_368), .o(n_2913) );
na02m02 TIMEBOOST_cell_42203 ( .a(n_9453), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q), .o(TIMEBOOST_net_13340) );
in01f02 g64060_u0 ( .a(n_2910), .o(n_3112) );
ao22f02 g64061_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_497), .c(n_3252), .d(configuration_pci_err_cs_bit_466), .o(n_2910) );
in01f02 g64062_u0 ( .a(n_2909), .o(n_3111) );
ao22f02 g64063_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_498), .c(n_3252), .d(configuration_pci_err_cs_bit_467), .o(n_2909) );
ao22s02 g64064_u0 ( .a(n_2699), .b(wbu_map_in_131), .c(n_2698), .d(wbu_map_in_132), .o(n_2700) );
ao22m02 g64065_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr), .c(configuration_wb_err_addr), .d(n_15445), .o(n_15435) );
ao22s02 g64066_u0 ( .a(n_2699), .b(wbu_pref_en_in_136), .c(n_2698), .d(wbu_pref_en_in_137), .o(n_2697) );
in01f02 g64067_u0 ( .a(n_2907), .o(n_3110) );
ao22f02 g64068_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_499), .c(n_3252), .d(configuration_pci_err_cs_bit_468), .o(n_2907) );
ao22f01 g64069_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_472), .c(configuration_interrupt_line_38), .d(n_3295), .o(n_3293) );
ao22m02 g64070_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_481), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_245), .o(n_2906) );
ao22s02 g64071_u0 ( .a(n_2699), .b(wbu_mrl_en_in_141), .c(n_2698), .d(wbu_mrl_en_in_142), .o(n_2696) );
ao22f02 g64072_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_482), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_246), .o(n_2905) );
ao22m02 g64073_u0 ( .a(n_3115), .b(configuration_icr_bit_2967), .c(configuration_wb_err_addr_534), .d(n_15444), .o(n_3109) );
ao22f02 g64074_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_483), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_247), .o(n_2904) );
ao22f02 g64075_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_484), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_248), .o(n_15434) );
ao22m02 g64076_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_496), .c(n_3252), .d(configuration_pci_err_cs_bit_465), .o(n_2902) );
ao22f02 g64077_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_485), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_249), .o(n_16852) );
in01s01 g64078_u0 ( .a(FE_OFN1077_n_4740), .o(g64078_sb) );
na02s01 TIMEBOOST_cell_16039 ( .a(TIMEBOOST_net_3276), .b(n_2515), .o(n_2516) );
na02s02 TIMEBOOST_cell_45222 ( .a(TIMEBOOST_net_14849), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_13265) );
na02s02 TIMEBOOST_cell_19163 ( .a(TIMEBOOST_net_4838), .b(g59093_sb), .o(TIMEBOOST_net_2409) );
in01s01 g64079_u0 ( .a(FE_OFN1046_n_16657), .o(g64079_sb) );
na02s02 TIMEBOOST_cell_39978 ( .a(TIMEBOOST_net_12227), .b(g63159_sb), .o(n_5819) );
na02s01 g64079_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__Q), .b(FE_OFN1046_n_16657), .o(g64079_db) );
na02m02 TIMEBOOST_cell_39980 ( .a(TIMEBOOST_net_12228), .b(g62416_sb), .o(n_6766) );
in01s01 g64080_u0 ( .a(FE_OFN1077_n_4740), .o(g64080_sb) );
na02s01 TIMEBOOST_cell_38476 ( .a(TIMEBOOST_net_11476), .b(g61899_sb), .o(n_7981) );
na02s01 g64080_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__12__Q), .b(FE_OFN1077_n_4740), .o(g64080_db) );
na02s01 TIMEBOOST_cell_18471 ( .a(TIMEBOOST_net_4492), .b(g63100_sb), .o(n_5054) );
in01s01 g64081_u0 ( .a(FE_OFN1075_n_4740), .o(g64081_sb) );
na02f02 TIMEBOOST_cell_44266 ( .a(TIMEBOOST_net_14371), .b(FE_OFN1405_n_8567), .o(TIMEBOOST_net_12831) );
na02s01 g64081_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__Q), .b(FE_OFN1075_n_4740), .o(g64081_db) );
na02f02 TIMEBOOST_cell_38802 ( .a(TIMEBOOST_net_11639), .b(FE_OFN2168_n_8567), .o(n_11555) );
in01s01 g64082_u0 ( .a(FE_OFN1077_n_4740), .o(g64082_sb) );
na02s02 TIMEBOOST_cell_38588 ( .a(TIMEBOOST_net_11532), .b(g60645_sb), .o(n_5682) );
na02s01 g64082_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__Q), .b(FE_OFN1077_n_4740), .o(g64082_db) );
na02s02 TIMEBOOST_cell_18475 ( .a(TIMEBOOST_net_4494), .b(g59372_sb), .o(n_7689) );
in01s01 g64083_u0 ( .a(FE_OFN1076_n_4740), .o(g64083_sb) );
na02s01 TIMEBOOST_cell_18109 ( .a(TIMEBOOST_net_4311), .b(g63089_sb), .o(n_5076) );
na02s01 g64083_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__Q), .b(FE_OFN1076_n_4740), .o(g64083_db) );
na02s02 TIMEBOOST_cell_10377 ( .a(TIMEBOOST_net_1755), .b(g61829_sb), .o(n_8128) );
in01s01 g64084_u0 ( .a(FE_OFN1077_n_4740), .o(g64084_sb) );
na02s01 TIMEBOOST_cell_38478 ( .a(TIMEBOOST_net_11477), .b(g61922_db), .o(n_7977) );
na02s01 g64084_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__Q), .b(FE_OFN1077_n_4740), .o(g64084_db) );
na02s01 TIMEBOOST_cell_18477 ( .a(TIMEBOOST_net_4495), .b(g59378_sb), .o(n_7683) );
in01s01 g64085_u0 ( .a(FE_OFN906_n_4736), .o(g64085_sb) );
na02m02 TIMEBOOST_cell_44635 ( .a(n_9831), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__Q), .o(TIMEBOOST_net_14556) );
na02s01 g64085_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__Q), .b(FE_OFN906_n_4736), .o(g64085_db) );
na02s02 TIMEBOOST_cell_15909 ( .a(TIMEBOOST_net_3211), .b(n_3083), .o(TIMEBOOST_net_150) );
in01s01 g64086_u0 ( .a(FE_OFN1075_n_4740), .o(g64086_sb) );
na02s01 g64086_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__Q), .b(FE_OFN1077_n_4740), .o(g64086_db) );
na02s02 TIMEBOOST_cell_39982 ( .a(TIMEBOOST_net_12229), .b(g62560_sb), .o(n_6440) );
in01s01 g64087_u0 ( .a(FE_OFN906_n_4736), .o(g64087_sb) );
na03f02 TIMEBOOST_cell_36103 ( .a(FE_OFN1554_n_12104), .b(TIMEBOOST_net_10215), .c(FE_OCP_RBN1979_n_10273), .o(n_12597) );
na02s01 g64087_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__Q), .b(FE_OFN905_n_4736), .o(g64087_db) );
na02s02 TIMEBOOST_cell_43484 ( .a(TIMEBOOST_net_13980), .b(FE_OFN1233_n_6391), .o(TIMEBOOST_net_12175) );
in01s01 g64088_u0 ( .a(FE_OFN1075_n_4740), .o(g64088_sb) );
na03s02 TIMEBOOST_cell_43323 ( .a(n_4491), .b(FE_OFN1273_n_4096), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__Q), .o(TIMEBOOST_net_13900) );
na02s01 g64088_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__Q), .b(FE_OFN1075_n_4740), .o(g64088_db) );
na02s02 TIMEBOOST_cell_38480 ( .a(TIMEBOOST_net_11478), .b(FE_OFN1697_n_5751), .o(TIMEBOOST_net_4832) );
in01s01 g64089_u0 ( .a(FE_OFN1077_n_4740), .o(g64089_sb) );
na02m02 TIMEBOOST_cell_44197 ( .a(n_9512), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__Q), .o(TIMEBOOST_net_14337) );
na02s01 g64089_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__Q), .b(FE_OFN1077_n_4740), .o(g64089_db) );
na02f04 TIMEBOOST_cell_39028 ( .a(TIMEBOOST_net_11752), .b(FE_OFN2242_g52675_p), .o(TIMEBOOST_net_10754) );
in01s01 g64090_u0 ( .a(FE_OFN1046_n_16657), .o(g64090_sb) );
na02s01 TIMEBOOST_cell_42624 ( .a(TIMEBOOST_net_13550), .b(g64799_db), .o(n_3757) );
na02s01 g64090_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__Q), .b(FE_OFN1046_n_16657), .o(g64090_db) );
in01s01 g64091_u0 ( .a(FE_OFN1051_n_16657), .o(g64091_sb) );
na02s01 g64091_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__13__Q), .b(FE_OFN1051_n_16657), .o(g64091_db) );
na02s02 TIMEBOOST_cell_39984 ( .a(TIMEBOOST_net_12230), .b(g62407_sb), .o(n_6785) );
in01s01 g64092_u0 ( .a(FE_OFN1075_n_4740), .o(g64092_sb) );
na02f02 TIMEBOOST_cell_10386 ( .a(FE_OFN2128_n_16497), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_12__Q), .o(TIMEBOOST_net_1760) );
na02s01 g64092_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__Q), .b(FE_OFN1075_n_4740), .o(g64092_db) );
na02f02 TIMEBOOST_cell_18455 ( .a(TIMEBOOST_net_4484), .b(n_3440), .o(TIMEBOOST_net_530) );
in01s01 g64093_u0 ( .a(FE_OFN1049_n_16657), .o(g64093_sb) );
na02s01 g64093_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_127), .b(g64093_sb), .o(g64093_da) );
na02s01 g64093_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__Q), .b(FE_OFN1049_n_16657), .o(g64093_db) );
na02s02 TIMEBOOST_cell_38583 ( .a(TIMEBOOST_net_9932), .b(FE_OFN1181_n_3476), .o(TIMEBOOST_net_11530) );
in01s01 g64094_u0 ( .a(FE_OFN1074_n_4740), .o(g64094_sb) );
na02s01 TIMEBOOST_cell_17130 ( .a(FE_OFN217_n_9889), .b(FE_OFN572_n_9502), .o(TIMEBOOST_net_3822) );
na02s01 g64094_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__Q), .b(FE_OFN1074_n_4740), .o(g64094_db) );
na02s01 TIMEBOOST_cell_17131 ( .a(TIMEBOOST_net_3822), .b(TIMEBOOST_net_1405), .o(n_9499) );
in01s01 g64095_u0 ( .a(FE_OFN905_n_4736), .o(g64095_sb) );
na02f02 TIMEBOOST_cell_40885 ( .a(n_9813), .b(g57115_sb), .o(TIMEBOOST_net_12681) );
na02s01 g64095_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__Q), .b(FE_OFN905_n_4736), .o(g64095_db) );
na02s01 TIMEBOOST_cell_42919 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__Q), .b(FE_OFN580_n_9531), .o(TIMEBOOST_net_13698) );
in01s01 g64096_u0 ( .a(FE_OFN905_n_4736), .o(g64096_sb) );
na02s01 g64096_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_142), .b(g64096_sb), .o(g64096_da) );
na02s01 g64096_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__22__Q), .b(FE_OFN905_n_4736), .o(g64096_db) );
in01s01 g64097_u0 ( .a(FE_OFN1049_n_16657), .o(g64097_sb) );
na02s01 TIMEBOOST_cell_9884 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__Q), .b(g58284_sb), .o(TIMEBOOST_net_1509) );
na02s01 g64097_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__Q), .b(FE_OFN1049_n_16657), .o(g64097_db) );
na02s01 TIMEBOOST_cell_9885 ( .a(TIMEBOOST_net_1509), .b(g58284_db), .o(n_9518) );
in01s01 g64098_u0 ( .a(FE_OFN1049_n_16657), .o(g64098_sb) );
na02s02 TIMEBOOST_cell_45200 ( .a(TIMEBOOST_net_14838), .b(FE_OFN1264_n_4095), .o(TIMEBOOST_net_12101) );
na02s01 g64098_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__Q), .b(FE_OFN1049_n_16657), .o(g64098_db) );
na02s02 TIMEBOOST_cell_39986 ( .a(TIMEBOOST_net_12231), .b(g62660_sb), .o(n_6223) );
in01s01 g64099_u0 ( .a(FE_OFN1049_n_16657), .o(g64099_sb) );
na02s02 TIMEBOOST_cell_45157 ( .a(n_4238), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__Q), .o(TIMEBOOST_net_14817) );
na02s01 g64099_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__Q), .b(FE_OFN1049_n_16657), .o(g64099_db) );
na02m02 TIMEBOOST_cell_39988 ( .a(TIMEBOOST_net_12232), .b(g62968_sb), .o(n_5946) );
in01s01 g64100_u0 ( .a(FE_OFN1076_n_4740), .o(g64100_sb) );
na02f02 TIMEBOOST_cell_17132 ( .a(configuration_pci_err_data_513), .b(n_16429), .o(TIMEBOOST_net_3823) );
na02s01 g64100_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__Q), .b(FE_OFN1076_n_4740), .o(g64100_db) );
na02s02 TIMEBOOST_cell_45158 ( .a(TIMEBOOST_net_14817), .b(FE_OFN1248_n_4093), .o(TIMEBOOST_net_12651) );
oa12s01 g64101_u0 ( .a(n_1815), .b(FE_OFN923_n_4740), .c(pci_target_unit_fifos_pciw_control_in), .o(n_4528) );
in01s01 g64102_u0 ( .a(FE_OFN905_n_4736), .o(g64102_sb) );
na02s01 g64102_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_141), .b(g64102_sb), .o(g64102_da) );
na02s01 g64102_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__Q), .b(FE_OFN905_n_4736), .o(g64102_db) );
na02s02 TIMEBOOST_cell_45098 ( .a(TIMEBOOST_net_14787), .b(FE_OFN1812_n_7845), .o(TIMEBOOST_net_11387) );
in01s01 g64103_u0 ( .a(FE_OFN1076_n_4740), .o(g64103_sb) );
na02s01 g64103_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__Q), .b(FE_OFN1076_n_4740), .o(g64103_db) );
na02s02 TIMEBOOST_cell_39990 ( .a(TIMEBOOST_net_12233), .b(g62561_sb), .o(n_6438) );
oa12s01 g64104_u0 ( .a(n_1795), .b(FE_OFN1046_n_16657), .c(pci_target_unit_fifos_pciw_control_in), .o(n_4527) );
in01s01 g64105_u0 ( .a(FE_OFN904_n_4736), .o(g64105_sb) );
na02s01 g64105_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_150), .b(g64105_sb), .o(g64105_da) );
na02s01 g64105_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__Q), .b(FE_OFN904_n_4736), .o(g64105_db) );
na02s01 TIMEBOOST_cell_44972 ( .a(TIMEBOOST_net_14724), .b(FE_OFN1801_n_9690), .o(TIMEBOOST_net_11012) );
in01s01 g64106_u0 ( .a(FE_OFN1046_n_16657), .o(g64106_sb) );
na02s01 g64106_u1 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(g64106_sb), .o(g64106_da) );
na02s01 g64106_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__Q), .b(FE_OFN1046_n_16657), .o(g64106_db) );
na02s01 TIMEBOOST_cell_38585 ( .a(TIMEBOOST_net_4789), .b(FE_OFN1183_n_3476), .o(TIMEBOOST_net_11531) );
in01s01 g64107_u0 ( .a(FE_OFN1049_n_16657), .o(g64107_sb) );
na02s01 TIMEBOOST_cell_9890 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__Q), .b(g65360_sb), .o(TIMEBOOST_net_1512) );
na02s01 g64107_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__Q), .b(FE_OFN1049_n_16657), .o(g64107_db) );
na02s01 TIMEBOOST_cell_9891 ( .a(TIMEBOOST_net_1512), .b(g65360_db), .o(n_3537) );
in01s01 g64108_u0 ( .a(FE_OFN1046_n_16657), .o(g64108_sb) );
na02s01 g64108_u1 ( .a(pci_target_unit_fifos_pciw_cbe_in_153), .b(g64108_sb), .o(g64108_da) );
na02s01 g64108_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__Q), .b(FE_OFN1046_n_16657), .o(g64108_db) );
na02s02 TIMEBOOST_cell_43626 ( .a(TIMEBOOST_net_14051), .b(FE_OFN1314_n_6624), .o(TIMEBOOST_net_12237) );
in01s01 g64109_u0 ( .a(FE_OFN1076_n_4740), .o(g64109_sb) );
na02s02 TIMEBOOST_cell_45159 ( .a(n_4233), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__Q), .o(TIMEBOOST_net_14818) );
na02s01 g64109_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__Q), .b(FE_OFN1076_n_4740), .o(g64109_db) );
na02s02 TIMEBOOST_cell_39992 ( .a(TIMEBOOST_net_12234), .b(g62593_sb), .o(n_6366) );
in01s01 g64110_u0 ( .a(FE_OFN1046_n_16657), .o(g64110_sb) );
na02s02 TIMEBOOST_cell_45160 ( .a(TIMEBOOST_net_14818), .b(FE_OFN1194_n_6935), .o(TIMEBOOST_net_12650) );
na02s01 g64110_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__Q), .b(FE_OFN1046_n_16657), .o(g64110_db) );
na02m02 TIMEBOOST_cell_39994 ( .a(TIMEBOOST_net_12235), .b(g62983_sb), .o(n_5916) );
in01s01 g64111_u0 ( .a(FE_OFN1074_n_4740), .o(g64111_sb) );
na02s01 TIMEBOOST_cell_39285 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(g65799_sb), .o(TIMEBOOST_net_11881) );
na02s01 g64111_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__Q), .b(FE_OFN1074_n_4740), .o(g64111_db) );
na02s01 TIMEBOOST_cell_39272 ( .a(TIMEBOOST_net_11874), .b(g64270_db), .o(n_3903) );
in01s01 g64112_u0 ( .a(FE_OFN1077_n_4740), .o(g64112_sb) );
na03s02 TIMEBOOST_cell_33910 ( .a(n_2559), .b(TIMEBOOST_net_905), .c(TIMEBOOST_net_471), .o(n_4892) );
na02s01 g64112_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__16__Q), .b(FE_OFN1077_n_4740), .o(g64112_db) );
na02s01 TIMEBOOST_cell_42896 ( .a(TIMEBOOST_net_13686), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_11156) );
in01s01 g64113_u0 ( .a(FE_OFN1046_n_16657), .o(g64113_sb) );
na02m04 TIMEBOOST_cell_17924 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__Q), .b(FE_OFN2059_n_13447), .o(TIMEBOOST_net_4219) );
na02s01 g64113_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__Q), .b(FE_OFN1049_n_16657), .o(g64113_db) );
na02f04 TIMEBOOST_cell_17925 ( .a(TIMEBOOST_net_4219), .b(FE_OFN1151_n_13249), .o(TIMEBOOST_net_1834) );
in01s01 g64114_u0 ( .a(FE_OFN937_n_2292), .o(g64114_sb) );
na02s01 g64114_u1 ( .a(pci_target_unit_fifos_pcir_control_in_192), .b(g64114_sb), .o(g64114_da) );
na02s01 g64114_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__Q), .b(FE_OFN937_n_2292), .o(g64114_db) );
na02s01 g64114_u3 ( .a(g64114_da), .b(g64114_db), .o(n_4525) );
in01s01 g64115_u0 ( .a(FE_OFN1076_n_4740), .o(g64115_sb) );
na02s02 TIMEBOOST_cell_42366 ( .a(TIMEBOOST_net_13421), .b(g54357_sb), .o(n_13085) );
na02s01 g64115_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__Q), .b(FE_OFN1076_n_4740), .o(g64115_db) );
na02s01 TIMEBOOST_cell_42907 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q), .b(FE_OFN580_n_9531), .o(TIMEBOOST_net_13692) );
in01s01 g64116_u0 ( .a(FE_OFN1049_n_16657), .o(g64116_sb) );
na02s01 TIMEBOOST_cell_18286 ( .a(g61943_sb), .b(g61943_db), .o(TIMEBOOST_net_4400) );
na02s01 g64116_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__Q), .b(FE_OFN1049_n_16657), .o(g64116_db) );
na02f06 TIMEBOOST_cell_38482 ( .a(TIMEBOOST_net_11479), .b(g54319_da), .o(n_13289) );
in01s01 g64117_u0 ( .a(FE_OFN1075_n_4740), .o(g64117_sb) );
na02f02 TIMEBOOST_cell_42953 ( .a(TIMEBOOST_net_9656), .b(FE_OFN1149_n_13249), .o(TIMEBOOST_net_13715) );
na02s01 g64117_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__Q), .b(FE_OFN1075_n_4740), .o(g64117_db) );
na02s02 TIMEBOOST_cell_41892 ( .a(TIMEBOOST_net_13184), .b(n_8757), .o(g52396_db) );
in01s01 g64118_u0 ( .a(FE_OFN908_n_4734), .o(g64118_sb) );
na02s01 TIMEBOOST_cell_31238 ( .a(n_3785), .b(g64950_sb), .o(TIMEBOOST_net_9530) );
na02s01 g64118_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__Q), .b(FE_OFN908_n_4734), .o(g64118_db) );
na02s01 TIMEBOOST_cell_31237 ( .a(TIMEBOOST_net_9529), .b(g64949_db), .o(n_3667) );
in01s01 g64119_u0 ( .a(FE_OFN906_n_4736), .o(g64119_sb) );
na02s01 g64119_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_149), .b(g64119_sb), .o(g64119_da) );
na02s01 g64119_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__Q), .b(FE_OFN906_n_4736), .o(g64119_db) );
na02s02 TIMEBOOST_cell_45099 ( .a(n_2152), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__Q), .o(TIMEBOOST_net_14788) );
in01s01 g64120_u0 ( .a(FE_OFN904_n_4736), .o(g64120_sb) );
na02s01 g64120_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_125), .b(g64120_sb), .o(g64120_da) );
na02s01 g64120_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__Q), .b(FE_OFN904_n_4736), .o(g64120_db) );
na02s02 TIMEBOOST_cell_45100 ( .a(TIMEBOOST_net_14788), .b(FE_OFN1812_n_7845), .o(TIMEBOOST_net_11381) );
oa12s01 g64121_u0 ( .a(n_1804), .b(FE_OFN903_n_4736), .c(pci_target_unit_fifos_pciw_control_in), .o(n_4524) );
in01s01 g64122_u0 ( .a(FE_OFN902_n_4736), .o(g64122_sb) );
na03f02 TIMEBOOST_cell_36104 ( .a(FE_OFN1554_n_12104), .b(TIMEBOOST_net_10212), .c(FE_OFN1513_n_14987), .o(n_12738) );
na02s01 g64122_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__Q), .b(FE_OFN902_n_4736), .o(g64122_db) );
na02s02 TIMEBOOST_cell_38716 ( .a(TIMEBOOST_net_11596), .b(g62633_sb), .o(n_6286) );
in01s01 g64123_u0 ( .a(FE_OFN904_n_4736), .o(g64123_sb) );
na02s01 g64123_u1 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(g64123_sb), .o(g64123_da) );
na02s01 g64123_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__Q), .b(FE_OFN904_n_4736), .o(g64123_db) );
na02s02 TIMEBOOST_cell_45101 ( .a(n_1863), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__Q), .o(TIMEBOOST_net_14789) );
no02s02 g64124_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_4_), .b(n_1176), .o(g64124_p) );
ao12s02 g64124_u1 ( .a(g64124_p), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_4_), .c(n_1176), .o(n_1750) );
in01s01 g64125_u0 ( .a(FE_OFN923_n_4740), .o(g64125_sb) );
na02s01 TIMEBOOST_cell_41693 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_71), .b(wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_13085) );
na02s01 g64125_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__Q), .b(FE_OFN923_n_4740), .o(g64125_db) );
na02s01 TIMEBOOST_cell_41928 ( .a(TIMEBOOST_net_13202), .b(g57895_db), .o(n_9229) );
in01s01 g64126_u0 ( .a(FE_OFN905_n_4736), .o(g64126_sb) );
na02s01 g64126_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_135), .b(g64126_sb), .o(g64126_da) );
na02s01 g64126_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q), .b(FE_OFN905_n_4736), .o(g64126_db) );
in01s01 g64127_u0 ( .a(FE_OFN1049_n_16657), .o(g64127_sb) );
na02f02 TIMEBOOST_cell_17926 ( .a(n_16452), .b(wishbone_slave_unit_wbs_sm_wbr_control_in_190), .o(TIMEBOOST_net_4220) );
na02s01 g64127_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__Q), .b(FE_OFN1049_n_16657), .o(g64127_db) );
na02f02 TIMEBOOST_cell_17927 ( .a(TIMEBOOST_net_4220), .b(n_7725), .o(TIMEBOOST_net_539) );
in01s01 g64128_u0 ( .a(FE_OFN905_n_4736), .o(g64128_sb) );
na02m02 TIMEBOOST_cell_32148 ( .a(FE_OFN2072_n_15978), .b(g53937_sb), .o(TIMEBOOST_net_9985) );
na02s01 g64128_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__Q), .b(FE_OFN905_n_4736), .o(g64128_db) );
na02f06 TIMEBOOST_cell_32147 ( .a(TIMEBOOST_net_9984), .b(n_16165), .o(TIMEBOOST_net_624) );
in01s01 g64129_u0 ( .a(FE_OFN1010_n_4734), .o(g64129_sb) );
na02s01 g64129_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_127), .b(g64129_sb), .o(g64129_da) );
na02s01 g64129_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__Q), .b(FE_OFN1010_n_4734), .o(g64129_db) );
na02s01 g64129_u3 ( .a(g64129_da), .b(g64129_db), .o(n_4033) );
in01s01 g64130_u0 ( .a(FE_OFN1013_n_4734), .o(g64130_sb) );
na02s01 TIMEBOOST_cell_31236 ( .a(n_3741), .b(g64949_sb), .o(TIMEBOOST_net_9529) );
na02s01 g64130_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__Q), .b(FE_OFN1013_n_4734), .o(g64130_db) );
na02s02 TIMEBOOST_cell_31235 ( .a(TIMEBOOST_net_9528), .b(g64945_db), .o(n_4381) );
in01s01 g64131_u0 ( .a(FE_OFN1046_n_16657), .o(g64131_sb) );
na02s01 g64131_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(g64131_sb), .o(g64131_da) );
na02s01 g64131_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__Q), .b(FE_OFN1046_n_16657), .o(g64131_db) );
na03s02 TIMEBOOST_cell_38577 ( .a(wishbone_slave_unit_pcim_sm_last_in), .b(n_4936), .c(n_7538), .o(TIMEBOOST_net_11527) );
in01s01 g64132_u0 ( .a(FE_OFN908_n_4734), .o(g64132_sb) );
na02s01 g64132_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_128), .b(g64132_sb), .o(g64132_da) );
na02s01 g64132_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__Q), .b(FE_OFN908_n_4734), .o(g64132_db) );
na02s01 g64132_u3 ( .a(g64132_da), .b(g64132_db), .o(n_4030) );
in01s01 g64133_u0 ( .a(FE_OFN1046_n_16657), .o(g64133_sb) );
na02s02 TIMEBOOST_cell_39996 ( .a(TIMEBOOST_net_12236), .b(g62481_sb), .o(n_6626) );
na02s01 g64133_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__Q), .b(FE_OFN1046_n_16657), .o(g64133_db) );
na02s02 TIMEBOOST_cell_39998 ( .a(TIMEBOOST_net_12237), .b(g62666_sb), .o(n_6206) );
in01s01 g64134_u0 ( .a(FE_OFN1049_n_16657), .o(g64134_sb) );
na02m02 TIMEBOOST_cell_40000 ( .a(TIMEBOOST_net_12238), .b(g62451_sb), .o(n_6695) );
na02s01 g64134_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__Q), .b(FE_OFN1049_n_16657), .o(g64134_db) );
na02s02 TIMEBOOST_cell_40002 ( .a(TIMEBOOST_net_12239), .b(g62425_sb), .o(n_6747) );
in01s01 g64135_u0 ( .a(FE_OFN906_n_4736), .o(g64135_sb) );
na02f02 TIMEBOOST_cell_44536 ( .a(TIMEBOOST_net_14506), .b(FE_OFN2188_n_8567), .o(TIMEBOOST_net_13459) );
na02s01 g64135_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__14__Q), .b(FE_OFN906_n_4736), .o(g64135_db) );
na02s01 TIMEBOOST_cell_32145 ( .a(TIMEBOOST_net_9983), .b(g62012_sb), .o(n_7871) );
in01s01 g64136_u0 ( .a(FE_OFN1076_n_4740), .o(g64136_sb) );
na02f08 TIMEBOOST_cell_36280 ( .a(TIMEBOOST_net_10378), .b(FE_RN_305_0), .o(TIMEBOOST_net_213) );
na02s01 TIMEBOOST_cell_18288 ( .a(g61923_sb), .b(g61968_db), .o(TIMEBOOST_net_4401) );
na02m08 TIMEBOOST_cell_36281 ( .a(n_3083), .b(TIMEBOOST_net_9297), .o(TIMEBOOST_net_10379) );
in01s01 g64137_u0 ( .a(FE_OFN1049_n_16657), .o(g64137_sb) );
na02s01 TIMEBOOST_cell_36507 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__Q), .b(FE_OFN205_n_9140), .o(TIMEBOOST_net_10492) );
na02s01 g64137_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__Q), .b(FE_OFN1049_n_16657), .o(g64137_db) );
na02s01 TIMEBOOST_cell_9903 ( .a(TIMEBOOST_net_1518), .b(FE_OFN235_n_9834), .o(n_9759) );
in01s01 g64138_u0 ( .a(FE_OFN904_n_4736), .o(g64138_sb) );
na02f02 TIMEBOOST_cell_44186 ( .a(TIMEBOOST_net_14331), .b(FE_OFN1399_n_8567), .o(TIMEBOOST_net_12767) );
na02s01 g64138_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__Q), .b(FE_OFN904_n_4736), .o(g64138_db) );
na02f02 TIMEBOOST_cell_38816 ( .a(TIMEBOOST_net_11646), .b(n_10256), .o(TIMEBOOST_net_10694) );
in01s01 g64139_u0 ( .a(FE_OFN905_n_4736), .o(g64139_sb) );
na02s01 g64139_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q), .b(FE_OFN905_n_4736), .o(g64139_db) );
na02s01 TIMEBOOST_cell_42642 ( .a(TIMEBOOST_net_13559), .b(g58172_db), .o(n_9062) );
in01s01 g64140_u0 ( .a(FE_OFN923_n_4740), .o(g64140_sb) );
na02f02 TIMEBOOST_cell_41686 ( .a(n_11898), .b(TIMEBOOST_net_13081), .o(n_12485) );
na02s01 g64140_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__Q), .b(FE_OFN923_n_4740), .o(g64140_db) );
na02s01 TIMEBOOST_cell_41929 ( .a(FE_OFN201_n_9230), .b(g57900_sb), .o(TIMEBOOST_net_13203) );
in01s01 g64141_u0 ( .a(FE_OFN906_n_4736), .o(g64141_sb) );
na02s01 g64141_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_145), .b(g64141_sb), .o(g64141_da) );
na02s01 g64141_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__Q), .b(FE_OFN906_n_4736), .o(g64141_db) );
na02s02 TIMEBOOST_cell_44973 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__Q), .b(FE_OFN207_n_9865), .o(TIMEBOOST_net_14725) );
in01s01 g64142_u0 ( .a(FE_OFN953_n_2055), .o(g64142_sb) );
na02m02 TIMEBOOST_cell_41798 ( .a(n_3351), .b(TIMEBOOST_net_13137), .o(TIMEBOOST_net_11686) );
na02s01 g64142_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__Q), .b(FE_OFN953_n_2055), .o(g64142_db) );
na02s01 TIMEBOOST_cell_42590 ( .a(TIMEBOOST_net_13533), .b(g57902_db), .o(n_9137) );
in01s01 g64143_u0 ( .a(FE_OFN908_n_4734), .o(g64143_sb) );
na02s01 g64143_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(g64143_sb), .o(g64143_da) );
na02s01 g64143_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__Q), .b(FE_OFN908_n_4734), .o(g64143_db) );
na02s01 g64143_u3 ( .a(g64143_da), .b(g64143_db), .o(n_4021) );
in01s01 g64144_u0 ( .a(FE_OFN1013_n_4734), .o(g64144_sb) );
na02s02 TIMEBOOST_cell_31234 ( .a(n_4447), .b(g64945_sb), .o(TIMEBOOST_net_9528) );
na02s01 g64144_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__Q), .b(FE_OFN1013_n_4734), .o(g64144_db) );
na02s01 TIMEBOOST_cell_31233 ( .a(TIMEBOOST_net_9527), .b(g64942_db), .o(n_3673) );
in01s01 g64145_u0 ( .a(FE_OFN2109_n_2047), .o(g64145_sb) );
na02s01 TIMEBOOST_cell_9078 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__Q), .o(TIMEBOOST_net_1106) );
na02s01 g64145_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__Q), .b(FE_OFN2109_n_2047), .o(g64145_db) );
na02s01 TIMEBOOST_cell_9079 ( .a(TIMEBOOST_net_1106), .b(n_4725), .o(TIMEBOOST_net_155) );
in01s01 g64146_u0 ( .a(FE_OFN1010_n_4734), .o(g64146_sb) );
na03s02 TIMEBOOST_cell_33981 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__Q), .b(FE_OFN881_g64577_p), .c(g62720_sb), .o(TIMEBOOST_net_9856) );
na02s01 g64146_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q), .b(FE_OFN1010_n_4734), .o(g64146_db) );
na02s01 TIMEBOOST_cell_36477 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(g65769_sb), .o(TIMEBOOST_net_10477) );
in01s01 g64147_u0 ( .a(FE_OFN906_n_4736), .o(g64147_sb) );
na02s01 g64147_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(g64147_sb), .o(g64147_da) );
na02s01 g64147_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__28__Q), .b(FE_OFN906_n_4736), .o(g64147_db) );
na02s01 TIMEBOOST_cell_44974 ( .a(TIMEBOOST_net_14725), .b(FE_OFN1801_n_9690), .o(TIMEBOOST_net_11016) );
in01s01 g64148_u0 ( .a(FE_OFN906_n_4736), .o(g64148_sb) );
na02s01 g64148_u1 ( .a(pci_target_unit_fifos_pciw_cbe_in_152), .b(g64148_sb), .o(g64148_da) );
na02s01 g64148_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__Q), .b(FE_OFN906_n_4736), .o(g64148_db) );
na02s02 TIMEBOOST_cell_45102 ( .a(TIMEBOOST_net_14789), .b(FE_OFN1812_n_7845), .o(TIMEBOOST_net_11382) );
in01s01 g64149_u0 ( .a(FE_OFN1074_n_4740), .o(g64149_sb) );
na02s02 TIMEBOOST_cell_43041 ( .a(TIMEBOOST_net_9870), .b(FE_OFN1671_n_9477), .o(TIMEBOOST_net_13759) );
na02s01 g64149_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__Q), .b(FE_OFN1074_n_4740), .o(g64149_db) );
na02s01 TIMEBOOST_cell_41930 ( .a(TIMEBOOST_net_13203), .b(g57900_db), .o(n_9225) );
in01s01 g64150_u0 ( .a(FE_OFN1011_n_4734), .o(g64150_sb) );
na02s01 TIMEBOOST_cell_31232 ( .a(n_3777), .b(g64942_sb), .o(TIMEBOOST_net_9527) );
na02s01 g64150_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__16__Q), .b(FE_OFN1011_n_4734), .o(g64150_db) );
na03f02 TIMEBOOST_cell_36117 ( .a(n_15591), .b(n_15593), .c(n_15586), .o(n_15594) );
in01s01 g64151_u0 ( .a(FE_OFN1011_n_4734), .o(g64151_sb) );
na02s01 TIMEBOOST_cell_43477 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__Q), .b(n_4477), .o(TIMEBOOST_net_13977) );
na02s01 g64151_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__13__Q), .b(FE_OFN1011_n_4734), .o(g64151_db) );
na02s01 TIMEBOOST_cell_16566 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(g65888_sb), .o(TIMEBOOST_net_3540) );
in01s01 g64152_u0 ( .a(FE_OFN1010_n_4734), .o(g64152_sb) );
na02s01 g64152_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_135), .b(g64152_sb), .o(g64152_da) );
na02s01 g64152_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q), .b(FE_OFN1010_n_4734), .o(g64152_db) );
na02s01 g64152_u3 ( .a(g64152_da), .b(g64152_db), .o(n_4013) );
in01s01 g64153_u0 ( .a(FE_OFN1013_n_4734), .o(g64153_sb) );
na02s02 TIMEBOOST_cell_45723 ( .a(n_4900), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q), .o(TIMEBOOST_net_15100) );
na02s01 g64153_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__Q), .b(FE_OFN1013_n_4734), .o(g64153_db) );
na02s02 TIMEBOOST_cell_45724 ( .a(TIMEBOOST_net_15100), .b(FE_OFN1274_n_4096), .o(TIMEBOOST_net_12612) );
in01s01 g64154_u0 ( .a(FE_OFN1010_n_4734), .o(g64154_sb) );
na02s01 TIMEBOOST_cell_17838 ( .a(n_3785), .b(g64763_sb), .o(TIMEBOOST_net_4176) );
na02s01 g64154_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__14__Q), .b(FE_OFN1010_n_4734), .o(g64154_db) );
na02s02 TIMEBOOST_cell_38453 ( .a(TIMEBOOST_net_9853), .b(FE_OFN1084_n_13221), .o(TIMEBOOST_net_11465) );
in01s01 g64155_u0 ( .a(FE_OFN1010_n_4734), .o(g64155_sb) );
na02s02 TIMEBOOST_cell_45725 ( .a(n_3634), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__Q), .o(TIMEBOOST_net_15101) );
na02s01 g64155_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q), .b(FE_OFN1010_n_4734), .o(g64155_db) );
na03f02 TIMEBOOST_cell_36082 ( .a(n_11900), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__Q), .c(FE_OFN1747_n_12004), .o(n_12622) );
in01s01 g64156_u0 ( .a(FE_OFN1012_n_4734), .o(g64156_sb) );
na02s02 TIMEBOOST_cell_45726 ( .a(TIMEBOOST_net_15101), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_13263) );
na02s01 g64156_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__Q), .b(FE_OFN1012_n_4734), .o(g64156_db) );
na02s01 TIMEBOOST_cell_45733 ( .a(n_3633), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__Q), .o(TIMEBOOST_net_15105) );
in01s01 g64157_u0 ( .a(FE_OFN1075_n_4740), .o(g64157_sb) );
na02m02 TIMEBOOST_cell_42153 ( .a(n_9837), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__Q), .o(TIMEBOOST_net_13315) );
na02s01 g64157_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__Q), .b(FE_OFN1075_n_4740), .o(g64157_db) );
na02s01 TIMEBOOST_cell_42908 ( .a(TIMEBOOST_net_13692), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_11158) );
in01s01 g64158_u0 ( .a(FE_OFN1011_n_4734), .o(g64158_sb) );
na02s01 g64158_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_132), .b(g64158_sb), .o(g64158_da) );
na02s01 g64158_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q), .b(FE_OFN1011_n_4734), .o(g64158_db) );
na02s01 g64158_u3 ( .a(g64158_da), .b(g64158_db), .o(n_4007) );
in01s01 g64159_u0 ( .a(FE_OFN1013_n_4734), .o(g64159_sb) );
na02s01 g64159_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__Q), .b(FE_OFN1013_n_4734), .o(g64159_db) );
na03f02 TIMEBOOST_cell_36086 ( .a(n_12041), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__Q), .c(n_12313), .o(n_12748) );
in01s01 g64160_u0 ( .a(FE_OFN1010_n_4734), .o(g64160_sb) );
na02s02 TIMEBOOST_cell_17840 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__Q), .b(g65906_sb), .o(TIMEBOOST_net_4177) );
na02s01 g64160_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__Q), .b(FE_OFN1010_n_4734), .o(g64160_db) );
na02s02 TIMEBOOST_cell_17841 ( .a(TIMEBOOST_net_4177), .b(g65906_db), .o(n_1856) );
in01s01 g64161_u0 ( .a(FE_OFN1011_n_4734), .o(g64161_sb) );
na02s01 TIMEBOOST_cell_16567 ( .a(TIMEBOOST_net_3540), .b(g65888_db), .o(n_1861) );
na02s01 g64161_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__Q), .b(FE_OFN1011_n_4734), .o(g64161_db) );
na02s01 TIMEBOOST_cell_42933 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__Q), .b(FE_OFN535_n_9823), .o(TIMEBOOST_net_13705) );
in01s01 g64162_u0 ( .a(FE_OFN908_n_4734), .o(g64162_sb) );
na02s01 TIMEBOOST_cell_31220 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__Q), .o(TIMEBOOST_net_9521) );
na02s01 g64162_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q), .b(FE_OFN908_n_4734), .o(g64162_db) );
na02s01 TIMEBOOST_cell_31219 ( .a(TIMEBOOST_net_9520), .b(g65289_db), .o(n_3579) );
in01s01 g64163_u0 ( .a(FE_OFN1011_n_4734), .o(g64163_sb) );
na02s01 TIMEBOOST_cell_31218 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__Q), .b(g65289_sb), .o(TIMEBOOST_net_9520) );
na02s01 g64163_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__Q), .b(FE_OFN1011_n_4734), .o(g64163_db) );
na02s01 TIMEBOOST_cell_45718 ( .a(TIMEBOOST_net_15097), .b(g62572_sb), .o(n_6410) );
in01s01 g64164_u0 ( .a(FE_OFN1010_n_4734), .o(g64164_sb) );
na02s01 g64164_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(g64164_sb), .o(g64164_da) );
na02s01 g64164_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__Q), .b(FE_OFN1010_n_4734), .o(g64164_db) );
na02s02 TIMEBOOST_cell_36640 ( .a(TIMEBOOST_net_10558), .b(g52641_db), .o(n_14749) );
in01s01 g64165_u0 ( .a(FE_OFN1074_n_4740), .o(g64165_sb) );
na02f02 TIMEBOOST_cell_42154 ( .a(TIMEBOOST_net_13315), .b(FE_OFN1419_n_8567), .o(TIMEBOOST_net_12280) );
na02s01 g64165_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__Q), .b(FE_OFN1074_n_4740), .o(g64165_db) );
na02s01 TIMEBOOST_cell_41893 ( .a(g64352_da), .b(g64352_db), .o(TIMEBOOST_net_13185) );
in01s01 g64166_u0 ( .a(FE_OFN1013_n_4734), .o(g64166_sb) );
na03f02 TIMEBOOST_cell_35932 ( .a(TIMEBOOST_net_10092), .b(g58600_sb), .c(g58600_db), .o(n_9239) );
na02s01 g64166_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q), .b(FE_OFN1013_n_4734), .o(g64166_db) );
na03f02 TIMEBOOST_cell_35935 ( .a(TIMEBOOST_net_10096), .b(FE_OFN1472_g52675_p), .c(g52509_sb), .o(n_13744) );
in01s01 g64167_u0 ( .a(FE_OFN905_n_4736), .o(g64167_sb) );
na02s01 g64167_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_139), .b(g64167_sb), .o(g64167_da) );
na02s01 g64167_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__Q), .b(FE_OFN905_n_4736), .o(g64167_db) );
na02s02 TIMEBOOST_cell_45161 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__Q), .b(n_3523), .o(TIMEBOOST_net_14819) );
in01s01 g64168_u0 ( .a(FE_OFN1012_n_4734), .o(g64168_sb) );
na03f02 TIMEBOOST_cell_35934 ( .a(TIMEBOOST_net_10097), .b(FE_OFN1472_g52675_p), .c(g52528_sb), .o(n_13693) );
na02s01 g64168_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__Q), .b(FE_OFN1012_n_4734), .o(g64168_db) );
in01s01 g64169_u0 ( .a(FE_OFN906_n_4736), .o(g64169_sb) );
na02s01 g64169_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_146), .b(g64169_sb), .o(g64169_da) );
na02s01 g64169_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__Q), .b(FE_OFN906_n_4736), .o(g64169_db) );
na02s02 TIMEBOOST_cell_43542 ( .a(TIMEBOOST_net_14009), .b(FE_OFN1316_n_6624), .o(TIMEBOOST_net_12676) );
in01s01 g64170_u0 ( .a(FE_OFN923_n_4740), .o(g64170_sb) );
na02s01 TIMEBOOST_cell_39273 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__16__Q), .b(g64275_sb), .o(TIMEBOOST_net_11875) );
na02s01 g64170_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__Q), .b(FE_OFN923_n_4740), .o(g64170_db) );
na02s01 TIMEBOOST_cell_39274 ( .a(TIMEBOOST_net_11875), .b(g64275_db), .o(n_3898) );
in01s01 g64171_u0 ( .a(FE_OFN1010_n_4734), .o(g64171_sb) );
na02m02 TIMEBOOST_cell_40004 ( .a(TIMEBOOST_net_12240), .b(g63160_sb), .o(n_5816) );
na02s01 g64171_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__Q), .b(FE_OFN1010_n_4734), .o(g64171_db) );
na02s01 TIMEBOOST_cell_37576 ( .a(TIMEBOOST_net_11026), .b(g65927_db), .o(n_2584) );
in01s01 g64172_u0 ( .a(FE_OFN904_n_4736), .o(g64172_sb) );
na02m02 TIMEBOOST_cell_38817 ( .a(n_1680), .b(wbu_addr_in_253), .o(TIMEBOOST_net_11647) );
na02s01 g64172_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__Q), .b(FE_OFN904_n_4736), .o(g64172_db) );
na02f02 TIMEBOOST_cell_38818 ( .a(TIMEBOOST_net_11647), .b(n_10256), .o(TIMEBOOST_net_10696) );
in01s01 g64173_u0 ( .a(FE_OFN1050_n_16657), .o(g64173_sb) );
na02f02 TIMEBOOST_cell_39101 ( .a(FE_RN_221_0), .b(n_10656), .o(TIMEBOOST_net_11789) );
na02s01 g64173_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__Q), .b(FE_OFN1050_n_16657), .o(g64173_db) );
na02f04 TIMEBOOST_cell_39030 ( .a(TIMEBOOST_net_11753), .b(FE_OFN2241_g52675_p), .o(TIMEBOOST_net_10748) );
oa12s01 g64174_u0 ( .a(n_1803), .b(FE_OFN1012_n_4734), .c(pci_target_unit_fifos_pciw_control_in), .o(n_4521) );
in01s01 g64175_u0 ( .a(FE_OFN1013_n_4734), .o(g64175_sb) );
na02s01 g64175_u1 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(g64175_sb), .o(g64175_da) );
na02s01 g64175_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__Q), .b(FE_OFN1013_n_4734), .o(g64175_db) );
na02m04 TIMEBOOST_cell_39031 ( .a(wbs_wbb3_2_wbb2_dat_o_i_117), .b(wbs_dat_o_18_), .o(TIMEBOOST_net_11754) );
in01s01 g64176_u0 ( .a(FE_OFN1012_n_4734), .o(g64176_sb) );
na02s01 g64176_u1 ( .a(pci_target_unit_fifos_pciw_cbe_in_153), .b(g64176_sb), .o(g64176_da) );
na02s01 g64176_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__Q), .b(FE_OFN1012_n_4734), .o(g64176_db) );
na02f02 TIMEBOOST_cell_39487 ( .a(n_3238), .b(n_2768), .o(TIMEBOOST_net_11982) );
in01s01 g64177_u0 ( .a(FE_OFN906_n_4736), .o(g64177_sb) );
na02s01 g64177_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_143), .b(g64177_sb), .o(g64177_da) );
na02s01 g64177_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__Q), .b(FE_OFN906_n_4736), .o(g64177_db) );
na02s02 TIMEBOOST_cell_44975 ( .a(FE_OFN213_n_9124), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__Q), .o(TIMEBOOST_net_14726) );
in01s01 g64178_u0 ( .a(FE_OFN908_n_4734), .o(g64178_sb) );
na02s01 TIMEBOOST_cell_45717 ( .a(TIMEBOOST_net_4811), .b(FE_OFN1200_n_4090), .o(TIMEBOOST_net_15097) );
na02s01 g64178_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__Q), .b(FE_OFN908_n_4734), .o(g64178_db) );
na03f03 TIMEBOOST_cell_36005 ( .a(n_16967), .b(n_16970), .c(n_16974), .o(n_13674) );
in01s01 g64179_u0 ( .a(FE_OFN1049_n_16657), .o(g64179_sb) );
na02s01 TIMEBOOST_cell_9906 ( .a(FE_OFN211_n_9858), .b(FE_OFN572_n_9502), .o(TIMEBOOST_net_1520) );
na02s01 g64179_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__Q), .b(FE_OFN1049_n_16657), .o(g64179_db) );
na02s01 TIMEBOOST_cell_9907 ( .a(TIMEBOOST_net_1520), .b(g58311_da), .o(n_9500) );
in01s01 g64180_u0 ( .a(FE_OFN1011_n_4734), .o(g64180_sb) );
na02s01 g64180_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__Q), .b(FE_OFN1011_n_4734), .o(g64180_db) );
na02s01 TIMEBOOST_cell_44784 ( .a(TIMEBOOST_net_14630), .b(g58083_sb), .o(TIMEBOOST_net_13162) );
in01s01 g64181_u0 ( .a(FE_OFN908_n_4734), .o(g64181_sb) );
na02s01 TIMEBOOST_cell_42893 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__Q), .b(FE_OFN593_n_9694), .o(TIMEBOOST_net_13685) );
na02s01 g64181_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__Q), .b(FE_OFN908_n_4734), .o(g64181_db) );
na02s01 TIMEBOOST_cell_31208 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__Q), .b(pci_target_unit_fifos_pcir_data_in_182), .o(TIMEBOOST_net_9515) );
in01s01 g64182_u0 ( .a(FE_OFN1011_n_4734), .o(g64182_sb) );
na02s01 g64182_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_142), .b(g64182_sb), .o(g64182_da) );
na02s01 g64182_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__Q), .b(FE_OFN1011_n_4734), .o(g64182_db) );
na02s01 g64182_u3 ( .a(g64182_da), .b(g64182_db), .o(n_3984) );
in01s01 g64183_u0 ( .a(FE_OFN1049_n_16657), .o(g64183_sb) );
na02s01 TIMEBOOST_cell_45067 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__Q), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_14772) );
na02s01 g64183_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q), .b(FE_OFN1049_n_16657), .o(g64183_db) );
na02s01 TIMEBOOST_cell_38690 ( .a(TIMEBOOST_net_11583), .b(g62808_db), .o(n_5363) );
in01s01 g64184_u0 ( .a(FE_OFN1011_n_4734), .o(g64184_sb) );
na03f04 TIMEBOOST_cell_36009 ( .a(FE_OCP_RBN2016_n_16970), .b(n_14939), .c(n_16205), .o(n_13701) );
na02s01 g64184_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN1011_n_4734), .o(g64184_db) );
na02s02 TIMEBOOST_cell_41867 ( .a(TIMEBOOST_net_327), .b(g61894_sb), .o(TIMEBOOST_net_13172) );
in01s01 g64185_u0 ( .a(FE_OFN908_n_4734), .o(g64185_sb) );
na02s01 g64185_u1 ( .a(pci_target_unit_fifos_pciw_cbe_in_152), .b(g64185_sb), .o(g64185_da) );
na02s01 g64185_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__Q), .b(FE_OFN908_n_4734), .o(g64185_db) );
na02s01 g64185_u3 ( .a(g64185_da), .b(g64185_db), .o(n_3981) );
in01s01 g64186_u0 ( .a(FE_OFN1013_n_4734), .o(g64186_sb) );
na03f02 TIMEBOOST_cell_36010 ( .a(n_10904), .b(FE_RN_477_0), .c(n_12569), .o(n_12831) );
na02s01 g64186_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q), .b(FE_OFN1013_n_4734), .o(g64186_db) );
na02s01 TIMEBOOST_cell_31204 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__Q), .b(pci_target_unit_fifos_pcir_data_in_174), .o(TIMEBOOST_net_9513) );
in01s01 g64187_u0 ( .a(FE_OFN1051_n_16657), .o(g64187_sb) );
na02s02 TIMEBOOST_cell_43377 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__Q), .b(n_4255), .o(TIMEBOOST_net_13927) );
na02s01 TIMEBOOST_cell_9080 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__Q), .o(TIMEBOOST_net_1107) );
na02m02 TIMEBOOST_cell_40006 ( .a(TIMEBOOST_net_12241), .b(g62636_sb), .o(n_6278) );
in01s01 g64188_u0 ( .a(FE_OFN906_n_4736), .o(g64188_sb) );
na02s01 g64188_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(g64188_sb), .o(g64188_da) );
na02s01 g64188_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__Q), .b(FE_OFN906_n_4736), .o(g64188_db) );
na02s02 TIMEBOOST_cell_45162 ( .a(TIMEBOOST_net_14819), .b(FE_OFN1204_n_4090), .o(TIMEBOOST_net_12597) );
in01s01 g64189_u0 ( .a(FE_OFN905_n_4736), .o(g64189_sb) );
na02s01 g64189_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(g64189_sb), .o(g64189_da) );
na02s01 g64189_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__Q), .b(FE_OFN905_n_4736), .o(g64189_db) );
na02s01 TIMEBOOST_cell_45068 ( .a(TIMEBOOST_net_14772), .b(FE_OFN587_n_9692), .o(TIMEBOOST_net_11174) );
in01s01 g64190_u0 ( .a(FE_OFN1785_n_1699), .o(g64190_sb) );
na02s01 g64190_u1 ( .a(pci_target_unit_fifos_pcir_control_in_192), .b(g64190_sb), .o(g64190_da) );
na02s01 g64190_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__Q), .b(FE_OFN1785_n_1699), .o(g64190_db) );
na02s01 g64190_u3 ( .a(g64190_da), .b(g64190_db), .o(n_4520) );
in01s01 g64191_u0 ( .a(FE_OFN905_n_4736), .o(g64191_sb) );
na02s01 g64191_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_132), .b(g64191_sb), .o(g64191_da) );
na02s01 g64191_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q), .b(FE_OFN905_n_4736), .o(g64191_db) );
na02m04 TIMEBOOST_cell_40223 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__Q), .o(TIMEBOOST_net_12350) );
in01s01 g64192_u0 ( .a(FE_OFN1051_n_16657), .o(g64192_sb) );
na02s01 g64192_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(g64192_sb), .o(g64192_da) );
na02s01 g64192_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__Q), .b(FE_OFN1051_n_16657), .o(g64192_db) );
na02s02 TIMEBOOST_cell_43627 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__Q), .b(n_4483), .o(TIMEBOOST_net_14052) );
in01s01 g64193_u0 ( .a(FE_OFN1051_n_16657), .o(g64193_sb) );
na02s01 g64193_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_135), .b(g64193_sb), .o(g64193_da) );
na02s01 g64193_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__15__Q), .b(FE_OFN1051_n_16657), .o(g64193_db) );
na02s02 TIMEBOOST_cell_43628 ( .a(TIMEBOOST_net_14052), .b(FE_OFN1311_n_6624), .o(TIMEBOOST_net_12239) );
no02s01 g64194_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_3_), .b(n_1437), .o(g64194_p) );
ao12s01 g64194_u1 ( .a(g64194_p), .b(pci_target_unit_wishbone_master_rty_counter_3_), .c(n_1437), .o(n_1662) );
in01s01 g64195_u0 ( .a(FE_OFN1051_n_16657), .o(g64195_sb) );
na02m06 TIMEBOOST_cell_17928 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_395), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__Q), .o(TIMEBOOST_net_4221) );
na02s01 g64195_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__16__Q), .b(FE_OFN1051_n_16657), .o(g64195_db) );
na02s01 TIMEBOOST_cell_45069 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__Q), .b(FE_OFN553_n_9864), .o(TIMEBOOST_net_14773) );
in01s01 g64196_u0 ( .a(FE_OFN903_n_4736), .o(g64196_sb) );
na02s01 g64196_u1 ( .a(pci_target_unit_fifos_pciw_cbe_in_153), .b(g64196_sb), .o(g64196_da) );
na02s01 g64196_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__Q), .b(FE_OFN903_n_4736), .o(g64196_db) );
na02s01 TIMEBOOST_cell_45070 ( .a(TIMEBOOST_net_14773), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_11175) );
in01s01 g64197_u0 ( .a(FE_OFN906_n_4736), .o(g64197_sb) );
na02f02 TIMEBOOST_cell_32143 ( .a(TIMEBOOST_net_9982), .b(n_3456), .o(n_14812) );
na02s01 g64197_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__Q), .b(FE_OFN906_n_4736), .o(g64197_db) );
na02f02 TIMEBOOST_cell_32142 ( .a(g52440_sb), .b(g52440_db), .o(TIMEBOOST_net_9982) );
in01s01 g64198_u0 ( .a(FE_OFN1011_n_4734), .o(g64198_sb) );
na02s01 TIMEBOOST_cell_41896 ( .a(TIMEBOOST_net_13186), .b(g62127_sb), .o(TIMEBOOST_net_11976) );
na02s01 g64198_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__Q), .b(FE_OFN1011_n_4734), .o(g64198_db) );
na02s01 TIMEBOOST_cell_31202 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__Q), .b(pci_target_unit_fifos_pcir_data_in_173), .o(TIMEBOOST_net_9512) );
in01s01 g64199_u0 ( .a(FE_OFN906_n_4736), .o(g64199_sb) );
na02m02 TIMEBOOST_cell_15912 ( .a(n_1724), .b(pci_target_unit_pci_target_sm_rd_from_fifo), .o(TIMEBOOST_net_3213) );
na02s01 g64199_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__Q), .b(FE_OFN906_n_4736), .o(g64199_db) );
na03s02 TIMEBOOST_cell_38077 ( .a(TIMEBOOST_net_4242), .b(g64214_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q), .o(TIMEBOOST_net_11277) );
in01s01 g64200_u0 ( .a(FE_OFN1051_n_16657), .o(g64200_sb) );
na02s01 g64200_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(g64200_sb), .o(g64200_da) );
na02s01 g64200_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q), .b(FE_OFN1051_n_16657), .o(g64200_db) );
na02s02 TIMEBOOST_cell_40008 ( .a(TIMEBOOST_net_12242), .b(g62401_sb), .o(n_6797) );
in01s01 g64201_u0 ( .a(FE_OFN906_n_4736), .o(g64201_sb) );
na02s01 g64201_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_128), .b(g64201_sb), .o(g64201_da) );
na02s01 g64201_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__Q), .b(FE_OFN906_n_4736), .o(g64201_db) );
na02s02 TIMEBOOST_cell_44976 ( .a(TIMEBOOST_net_14726), .b(FE_OFN1634_n_9531), .o(TIMEBOOST_net_11015) );
in01s01 g64202_u0 ( .a(FE_OFN905_n_4736), .o(g64202_sb) );
na02m02 TIMEBOOST_cell_32140 ( .a(FE_OFN1189_n_5742), .b(wishbone_slave_unit_wishbone_slave_del_addr_hit), .o(TIMEBOOST_net_9981) );
na02s01 g64202_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__Q), .b(FE_OFN905_n_4736), .o(g64202_db) );
na02s02 TIMEBOOST_cell_43601 ( .a(n_4292), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__Q), .o(TIMEBOOST_net_14039) );
in01s01 g64203_u0 ( .a(FE_OFN906_n_4736), .o(g64203_sb) );
na02s01 g64203_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_127), .b(g64203_sb), .o(g64203_da) );
na02s01 g64203_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__Q), .b(FE_OFN906_n_4736), .o(g64203_db) );
na02f02 TIMEBOOST_cell_44706 ( .a(TIMEBOOST_net_14591), .b(TIMEBOOST_net_6359), .o(n_14284) );
in01s01 g64204_u0 ( .a(FE_OFN1051_n_16657), .o(g64204_sb) );
na02s01 TIMEBOOST_cell_38691 ( .a(n_3982), .b(g62835_sb), .o(TIMEBOOST_net_11584) );
na02s01 g64204_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__Q), .b(FE_OFN1051_n_16657), .o(g64204_db) );
na02s01 TIMEBOOST_cell_38692 ( .a(TIMEBOOST_net_11584), .b(g62835_db), .o(n_5303) );
in01s01 g64205_u0 ( .a(FE_OFN1075_n_4740), .o(g64205_sb) );
na02m04 TIMEBOOST_cell_39029 ( .a(wbs_wbb3_2_wbb2_dat_o_i_122), .b(wbs_dat_o_23_), .o(TIMEBOOST_net_11753) );
na02s01 g64205_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__Q), .b(FE_OFN1075_n_4740), .o(g64205_db) );
na02m02 TIMEBOOST_cell_38484 ( .a(TIMEBOOST_net_11480), .b(n_3305), .o(TIMEBOOST_net_5429) );
in01s01 g64206_u0 ( .a(FE_OFN1049_n_16657), .o(g64206_sb) );
na02s01 g64206_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(g64206_sb), .o(g64206_da) );
na02s01 g64206_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__Q), .b(FE_OFN1049_n_16657), .o(g64206_db) );
na02f02 TIMEBOOST_cell_38570 ( .a(TIMEBOOST_net_11523), .b(n_3039), .o(TIMEBOOST_net_637) );
in01s01 g64207_u0 ( .a(FE_OFN905_n_4736), .o(g64207_sb) );
na02s01 g64207_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_136), .b(g64207_sb), .o(g64207_da) );
na02s01 g64207_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__16__Q), .b(FE_OFN905_n_4736), .o(g64207_db) );
na02s02 TIMEBOOST_cell_45163 ( .a(n_263), .b(n_4902), .o(TIMEBOOST_net_14820) );
in01s01 g64208_u0 ( .a(FE_OFN1049_n_16657), .o(g64208_sb) );
na02s01 TIMEBOOST_cell_9914 ( .a(n_4084), .b(FE_OFN2121_n_2687), .o(TIMEBOOST_net_1524) );
na02s01 g64208_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__Q), .b(FE_OFN1049_n_16657), .o(g64208_db) );
na02s01 TIMEBOOST_cell_9915 ( .a(TIMEBOOST_net_1524), .b(FE_OFN2052_n_6965), .o(TIMEBOOST_net_808) );
in01s01 g64209_u0 ( .a(FE_OFN1075_n_4740), .o(g64209_sb) );
na02s01 TIMEBOOST_cell_38485 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_0__Q), .b(FE_OFN1082_n_13221), .o(TIMEBOOST_net_11481) );
na02s01 g64209_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__Q), .b(FE_OFN1075_n_4740), .o(g64209_db) );
na02s02 TIMEBOOST_cell_38486 ( .a(TIMEBOOST_net_11481), .b(TIMEBOOST_net_9875), .o(n_13497) );
in01s01 g64210_u0 ( .a(FE_OFN1051_n_16657), .o(g64210_sb) );
na02s01 g64210_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_143), .b(g64210_sb), .o(g64210_da) );
na02s01 g64210_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__Q), .b(FE_OFN1051_n_16657), .o(g64210_db) );
na02m02 TIMEBOOST_cell_43629 ( .a(n_4337), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__Q), .o(TIMEBOOST_net_14053) );
in01s01 g64211_u0 ( .a(FE_OFN1077_n_4740), .o(g64211_sb) );
na02f02 TIMEBOOST_cell_44394 ( .a(TIMEBOOST_net_14435), .b(FE_OFN1414_n_8567), .o(TIMEBOOST_net_12781) );
na02s01 g64211_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q), .b(FE_OFN1077_n_4740), .o(g64211_db) );
na02m02 TIMEBOOST_cell_44537 ( .a(n_9588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__Q), .o(TIMEBOOST_net_14507) );
in01s01 g64212_u0 ( .a(FE_OFN923_n_4740), .o(g64212_sb) );
na02m02 TIMEBOOST_cell_44127 ( .a(n_9568), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__Q), .o(TIMEBOOST_net_14302) );
na02s01 g64212_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__28__Q), .b(FE_OFN923_n_4740), .o(g64212_db) );
na02s02 TIMEBOOST_cell_38488 ( .a(TIMEBOOST_net_11482), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_10663) );
in01s01 g64213_u0 ( .a(FE_OFN1051_n_16657), .o(g64213_sb) );
na02m02 TIMEBOOST_cell_9916 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_27__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_792), .o(TIMEBOOST_net_1525) );
na02s01 g64213_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__Q), .b(FE_OFN1051_n_16657), .o(g64213_db) );
na02f02 TIMEBOOST_cell_9917 ( .a(TIMEBOOST_net_1525), .b(FE_OFN2127_n_16497), .o(TIMEBOOST_net_528) );
in01s01 g64214_u0 ( .a(FE_OFN1076_n_4740), .o(g64214_sb) );
na02s01 TIMEBOOST_cell_38489 ( .a(configuration_pci_err_data_527), .b(wbm_dat_o_26_), .o(TIMEBOOST_net_11483) );
na02s01 g64214_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q), .b(FE_OFN1076_n_4740), .o(g64214_db) );
na02s02 TIMEBOOST_cell_38490 ( .a(TIMEBOOST_net_11483), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_10664) );
in01s01 g64215_u0 ( .a(FE_OFN1050_n_16657), .o(g64215_sb) );
na02m02 TIMEBOOST_cell_9918 ( .a(n_7822), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_7__Q), .o(TIMEBOOST_net_1526) );
na02s01 g64215_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__Q), .b(FE_OFN1050_n_16657), .o(g64215_db) );
na02f02 TIMEBOOST_cell_9919 ( .a(TIMEBOOST_net_1526), .b(FE_OFN2127_n_16497), .o(TIMEBOOST_net_467) );
in01s01 g64216_u0 ( .a(FE_OFN905_n_4736), .o(g64216_sb) );
na02s02 TIMEBOOST_cell_38492 ( .a(TIMEBOOST_net_11484), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_10665) );
na02s01 g64216_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__Q), .b(FE_OFN905_n_4736), .o(g64216_db) );
na02s01 TIMEBOOST_cell_32137 ( .a(TIMEBOOST_net_9979), .b(g62515_sb), .o(TIMEBOOST_net_5279) );
in01s01 g64217_u0 ( .a(FE_OFN1051_n_16657), .o(g64217_sb) );
na02s02 TIMEBOOST_cell_9920 ( .a(conf_wb_err_addr_in_953), .b(FE_OFN2071_n_15978), .o(TIMEBOOST_net_1527) );
na02s01 g64217_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q), .b(FE_OFN1051_n_16657), .o(g64217_db) );
na02s02 TIMEBOOST_cell_9921 ( .a(TIMEBOOST_net_1527), .b(FE_OFN1143_n_15261), .o(TIMEBOOST_net_607) );
in01s01 g64218_u0 ( .a(FE_OFN1077_n_4740), .o(g64218_sb) );
na02s02 TIMEBOOST_cell_43473 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__23__Q), .b(n_3742), .o(TIMEBOOST_net_13975) );
na02s01 g64218_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__Q), .b(FE_OFN1077_n_4740), .o(g64218_db) );
na02s02 TIMEBOOST_cell_38494 ( .a(TIMEBOOST_net_11485), .b(g59122_sb), .o(n_8585) );
in01s01 g64219_u0 ( .a(FE_OFN903_n_4736), .o(g64219_sb) );
na02s01 g64219_u1 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(g64219_sb), .o(g64219_da) );
na02s01 g64219_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__Q), .b(FE_OFN903_n_4736), .o(g64219_db) );
na02s01 TIMEBOOST_cell_45071 ( .a(FE_OFN270_n_9836), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__Q), .o(TIMEBOOST_net_14774) );
in01s01 g64220_u0 ( .a(FE_OFN1076_n_4740), .o(g64220_sb) );
na02s01 TIMEBOOST_cell_38491 ( .a(configuration_pci_err_data_508), .b(wbm_dat_o_7_), .o(TIMEBOOST_net_11484) );
na02s01 g64220_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__14__Q), .b(FE_OFN1076_n_4740), .o(g64220_db) );
na02s01 TIMEBOOST_cell_38496 ( .a(TIMEBOOST_net_11486), .b(FE_OFN1219_n_6886), .o(TIMEBOOST_net_5193) );
in01s01 g64221_u0 ( .a(FE_OFN1076_n_4740), .o(g64221_sb) );
na02f04 TIMEBOOST_cell_39032 ( .a(TIMEBOOST_net_11754), .b(FE_OFN2243_g52675_p), .o(TIMEBOOST_net_10745) );
na02s01 g64221_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__Q), .b(FE_OFN1076_n_4740), .o(g64221_db) );
na02s01 TIMEBOOST_cell_18599 ( .a(TIMEBOOST_net_4556), .b(g62797_sb), .o(n_5391) );
in01s01 g64222_u0 ( .a(FE_OFN1074_n_4740), .o(g64222_sb) );
na03s02 TIMEBOOST_cell_38495 ( .a(TIMEBOOST_net_4184), .b(g65352_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__1__Q), .o(TIMEBOOST_net_11486) );
na02s01 g64222_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__Q), .b(FE_OFN1074_n_4740), .o(g64222_db) );
na02s02 TIMEBOOST_cell_39342 ( .a(TIMEBOOST_net_11909), .b(g65949_sb), .o(n_1562) );
in01s01 g64223_u0 ( .a(FE_OFN1051_n_16657), .o(g64223_sb) );
na02s02 TIMEBOOST_cell_9922 ( .a(conf_wb_err_addr_in_952), .b(FE_OFN2069_n_15978), .o(TIMEBOOST_net_1528) );
na02s01 g64223_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__Q), .b(FE_OFN1051_n_16657), .o(g64223_db) );
na02s02 TIMEBOOST_cell_9923 ( .a(TIMEBOOST_net_1528), .b(FE_OFN1142_n_15261), .o(TIMEBOOST_net_890) );
in01s01 g64224_u0 ( .a(FE_OFN1016_n_2053), .o(g64224_sb) );
na02s01 TIMEBOOST_cell_40269 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__Q), .b(n_8069), .o(TIMEBOOST_net_12373) );
na02s01 g64224_u2 ( .a(pci_target_unit_fifos_pcir_control_in_192), .b(FE_OFN1016_n_2053), .o(g64224_db) );
na02s01 TIMEBOOST_cell_16906 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__Q), .b(g65855_sb), .o(TIMEBOOST_net_3710) );
in01s01 g64225_u0 ( .a(FE_OFN2111_n_2248), .o(g64225_sb) );
na02s01 g64225_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__Q), .b(g64225_sb), .o(g64225_da) );
na02s01 g64225_u2 ( .a(pci_target_unit_fifos_pcir_control_in_192), .b(FE_OFN2111_n_2248), .o(g64225_db) );
na02s01 TIMEBOOST_cell_39559 ( .a(n_7078), .b(wishbone_slave_unit_pci_initiator_if_read_count_0_), .o(TIMEBOOST_net_12018) );
in01s01 g64226_u0 ( .a(FE_OFN1042_n_2037), .o(g64226_sb) );
na02s01 g64226_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__Q), .b(g64226_sb), .o(g64226_da) );
na02s01 g64226_u2 ( .a(pci_target_unit_fifos_pcir_control_in_192), .b(FE_OFN1042_n_2037), .o(g64226_db) );
na02f02 TIMEBOOST_cell_37072 ( .a(TIMEBOOST_net_10774), .b(FE_OFN1589_n_13736), .o(n_16259) );
in01s01 g64227_u0 ( .a(FE_OFN918_n_4725), .o(g64227_sb) );
na02s01 TIMEBOOST_cell_16263 ( .a(TIMEBOOST_net_3388), .b(g65668_db), .o(n_1960) );
na02s01 g64227_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_145), .b(FE_OFN918_n_4725), .o(g64227_db) );
na02m02 TIMEBOOST_cell_40535 ( .a(FE_OFN1084_n_13221), .b(TIMEBOOST_net_1837), .o(TIMEBOOST_net_12506) );
in01s01 g64228_u0 ( .a(FE_OFN912_n_4727), .o(g64228_sb) );
na02m04 TIMEBOOST_cell_39027 ( .a(wbs_wbb3_2_wbb2_dat_o_i_124), .b(wbs_dat_o_25_), .o(TIMEBOOST_net_11752) );
na02s01 g64228_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_130), .b(FE_OFN912_n_4727), .o(g64228_db) );
na02s02 TIMEBOOST_cell_38498 ( .a(TIMEBOOST_net_11487), .b(g58352_db), .o(n_9469) );
in01s01 g64229_u0 ( .a(FE_OFN1056_n_4727), .o(g64229_sb) );
na03s02 TIMEBOOST_cell_38499 ( .a(TIMEBOOST_net_9645), .b(g64760_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__Q), .o(TIMEBOOST_net_11488) );
na02s01 g64229_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_132), .b(FE_OFN1056_n_4727), .o(g64229_db) );
na02s02 TIMEBOOST_cell_38500 ( .a(TIMEBOOST_net_11488), .b(FE_OFN1258_n_4143), .o(TIMEBOOST_net_5235) );
in01s01 g64230_u0 ( .a(FE_OFN1056_n_4727), .o(g64230_sb) );
na02s02 TIMEBOOST_cell_38501 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__Q), .b(g58289_sb), .o(TIMEBOOST_net_11489) );
na02s01 g64230_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(FE_OFN1056_n_4727), .o(g64230_db) );
na02s01 TIMEBOOST_cell_39190 ( .a(TIMEBOOST_net_11833), .b(n_2159), .o(TIMEBOOST_net_11232) );
in01s01 g64231_u0 ( .a(FE_OFN1035_n_4732), .o(g64231_sb) );
na02s02 TIMEBOOST_cell_17930 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__Q), .b(n_504), .o(TIMEBOOST_net_4222) );
na02s01 g64231_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_145), .b(FE_OFN1031_n_4732), .o(g64231_db) );
na02s02 TIMEBOOST_cell_17931 ( .a(TIMEBOOST_net_4222), .b(FE_OFN1147_n_13249), .o(TIMEBOOST_net_489) );
in01s01 g64232_u0 ( .a(FE_OFN1055_n_4727), .o(g64232_sb) );
na02m02 TIMEBOOST_cell_38838 ( .a(TIMEBOOST_net_11657), .b(g58478_sb), .o(n_9361) );
na02s01 g64232_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(FE_OFN1055_n_4727), .o(g64232_db) );
na02s02 TIMEBOOST_cell_17679 ( .a(TIMEBOOST_net_4096), .b(g61753_sb), .o(n_8309) );
in01s01 g64233_u0 ( .a(FE_OFN1055_n_4727), .o(g64233_sb) );
na02s01 TIMEBOOST_cell_39344 ( .a(TIMEBOOST_net_11910), .b(g64266_db), .o(n_3907) );
na02s01 g64233_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_135), .b(FE_OFN1055_n_4727), .o(g64233_db) );
na02s01 TIMEBOOST_cell_17681 ( .a(TIMEBOOST_net_4097), .b(g61758_sb), .o(n_8297) );
in01s01 g64234_u0 ( .a(FE_OFN1056_n_4727), .o(g64234_sb) );
na02m02 TIMEBOOST_cell_40010 ( .a(TIMEBOOST_net_12243), .b(g62444_sb), .o(n_6707) );
na02s01 g64234_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_136), .b(FE_OFN1056_n_4727), .o(g64234_db) );
na02s01 TIMEBOOST_cell_17683 ( .a(TIMEBOOST_net_4098), .b(g61792_sb), .o(n_8215) );
in01s01 g64235_u0 ( .a(FE_OFN1034_n_4732), .o(g64235_sb) );
na02s02 TIMEBOOST_cell_38497 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__Q), .b(g58352_sb), .o(TIMEBOOST_net_11487) );
na02s01 g64235_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_128), .b(FE_OFN1034_n_4732), .o(g64235_db) );
na02s02 TIMEBOOST_cell_38502 ( .a(TIMEBOOST_net_11489), .b(g58289_db), .o(n_9515) );
in01s01 g64236_u0 ( .a(FE_OFN1033_n_4732), .o(g64236_sb) );
na02s01 TIMEBOOST_cell_38487 ( .a(configuration_pci_err_data), .b(wbm_dat_o_0_), .o(TIMEBOOST_net_11482) );
na02s01 g64236_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_124), .b(FE_OFN1033_n_4732), .o(g64236_db) );
na02f02 TIMEBOOST_cell_38840 ( .a(TIMEBOOST_net_11658), .b(g58460_sb), .o(n_8986) );
in01s01 g64237_u0 ( .a(FE_OFN1055_n_4727), .o(g64237_sb) );
na02m02 TIMEBOOST_cell_40012 ( .a(TIMEBOOST_net_12244), .b(g63008_sb), .o(n_5866) );
na02s01 g64237_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(FE_OFN1055_n_4727), .o(g64237_db) );
na02s02 TIMEBOOST_cell_17685 ( .a(TIMEBOOST_net_4099), .b(g61947_sb), .o(n_7931) );
in01s01 g64238_u0 ( .a(FE_OFN1056_n_4727), .o(g64238_sb) );
na02s02 TIMEBOOST_cell_45103 ( .a(n_1562), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__Q), .o(TIMEBOOST_net_14790) );
na02s01 g64238_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(FE_OFN1056_n_4727), .o(g64238_db) );
na02s02 TIMEBOOST_cell_40014 ( .a(TIMEBOOST_net_12245), .b(g62988_sb), .o(n_5906) );
in01s01 g64239_u0 ( .a(FE_OFN1032_n_4732), .o(g64239_sb) );
na02s01 g64239_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__Q), .b(g64239_sb), .o(g64239_da) );
na02s01 g64239_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_143), .b(FE_OFN1032_n_4732), .o(g64239_db) );
na03s02 TIMEBOOST_cell_38369 ( .a(n_3999), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q), .c(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_11423) );
in01s01 g64240_u0 ( .a(FE_OFN1055_n_4727), .o(g64240_sb) );
na02s01 TIMEBOOST_cell_17932 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__Q), .b(g61943_sb), .o(TIMEBOOST_net_4223) );
na02s01 g64240_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_139), .b(FE_OFN1055_n_4727), .o(g64240_db) );
na02s02 TIMEBOOST_cell_17933 ( .a(TIMEBOOST_net_4223), .b(FE_OFN2021_n_4778), .o(TIMEBOOST_net_859) );
in01s01 g64241_u0 ( .a(FE_OFN917_n_4725), .o(g64241_sb) );
na02s01 g64241_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__21__Q), .b(g64241_sb), .o(g64241_da) );
na02s01 g64241_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_141), .b(FE_OFN917_n_4725), .o(g64241_db) );
na02s01 g64241_u3 ( .a(g64241_da), .b(g64241_db), .o(n_3931) );
in01s01 g64242_u0 ( .a(FE_OFN1056_n_4727), .o(g64242_sb) );
na02s02 TIMEBOOST_cell_43324 ( .a(TIMEBOOST_net_13900), .b(g62358_sb), .o(n_6883) );
na02s01 TIMEBOOST_cell_36301 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__Q), .b(pci_target_unit_fifos_pcir_data_in_174), .o(TIMEBOOST_net_10389) );
na02s01 TIMEBOOST_cell_39366 ( .a(TIMEBOOST_net_11921), .b(g65820_sb), .o(n_1896) );
in01s01 g64243_u0 ( .a(FE_OFN1056_n_4727), .o(g64243_sb) );
na02s01 TIMEBOOST_cell_17934 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__Q), .b(g61943_sb), .o(TIMEBOOST_net_4224) );
na02s01 g64243_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_142), .b(FE_OFN1056_n_4727), .o(g64243_db) );
na02s02 TIMEBOOST_cell_17935 ( .a(TIMEBOOST_net_4224), .b(FE_OFN2021_n_4778), .o(TIMEBOOST_net_858) );
in01s01 g64244_u0 ( .a(FE_OFN1055_n_4727), .o(g64244_sb) );
na02s01 TIMEBOOST_cell_17936 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__Q), .b(g61943_sb), .o(TIMEBOOST_net_4225) );
na02s01 g64244_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_143), .b(FE_OFN1055_n_4727), .o(g64244_db) );
na02s01 TIMEBOOST_cell_17937 ( .a(TIMEBOOST_net_4225), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_861) );
in01s01 g64245_u0 ( .a(FE_OFN1057_n_4727), .o(g64245_sb) );
na02s01 TIMEBOOST_cell_17938 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__Q), .b(g61943_sb), .o(TIMEBOOST_net_4226) );
na02s01 g64245_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_145), .b(FE_OFN1057_n_4727), .o(g64245_db) );
na02s02 TIMEBOOST_cell_17939 ( .a(TIMEBOOST_net_4226), .b(FE_OFN2021_n_4778), .o(TIMEBOOST_net_862) );
in01s01 g64246_u0 ( .a(FE_OFN1055_n_4727), .o(g64246_sb) );
na02m02 TIMEBOOST_cell_17940 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__Q), .b(g53892_sb), .o(TIMEBOOST_net_4227) );
na02s01 g64246_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_146), .b(FE_OFN1055_n_4727), .o(g64246_db) );
na02m02 TIMEBOOST_cell_17941 ( .a(FE_OFN1147_n_13249), .b(TIMEBOOST_net_4227), .o(TIMEBOOST_net_501) );
in01s01 g64247_u0 ( .a(FE_OFN1032_n_4732), .o(g64247_sb) );
na02s01 g64247_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__21__Q), .b(g64247_sb), .o(g64247_da) );
na02s01 g64247_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_141), .b(FE_OFN1032_n_4732), .o(g64247_db) );
na03s02 TIMEBOOST_cell_38145 ( .a(TIMEBOOST_net_4041), .b(g64323_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__Q), .o(TIMEBOOST_net_11311) );
in01s01 g64248_u0 ( .a(FE_OFN1056_n_4727), .o(g64248_sb) );
na02f02 TIMEBOOST_cell_38903 ( .a(n_2695), .b(wbu_addr_in_260), .o(TIMEBOOST_net_11690) );
na02s01 g64248_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_147), .b(FE_OFN1056_n_4727), .o(g64248_db) );
na02f02 TIMEBOOST_cell_38694 ( .a(TIMEBOOST_net_11585), .b(n_7213), .o(TIMEBOOST_net_5590) );
oa12s01 g64249_u0 ( .a(n_3805), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_2__231), .c(FE_OFN1036_n_4732), .o(n_4733) );
in01s01 g64250_u0 ( .a(FE_OFN912_n_4727), .o(g64250_sb) );
na02s02 TIMEBOOST_cell_39398 ( .a(TIMEBOOST_net_11937), .b(g58200_sb), .o(n_9585) );
na02s01 g64250_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(FE_OFN912_n_4727), .o(g64250_db) );
na02m02 TIMEBOOST_cell_44217 ( .a(n_9440), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__Q), .o(TIMEBOOST_net_14347) );
in01s01 g64251_u0 ( .a(FE_OFN1057_n_4727), .o(g64251_sb) );
na02s02 TIMEBOOST_cell_45129 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__Q), .b(n_4002), .o(TIMEBOOST_net_14803) );
na02s01 g64251_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_149), .b(FE_OFN1057_n_4727), .o(g64251_db) );
na02m02 TIMEBOOST_cell_38696 ( .a(TIMEBOOST_net_11586), .b(g59809_sb), .o(n_7614) );
in01s01 g64252_u0 ( .a(FE_OFN912_n_4727), .o(g64252_sb) );
na02s01 TIMEBOOST_cell_39192 ( .a(TIMEBOOST_net_11834), .b(g65734_sb), .o(n_1909) );
na02s01 g64252_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(FE_OFN912_n_4727), .o(g64252_db) );
na02s01 TIMEBOOST_cell_37165 ( .a(n_1992), .b(n_245), .o(TIMEBOOST_net_10821) );
in01s01 g64253_u0 ( .a(FE_OFN1033_n_4732), .o(g64253_sb) );
na02s01 g64253_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__Q), .b(g64253_sb), .o(g64253_da) );
na02s01 g64253_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(FE_OFN1033_n_4732), .o(g64253_db) );
na02s01 TIMEBOOST_cell_37456 ( .a(TIMEBOOST_net_10966), .b(FE_OFN775_n_15366), .o(TIMEBOOST_net_10566) );
in01s01 g64254_u0 ( .a(FE_OFN918_n_4725), .o(g64254_sb) );
na02f02 TIMEBOOST_cell_37049 ( .a(TIMEBOOST_net_10131), .b(n_13901), .o(TIMEBOOST_net_10763) );
na02s01 g64254_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_139), .b(FE_OFN918_n_4725), .o(g64254_db) );
na02f02 TIMEBOOST_cell_37048 ( .a(TIMEBOOST_net_10762), .b(FE_OFN1768_n_14054), .o(g53262_p) );
in01s01 g64255_u0 ( .a(FE_OFN912_n_4727), .o(g64255_sb) );
na03s02 TIMEBOOST_cell_38121 ( .a(g64169_da), .b(g64169_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__Q), .o(TIMEBOOST_net_11299) );
na02s02 TIMEBOOST_cell_40016 ( .a(TIMEBOOST_net_12246), .b(g62562_sb), .o(n_6435) );
na02s01 TIMEBOOST_cell_19873 ( .a(TIMEBOOST_net_5193), .b(g62984_sb), .o(n_5914) );
in01s01 g64256_u0 ( .a(FE_OFN912_n_4727), .o(g64256_sb) );
na02s02 TIMEBOOST_cell_44426 ( .a(TIMEBOOST_net_14451), .b(FE_OFN1305_n_13124), .o(TIMEBOOST_net_13426) );
na02s01 g64256_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in_153), .b(FE_OFN912_n_4727), .o(g64256_db) );
na02m02 TIMEBOOST_cell_38698 ( .a(TIMEBOOST_net_11587), .b(g62960_sb), .o(n_5962) );
in01s01 g64257_u0 ( .a(FE_OFN1057_n_4727), .o(g64257_sb) );
na02f02 TIMEBOOST_cell_43796 ( .a(TIMEBOOST_net_14136), .b(FE_OFN1370_n_8567), .o(TIMEBOOST_net_12687) );
na02s01 g64257_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(FE_OFN1057_n_4727), .o(g64257_db) );
na02s02 TIMEBOOST_cell_38768 ( .a(TIMEBOOST_net_11622), .b(g53923_sb), .o(n_13521) );
in01s01 g64258_u0 ( .a(FE_OFN1032_n_4732), .o(g64258_sb) );
na02s01 TIMEBOOST_cell_18290 ( .a(g61923_sb), .b(g61973_db), .o(TIMEBOOST_net_4402) );
na02s01 g64258_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_139), .b(FE_OFN1032_n_4732), .o(g64258_db) );
na02s02 TIMEBOOST_cell_38504 ( .a(TIMEBOOST_net_11490), .b(g58292_db), .o(n_9512) );
in01s01 g64259_u0 ( .a(FE_OFN1057_n_4727), .o(g64259_sb) );
na02s01 TIMEBOOST_cell_9834 ( .a(wbu_latency_tim_val_in_249), .b(n_6986), .o(TIMEBOOST_net_1484) );
na02s01 g64259_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_123), .b(FE_OFN1057_n_4727), .o(g64259_db) );
na02s01 TIMEBOOST_cell_9835 ( .a(TIMEBOOST_net_1484), .b(g58611_sb), .o(TIMEBOOST_net_905) );
in01s01 g64260_u0 ( .a(FE_OFN1055_n_4727), .o(g64260_sb) );
na02m02 TIMEBOOST_cell_43797 ( .a(n_9838), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__Q), .o(TIMEBOOST_net_14137) );
na02s01 g64260_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_124), .b(FE_OFN1055_n_4727), .o(g64260_db) );
na02s02 TIMEBOOST_cell_38770 ( .a(TIMEBOOST_net_11623), .b(g53902_sb), .o(n_13539) );
in01s01 g64261_u0 ( .a(FE_OFN1057_n_4727), .o(g64261_sb) );
na02s01 g64261_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__Q), .b(g64261_sb), .o(g64261_da) );
na02s01 g64261_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_125), .b(FE_OFN1057_n_4727), .o(g64261_db) );
na02s02 TIMEBOOST_cell_38506 ( .a(TIMEBOOST_net_11491), .b(g58358_db), .o(n_9465) );
in01s01 g64262_u0 ( .a(FE_OFN1058_n_4727), .o(g64262_sb) );
na02s01 g64262_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__6__Q), .b(g64262_sb), .o(g64262_da) );
na02s01 g64262_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(FE_OFN1058_n_4727), .o(g64262_db) );
na02s02 TIMEBOOST_cell_40018 ( .a(TIMEBOOST_net_12247), .b(g62956_sb), .o(n_5969) );
in01s01 g64263_u0 ( .a(FE_OFN1055_n_4727), .o(g64263_sb) );
na02f02 TIMEBOOST_cell_43798 ( .a(TIMEBOOST_net_14137), .b(FE_OFN1414_n_8567), .o(TIMEBOOST_net_12881) );
na02s01 g64263_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_127), .b(FE_OFN1055_n_4727), .o(g64263_db) );
na02f02 TIMEBOOST_cell_38900 ( .a(TIMEBOOST_net_11688), .b(FE_OFN2200_n_10256), .o(TIMEBOOST_net_10707) );
in01s01 g64264_u0 ( .a(FE_OFN912_n_4727), .o(g64264_sb) );
na02s01 TIMEBOOST_cell_17580 ( .a(FE_OFN1780_parchk_pci_ad_reg_in_1221), .b(g65813_sb), .o(TIMEBOOST_net_4047) );
na02s01 g64264_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_128), .b(FE_OFN912_n_4727), .o(g64264_db) );
na02s01 TIMEBOOST_cell_17581 ( .a(TIMEBOOST_net_4047), .b(g65968_db), .o(n_2570) );
in01s01 g64265_u0 ( .a(FE_OFN1055_n_4727), .o(g64265_sb) );
na02f02 TIMEBOOST_cell_38901 ( .a(n_3471), .b(wbu_addr_in_277), .o(TIMEBOOST_net_11689) );
na02s01 g64265_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(FE_OFN1055_n_4727), .o(g64265_db) );
na02s02 TIMEBOOST_cell_39400 ( .a(TIMEBOOST_net_11938), .b(FE_OFN266_n_9884), .o(n_9676) );
in01s01 g64266_u0 ( .a(FE_OFN1037_n_4732), .o(g64266_sb) );
na02s02 TIMEBOOST_cell_37430 ( .a(TIMEBOOST_net_10953), .b(n_4672), .o(TIMEBOOST_net_5436) );
na02s01 g64266_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_136), .b(FE_OFN1037_n_4732), .o(g64266_db) );
na02s01 TIMEBOOST_cell_37431 ( .a(TIMEBOOST_net_9401), .b(FE_OFN2108_n_2047), .o(TIMEBOOST_net_10954) );
in01s01 g64267_u0 ( .a(FE_OFN1036_n_4732), .o(g64267_sb) );
na02s01 g64267_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__Q), .b(g64267_sb), .o(g64267_da) );
na02s01 g64267_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in_153), .b(FE_OFN1036_n_4732), .o(g64267_db) );
na02m02 TIMEBOOST_cell_38307 ( .a(TIMEBOOST_net_1822), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_408), .o(TIMEBOOST_net_11392) );
in01s01 g64268_u0 ( .a(FE_OFN928_n_4730), .o(g64268_sb) );
na02s01 TIMEBOOST_cell_16907 ( .a(TIMEBOOST_net_3710), .b(g65855_db), .o(n_1873) );
na02s01 g64268_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_130), .b(FE_OFN928_n_4730), .o(g64268_db) );
na02s01 TIMEBOOST_cell_16908 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q), .b(g64289_sb), .o(TIMEBOOST_net_3711) );
in01s01 g64269_u0 ( .a(FE_OFN928_n_4730), .o(g64269_sb) );
na02s01 g64269_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__Q), .b(g64269_sb), .o(g64269_da) );
na02s01 g64269_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(FE_OFN928_n_4730), .o(g64269_db) );
na02s01 TIMEBOOST_cell_36642 ( .a(TIMEBOOST_net_10559), .b(g65947_db), .o(n_2574) );
in01s01 g64270_u0 ( .a(FE_OFN928_n_4730), .o(g64270_sb) );
na02s01 TIMEBOOST_cell_36644 ( .a(TIMEBOOST_net_10560), .b(g65945_db), .o(n_2576) );
na02s01 g64270_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_132), .b(FE_OFN928_n_4730), .o(g64270_db) );
na02m02 TIMEBOOST_cell_40020 ( .a(TIMEBOOST_net_12248), .b(g62558_sb), .o(n_6446) );
in01s01 g64271_u0 ( .a(FE_OFN928_n_4730), .o(g64271_sb) );
na02s01 TIMEBOOST_cell_45164 ( .a(TIMEBOOST_net_14820), .b(FE_OFN1252_n_4143), .o(TIMEBOOST_net_12031) );
na02s01 g64271_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(FE_OFN928_n_4730), .o(g64271_db) );
na02s02 TIMEBOOST_cell_40022 ( .a(TIMEBOOST_net_12249), .b(g62612_sb), .o(n_6333) );
in01s01 g64272_u0 ( .a(FE_OFN1032_n_4732), .o(g64272_sb) );
na02s01 g64272_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__Q), .b(g64272_sb), .o(g64272_da) );
na02s01 g64272_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_135), .b(FE_OFN1032_n_4732), .o(g64272_db) );
na03s02 TIMEBOOST_cell_38345 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__Q), .b(FE_OFN1128_g64577_p), .c(n_3588), .o(TIMEBOOST_net_11411) );
in01s01 g64273_u0 ( .a(FE_OFN928_n_4730), .o(g64273_sb) );
na02s01 g64273_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__14__Q), .b(g64273_sb), .o(g64273_da) );
na02s01 g64273_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(FE_OFN928_n_4730), .o(g64273_db) );
na02s01 TIMEBOOST_cell_44977 ( .a(FE_OFN211_n_9858), .b(g57981_sb), .o(TIMEBOOST_net_14727) );
in01s01 g64274_u0 ( .a(FE_OFN928_n_4730), .o(g64274_sb) );
na02s01 g64274_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__15__Q), .b(g64274_sb), .o(g64274_da) );
na02s01 g64274_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_135), .b(FE_OFN928_n_4730), .o(g64274_db) );
na02m02 TIMEBOOST_cell_44187 ( .a(n_9591), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__Q), .o(TIMEBOOST_net_14332) );
in01s01 g64275_u0 ( .a(FE_OFN928_n_4730), .o(g64275_sb) );
na02s01 TIMEBOOST_cell_16912 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__Q), .b(g65288_sb), .o(TIMEBOOST_net_3713) );
na02s01 g64275_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_136), .b(FE_OFN928_n_4730), .o(g64275_db) );
na02s01 TIMEBOOST_cell_16913 ( .a(TIMEBOOST_net_3713), .b(g65288_db), .o(n_3580) );
in01s01 g64276_u0 ( .a(FE_OFN928_n_4730), .o(g64276_sb) );
na02s01 TIMEBOOST_cell_16914 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__Q), .b(g65398_sb), .o(TIMEBOOST_net_3714) );
na02s01 g64276_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(FE_OFN928_n_4730), .o(g64276_db) );
na02s02 TIMEBOOST_cell_40024 ( .a(TIMEBOOST_net_12250), .b(g62569_sb), .o(n_6417) );
in01s01 g64277_u0 ( .a(FE_OFN930_n_4730), .o(g64277_sb) );
na02s01 g64277_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__18__Q), .b(g64277_sb), .o(g64277_da) );
na02s01 g64277_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(FE_OFN930_n_4730), .o(g64277_db) );
na02f02 TIMEBOOST_cell_38813 ( .a(n_3006), .b(wbu_addr_in_259), .o(TIMEBOOST_net_11645) );
in01s01 g64278_u0 ( .a(FE_OFN917_n_4725), .o(g64278_sb) );
na02s01 g64278_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__Q), .b(g64278_sb), .o(g64278_da) );
na02s01 g64278_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(FE_OFN917_n_4725), .o(g64278_db) );
na02s01 TIMEBOOST_cell_44978 ( .a(TIMEBOOST_net_14727), .b(g57981_db), .o(n_9818) );
in01s01 g64279_u0 ( .a(FE_OFN930_n_4730), .o(g64279_sb) );
na02s02 TIMEBOOST_cell_40026 ( .a(TIMEBOOST_net_12251), .b(g62947_sb), .o(n_5987) );
na02s01 g64279_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_139), .b(FE_OFN930_n_4730), .o(g64279_db) );
na02s02 TIMEBOOST_cell_39549 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__Q), .b(g58363_sb), .o(TIMEBOOST_net_12013) );
in01s01 g64280_u0 ( .a(FE_OFN928_n_4730), .o(g64280_sb) );
na02s02 TIMEBOOST_cell_40028 ( .a(TIMEBOOST_net_12252), .b(g63178_sb), .o(n_5792) );
na02s01 g64280_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_140), .b(FE_OFN928_n_4730), .o(g64280_db) );
na02s02 TIMEBOOST_cell_42867 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__Q), .b(FE_OFN1654_n_9502), .o(TIMEBOOST_net_13672) );
in01s01 g64281_u0 ( .a(FE_OFN930_n_4730), .o(g64281_sb) );
na02s01 g64281_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__21__Q), .b(g64281_sb), .o(g64281_da) );
na02s01 g64281_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_141), .b(FE_OFN930_n_4730), .o(g64281_db) );
na02f02 TIMEBOOST_cell_38815 ( .a(n_3139), .b(wbu_addr_in_269), .o(TIMEBOOST_net_11646) );
in01s01 g64282_u0 ( .a(FE_OFN928_n_4730), .o(g64282_sb) );
na02s02 TIMEBOOST_cell_40030 ( .a(TIMEBOOST_net_12253), .b(g63004_sb), .o(n_5874) );
na02s01 g64282_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_142), .b(FE_OFN928_n_4730), .o(g64282_db) );
na02s02 TIMEBOOST_cell_45165 ( .a(n_4407), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__Q), .o(TIMEBOOST_net_14821) );
in01s01 g64283_u0 ( .a(FE_OFN1037_n_4732), .o(g64283_sb) );
na02s02 TIMEBOOST_cell_37432 ( .a(TIMEBOOST_net_10954), .b(g65690_sb), .o(n_1953) );
na02s01 g64283_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(FE_OFN1037_n_4732), .o(g64283_db) );
na02s02 TIMEBOOST_cell_37433 ( .a(TIMEBOOST_net_9404), .b(FE_OFN1797_n_2299), .o(TIMEBOOST_net_10955) );
in01s01 g64284_u0 ( .a(FE_OFN928_n_4730), .o(g64284_sb) );
na02s01 g64284_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__Q), .b(g64284_sb), .o(g64284_da) );
na02s01 g64284_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_143), .b(FE_OFN928_n_4730), .o(g64284_db) );
na02s02 TIMEBOOST_cell_44979 ( .a(n_2167), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__Q), .o(TIMEBOOST_net_14728) );
in01s01 g64285_u0 ( .a(FE_OFN930_n_4730), .o(g64285_sb) );
na02s02 TIMEBOOST_cell_45166 ( .a(TIMEBOOST_net_14821), .b(FE_OFN1283_n_4097), .o(TIMEBOOST_net_12032) );
na02s01 g64285_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_144), .b(FE_OFN930_n_4730), .o(g64285_db) );
na02s01 TIMEBOOST_cell_16876 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__Q), .b(g64292_sb), .o(TIMEBOOST_net_3695) );
in01s01 g64286_u0 ( .a(FE_OFN927_n_4730), .o(g64286_sb) );
na02s02 TIMEBOOST_cell_45683 ( .a(n_3565), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__Q), .o(TIMEBOOST_net_15080) );
na03s02 TIMEBOOST_cell_43325 ( .a(n_4402), .b(FE_OFN1223_n_6391), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__Q), .o(TIMEBOOST_net_13901) );
na02f02 TIMEBOOST_cell_42488 ( .a(TIMEBOOST_net_13482), .b(g57485_sb), .o(n_10332) );
in01s01 g64287_u0 ( .a(FE_OFN928_n_4730), .o(g64287_sb) );
na02s01 TIMEBOOST_cell_16877 ( .a(TIMEBOOST_net_3695), .b(g64292_db), .o(n_3881) );
na02s01 g64287_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_147), .b(FE_OFN928_n_4730), .o(g64287_db) );
na02s02 TIMEBOOST_cell_40670 ( .a(TIMEBOOST_net_12573), .b(g62450_sb), .o(n_6697) );
in01s01 g64288_u0 ( .a(FE_OFN1031_n_4732), .o(g64288_sb) );
na02s01 g64288_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__Q), .b(g64288_sb), .o(g64288_da) );
na02s01 g64288_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_150), .b(FE_OFN1031_n_4732), .o(g64288_db) );
in01s01 TIMEBOOST_cell_45934 ( .a(TIMEBOOST_net_15240), .o(TIMEBOOST_net_15241) );
in01s01 g64289_u0 ( .a(FE_OFN927_n_4730), .o(g64289_sb) );
na02s01 TIMEBOOST_cell_42934 ( .a(TIMEBOOST_net_13705), .b(FE_OFN270_n_9836), .o(TIMEBOOST_net_11932) );
na02s01 g64289_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(FE_OFN927_n_4730), .o(g64289_db) );
na03s02 TIMEBOOST_cell_42909 ( .a(g64293_da), .b(g64293_db), .c(g63077_sb), .o(TIMEBOOST_net_13693) );
in01s01 g64290_u0 ( .a(FE_OFN927_n_4730), .o(g64290_sb) );
na02s01 g64290_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__Q), .b(g64290_sb), .o(g64290_da) );
na02s01 g64290_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(FE_OFN927_n_4730), .o(g64290_db) );
na02s02 TIMEBOOST_cell_45197 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__Q), .b(n_3597), .o(TIMEBOOST_net_14837) );
in01s01 g64291_u0 ( .a(FE_OFN929_n_4730), .o(g64291_sb) );
na02s01 g64291_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__Q), .b(g64291_sb), .o(g64291_da) );
na02s01 g64291_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_150), .b(FE_OFN929_n_4730), .o(g64291_db) );
na02m02 TIMEBOOST_cell_44195 ( .a(n_9456), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__Q), .o(TIMEBOOST_net_14336) );
in01s01 g64292_u0 ( .a(FE_OFN927_n_4730), .o(g64292_sb) );
na02s02 TIMEBOOST_cell_41894 ( .a(TIMEBOOST_net_13185), .b(TIMEBOOST_net_4332), .o(n_4965) );
na02s01 g64292_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_151), .b(FE_OFN927_n_4730), .o(g64292_db) );
na02s01 TIMEBOOST_cell_30966 ( .a(n_3749), .b(g64929_sb), .o(TIMEBOOST_net_9394) );
in01s01 g64293_u0 ( .a(FE_OFN929_n_4730), .o(g64293_sb) );
na02s01 g64293_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q), .b(g64293_sb), .o(g64293_da) );
na02s01 g64293_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in), .b(FE_OFN929_n_4730), .o(g64293_db) );
na02s01 TIMEBOOST_cell_16924 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__Q), .b(g65410_sb), .o(TIMEBOOST_net_3719) );
na02s02 TIMEBOOST_cell_43013 ( .a(n_3864), .b(g63101_db), .o(TIMEBOOST_net_13745) );
na02s02 TIMEBOOST_cell_43056 ( .a(TIMEBOOST_net_13766), .b(FE_OFN1268_n_4095), .o(TIMEBOOST_net_12139) );
na02f02 TIMEBOOST_cell_42204 ( .a(TIMEBOOST_net_13340), .b(FE_OFN1407_n_8567), .o(TIMEBOOST_net_12292) );
in01s01 g64295_u0 ( .a(FE_OFN927_n_4730), .o(g64295_sb) );
na02s01 g64295_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__Q), .b(g64295_sb), .o(g64295_da) );
na02s01 g64295_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in_153), .b(FE_OFN927_n_4730), .o(g64295_db) );
na02m02 TIMEBOOST_cell_43799 ( .a(n_9805), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__Q), .o(TIMEBOOST_net_14138) );
in01s01 g64296_u0 ( .a(FE_OFN917_n_4725), .o(g64296_sb) );
na02s01 TIMEBOOST_cell_40526 ( .a(TIMEBOOST_net_12501), .b(FE_OFN1301_n_5763), .o(TIMEBOOST_net_11499) );
na02s01 g64296_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_132), .b(FE_OFN917_n_4725), .o(g64296_db) );
na02f02 TIMEBOOST_cell_37051 ( .a(TIMEBOOST_net_10129), .b(n_13891), .o(TIMEBOOST_net_10764) );
in01s01 g64297_u0 ( .a(FE_OFN1034_n_4732), .o(g64297_sb) );
na02s01 TIMEBOOST_cell_18146 ( .a(g63561_sb), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_), .o(TIMEBOOST_net_4330) );
na02s01 g64297_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_130), .b(FE_OFN1034_n_4732), .o(g64297_db) );
na02s01 TIMEBOOST_cell_18147 ( .a(TIMEBOOST_net_4330), .b(g63561_db), .o(n_4113) );
in01s01 g64298_u0 ( .a(FE_OFN929_n_4730), .o(g64298_sb) );
na02s02 TIMEBOOST_cell_42944 ( .a(TIMEBOOST_net_13710), .b(g63141_sb), .o(TIMEBOOST_net_4332) );
na02s01 g64298_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(FE_OFN929_n_4730), .o(g64298_db) );
na03f02 TIMEBOOST_cell_8797 ( .a(n_11839), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__Q), .c(FE_OCPN1866_n_12377), .o(n_12742) );
oa12s01 g64299_u0 ( .a(n_3807), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_1__192), .c(n_4730), .o(n_4729) );
in01s01 g64300_u0 ( .a(FE_OFN1031_n_4732), .o(g64300_sb) );
na02s02 TIMEBOOST_cell_38503 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__Q), .b(g58292_sb), .o(TIMEBOOST_net_11490) );
na02s01 g64300_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_123), .b(FE_OFN1031_n_4732), .o(g64300_db) );
na02s01 TIMEBOOST_cell_38508 ( .a(TIMEBOOST_net_11492), .b(FE_OFN1279_n_4097), .o(TIMEBOOST_net_5199) );
in01s01 g64301_u0 ( .a(FE_OFN929_n_4730), .o(g64301_sb) );
na03f02 TIMEBOOST_cell_36056 ( .a(FE_OFN1601_n_13995), .b(TIMEBOOST_net_10174), .c(FE_OFN1605_n_13997), .o(n_14512) );
na02s01 g64301_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_123), .b(FE_OFN929_n_4730), .o(g64301_db) );
na02s01 TIMEBOOST_cell_16898 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q), .b(g64271_sb), .o(TIMEBOOST_net_3706) );
in01s01 g64302_u0 ( .a(FE_OFN929_n_4730), .o(g64302_sb) );
na02s01 g64302_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__Q), .b(g64302_sb), .o(g64302_da) );
na02s01 g64302_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_125), .b(FE_OFN929_n_4730), .o(g64302_db) );
na02s02 TIMEBOOST_cell_36772 ( .a(TIMEBOOST_net_10624), .b(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_4693) );
na02f02 TIMEBOOST_cell_21993 ( .a(TIMEBOOST_net_6253), .b(FE_OFN1774_n_13800), .o(n_14479) );
na02s02 TIMEBOOST_cell_45684 ( .a(TIMEBOOST_net_15080), .b(FE_OFN1275_n_4096), .o(TIMEBOOST_net_13271) );
na02s02 TIMEBOOST_cell_40032 ( .a(TIMEBOOST_net_12254), .b(g62535_sb), .o(n_6501) );
in01s01 g64304_u0 ( .a(FE_OFN928_n_4730), .o(g64304_sb) );
na02s01 TIMEBOOST_cell_42935 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__Q), .b(FE_OFN533_n_9823), .o(TIMEBOOST_net_13706) );
na02s01 g64304_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_127), .b(FE_OFN928_n_4730), .o(g64304_db) );
na02s02 TIMEBOOST_cell_43265 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__Q), .b(n_4484), .o(TIMEBOOST_net_13871) );
na02m02 TIMEBOOST_cell_39194 ( .a(TIMEBOOST_net_11835), .b(wbu_addr_in_252), .o(n_9828) );
na03s02 TIMEBOOST_cell_40727 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__Q), .b(n_3567), .c(FE_OFN1207_n_6356), .o(TIMEBOOST_net_12602) );
na02s01 TIMEBOOST_cell_17245 ( .a(TIMEBOOST_net_3879), .b(g65424_da), .o(n_4224) );
in01s01 g64306_u0 ( .a(FE_OFN928_n_4730), .o(g64306_sb) );
na02s01 g64306_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__Q), .b(g64306_sb), .o(g64306_da) );
na02s01 g64306_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(FE_OFN928_n_4730), .o(g64306_db) );
na02s01 TIMEBOOST_cell_9850 ( .a(n_272), .b(FE_OCP_RBN1917_wbs_cti_i_1_), .o(TIMEBOOST_net_1492) );
in01s01 g64307_u0 ( .a(FE_OFN1033_n_4732), .o(g64307_sb) );
na02s01 g64307_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__Q), .b(g64307_sb), .o(g64307_da) );
na02s01 g64307_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(FE_OFN1033_n_4732), .o(g64307_db) );
na02s01 TIMEBOOST_cell_39333 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__Q), .b(g64243_sb), .o(TIMEBOOST_net_11905) );
in01s01 g64308_u0 ( .a(FE_OFN1037_n_4732), .o(g64308_sb) );
na02s02 TIMEBOOST_cell_44839 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__Q), .b(FE_OFN1642_n_4671), .o(TIMEBOOST_net_14658) );
na02s01 g64308_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_132), .b(FE_OFN1037_n_4732), .o(g64308_db) );
na02s02 TIMEBOOST_cell_40034 ( .a(TIMEBOOST_net_12255), .b(g63161_sb), .o(n_5814) );
in01s01 g64309_u0 ( .a(FE_OFN1032_n_4732), .o(g64309_sb) );
na02s01 g64309_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__Q), .b(g64309_sb), .o(g64309_da) );
na02s01 g64309_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(FE_OFN1032_n_4732), .o(g64309_db) );
na02m02 TIMEBOOST_cell_38975 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_5__Q), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__Q), .o(TIMEBOOST_net_11726) );
in01s01 g64310_u0 ( .a(FE_OFN1032_n_4732), .o(g64310_sb) );
na02s01 g64310_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__Q), .b(g64310_sb), .o(g64310_da) );
na02s01 g64310_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(FE_OFN1032_n_4732), .o(g64310_db) );
na03s02 TIMEBOOST_cell_38115 ( .a(g64119_da), .b(g64119_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__Q), .o(TIMEBOOST_net_11296) );
in01s01 g64311_u0 ( .a(FE_OFN1032_n_4732), .o(g64311_sb) );
na02s01 TIMEBOOST_cell_18152 ( .a(g63573_sb), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_), .o(TIMEBOOST_net_4333) );
na02s01 g64311_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(FE_OFN1032_n_4732), .o(g64311_db) );
na02s01 TIMEBOOST_cell_18153 ( .a(TIMEBOOST_net_4333), .b(g63573_db), .o(n_4108) );
in01s01 g64312_u0 ( .a(FE_OFN1037_n_4732), .o(g64312_sb) );
na03s01 TIMEBOOST_cell_38509 ( .a(g65377_da), .b(g65377_db), .c(n_14), .o(TIMEBOOST_net_11493) );
na02s01 g64312_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_140), .b(FE_OFN1037_n_4732), .o(g64312_db) );
na02s01 TIMEBOOST_cell_38510 ( .a(TIMEBOOST_net_11493), .b(FE_OFN1226_n_6391), .o(TIMEBOOST_net_5231) );
in01s01 g64313_u0 ( .a(FE_OFN1037_n_4732), .o(g64313_sb) );
na02s01 TIMEBOOST_cell_43098 ( .a(TIMEBOOST_net_13787), .b(FE_OFN1223_n_6391), .o(TIMEBOOST_net_13250) );
na02s01 g64313_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_142), .b(FE_OFN1037_n_4732), .o(g64313_db) );
na02s02 TIMEBOOST_cell_18157 ( .a(TIMEBOOST_net_4335), .b(g58341_sb), .o(n_9479) );
in01s01 g64314_u0 ( .a(FE_OFN1034_n_4732), .o(g64314_sb) );
na02s02 TIMEBOOST_cell_43099 ( .a(n_3575), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__Q), .o(TIMEBOOST_net_13788) );
na02s01 g64314_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_144), .b(FE_OFN1034_n_4732), .o(g64314_db) );
na02s02 TIMEBOOST_cell_42857 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__Q), .b(n_2154), .o(TIMEBOOST_net_13667) );
in01s01 g64315_u0 ( .a(FE_OFN959_n_2299), .o(g64315_sb) );
na03s02 TIMEBOOST_cell_36775 ( .a(g64348_da), .b(g64348_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__Q), .o(TIMEBOOST_net_10626) );
na02s01 g64315_u2 ( .a(pci_target_unit_fifos_pcir_control_in_192), .b(FE_OFN959_n_2299), .o(g64315_db) );
na02s02 TIMEBOOST_cell_44980 ( .a(TIMEBOOST_net_14728), .b(FE_OFN706_n_8119), .o(TIMEBOOST_net_11049) );
in01s01 g64316_u0 ( .a(FE_OFN1033_n_4732), .o(g64316_sb) );
na02s01 g64316_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__Q), .b(g64316_sb), .o(g64316_da) );
na02s01 g64316_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_146), .b(FE_OFN1033_n_4732), .o(g64316_db) );
na02s01 TIMEBOOST_cell_38477 ( .a(n_1709), .b(g61746_sb), .o(TIMEBOOST_net_11477) );
in01s01 g64317_u0 ( .a(FE_OFN930_n_4730), .o(g64317_sb) );
na02s01 g64317_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_124), .b(FE_OFN930_n_4730), .o(g64317_db) );
na02s02 TIMEBOOST_cell_40036 ( .a(TIMEBOOST_net_12256), .b(g62902_sb), .o(n_6073) );
in01s01 g64318_u0 ( .a(FE_OFN1037_n_4732), .o(g64318_sb) );
na02s02 TIMEBOOST_cell_45685 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__Q), .b(n_4345), .o(TIMEBOOST_net_15081) );
na02s01 g64318_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_147), .b(FE_OFN1037_n_4732), .o(g64318_db) );
na03s02 TIMEBOOST_cell_38149 ( .a(TIMEBOOST_net_3550), .b(g64360_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__Q), .o(TIMEBOOST_net_11313) );
in01s01 g64319_u0 ( .a(FE_OFN1034_n_4732), .o(g64319_sb) );
na02f02 TIMEBOOST_cell_42490 ( .a(TIMEBOOST_net_13483), .b(g57093_sb), .o(n_11648) );
na02s01 g64319_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(FE_OFN1034_n_4732), .o(g64319_db) );
na02f02 TIMEBOOST_cell_44702 ( .a(TIMEBOOST_net_14589), .b(g52516_sb), .o(n_13709) );
in01s01 g64320_u0 ( .a(FE_OFN1031_n_4732), .o(g64320_sb) );
na02s01 g64320_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__Q), .b(g64320_sb), .o(g64320_da) );
na02s01 g64320_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_149), .b(FE_OFN1031_n_4732), .o(g64320_db) );
in01s01 TIMEBOOST_cell_45935 ( .a(wbm_dat_i_26_), .o(TIMEBOOST_net_15242) );
in01s01 g64321_u0 ( .a(FE_OFN1033_n_4732), .o(g64321_sb) );
na02s01 g64321_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__Q), .b(g64321_sb), .o(g64321_da) );
na02s01 g64321_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_127), .b(FE_OFN1033_n_4732), .o(g64321_db) );
na02s02 TIMEBOOST_cell_43595 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__26__Q), .b(n_4335), .o(TIMEBOOST_net_14036) );
in01s01 g64322_u0 ( .a(FE_OFN1034_n_4732), .o(g64322_sb) );
na02f02 TIMEBOOST_cell_38902 ( .a(TIMEBOOST_net_11689), .b(FE_OFN2200_n_10256), .o(TIMEBOOST_net_10708) );
na02s01 g64322_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(FE_OFN1034_n_4732), .o(g64322_db) );
na02m02 TIMEBOOST_cell_18165 ( .a(TIMEBOOST_net_4339), .b(g54161_sb), .o(n_13554) );
in01s01 g64323_u0 ( .a(FE_OFN1034_n_4732), .o(g64323_sb) );
na03s02 TIMEBOOST_cell_38393 ( .a(n_4032), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__Q), .c(FE_OFN1119_g64577_p), .o(TIMEBOOST_net_11435) );
na02s01 g64323_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_151), .b(FE_OFN1034_n_4732), .o(g64323_db) );
na02s02 TIMEBOOST_cell_38512 ( .a(TIMEBOOST_net_11494), .b(g58359_db), .o(n_9464) );
in01s01 g64324_u0 ( .a(FE_OFN1034_n_4732), .o(g64324_sb) );
na02s01 g64324_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__Q), .b(g64324_sb), .o(g64324_da) );
na02s01 g64324_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in_152), .b(FE_OFN1034_n_4732), .o(g64324_db) );
na03s02 TIMEBOOST_cell_38513 ( .a(TIMEBOOST_net_4176), .b(g64763_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__Q), .o(TIMEBOOST_net_11495) );
in01s01 g64325_u0 ( .a(FE_OFN1031_n_4732), .o(g64325_sb) );
na02s01 TIMEBOOST_cell_38455 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__Q), .b(g58409_sb), .o(TIMEBOOST_net_11466) );
na02s01 g64325_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(FE_OFN1031_n_4732), .o(g64325_db) );
na02s02 TIMEBOOST_cell_38514 ( .a(TIMEBOOST_net_11495), .b(FE_OFN1261_n_4143), .o(TIMEBOOST_net_5234) );
in01s01 g64326_u0 ( .a(FE_OFN1035_n_4732), .o(g64326_sb) );
na02f04 TIMEBOOST_cell_45520 ( .a(TIMEBOOST_net_14998), .b(g54340_sb), .o(n_12976) );
na02s01 g64326_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(FE_OFN1035_n_4732), .o(g64326_db) );
na02m02 TIMEBOOST_cell_18171 ( .a(TIMEBOOST_net_4342), .b(TIMEBOOST_net_501), .o(n_13553) );
in01s01 g64327_u0 ( .a(FE_OFN916_n_4725), .o(g64327_sb) );
na02s01 TIMEBOOST_cell_40527 ( .a(wishbone_slave_unit_pcim_sm_data_in_645), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__Q), .o(TIMEBOOST_net_12502) );
na02s01 g64327_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_130), .b(FE_OFN916_n_4725), .o(g64327_db) );
na02s01 TIMEBOOST_cell_40528 ( .a(TIMEBOOST_net_12502), .b(FE_OFN1301_n_5763), .o(TIMEBOOST_net_11517) );
in01s01 g64328_u0 ( .a(FE_OFN917_n_4725), .o(g64328_sb) );
na02s01 TIMEBOOST_cell_40529 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__Q), .b(wishbone_slave_unit_pcim_sm_data_in_639), .o(TIMEBOOST_net_12503) );
na02f02 TIMEBOOST_cell_44188 ( .a(TIMEBOOST_net_14332), .b(FE_OFN1370_n_8567), .o(TIMEBOOST_net_13400) );
na02f02 TIMEBOOST_cell_37050 ( .a(FE_OFN1593_n_13741), .b(TIMEBOOST_net_10763), .o(g53243_p) );
in01s01 g64329_u0 ( .a(FE_OFN917_n_4725), .o(g64329_sb) );
na02s01 g64329_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__Q), .b(g64329_sb), .o(g64329_da) );
na02s01 g64329_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_135), .b(FE_OFN917_n_4725), .o(g64329_db) );
na02s02 TIMEBOOST_cell_45104 ( .a(TIMEBOOST_net_14790), .b(FE_OFN1812_n_7845), .o(TIMEBOOST_net_11389) );
in01s01 g64330_u0 ( .a(FE_OFN917_n_4725), .o(g64330_sb) );
na02s01 g64330_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__16__Q), .b(g64330_sb), .o(g64330_da) );
na02s01 g64330_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_136), .b(FE_OFN917_n_4725), .o(g64330_db) );
na02s01 TIMEBOOST_cell_9194 ( .a(pci_target_unit_fifos_pcir_data_in), .b(g65712_sb), .o(TIMEBOOST_net_1164) );
in01s01 g64331_u0 ( .a(FE_OFN917_n_4725), .o(g64331_sb) );
na02s01 g64331_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__Q), .b(g64331_sb), .o(g64331_da) );
na02s01 g64331_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(FE_OFN917_n_4725), .o(g64331_db) );
in01s01 g64332_u0 ( .a(FE_OFN1057_n_4727), .o(g64332_sb) );
na02s01 TIMEBOOST_cell_17956 ( .a(n_4452), .b(FE_OFN1680_n_4655), .o(TIMEBOOST_net_4235) );
na02s01 g64332_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in), .b(FE_OFN1057_n_4727), .o(g64332_db) );
na02s01 TIMEBOOST_cell_17957 ( .a(TIMEBOOST_net_4235), .b(g65396_da), .o(n_4239) );
in01s01 g64333_u0 ( .a(FE_OFN917_n_4725), .o(g64333_sb) );
na02s02 TIMEBOOST_cell_40672 ( .a(TIMEBOOST_net_12574), .b(g62904_sb), .o(n_6069) );
na02s01 g64333_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_140), .b(FE_OFN917_n_4725), .o(g64333_db) );
na02s01 TIMEBOOST_cell_37459 ( .a(pci_target_unit_del_sync_addr_in_233), .b(n_2509), .o(TIMEBOOST_net_10968) );
in01s01 g64334_u0 ( .a(FE_OFN917_n_4725), .o(g64334_sb) );
na02s01 TIMEBOOST_cell_37458 ( .a(TIMEBOOST_net_10967), .b(FE_OFN775_n_15366), .o(TIMEBOOST_net_10567) );
na02s01 g64334_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_144), .b(FE_OFN917_n_4725), .o(g64334_db) );
na03s02 TIMEBOOST_cell_40673 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__Q), .b(n_4358), .c(FE_OFN1243_n_4092), .o(TIMEBOOST_net_12575) );
in01s01 g64335_u0 ( .a(FE_OFN917_n_4725), .o(g64335_sb) );
na02s02 TIMEBOOST_cell_40674 ( .a(TIMEBOOST_net_12575), .b(g62509_sb), .o(n_6561) );
na02s01 g64335_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_147), .b(FE_OFN916_n_4725), .o(g64335_db) );
in01s01 g64336_u0 ( .a(FE_OFN916_n_4725), .o(g64336_sb) );
na02s01 TIMEBOOST_cell_40530 ( .a(TIMEBOOST_net_12503), .b(FE_OFN1300_n_5763), .o(TIMEBOOST_net_11509) );
na02s01 g64336_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(FE_OFN916_n_4725), .o(g64336_db) );
in01s01 g64337_u0 ( .a(FE_OFN912_n_4727), .o(g64337_sb) );
na02s01 TIMEBOOST_cell_17958 ( .a(n_4488), .b(FE_OFN1676_n_4655), .o(TIMEBOOST_net_4236) );
na02s01 g64337_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_151), .b(FE_OFN912_n_4727), .o(g64337_db) );
na02s01 TIMEBOOST_cell_17959 ( .a(TIMEBOOST_net_4236), .b(g65347_da), .o(n_4259) );
oa12s01 g64338_u0 ( .a(n_3797), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_3__270), .c(n_4725), .o(n_4726) );
in01s01 g64339_u0 ( .a(FE_OFN1057_n_4727), .o(g64339_sb) );
na02f02 TIMEBOOST_cell_42252 ( .a(TIMEBOOST_net_13364), .b(FE_OFN1399_n_8567), .o(TIMEBOOST_net_12322) );
na02s01 g64339_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_150), .b(FE_OFN1057_n_4727), .o(g64339_db) );
na02s02 TIMEBOOST_cell_40038 ( .a(TIMEBOOST_net_12257), .b(g62574_sb), .o(n_6405) );
in01s01 g64340_u0 ( .a(FE_OFN918_n_4725), .o(g64340_sb) );
na02s01 g64340_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__Q), .b(g64340_sb), .o(g64340_da) );
na02s01 g64340_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(FE_OFN918_n_4725), .o(g64340_db) );
na02s02 TIMEBOOST_cell_45072 ( .a(TIMEBOOST_net_14774), .b(FE_OFN1635_n_9531), .o(TIMEBOOST_net_11170) );
in01s01 g64341_u0 ( .a(FE_OFN1056_n_4727), .o(g64341_sb) );
na02s02 TIMEBOOST_cell_45167 ( .a(n_4383), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__Q), .o(TIMEBOOST_net_14822) );
na02s01 g64341_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_144), .b(FE_OFN1056_n_4727), .o(g64341_db) );
na03s02 TIMEBOOST_cell_38363 ( .a(n_3942), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q), .c(FE_OFN2104_g64577_p), .o(TIMEBOOST_net_11420) );
in01s01 g64342_u0 ( .a(FE_OFN1056_n_4727), .o(g64342_sb) );
na02s01 TIMEBOOST_cell_18006 ( .a(pci_target_unit_fifos_pciw_addr_data_in_151), .b(g64082_sb), .o(TIMEBOOST_net_4260) );
na02s01 g64342_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_140), .b(FE_OFN1056_n_4727), .o(g64342_db) );
na02m02 TIMEBOOST_cell_44189 ( .a(n_9083), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q), .o(TIMEBOOST_net_14333) );
in01s01 g64343_u0 ( .a(FE_OFN918_n_4725), .o(g64343_sb) );
na02s01 g64343_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__Q), .b(g64343_sb), .o(g64343_da) );
na02s01 g64343_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_149), .b(FE_OFN918_n_4725), .o(g64343_db) );
na02s01 TIMEBOOST_cell_45073 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q), .b(FE_OFN1650_n_9428), .o(TIMEBOOST_net_14775) );
in01s01 g64344_u0 ( .a(FE_OFN917_n_4725), .o(g64344_sb) );
na02s01 TIMEBOOST_cell_44981 ( .a(g61962_sb), .b(g61984_db), .o(TIMEBOOST_net_14729) );
na02s01 g64344_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_142), .b(FE_OFN917_n_4725), .o(g64344_db) );
na02s02 TIMEBOOST_cell_40040 ( .a(TIMEBOOST_net_12258), .b(g62431_sb), .o(n_6735) );
in01s01 g64345_u0 ( .a(FE_OFN918_n_4725), .o(g64345_sb) );
na02s01 g64345_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__Q), .b(g64345_sb), .o(g64345_da) );
na02s01 g64345_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(FE_OFN918_n_4725), .o(g64345_db) );
na02s01 g64345_u3 ( .a(g64345_da), .b(g64345_db), .o(n_3833) );
in01s01 g64346_u0 ( .a(FE_OFN930_n_4730), .o(g64346_sb) );
na02f02 TIMEBOOST_cell_41114 ( .a(TIMEBOOST_net_12795), .b(g57499_sb), .o(n_11239) );
na02s01 g64346_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_149), .b(FE_OFN930_n_4730), .o(g64346_db) );
na02s02 TIMEBOOST_cell_45521 ( .a(TIMEBOOST_net_5436), .b(FE_OFN1312_n_6624), .o(TIMEBOOST_net_14999) );
in01s01 g64347_u0 ( .a(FE_OFN1055_n_4727), .o(g64347_sb) );
na02f02 TIMEBOOST_cell_38693 ( .a(TIMEBOOST_net_2028), .b(n_13127), .o(TIMEBOOST_net_11585) );
na02s01 g64347_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(FE_OFN1055_n_4727), .o(g64347_db) );
na02s02 TIMEBOOST_cell_38700 ( .a(TIMEBOOST_net_11588), .b(g62906_sb), .o(n_6065) );
in01s01 g64348_u0 ( .a(FE_OFN917_n_4725), .o(g64348_sb) );
na02s01 g64348_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__Q), .b(g64348_sb), .o(g64348_da) );
na02s01 g64348_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_143), .b(FE_OFN917_n_4725), .o(g64348_db) );
in01s01 g64349_u0 ( .a(FE_OFN1031_n_4732), .o(g64349_sb) );
na02s01 g64349_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__Q), .b(g64349_sb), .o(g64349_da) );
na02s01 g64349_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in), .b(FE_OFN1031_n_4732), .o(g64349_db) );
na03s02 TIMEBOOST_cell_38233 ( .a(TIMEBOOST_net_3685), .b(g64285_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__Q), .o(TIMEBOOST_net_11355) );
in01s01 g64350_u0 ( .a(FE_OFN930_n_4730), .o(g64350_sb) );
na02s01 g64350_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__Q), .b(g64350_sb), .o(g64350_da) );
na02s01 g64350_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_146), .b(FE_OFN930_n_4730), .o(g64350_db) );
na02s02 TIMEBOOST_cell_38725 ( .a(n_1845), .b(g61864_sb), .o(TIMEBOOST_net_11601) );
in01s01 g64351_u0 ( .a(FE_OFN917_n_4725), .o(g64351_sb) );
na02s02 TIMEBOOST_cell_45212 ( .a(TIMEBOOST_net_14844), .b(FE_OFN1244_n_4092), .o(TIMEBOOST_net_12121) );
na02s01 TIMEBOOST_cell_17518 ( .a(pci_target_unit_fifos_pciw_addr_data_in_141), .b(g64217_sb), .o(TIMEBOOST_net_4016) );
na02m02 TIMEBOOST_cell_40042 ( .a(TIMEBOOST_net_12259), .b(g58622_db), .o(n_8854) );
in01s01 g64352_u0 ( .a(FE_OFN918_n_4725), .o(g64352_sb) );
na02s01 g64352_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__Q), .b(g64352_sb), .o(g64352_da) );
na02s01 g64352_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(FE_OFN918_n_4725), .o(g64352_db) );
na02s01 TIMEBOOST_cell_45105 ( .a(n_2199), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__Q), .o(TIMEBOOST_net_14791) );
in01s01 g64353_u0 ( .a(FE_OFN916_n_4725), .o(g64353_sb) );
no02f06 TIMEBOOST_cell_40043 ( .a(FE_RN_153_0), .b(n_2250), .o(TIMEBOOST_net_12260) );
na02s01 g64353_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_128), .b(FE_OFN916_n_4725), .o(g64353_db) );
no02f06 TIMEBOOST_cell_40044 ( .a(TIMEBOOST_net_12260), .b(n_3466), .o(TIMEBOOST_net_5448) );
in01s01 g64354_u0 ( .a(FE_OFN918_n_4725), .o(g64354_sb) );
na02s01 g64354_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__Q), .b(g64354_sb), .o(g64354_da) );
na02s01 g64354_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_125), .b(FE_OFN918_n_4725), .o(g64354_db) );
na02m02 TIMEBOOST_cell_36264 ( .a(TIMEBOOST_net_10370), .b(n_3194), .o(TIMEBOOST_net_482) );
in01s01 g64355_u0 ( .a(FE_OFN916_n_4725), .o(g64355_sb) );
na02s01 TIMEBOOST_cell_40532 ( .a(TIMEBOOST_net_12504), .b(FE_OFN1301_n_5763), .o(TIMEBOOST_net_11507) );
na02s01 TIMEBOOST_cell_42643 ( .a(n_3739), .b(g64855_sb), .o(TIMEBOOST_net_13560) );
na02s01 TIMEBOOST_cell_9253 ( .a(TIMEBOOST_net_1193), .b(g65677_db), .o(n_2212) );
in01s01 g64356_u0 ( .a(FE_OFN916_n_4725), .o(g64356_sb) );
na02s01 g64356_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__Q), .b(g64356_sb), .o(g64356_da) );
na02s01 g64356_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in_152), .b(FE_OFN916_n_4725), .o(g64356_db) );
na02s02 TIMEBOOST_cell_45195 ( .a(n_4262), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__Q), .o(TIMEBOOST_net_14836) );
in01s01 g64357_u0 ( .a(FE_OFN918_n_4725), .o(g64357_sb) );
na02s01 TIMEBOOST_cell_16280 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__Q), .o(TIMEBOOST_net_3397) );
na02s01 g64357_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_124), .b(FE_OFN918_n_4725), .o(g64357_db) );
na02f02 TIMEBOOST_cell_40045 ( .a(n_9775), .b(g57148_sb), .o(TIMEBOOST_net_12261) );
in01s01 g64358_u0 ( .a(FE_OFN918_n_4725), .o(g64358_sb) );
na02s01 g64358_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__Q), .b(g64358_sb), .o(g64358_da) );
na02s01 g64358_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in), .b(FE_OFN918_n_4725), .o(g64358_db) );
na02s01 TIMEBOOST_cell_9196 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(g65772_sb), .o(TIMEBOOST_net_1165) );
in01s01 g64359_u0 ( .a(FE_OFN918_n_4725), .o(g64359_sb) );
na02s01 TIMEBOOST_cell_44982 ( .a(TIMEBOOST_net_14729), .b(g63607_db), .o(TIMEBOOST_net_13152) );
na02s01 g64359_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_123), .b(FE_OFN918_n_4725), .o(g64359_db) );
na02f02 TIMEBOOST_cell_40046 ( .a(TIMEBOOST_net_12261), .b(g57148_db), .o(n_11602) );
in01s01 g64360_u0 ( .a(FE_OFN916_n_4725), .o(g64360_sb) );
na02s01 TIMEBOOST_cell_40534 ( .a(TIMEBOOST_net_12505), .b(TIMEBOOST_net_9879), .o(n_13496) );
na02s01 g64360_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_151), .b(FE_OFN916_n_4725), .o(g64360_db) );
na02s01 TIMEBOOST_cell_16286 ( .a(wishbone_slave_unit_pci_initiator_if_data_source), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_3400) );
in01s01 g64361_u0 ( .a(FE_OFN918_n_4725), .o(g64361_sb) );
na02s01 TIMEBOOST_cell_16287 ( .a(TIMEBOOST_net_3400), .b(g53940_sb), .o(TIMEBOOST_net_829) );
na02s01 g64361_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_127), .b(FE_OFN918_n_4725), .o(g64361_db) );
na02f02 TIMEBOOST_cell_40047 ( .a(n_9759), .b(g57160_sb), .o(TIMEBOOST_net_12262) );
in01s01 g64362_u0 ( .a(FE_OFN918_n_4725), .o(g64362_sb) );
na02f02 TIMEBOOST_cell_40048 ( .a(TIMEBOOST_net_12262), .b(g57160_db), .o(n_11589) );
na02s01 g64362_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_150), .b(FE_OFN918_n_4725), .o(g64362_db) );
na03s02 TIMEBOOST_cell_16290 ( .a(n_2580), .b(n_2172), .c(n_1848), .o(TIMEBOOST_net_3402) );
in01s01 g64363_u0 ( .a(FE_OFN916_n_4725), .o(g64363_sb) );
na02s02 TIMEBOOST_cell_16291 ( .a(TIMEBOOST_net_3402), .b(n_2377), .o(n_3298) );
na02s01 g64363_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(FE_OFN916_n_4725), .o(g64363_db) );
na02f02 TIMEBOOST_cell_40049 ( .a(n_9746), .b(g57178_sb), .o(TIMEBOOST_net_12263) );
oa12s01 g64364_u0 ( .a(n_3808), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_0__153), .c(FE_OFN1059_n_4727), .o(n_4722) );
na02s02 TIMEBOOST_cell_10581 ( .a(TIMEBOOST_net_1857), .b(g65400_db), .o(n_4237) );
na02s02 TIMEBOOST_cell_45522 ( .a(TIMEBOOST_net_14999), .b(g62673_sb), .o(n_6193) );
na02s01 TIMEBOOST_cell_39196 ( .a(TIMEBOOST_net_11836), .b(g65710_sb), .o(n_1907) );
in01s01 g64366_u0 ( .a(FE_OFN1033_n_4732), .o(g64366_sb) );
na02s01 g64366_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__Q), .b(g64366_sb), .o(g64366_da) );
na02s01 g64366_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_125), .b(FE_OFN1033_n_4732), .o(g64366_db) );
na02s01 g64366_u3 ( .a(g64366_da), .b(g64366_db), .o(n_3814) );
in01s01 g64367_u0 ( .a(FE_OFN918_n_4725), .o(g64367_sb) );
na02s01 g64367_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__Q), .b(g64367_sb), .o(g64367_da) );
na02s01 g64367_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_146), .b(FE_OFN918_n_4725), .o(g64367_db) );
na02s02 TIMEBOOST_cell_45106 ( .a(TIMEBOOST_net_14791), .b(FE_OFN1812_n_7845), .o(TIMEBOOST_net_11388) );
no02s01 g64368_u0 ( .a(wbu_addr_in_260), .b(n_2694), .o(g64368_p) );
ao12s02 g64368_u1 ( .a(g64368_p), .b(wbu_addr_in_260), .c(n_2694), .o(n_2695) );
no02s01 g64369_u0 ( .a(n_2419), .b(wbm_adr_o_11_), .o(g64369_p) );
ao12m01 g64369_u1 ( .a(g64369_p), .b(wbm_adr_o_11_), .c(n_2419), .o(n_2693) );
no02s02 g64370_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_9_), .b(n_1633), .o(g64370_p) );
ao12s02 g64370_u1 ( .a(g64370_p), .b(pci_target_unit_del_sync_comp_cycle_count_9_), .c(n_1633), .o(n_2423) );
no02s02 g64371_u0 ( .a(n_1992), .b(n_1631), .o(g64371_p) );
ao12s02 g64371_u1 ( .a(g64371_p), .b(n_1992), .c(n_1631), .o(n_2422) );
in01s01 g64372_u0 ( .a(n_1669), .o(n_1463) );
in01s01 g64373_u0 ( .a(n_1438), .o(n_1190) );
in01s01 g64374_u0 ( .a(n_1476), .o(n_1213) );
no02m01 g64375_u0 ( .a(n_2691), .b(conf_wb_err_addr_in_952), .o(g64375_p) );
ao12m01 g64375_u1 ( .a(g64375_p), .b(conf_wb_err_addr_in_952), .c(n_2691), .o(n_2692) );
no02s01 g64376_u0 ( .a(conf_wb_err_addr_in_949), .b(n_2260), .o(g64376_p) );
ao12s01 g64376_u1 ( .a(g64376_p), .b(conf_wb_err_addr_in_949), .c(n_2260), .o(n_2261) );
no02s01 g64377_u0 ( .a(wbm_adr_o_8_), .b(n_2258), .o(g64377_p) );
ao12s01 g64377_u1 ( .a(g64377_p), .b(wbm_adr_o_8_), .c(n_2258), .o(n_2259) );
no02s01 g64378_u0 ( .a(wbu_addr_in_257), .b(n_2256), .o(g64378_p) );
ao12s01 g64378_u1 ( .a(g64378_p), .b(wbu_addr_in_257), .c(n_2256), .o(n_2257) );
no02f02 g64379_u0 ( .a(n_1396), .b(n_1395), .o(g64379_p) );
ao12f02 g64379_u1 ( .a(g64379_p), .b(n_1396), .c(n_1395), .o(n_2255) );
no02f02 g64380_u0 ( .a(n_1393), .b(n_1404), .o(g64380_p) );
ao12f02 g64380_u1 ( .a(g64380_p), .b(n_1393), .c(n_1404), .o(n_2254) );
na02s01 TIMEBOOST_cell_17208 ( .a(pci_target_unit_fifos_pcir_data_in_187), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__Q), .o(TIMEBOOST_net_3861) );
no02f02 g64382_u0 ( .a(n_1400), .b(n_1398), .o(g64382_p) );
ao12f02 g64382_u1 ( .a(g64382_p), .b(n_1400), .c(n_1398), .o(n_2252) );
no02f03 g64383_u0 ( .a(n_1449), .b(n_1405), .o(g64383_p) );
ao12f02 g64383_u1 ( .a(g64383_p), .b(n_1449), .c(n_1405), .o(n_2251) );
no02f02 g64384_u0 ( .a(n_1402), .b(n_1401), .o(g64384_p) );
ao12f04 g64384_u1 ( .a(g64384_p), .b(n_1402), .c(n_1401), .o(n_2250) );
no02f02 g64385_u0 ( .a(n_1394), .b(n_1439), .o(g64385_p) );
ao12f02 g64385_u1 ( .a(g64385_p), .b(n_1394), .c(n_1439), .o(n_2249) );
na02s04 g64450_u0 ( .a(n_2219), .b(pci_gnt_i), .o(n_3126) );
na02s02 TIMEBOOST_cell_45686 ( .a(TIMEBOOST_net_15081), .b(FE_OFN1214_n_4151), .o(TIMEBOOST_net_12604) );
na02f02 g64452_u0 ( .a(n_3290), .b(pciu_bar0_in_364), .o(n_3292) );
na02s01 g64454_u0 ( .a(n_4718), .b(n_3314), .o(g64454_p) );
in01s01 g64454_u1 ( .a(g64454_p), .o(n_3289) );
na02s01 TIMEBOOST_cell_37265 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__Q), .b(n_3747), .o(TIMEBOOST_net_10871) );
na02s01 g64456_u0 ( .a(n_4512), .b(n_4669), .o(n_4514) );
na02s02 TIMEBOOST_cell_37171 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_413), .b(wishbone_slave_unit_del_sync_addr_out_reg_30__Q), .o(TIMEBOOST_net_10824) );
na02s02 TIMEBOOST_cell_38590 ( .a(TIMEBOOST_net_11533), .b(g60643_sb), .o(n_5686) );
no02s01 g64459_u0 ( .a(n_2726), .b(n_3023), .o(n_3812) );
na02s01 g64460_u0 ( .a(n_4512), .b(n_4677), .o(n_4513) );
no02s01 g64461_u0 ( .a(n_1621), .b(n_2248), .o(g64461_p) );
in01s01 g64461_u1 ( .a(g64461_p), .o(n_7835) );
na02s01 g64462_u0 ( .a(n_4512), .b(FE_OFN1678_n_4655), .o(n_4511) );
na02s01 g64463_u0 ( .a(n_4512), .b(FE_OFN1640_n_4671), .o(n_4510) );
no02f06 g64464_u0 ( .a(n_15324), .b(n_2308), .o(n_2897) );
no02f02 g64465_u0 ( .a(n_3016), .b(n_2449), .o(g64465_p) );
in01f02 g64465_u1 ( .a(g64465_p), .o(n_3390) );
no02s01 g64466_u0 ( .a(n_1623), .b(n_4725), .o(g64466_p) );
in01s01 g64466_u1 ( .a(g64466_p), .o(n_2247) );
na02f02 g64467_u0 ( .a(n_3290), .b(pciu_bar0_in_378), .o(n_3285) );
na02f06 g64577_u0 ( .a(n_2399), .b(pci_target_unit_fifos_pciw_wenable_in), .o(g64577_p) );
na02m04 g64578_u0 ( .a(n_2691), .b(n_1482), .o(g64578_p) );
in01m02 g64578_u1 ( .a(g64578_p), .o(n_3130) );
na02s02 TIMEBOOST_cell_38592 ( .a(TIMEBOOST_net_11534), .b(g60646_sb), .o(n_5681) );
na02s01 g64580_u0 ( .a(n_4512), .b(FE_OFN651_n_4508), .o(n_4509) );
na02m04 g64581_u0 ( .a(n_2260), .b(n_1388), .o(g64581_p) );
in01m04 g64581_u1 ( .a(g64581_p), .o(n_2722) );
na02s02 g64582_u0 ( .a(n_1437), .b(pci_target_unit_wishbone_master_rty_counter_3_), .o(g64582_p) );
in01s02 g64582_u1 ( .a(g64582_p), .o(n_1273) );
na02f04 g64583_u0 ( .a(n_3023), .b(FE_OFN2121_n_2687), .o(n_6986) );
in01s01 g64584_u0 ( .a(n_3313), .o(n_2888) );
na02f06 g64585_u0 ( .a(n_4718), .b(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(g64585_p) );
in01f04 g64585_u1 ( .a(g64585_p), .o(n_3313) );
na02s02 TIMEBOOST_cell_43645 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__Q), .b(n_3601), .o(TIMEBOOST_net_14061) );
no02m02 g64587_u0 ( .a(FE_OFN2100_n_3281), .b(n_3280), .o(g64587_p) );
in01m02 g64587_u1 ( .a(g64587_p), .o(n_3282) );
in01s01 g64588_u0 ( .a(n_2245), .o(n_2246) );
no02m06 g64589_u0 ( .a(n_3395), .b(FE_OFN999_n_15978), .o(n_2245) );
na02m02 g64590_u0 ( .a(n_3089), .b(n_2308), .o(n_3090) );
no02s01 g64591_u0 ( .a(n_3388), .b(n_3275), .o(n_3389) );
no02s01 g64592_u0 ( .a(n_3388), .b(n_3265), .o(n_3387) );
no02s01 g64593_u0 ( .a(n_3278), .b(n_3277), .o(n_3279) );
na02m02 g64595_u0 ( .a(n_4718), .b(n_2685), .o(g64595_p) );
in01f02 g64595_u1 ( .a(g64595_p), .o(n_3119) );
na02f02 g64596_u0 ( .a(n_1282), .b(n_2256), .o(g64596_p) );
in01f02 g64596_u1 ( .a(g64596_p), .o(n_2437) );
na02m04 g64597_u0 ( .a(n_2419), .b(n_1373), .o(g64597_p) );
in01m04 g64597_u1 ( .a(g64597_p), .o(n_2931) );
oa12s01 g64598_u0 ( .a(n_2406), .b(n_990), .c(n_691), .o(n_2418) );
na02s01 g64599_u0 ( .a(n_3810), .b(n_4084), .o(n_3811) );
na02f02 TIMEBOOST_cell_40050 ( .a(TIMEBOOST_net_12263), .b(g57178_db), .o(n_11577) );
no02s01 g64601_u0 ( .a(n_3278), .b(n_3275), .o(n_3276) );
no02f03 g64602_u0 ( .a(pci_target_unit_pci_target_sm_state_transfere_reg), .b(n_532), .o(n_2887) );
in01s01 g64603_u0 ( .a(n_4533), .o(n_3809) );
na02f02 TIMEBOOST_cell_41054 ( .a(TIMEBOOST_net_12765), .b(g57302_sb), .o(n_10407) );
na02s01 g64605_u0 ( .a(FE_OFN1059_n_4727), .b(n_3806), .o(n_3808) );
no02s01 g64606_u0 ( .a(n_3386), .b(n_3395), .o(n_3385) );
no02s01 g64607_u0 ( .a(n_3388), .b(n_3273), .o(n_3384) );
no02s01 g64608_u0 ( .a(n_3278), .b(n_3273), .o(n_3274) );
na02s01 g64609_u0 ( .a(n_4730), .b(n_3806), .o(n_3807) );
no02f01 g64610_u0 ( .a(n_13820), .b(n_2415), .o(g64610_p) );
in01m02 g64610_u1 ( .a(g64610_p), .o(n_2416) );
na02s01 g64611_u0 ( .a(FE_OFN1036_n_4732), .b(n_3806), .o(n_3805) );
na02m02 TIMEBOOST_cell_42205 ( .a(n_9798), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__Q), .o(TIMEBOOST_net_13341) );
na02m02 TIMEBOOST_cell_44263 ( .a(n_9840), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__Q), .o(TIMEBOOST_net_14370) );
na02s01 TIMEBOOST_cell_42769 ( .a(FE_OFN252_n_9868), .b(g57944_sb), .o(TIMEBOOST_net_13623) );
in01s01 g64630_u3 ( .a(g64630_p), .o(n_1995) );
na02s02 g64631_u0 ( .a(n_3089), .b(n_2742), .o(g64631_p) );
in01s02 g64631_u1 ( .a(g64631_p), .o(n_3271) );
no02s01 g64632_u0 ( .a(n_3798), .b(n_2464), .o(g64632_p) );
in01s01 g64632_u1 ( .a(g64632_p), .o(n_3800) );
na02f04 g64633_u0 ( .a(n_2694), .b(n_1479), .o(g64633_p) );
in01f04 g64633_u1 ( .a(g64633_p), .o(n_3132) );
na02m02 TIMEBOOST_cell_42155 ( .a(n_9571), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__Q), .o(TIMEBOOST_net_13316) );
no02s02 g64639_u0 ( .a(n_3278), .b(n_3030), .o(g64639_p) );
in01s02 g64639_u1 ( .a(g64639_p), .o(n_4630) );
na02f02 TIMEBOOST_cell_40052 ( .a(TIMEBOOST_net_12264), .b(g57565_db), .o(n_11187) );
no02s02 g64641_u0 ( .a(n_3798), .b(n_2319), .o(n_3799) );
no02s02 g64642_u0 ( .a(n_4720), .b(n_3280), .o(n_4721) );
na02m02 g64643_u0 ( .a(n_2258), .b(n_1241), .o(g64643_p) );
in01m02 g64643_u1 ( .a(g64643_p), .o(n_2441) );
no02f10 g64644_u0 ( .a(n_842), .b(n_938), .o(n_1434) );
no02s02 g64645_u0 ( .a(n_1987), .b(n_1974), .o(n_2414) );
no02s01 g64646_u0 ( .a(n_4718), .b(n_691), .o(g64646_p) );
in01s01 g64646_u1 ( .a(g64646_p), .o(n_3087) );
na02s01 g64647_u0 ( .a(n_4725), .b(n_3806), .o(n_3797) );
na02s01 g64648_u0 ( .a(n_2799), .b(n_12179), .o(n_3269) );
na02s01 g64649_u0 ( .a(n_3267), .b(n_2966), .o(n_3268) );
no02f08 g64650_u0 ( .a(n_3395), .b(n_1514), .o(n_2443) );
no02s01 g64651_u0 ( .a(n_3278), .b(n_3265), .o(n_3266) );
no02s01 g64652_u0 ( .a(n_3388), .b(n_3277), .o(n_3381) );
in01f06 g64667_u0 ( .a(n_15260), .o(n_13249) );
na02s02 g64670_u0 ( .a(n_1961), .b(n_2337), .o(n_4152) );
no02s02 g64671_u0 ( .a(n_3388), .b(n_3030), .o(g64671_p) );
in01s02 g64671_u1 ( .a(g64671_p), .o(n_4783) );
in01s01 g64676_u0 ( .a(n_2727), .o(n_2412) );
ao12f04 g64677_u0 ( .a(n_1588), .b(n_1211), .c(n_545), .o(n_2727) );
na02s02 g64678_u0 ( .a(n_3795), .b(n_1533), .o(g64678_p) );
in01s01 g64678_u1 ( .a(g64678_p), .o(n_3796) );
na02f02 TIMEBOOST_cell_40054 ( .a(TIMEBOOST_net_12265), .b(g57571_sb), .o(n_11180) );
na02f02 TIMEBOOST_cell_42206 ( .a(TIMEBOOST_net_13341), .b(FE_OFN1419_n_8567), .o(TIMEBOOST_net_12279) );
na02s03 TIMEBOOST_cell_45778 ( .a(TIMEBOOST_net_15127), .b(g62520_sb), .o(n_6536) );
na02s02 TIMEBOOST_cell_45687 ( .a(n_4243), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__Q), .o(TIMEBOOST_net_15082) );
na02s02 TIMEBOOST_cell_43535 ( .a(n_27), .b(n_3641), .o(TIMEBOOST_net_14006) );
na02f04 TIMEBOOST_cell_39034 ( .a(TIMEBOOST_net_11755), .b(FE_OFN2243_g52675_p), .o(TIMEBOOST_net_10744) );
ao12s01 g64685_u0 ( .a(pci_target_unit_del_sync_req_comp_pending), .b(pci_target_unit_del_sync_req_rty_exp_reg), .c(pci_target_unit_del_sync_req_rty_exp_clr), .o(n_646) );
no02s01 g64687_u0 ( .a(n_2070), .b(n_3261), .o(g64687_p) );
in01s01 g64687_u1 ( .a(g64687_p), .o(n_3262) );
na02s02 TIMEBOOST_cell_42092 ( .a(TIMEBOOST_net_13284), .b(FE_OFN1230_n_6391), .o(TIMEBOOST_net_11568) );
ao12s01 g64689_u0 ( .a(n_152), .b(n_2765), .c(output_backup_trdy_out_reg_Q), .o(n_3380) );
na02s01 g64694_u0 ( .a(n_2303), .b(n_4718), .o(g64694_p) );
in01s01 g64694_u1 ( .a(g64694_p), .o(n_3081) );
oa12s01 g64695_u0 ( .a(n_2803), .b(n_15762), .c(n_3022), .o(n_2900) );
na02f01 g64696_u0 ( .a(n_2805), .b(FE_OFN2121_n_2687), .o(n_3260) );
na02s01 g64697_u0 ( .a(n_3481), .b(n_4718), .o(g64697_p) );
in01s01 g64697_u1 ( .a(g64697_p), .o(n_4719) );
ao22f02 g64698_u0 ( .a(n_2555), .b(n_14909), .c(n_2358), .d(n_2331), .o(n_3259) );
ao12s01 g64699_u0 ( .a(n_2086), .b(n_3123), .c(n_1554), .o(n_2878) );
na02s02 g64700_u0 ( .a(n_2065), .b(FE_OFN197_n_2683), .o(g64700_p) );
in01s01 g64700_u1 ( .a(g64700_p), .o(n_2684) );
no02s01 g64701_u0 ( .a(n_2072), .b(n_3261), .o(g64701_p) );
in01s01 g64701_u1 ( .a(g64701_p), .o(n_3258) );
no02s01 g64702_u0 ( .a(n_3261), .b(n_2068), .o(g64702_p) );
in01s01 g64702_u1 ( .a(g64702_p), .o(n_3257) );
ao12s01 g64703_u0 ( .a(n_2409), .b(n_8498), .c(pci_target_unit_pcit_if_req_req_pending_in), .o(n_2410) );
no02s01 g64704_u0 ( .a(n_3261), .b(n_8540), .o(g64704_p) );
in01s01 g64704_u1 ( .a(g64704_p), .o(n_3256) );
no02s01 g64705_u0 ( .a(n_2080), .b(n_3261), .o(g64705_p) );
in01s01 g64705_u1 ( .a(g64705_p), .o(n_3255) );
ao12s01 g64706_u0 ( .a(n_1659), .b(wishbone_slave_unit_pci_initiator_if_read_count_2_), .c(n_660), .o(n_1660) );
na02f02 g64707_u0 ( .a(n_3163), .b(n_3378), .o(g64707_p) );
in01f02 g64707_u1 ( .a(g64707_p), .o(n_3379) );
no02s02 g64708_u0 ( .a(n_1832), .b(n_1834), .o(n_8564) );
ao12s01 g64709_u0 ( .a(n_1178), .b(n_1011), .c(wishbone_slave_unit_pci_initiator_sm_latency_timer_2_), .o(n_1658) );
in01s01 g64710_u0 ( .a(n_2682), .o(n_2877) );
ao12s01 g64711_u0 ( .a(wishbone_slave_unit_del_sync_req_comp_pending), .b(wishbone_slave_unit_del_sync_req_rty_exp_reg), .c(wishbone_slave_unit_del_sync_req_rty_exp_clr), .o(n_2682) );
no02s01 g64712_u0 ( .a(n_2079), .b(n_3261), .o(g64712_p) );
in01s01 g64712_u1 ( .a(g64712_p), .o(n_3254) );
oa12s01 g64714_u0 ( .a(n_2406), .b(wishbone_slave_unit_pci_initiator_if_read_count_0_), .c(n_691), .o(n_2407) );
oa12s02 g64715_u0 ( .a(n_2406), .b(n_292), .c(n_692), .o(n_2405) );
ao12s01 g64716_u0 ( .a(n_2049), .b(wbu_cache_line_size_in_206), .c(n_691), .o(n_2234) );
na02s02 TIMEBOOST_cell_21951 ( .a(TIMEBOOST_net_6232), .b(n_10106), .o(n_11858) );
na02f02 TIMEBOOST_cell_44264 ( .a(TIMEBOOST_net_14370), .b(FE_OFN1414_n_8567), .o(TIMEBOOST_net_12754) );
na02s02 TIMEBOOST_cell_43536 ( .a(TIMEBOOST_net_14006), .b(FE_OFN1310_n_6624), .o(TIMEBOOST_net_12677) );
in01s01 TIMEBOOST_cell_45869 ( .a(n_11869), .o(TIMEBOOST_net_15176) );
in01s01 TIMEBOOST_cell_45870 ( .a(TIMEBOOST_net_15176), .o(TIMEBOOST_net_15177) );
na03s02 TIMEBOOST_cell_5783 ( .a(n_3774), .b(g64927_sb), .c(g64927_db), .o(n_3681) );
na02m02 TIMEBOOST_cell_42207 ( .a(n_8999), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__34__Q), .o(TIMEBOOST_net_13342) );
na02s01 TIMEBOOST_cell_41694 ( .a(TIMEBOOST_net_13085), .b(FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_1009) );
na02f04 g64727_u0 ( .a(n_2399), .b(n_1976), .o(g64727_p) );
in01f02 g64727_u1 ( .a(g64727_p), .o(n_3335) );
oa22s03 g64728_u0 ( .a(n_1809), .b(n_16168), .c(n_16160), .d(n_3250), .o(n_5751) );
ao12f01 g64729_u0 ( .a(n_3026), .b(n_16000), .c(n_3078), .o(n_3079) );
na02f02 TIMEBOOST_cell_45756 ( .a(TIMEBOOST_net_15116), .b(FE_OCPN1845_n_16427), .o(TIMEBOOST_net_632) );
na02f02 TIMEBOOST_cell_42208 ( .a(TIMEBOOST_net_13342), .b(FE_OFN1391_n_8567), .o(TIMEBOOST_net_12294) );
na02m02 TIMEBOOST_cell_45779 ( .a(n_3350), .b(TIMEBOOST_net_589), .o(TIMEBOOST_net_15128) );
na02s01 TIMEBOOST_cell_43326 ( .a(TIMEBOOST_net_13901), .b(g62605_sb), .o(n_6342) );
na02m02 TIMEBOOST_cell_43537 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__Q), .b(n_3626), .o(TIMEBOOST_net_14007) );
ao22f02 g64735_u0 ( .a(n_2339), .b(n_14910), .c(configuration_wb_err_data_572), .d(FE_OFN1071_n_15729), .o(n_3077) );
no02s01 g64736_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_5_), .b(n_1425), .o(g64736_p) );
ao12s01 g64736_u1 ( .a(g64736_p), .b(pci_target_unit_del_sync_comp_cycle_count_5_), .c(n_1425), .o(n_1701) );
ao22s01 g64738_u0 ( .a(n_547), .b(wishbone_slave_unit_pci_initiator_sm_decode_count_2_), .c(n_401), .d(n_1471), .o(n_1472) );
ao12s01 g64739_u0 ( .a(n_2806), .b(pci_target_unit_wishbone_master_read_count_1_), .c(n_3250), .o(n_3251) );
no02m01 g64740_u0 ( .a(n_1469), .b(pci_target_unit_wishbone_master_rty_counter_5_), .o(g64740_p) );
ao12m01 g64740_u1 ( .a(g64740_p), .b(pci_target_unit_wishbone_master_rty_counter_5_), .c(n_1469), .o(n_2291) );
oa12m01 g64741_u0 ( .a(n_2002), .b(n_2001), .c(pci_target_unit_wishbone_master_rty_counter_6_), .o(n_2396) );
ao22f02 g64742_u0 ( .a(configuration_isr_bit_631), .b(n_3246), .c(n_3248), .d(configuration_sync_command_bit0), .o(n_15436) );
in01s01 g64743_u0 ( .a(n_3377), .o(n_3794) );
na02f02 TIMEBOOST_cell_22425 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_6469), .o(TIMEBOOST_net_3084) );
ao22f02 g64745_u0 ( .a(configuration_command_bit), .b(n_3248), .c(n_3246), .d(configuration_isr_bit_618), .o(n_3247) );
no02s01 g64746_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_5_), .b(n_1426), .o(g64746_p) );
ao12s01 g64746_u1 ( .a(g64746_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_5_), .c(n_1426), .o(n_1656) );
no02f06 g64747_u0 ( .a(n_1279), .b(n_1081), .o(g64747_p) );
ao12f04 g64747_u1 ( .a(g64747_p), .b(n_1081), .c(n_1279), .o(n_2227) );
in01s01 g64748_u0 ( .a(FE_OFN672_n_4505), .o(g64748_sb) );
na02s01 TIMEBOOST_cell_31400 ( .a(g65023_sb), .b(g65023_db), .o(TIMEBOOST_net_9611) );
na02s01 g64748_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__Q), .b(FE_OFN672_n_4505), .o(g64748_db) );
na02s01 TIMEBOOST_cell_16370 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(g65673_sb), .o(TIMEBOOST_net_3442) );
in01s01 g64749_u0 ( .a(FE_OFN682_n_4460), .o(g64749_sb) );
na02f02 TIMEBOOST_cell_40056 ( .a(TIMEBOOST_net_12266), .b(g57219_sb), .o(n_11536) );
na02f02 TIMEBOOST_cell_44090 ( .a(TIMEBOOST_net_14283), .b(FE_OFN1390_n_8567), .o(TIMEBOOST_net_12909) );
na02s02 TIMEBOOST_cell_40057 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_767), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_2__Q), .o(TIMEBOOST_net_12267) );
in01s01 g64750_u0 ( .a(FE_OFN671_n_4505), .o(g64750_sb) );
na02s02 TIMEBOOST_cell_37772 ( .a(TIMEBOOST_net_11124), .b(g61921_sb), .o(n_7979) );
na02s01 TIMEBOOST_cell_40835 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__Q), .b(n_13548), .o(TIMEBOOST_net_12656) );
na02s02 TIMEBOOST_cell_37774 ( .a(TIMEBOOST_net_11125), .b(g61948_sb), .o(n_7929) );
in01s01 g64751_u0 ( .a(FE_OFN614_n_4501), .o(g64751_sb) );
na02s01 TIMEBOOST_cell_42763 ( .a(g63545_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__Q), .o(TIMEBOOST_net_13620) );
na02s01 g64751_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__Q), .b(FE_OFN614_n_4501), .o(g64751_db) );
in01s01 g64752_u0 ( .a(FE_OFN678_n_4460), .o(g64752_sb) );
na02m02 TIMEBOOST_cell_40058 ( .a(TIMEBOOST_net_12267), .b(FE_OFN1305_n_13124), .o(TIMEBOOST_net_11635) );
na02m02 TIMEBOOST_cell_44452 ( .a(TIMEBOOST_net_14464), .b(g54244_sb), .o(n_13146) );
na02s01 TIMEBOOST_cell_45074 ( .a(TIMEBOOST_net_14775), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_11154) );
in01s01 g64753_u0 ( .a(FE_OFN618_n_4490), .o(g64753_sb) );
na03f02 TIMEBOOST_cell_8628 ( .a(FE_OFN1602_n_13995), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__Q), .c(n_13949), .o(g53268_p) );
na02s01 g64753_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__30__Q), .b(FE_OFN618_n_4490), .o(g64753_db) );
na02s01 TIMEBOOST_cell_42625 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__Q), .b(FE_OFN1795_n_9904), .o(TIMEBOOST_net_13551) );
in01s01 g64754_u0 ( .a(FE_OFN672_n_4505), .o(g64754_sb) );
na02s02 TIMEBOOST_cell_40740 ( .a(TIMEBOOST_net_12608), .b(g62490_sb), .o(n_6605) );
na02s01 g64754_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__Q), .b(FE_OFN672_n_4505), .o(g64754_db) );
na03s02 TIMEBOOST_cell_43327 ( .a(n_3650), .b(FE_OFN1222_n_6391), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__Q), .o(TIMEBOOST_net_13902) );
in01s01 g64755_u0 ( .a(FE_OFN671_n_4505), .o(g64755_sb) );
na02s02 TIMEBOOST_cell_43461 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__Q), .b(n_3707), .o(TIMEBOOST_net_13969) );
na02s01 g64755_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__13__Q), .b(FE_OFN671_n_4505), .o(g64755_db) );
na02s01 TIMEBOOST_cell_16371 ( .a(TIMEBOOST_net_3442), .b(g65673_db), .o(n_1958) );
in01s01 g64756_u0 ( .a(FE_OFN619_n_4490), .o(g64756_sb) );
na02s01 TIMEBOOST_cell_16669 ( .a(TIMEBOOST_net_3591), .b(g64168_db), .o(n_3997) );
na02s01 g64756_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__Q), .b(FE_OFN619_n_4490), .o(g64756_db) );
na03s02 TIMEBOOST_cell_42811 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__Q), .b(FE_OFN699_n_7845), .c(n_1837), .o(TIMEBOOST_net_13644) );
in01s01 g64757_u0 ( .a(FE_OFN646_n_4497), .o(g64757_sb) );
na02s02 TIMEBOOST_cell_45107 ( .a(TIMEBOOST_net_4364), .b(g54199_sb), .o(TIMEBOOST_net_14792) );
na02s01 g64757_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__Q), .b(FE_OFN646_n_4497), .o(g64757_db) );
na02f02 TIMEBOOST_cell_40060 ( .a(TIMEBOOST_net_12268), .b(g57382_sb), .o(n_11363) );
in01s01 g64758_u0 ( .a(FE_OFN667_n_4495), .o(g64758_sb) );
na02s02 TIMEBOOST_cell_43462 ( .a(TIMEBOOST_net_13969), .b(FE_OFN1232_n_6391), .o(TIMEBOOST_net_12202) );
na02s01 g64758_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__Q), .b(FE_OFN667_n_4495), .o(g64758_db) );
na02s01 TIMEBOOST_cell_31397 ( .a(TIMEBOOST_net_9609), .b(g65035_db), .o(n_3625) );
in01s01 g64759_u0 ( .a(FE_OFN670_n_4505), .o(g64759_sb) );
na02s01 TIMEBOOST_cell_42707 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__Q), .b(g65952_sb), .o(TIMEBOOST_net_13592) );
na02s01 g64759_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q), .b(FE_OFN670_n_4505), .o(g64759_db) );
na02s01 TIMEBOOST_cell_38616 ( .a(TIMEBOOST_net_11546), .b(g63189_sb), .o(n_5776) );
in01s01 g64760_u0 ( .a(FE_OFN1806_n_4501), .o(g64760_sb) );
na02s01 TIMEBOOST_cell_45044 ( .a(TIMEBOOST_net_14760), .b(FE_OFN720_n_8060), .o(TIMEBOOST_net_11253) );
na02s01 g64760_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__Q), .b(FE_OFN1806_n_4501), .o(g64760_db) );
na02s02 TIMEBOOST_cell_38511 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__Q), .b(g58359_sb), .o(TIMEBOOST_net_11494) );
in01s01 g64761_u0 ( .a(FE_OFN669_n_4505), .o(g64761_sb) );
na02s01 TIMEBOOST_cell_31396 ( .a(n_3770), .b(g65035_sb), .o(TIMEBOOST_net_9609) );
na02s01 g64761_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__Q), .b(FE_OFN669_n_4505), .o(g64761_db) );
na02s01 TIMEBOOST_cell_40531 ( .a(wishbone_slave_unit_pcim_sm_data_in_641), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__Q), .o(TIMEBOOST_net_12504) );
in01s01 g64762_u0 ( .a(FE_OFN1663_n_4490), .o(g64762_sb) );
na02s01 TIMEBOOST_cell_31200 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__Q), .b(pci_target_unit_fifos_pcir_data_in_170), .o(TIMEBOOST_net_9511) );
na02s01 g64762_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__Q), .b(FE_OFN1663_n_4490), .o(g64762_db) );
na02s02 TIMEBOOST_cell_45730 ( .a(TIMEBOOST_net_15103), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_13264) );
in01s01 g64763_u0 ( .a(FE_OFN1806_n_4501), .o(g64763_sb) );
na02s01 TIMEBOOST_cell_39275 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q), .b(g64298_sb), .o(TIMEBOOST_net_11876) );
na02s01 g64763_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__Q), .b(FE_OFN1806_n_4501), .o(g64763_db) );
na02s01 TIMEBOOST_cell_39276 ( .a(TIMEBOOST_net_11876), .b(g64298_db), .o(n_3876) );
in01s01 g64764_u0 ( .a(FE_OFN1659_n_4490), .o(g64764_sb) );
na02s01 TIMEBOOST_cell_31198 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__Q), .b(pci_target_unit_fifos_pcir_data_in), .o(TIMEBOOST_net_9510) );
na02m02 TIMEBOOST_cell_44091 ( .a(n_9421), .b(n_15567), .o(TIMEBOOST_net_14284) );
na02m02 TIMEBOOST_cell_44323 ( .a(n_9416), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__Q), .o(TIMEBOOST_net_14400) );
in01s01 g64765_u0 ( .a(FE_OFN1660_n_4490), .o(g64765_sb) );
na02s01 TIMEBOOST_cell_42977 ( .a(TIMEBOOST_net_4245), .b(g64205_db), .o(TIMEBOOST_net_13727) );
na02s02 TIMEBOOST_cell_18129 ( .a(TIMEBOOST_net_4321), .b(g58281_sb), .o(n_9521) );
in01s01 g64766_u0 ( .a(FE_OFN666_n_4495), .o(g64766_sb) );
na02s01 TIMEBOOST_cell_16739 ( .a(TIMEBOOST_net_3626), .b(g65405_sb), .o(n_3518) );
na02s01 TIMEBOOST_cell_42755 ( .a(FE_OFN213_n_9124), .b(g57951_sb), .o(TIMEBOOST_net_13616) );
na03f02 TIMEBOOST_cell_35936 ( .a(TIMEBOOST_net_10095), .b(FE_OFN1472_g52675_p), .c(g52530_sb), .o(n_13793) );
in01s01 g64767_u0 ( .a(FE_OFN620_n_4490), .o(g64767_sb) );
na02s02 TIMEBOOST_cell_17283 ( .a(TIMEBOOST_net_3898), .b(g58043_sb), .o(n_9746) );
na02s01 g64767_u2 ( .a(n_95), .b(FE_OFN620_n_4490), .o(g64767_db) );
na02m02 TIMEBOOST_cell_40536 ( .a(TIMEBOOST_net_2024), .b(TIMEBOOST_net_12506), .o(n_13432) );
in01s01 g64768_u0 ( .a(FE_OFN1660_n_4490), .o(g64768_sb) );
na02s01 TIMEBOOST_cell_42910 ( .a(TIMEBOOST_net_13693), .b(g63077_db), .o(n_7121) );
na02s01 g64768_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__Q), .b(FE_OFN1660_n_4490), .o(g64768_db) );
na02s01 TIMEBOOST_cell_31196 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__Q), .b(pci_target_unit_fifos_pcir_data_in_158), .o(TIMEBOOST_net_9509) );
in01s01 g64769_u0 ( .a(FE_OFN670_n_4505), .o(g64769_sb) );
na02s02 TIMEBOOST_cell_40742 ( .a(TIMEBOOST_net_12609), .b(g62628_sb), .o(n_6298) );
na02s01 g64769_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__Q), .b(FE_OFN670_n_4505), .o(g64769_db) );
na02s02 TIMEBOOST_cell_40743 ( .a(wbm_adr_o_13_), .b(g59387_sb), .o(TIMEBOOST_net_12610) );
in01s01 g64770_u0 ( .a(FE_OFN671_n_4505), .o(g64770_sb) );
na03f02 TIMEBOOST_cell_35937 ( .a(TIMEBOOST_net_10094), .b(FE_OFN1472_g52675_p), .c(g52525_sb), .o(n_13734) );
na02s01 g64770_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__Q), .b(FE_OFN671_n_4505), .o(g64770_db) );
in01s01 g64771_u0 ( .a(FE_OFN671_n_4505), .o(g64771_sb) );
na02f04 TIMEBOOST_cell_39036 ( .a(TIMEBOOST_net_11756), .b(FE_OFN2243_g52675_p), .o(TIMEBOOST_net_10743) );
na02s02 TIMEBOOST_cell_40828 ( .a(TIMEBOOST_net_12652), .b(FE_OFN1331_n_13547), .o(TIMEBOOST_net_11617) );
na03s02 TIMEBOOST_cell_34038 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(g64220_sb), .c(g64220_db), .o(n_3949) );
in01s01 g64772_u0 ( .a(FE_OFN670_n_4505), .o(g64772_sb) );
na02s02 TIMEBOOST_cell_40744 ( .a(TIMEBOOST_net_12610), .b(TIMEBOOST_net_2305), .o(n_3482) );
na02s01 g64772_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__Q), .b(FE_OFN670_n_4505), .o(g64772_db) );
in01s01 g64773_u0 ( .a(FE_OFN670_n_4505), .o(g64773_sb) );
na02s01 TIMEBOOST_cell_9235 ( .a(TIMEBOOST_net_1184), .b(g65695_db), .o(n_2205) );
na02s01 TIMEBOOST_cell_40829 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__Q), .b(n_13175), .o(TIMEBOOST_net_12653) );
na02s02 TIMEBOOST_cell_40538 ( .a(TIMEBOOST_net_12507), .b(g58364_db), .o(n_9460) );
in01s01 g64774_u0 ( .a(FE_OFN670_n_4505), .o(g64774_sb) );
na03f02 TIMEBOOST_cell_35938 ( .a(TIMEBOOST_net_10093), .b(FE_OFN1472_g52675_p), .c(g52515_sb), .o(n_13806) );
na02s01 g64774_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__1__Q), .b(FE_OFN670_n_4505), .o(g64774_db) );
na02s01 TIMEBOOST_cell_42869 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__Q), .b(FE_OFN529_n_9899), .o(TIMEBOOST_net_13673) );
in01s01 g64775_u0 ( .a(FE_OFN672_n_4505), .o(g64775_sb) );
na02f04 TIMEBOOST_cell_39038 ( .a(TIMEBOOST_net_11757), .b(FE_OFN2242_g52675_p), .o(TIMEBOOST_net_10742) );
na02f02 TIMEBOOST_cell_42209 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__Q), .b(n_9657), .o(TIMEBOOST_net_13343) );
na02s01 TIMEBOOST_cell_42770 ( .a(TIMEBOOST_net_13623), .b(g57944_db), .o(n_9869) );
in01s01 g64776_u0 ( .a(FE_OFN671_n_4505), .o(g64776_sb) );
na02s02 TIMEBOOST_cell_40746 ( .a(TIMEBOOST_net_12611), .b(g62690_sb), .o(n_7364) );
na02s01 g64776_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__Q), .b(FE_OFN671_n_4505), .o(g64776_db) );
na03s02 TIMEBOOST_cell_38517 ( .a(TIMEBOOST_net_1558), .b(g65282_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__Q), .o(TIMEBOOST_net_11497) );
in01s01 g64777_u0 ( .a(FE_OFN671_n_4505), .o(g64777_sb) );
na02f02 TIMEBOOST_cell_40062 ( .a(TIMEBOOST_net_12269), .b(g57185_sb), .o(n_11568) );
na02s01 g64777_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__Q), .b(FE_OFN671_n_4505), .o(g64777_db) );
na02f02 TIMEBOOST_cell_42210 ( .a(TIMEBOOST_net_13343), .b(FE_OFN1404_n_8567), .o(TIMEBOOST_net_12296) );
in01s01 g64778_u0 ( .a(FE_OFN670_n_4505), .o(g64778_sb) );
na02s01 TIMEBOOST_cell_9279 ( .a(TIMEBOOST_net_1206), .b(g65425_db), .o(n_3510) );
na02s01 TIMEBOOST_cell_17656 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__Q), .b(g65404_sb), .o(TIMEBOOST_net_4085) );
in01s01 g64779_u0 ( .a(FE_OFN669_n_4505), .o(g64779_sb) );
na02s01 TIMEBOOST_cell_31395 ( .a(TIMEBOOST_net_9608), .b(g65045_db), .o(n_3622) );
na02s01 g64779_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q), .b(FE_OFN669_n_4505), .o(g64779_db) );
na02s01 TIMEBOOST_cell_31394 ( .a(n_3774), .b(g65045_sb), .o(TIMEBOOST_net_9608) );
in01s01 g64780_u0 ( .a(FE_OFN670_n_4505), .o(g64780_sb) );
na02s02 TIMEBOOST_cell_16765 ( .a(TIMEBOOST_net_3639), .b(n_4493), .o(n_4225) );
na02s01 g64780_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__Q), .b(FE_OFN670_n_4505), .o(g64780_db) );
na02f02 TIMEBOOST_cell_44092 ( .a(TIMEBOOST_net_14284), .b(FE_OFN1387_n_8567), .o(TIMEBOOST_net_12910) );
in01s01 g64781_u0 ( .a(FE_OFN672_n_4505), .o(g64781_sb) );
na02f02 TIMEBOOST_cell_45523 ( .a(FE_OFN2102_n_2834), .b(n_3505), .o(TIMEBOOST_net_15000) );
na02s01 g64781_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__Q), .b(FE_OFN672_n_4505), .o(g64781_db) );
na02s01 TIMEBOOST_cell_42644 ( .a(TIMEBOOST_net_13560), .b(g64855_db), .o(n_3721) );
in01s01 g64782_u0 ( .a(FE_OFN672_n_4505), .o(g64782_sb) );
na02s01 TIMEBOOST_cell_15926 ( .a(FE_OCPN1839_n_1238), .b(n_15856), .o(TIMEBOOST_net_3220) );
na02s01 g64782_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__Q), .b(FE_OFN672_n_4505), .o(g64782_db) );
na02s01 TIMEBOOST_cell_15927 ( .a(TIMEBOOST_net_3220), .b(n_4078), .o(TIMEBOOST_net_313) );
in01s01 g64783_u0 ( .a(FE_OFN669_n_4505), .o(g64783_sb) );
na02s01 g64783_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__Q), .b(FE_OFN669_n_4505), .o(g64783_db) );
na02s02 TIMEBOOST_cell_38516 ( .a(TIMEBOOST_net_11496), .b(g58374_db), .o(n_9455) );
in01s01 g64784_u0 ( .a(FE_OFN1660_n_4490), .o(g64784_sb) );
na02s01 TIMEBOOST_cell_41895 ( .a(configuration_wb_err_addr_558), .b(conf_wb_err_addr_in_967), .o(TIMEBOOST_net_13186) );
na02s01 g64784_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__Q), .b(FE_OFN1660_n_4490), .o(g64784_db) );
na02s01 TIMEBOOST_cell_31194 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__Q), .b(pci_target_unit_fifos_pcir_data_in_168), .o(TIMEBOOST_net_9508) );
in01s01 g64785_u0 ( .a(FE_OFN669_n_4505), .o(g64785_sb) );
na02s01 TIMEBOOST_cell_42645 ( .a(FE_OFN245_n_9114), .b(g57941_sb), .o(TIMEBOOST_net_13561) );
na02s01 g64785_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__Q), .b(FE_OFN669_n_4505), .o(g64785_db) );
na02s01 TIMEBOOST_cell_15930 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .b(n_1218), .o(TIMEBOOST_net_3222) );
in01s01 g64786_u0 ( .a(FE_OFN1659_n_4490), .o(g64786_sb) );
na02s01 TIMEBOOST_cell_42897 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q), .b(FE_OFN608_n_9904), .o(TIMEBOOST_net_13687) );
na02s01 g64786_u2 ( .a(n_3763), .b(FE_OFN1659_n_4490), .o(g64786_db) );
na02s01 TIMEBOOST_cell_31192 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__Q), .b(pci_target_unit_fifos_pcir_data_in_165), .o(TIMEBOOST_net_9507) );
in01s01 g64787_u0 ( .a(FE_OFN671_n_4505), .o(g64787_sb) );
na02s01 TIMEBOOST_cell_9283 ( .a(TIMEBOOST_net_1208), .b(g65873_db), .o(n_1576) );
na02f04 TIMEBOOST_cell_39040 ( .a(TIMEBOOST_net_11758), .b(FE_OFN2243_g52675_p), .o(TIMEBOOST_net_10753) );
na02f01 TIMEBOOST_cell_9285 ( .a(TIMEBOOST_net_1209), .b(n_15065), .o(n_2389) );
in01s01 g64788_u0 ( .a(FE_OFN667_n_4495), .o(g64788_sb) );
na02s01 TIMEBOOST_cell_37434 ( .a(TIMEBOOST_net_10955), .b(g65971_sb), .o(n_2153) );
na02s01 g64788_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__Q), .b(FE_OFN667_n_4495), .o(g64788_db) );
na02s01 TIMEBOOST_cell_40521 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__Q), .b(wishbone_slave_unit_pcim_sm_data_in_653), .o(TIMEBOOST_net_12499) );
in01s01 g64789_u0 ( .a(FE_OFN666_n_4495), .o(g64789_sb) );
na02s01 TIMEBOOST_cell_40540 ( .a(TIMEBOOST_net_12508), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_11558) );
na02s01 g64789_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__Q), .b(FE_OFN666_n_4495), .o(g64789_db) );
na02s01 TIMEBOOST_cell_31393 ( .a(TIMEBOOST_net_9607), .b(g64919_db), .o(n_3684) );
in01s01 g64790_u0 ( .a(FE_OFN669_n_4505), .o(g64790_sb) );
na02s01 TIMEBOOST_cell_44983 ( .a(g61943_sb), .b(g61967_db), .o(TIMEBOOST_net_14730) );
na02s01 g64790_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__Q), .b(FE_OFN669_n_4505), .o(g64790_db) );
na02f02 TIMEBOOST_cell_40064 ( .a(TIMEBOOST_net_12270), .b(g57204_sb), .o(n_10443) );
in01s01 g64791_u0 ( .a(FE_OFN667_n_4495), .o(g64791_sb) );
na02s01 TIMEBOOST_cell_42898 ( .a(TIMEBOOST_net_13687), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_11199) );
na02s01 g64791_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__Q), .b(FE_OFN667_n_4495), .o(g64791_db) );
na02s01 TIMEBOOST_cell_40542 ( .a(TIMEBOOST_net_12509), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_11560) );
in01s01 g64792_u0 ( .a(FE_OFN667_n_4495), .o(g64792_sb) );
na02s01 TIMEBOOST_cell_16376 ( .a(pci_target_unit_fifos_pcir_data_in), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__Q), .o(TIMEBOOST_net_3445) );
na02s01 g64792_u2 ( .a(n_28), .b(FE_OFN667_n_4495), .o(g64792_db) );
na02s01 TIMEBOOST_cell_16377 ( .a(TIMEBOOST_net_3445), .b(FE_OFN1017_n_2053), .o(TIMEBOOST_net_245) );
in01s01 g64793_u0 ( .a(FE_OFN667_n_4495), .o(g64793_sb) );
na02s01 TIMEBOOST_cell_31392 ( .a(n_3747), .b(g64919_sb), .o(TIMEBOOST_net_9607) );
na02s01 g64793_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__Q), .b(FE_OFN667_n_4495), .o(g64793_db) );
na02s01 TIMEBOOST_cell_16378 ( .a(n_3764), .b(n_4677), .o(TIMEBOOST_net_3446) );
in01s01 g64794_u0 ( .a(FE_OFN665_n_4495), .o(g64794_sb) );
na02s01 TIMEBOOST_cell_40543 ( .a(TIMEBOOST_net_984), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_2__Q), .o(TIMEBOOST_net_12510) );
na02s01 TIMEBOOST_cell_40544 ( .a(TIMEBOOST_net_12510), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_11561) );
in01s01 g64795_u0 ( .a(FE_OFN666_n_4495), .o(g64795_sb) );
na02s01 TIMEBOOST_cell_31391 ( .a(TIMEBOOST_net_9606), .b(n_4450), .o(n_4326) );
na02s01 g64795_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__Q), .b(FE_OFN666_n_4495), .o(g64795_db) );
na02s01 TIMEBOOST_cell_16379 ( .a(TIMEBOOST_net_3446), .b(g65290_da), .o(n_3578) );
in01s01 g64796_u0 ( .a(FE_OFN618_n_4490), .o(g64796_sb) );
na02f02 TIMEBOOST_cell_44093 ( .a(n_9075), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__Q), .o(TIMEBOOST_net_14285) );
na02s01 g64796_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__1__Q), .b(FE_OFN618_n_4490), .o(g64796_db) );
na02f02 TIMEBOOST_cell_40066 ( .a(TIMEBOOST_net_12271), .b(g57105_sb), .o(n_11640) );
in01s01 g64797_u0 ( .a(FE_OFN671_n_4505), .o(g64797_sb) );
na02m02 TIMEBOOST_cell_9287 ( .a(n_2397), .b(TIMEBOOST_net_1210), .o(TIMEBOOST_net_278) );
na02s01 TIMEBOOST_cell_15828 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_87), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3171) );
na02f02 TIMEBOOST_cell_44094 ( .a(TIMEBOOST_net_14285), .b(FE_OFN1397_n_8567), .o(TIMEBOOST_net_12911) );
in01s01 g64798_u0 ( .a(FE_OFN664_n_4495), .o(g64798_sb) );
na02s01 TIMEBOOST_cell_16116 ( .a(parchk_pci_ad_reg_in_1217), .b(pci_target_unit_del_sync_addr_in_216), .o(TIMEBOOST_net_3315) );
na02s01 g64798_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__Q), .b(FE_OFN664_n_4495), .o(g64798_db) );
na02s01 TIMEBOOST_cell_16117 ( .a(TIMEBOOST_net_3315), .b(FE_OFN2096_n_2520), .o(TIMEBOOST_net_1296) );
in01s01 g64799_u0 ( .a(FE_OFN664_n_4495), .o(g64799_sb) );
na02s01 TIMEBOOST_cell_16118 ( .a(parchk_pci_ad_reg_in_1225), .b(pci_target_unit_del_sync_addr_in_224), .o(TIMEBOOST_net_3316) );
na02s01 g64799_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__Q), .b(FE_OFN664_n_4495), .o(g64799_db) );
na02s01 TIMEBOOST_cell_16119 ( .a(TIMEBOOST_net_3316), .b(FE_OFN2096_n_2520), .o(TIMEBOOST_net_1298) );
in01s01 g64800_u0 ( .a(FE_OFN1663_n_4490), .o(g64800_sb) );
na02s01 TIMEBOOST_cell_42899 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__Q), .b(FE_OFN592_n_9694), .o(TIMEBOOST_net_13688) );
na02s01 g64800_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__5__Q), .b(FE_OFN1663_n_4490), .o(g64800_db) );
na02s01 TIMEBOOST_cell_42627 ( .a(FE_OFN219_n_9853), .b(g58176_sb), .o(TIMEBOOST_net_13552) );
in01s01 g64801_u0 ( .a(FE_OFN664_n_4495), .o(g64801_sb) );
na02s01 TIMEBOOST_cell_31390 ( .a(g65043_sb), .b(g65043_db), .o(TIMEBOOST_net_9606) );
na02s01 g64801_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__Q), .b(FE_OFN664_n_4495), .o(g64801_db) );
na02s02 TIMEBOOST_cell_45108 ( .a(TIMEBOOST_net_14792), .b(g54199_db), .o(n_13419) );
in01s01 g64802_u0 ( .a(FE_OFN664_n_4495), .o(g64802_sb) );
na02f02 TIMEBOOST_cell_40068 ( .a(TIMEBOOST_net_12272), .b(g57043_sb), .o(n_11691) );
na02s01 g64802_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q), .b(FE_OFN666_n_4495), .o(g64802_db) );
na03f02 TIMEBOOST_cell_44453 ( .a(n_3290), .b(pciu_bar0_in_375), .c(n_3050), .o(TIMEBOOST_net_14465) );
in01s01 g64803_u0 ( .a(FE_OFN671_n_4505), .o(g64803_sb) );
na02f02 TIMEBOOST_cell_40070 ( .a(TIMEBOOST_net_12273), .b(g57270_sb), .o(n_10417) );
na02s01 g64803_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q), .b(FE_OFN671_n_4505), .o(g64803_db) );
na02s01 TIMEBOOST_cell_31389 ( .a(TIMEBOOST_net_9605), .b(n_4450), .o(n_4391) );
in01s01 g64804_u0 ( .a(FE_OFN669_n_4505), .o(g64804_sb) );
na02m02 TIMEBOOST_cell_41637 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_13__Q), .b(FE_OFN211_n_9858), .o(TIMEBOOST_net_13057) );
na02s01 g64804_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__Q), .b(FE_OFN669_n_4505), .o(g64804_db) );
na02f02 TIMEBOOST_cell_44454 ( .a(TIMEBOOST_net_14465), .b(n_2842), .o(n_4647) );
in01s01 g64805_u0 ( .a(FE_OFN649_n_4497), .o(g64805_sb) );
na02s02 TIMEBOOST_cell_44455 ( .a(FE_OFN1398_n_8567), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .o(TIMEBOOST_net_14466) );
na02s01 g64805_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__20__Q), .b(FE_OFN649_n_4497), .o(g64805_db) );
na02f02 TIMEBOOST_cell_40072 ( .a(TIMEBOOST_net_12274), .b(g57202_sb), .o(n_11553) );
in01s01 g64806_u0 ( .a(FE_OFN670_n_4505), .o(g64806_sb) );
na02s01 TIMEBOOST_cell_40447 ( .a(parchk_pci_ad_out_in_1179), .b(configuration_wb_err_data_582), .o(TIMEBOOST_net_12462) );
na02s01 g64806_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__20__Q), .b(FE_OFN670_n_4505), .o(g64806_db) );
na02s02 TIMEBOOST_cell_45191 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__Q), .b(n_3549), .o(TIMEBOOST_net_14834) );
in01s01 g64807_u0 ( .a(FE_OFN614_n_4501), .o(g64807_sb) );
na02s01 TIMEBOOST_cell_31190 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__Q), .b(pci_target_unit_fifos_pcir_data_in_175), .o(TIMEBOOST_net_9506) );
na02s01 g64807_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q), .b(FE_OFN614_n_4501), .o(g64807_db) );
na02s01 TIMEBOOST_cell_41886 ( .a(TIMEBOOST_net_13181), .b(g57936_db), .o(n_9131) );
in01s01 g64808_u0 ( .a(FE_OFN664_n_4495), .o(g64808_sb) );
na02s01 TIMEBOOST_cell_16120 ( .a(parchk_pci_ad_reg_in_1232), .b(pci_target_unit_del_sync_addr_in_231), .o(TIMEBOOST_net_3317) );
na02s01 g64808_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__Q), .b(FE_OFN664_n_4495), .o(g64808_db) );
na02s01 TIMEBOOST_cell_16121 ( .a(TIMEBOOST_net_3317), .b(FE_OFN795_n_2520), .o(TIMEBOOST_net_1301) );
in01s01 g64809_u0 ( .a(FE_OFN672_n_4505), .o(g64809_sb) );
na02s01 TIMEBOOST_cell_40748 ( .a(TIMEBOOST_net_12612), .b(g62362_sb), .o(n_7392) );
na02s01 g64809_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__Q), .b(FE_OFN672_n_4505), .o(g64809_db) );
na02f02 TIMEBOOST_cell_45524 ( .a(TIMEBOOST_net_15000), .b(n_4826), .o(TIMEBOOST_net_646) );
in01s01 g64810_u0 ( .a(n_4460), .o(g64810_sb) );
na02s01 TIMEBOOST_cell_18715 ( .a(TIMEBOOST_net_4614), .b(g63107_sb), .o(n_5040) );
na02s01 g64810_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__Q), .b(n_4460), .o(g64810_db) );
na02s02 TIMEBOOST_cell_10587 ( .a(TIMEBOOST_net_1860), .b(g63050_sb), .o(n_5151) );
in01s01 g64811_u0 ( .a(FE_OFN681_n_4460), .o(g64811_sb) );
na02f02 TIMEBOOST_cell_44616 ( .a(TIMEBOOST_net_14546), .b(FE_OFN2188_n_8567), .o(TIMEBOOST_net_13004) );
na02m02 TIMEBOOST_cell_44095 ( .a(n_9576), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__Q), .o(TIMEBOOST_net_14286) );
na02s01 TIMEBOOST_cell_16768 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(g65931_sb), .o(TIMEBOOST_net_3641) );
in01s01 g64812_u0 ( .a(FE_OFN681_n_4460), .o(g64812_sb) );
na02s02 TIMEBOOST_cell_31387 ( .a(TIMEBOOST_net_9604), .b(n_4450), .o(n_4407) );
na02s01 g64812_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__Q), .b(FE_OFN681_n_4460), .o(g64812_db) );
na02f02 TIMEBOOST_cell_41624 ( .a(FE_OFN1441_n_9372), .b(TIMEBOOST_net_13050), .o(TIMEBOOST_net_11660) );
in01s01 g64813_u0 ( .a(n_4460), .o(g64813_sb) );
na02f02 TIMEBOOST_cell_10155 ( .a(TIMEBOOST_net_1644), .b(FE_OFN1149_n_13249), .o(TIMEBOOST_net_490) );
na02s01 g64813_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__Q), .b(n_4460), .o(g64813_db) );
na02s02 TIMEBOOST_cell_10157 ( .a(TIMEBOOST_net_1645), .b(FE_OFN1151_n_13249), .o(TIMEBOOST_net_503) );
in01s01 g64814_u0 ( .a(n_4460), .o(g64814_sb) );
na02s01 TIMEBOOST_cell_9239 ( .a(TIMEBOOST_net_1186), .b(g65701_db), .o(n_2201) );
na02s01 g64814_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__Q), .b(n_4460), .o(g64814_db) );
na02s01 TIMEBOOST_cell_9241 ( .a(TIMEBOOST_net_1187), .b(g65703_db), .o(n_2060) );
in01s01 g64815_u0 ( .a(n_4460), .o(g64815_sb) );
na02s01 TIMEBOOST_cell_17233 ( .a(TIMEBOOST_net_3873), .b(g65336_da), .o(n_4263) );
na02s01 g64815_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__Q), .b(n_4460), .o(g64815_db) );
na02f04 TIMEBOOST_cell_39042 ( .a(TIMEBOOST_net_11759), .b(FE_OFN2243_g52675_p), .o(TIMEBOOST_net_10741) );
in01s01 g64816_u0 ( .a(FE_OFN682_n_4460), .o(g64816_sb) );
na02s01 TIMEBOOST_cell_9291 ( .a(TIMEBOOST_net_1212), .b(TIMEBOOST_net_773), .o(n_2374) );
na02f02 TIMEBOOST_cell_44096 ( .a(TIMEBOOST_net_14286), .b(FE_OFN1376_n_8567), .o(TIMEBOOST_net_12912) );
in01s01 g64817_u0 ( .a(FE_OFN681_n_4460), .o(g64817_sb) );
na02s02 TIMEBOOST_cell_40676 ( .a(TIMEBOOST_net_12576), .b(g62937_sb), .o(n_6007) );
na02s01 g64817_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__23__Q), .b(FE_OFN681_n_4460), .o(g64817_db) );
in01s01 g64818_u0 ( .a(FE_OFN682_n_4460), .o(g64818_sb) );
na02s02 TIMEBOOST_cell_31385 ( .a(TIMEBOOST_net_9603), .b(g65064_db), .o(n_3610) );
na02s01 g64818_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__Q), .b(FE_OFN682_n_4460), .o(g64818_db) );
na02s02 TIMEBOOST_cell_31384 ( .a(n_3744), .b(g65064_sb), .o(TIMEBOOST_net_9603) );
in01s01 g64819_u0 ( .a(FE_OFN623_n_4409), .o(g64819_sb) );
na02m02 TIMEBOOST_cell_38519 ( .a(FE_OFN1700_n_5751), .b(wbm_adr_o_31_), .o(TIMEBOOST_net_11498) );
na02s01 g64819_u2 ( .a(n_3738), .b(FE_OFN623_n_4409), .o(g64819_db) );
na02f02 TIMEBOOST_cell_40902 ( .a(TIMEBOOST_net_12689), .b(g57138_sb), .o(n_11611) );
in01s01 g64820_u0 ( .a(FE_OFN682_n_4460), .o(g64820_sb) );
na02f02 TIMEBOOST_cell_40074 ( .a(TIMEBOOST_net_12275), .b(g57481_sb), .o(n_11255) );
na02s02 g64820_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__Q), .b(FE_OFN682_n_4460), .o(g64820_db) );
in01s01 g64821_u0 ( .a(n_4460), .o(g64821_sb) );
na02s01 TIMEBOOST_cell_39346 ( .a(TIMEBOOST_net_11911), .b(g64313_db), .o(n_3862) );
na02s01 g64821_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__Q), .b(n_4460), .o(g64821_db) );
na02f04 TIMEBOOST_cell_39044 ( .a(TIMEBOOST_net_11760), .b(FE_OFN2243_g52675_p), .o(TIMEBOOST_net_10740) );
in01s01 g64822_u0 ( .a(FE_OFN682_n_4460), .o(g64822_sb) );
na02f02 TIMEBOOST_cell_40076 ( .a(TIMEBOOST_net_12276), .b(g57253_sb), .o(n_11502) );
na02s01 g64822_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__Q), .b(FE_OFN682_n_4460), .o(g64822_db) );
na02s02 TIMEBOOST_cell_37920 ( .a(TIMEBOOST_net_11198), .b(FE_OFN270_n_9836), .o(n_9667) );
in01s01 g64823_u0 ( .a(FE_OFN682_n_4460), .o(g64823_sb) );
na02s02 TIMEBOOST_cell_45591 ( .a(TIMEBOOST_net_9375), .b(FE_OFN784_n_2678), .o(TIMEBOOST_net_15034) );
na02s01 g64823_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__Q), .b(FE_OFN682_n_4460), .o(g64823_db) );
na02s01 TIMEBOOST_cell_37268 ( .a(TIMEBOOST_net_10872), .b(FE_OFN682_n_4460), .o(TIMEBOOST_net_9405) );
in01s01 g64824_u0 ( .a(FE_OFN679_n_4460), .o(g64824_sb) );
na02s02 TIMEBOOST_cell_43600 ( .a(TIMEBOOST_net_14038), .b(FE_OFN1310_n_6624), .o(TIMEBOOST_net_12230) );
na02s01 g64824_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__Q), .b(FE_OFN679_n_4460), .o(g64824_db) );
na02s02 TIMEBOOST_cell_43111 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__Q), .b(n_4223), .o(TIMEBOOST_net_13794) );
in01s01 g64825_u0 ( .a(FE_OFN679_n_4460), .o(g64825_sb) );
na02s02 TIMEBOOST_cell_43112 ( .a(TIMEBOOST_net_13794), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_12090) );
na02s01 g64825_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__Q), .b(FE_OFN679_n_4460), .o(g64825_db) );
na02s02 TIMEBOOST_cell_44891 ( .a(pci_target_unit_fifos_pcir_data_in_185), .b(g65747_sb), .o(TIMEBOOST_net_14684) );
in01s01 g64826_u0 ( .a(FE_OFN629_n_4454), .o(g64826_sb) );
na03f02 TIMEBOOST_cell_36140 ( .a(FE_RN_227_0), .b(n_11730), .c(n_12568), .o(n_12830) );
na02s01 g64826_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__Q), .b(FE_OFN629_n_4454), .o(g64826_db) );
na02s02 TIMEBOOST_cell_44456 ( .a(TIMEBOOST_net_14466), .b(n_9341), .o(n_9343) );
in01s01 g64827_u0 ( .a(FE_OFN1810_n_4454), .o(g64827_sb) );
na02s01 TIMEBOOST_cell_17892 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__Q), .b(g61943_sb), .o(TIMEBOOST_net_4203) );
na02s01 TIMEBOOST_cell_17893 ( .a(TIMEBOOST_net_4203), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_860) );
in01s01 g64828_u0 ( .a(FE_OFN631_n_4454), .o(g64828_sb) );
na02s01 TIMEBOOST_cell_36647 ( .a(TIMEBOOST_net_9564), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_10562) );
na02s01 g64828_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__Q), .b(FE_OFN631_n_4454), .o(g64828_db) );
na02f02 TIMEBOOST_cell_40078 ( .a(TIMEBOOST_net_12277), .b(g57218_sb), .o(n_11538) );
in01s01 g64829_u0 ( .a(FE_OFN634_n_4454), .o(g64829_sb) );
na02s02 TIMEBOOST_cell_38518 ( .a(TIMEBOOST_net_11497), .b(FE_OFN1216_n_4151), .o(TIMEBOOST_net_5210) );
na02s01 g64829_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__Q), .b(FE_OFN634_n_4454), .o(g64829_db) );
na02f04 TIMEBOOST_cell_15936 ( .a(FE_RN_264_0), .b(n_16496), .o(TIMEBOOST_net_3225) );
in01s01 g64830_u0 ( .a(FE_OFN631_n_4454), .o(g64830_sb) );
na02s02 TIMEBOOST_cell_37776 ( .a(TIMEBOOST_net_11126), .b(g61950_sb), .o(n_7925) );
na02m02 TIMEBOOST_cell_43630 ( .a(TIMEBOOST_net_14053), .b(FE_OFN1316_n_6624), .o(TIMEBOOST_net_12228) );
na02m02 TIMEBOOST_cell_41638 ( .a(FE_OFN1439_n_9372), .b(TIMEBOOST_net_13057), .o(TIMEBOOST_net_11649) );
in01s01 g64831_u0 ( .a(FE_OFN1810_n_4454), .o(g64831_sb) );
na02s01 TIMEBOOST_cell_9738 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__Q), .b(g65821_sb), .o(TIMEBOOST_net_1436) );
na02s02 g64831_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__Q), .b(FE_OFN1810_n_4454), .o(g64831_db) );
na02s01 TIMEBOOST_cell_9739 ( .a(TIMEBOOST_net_1436), .b(g65821_db), .o(n_1895) );
in01s01 g64832_u0 ( .a(FE_OFN1810_n_4454), .o(g64832_sb) );
na02s01 TIMEBOOST_cell_9740 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__Q), .b(g65881_sb), .o(TIMEBOOST_net_1437) );
na02s02 g64832_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__Q), .b(FE_OFN1810_n_4454), .o(g64832_db) );
na02s01 TIMEBOOST_cell_9741 ( .a(TIMEBOOST_net_1437), .b(g65881_db), .o(n_1865) );
in01s01 g64833_u0 ( .a(FE_OFN633_n_4454), .o(g64833_sb) );
na02s01 TIMEBOOST_cell_40553 ( .a(TIMEBOOST_net_982), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_0__Q), .o(TIMEBOOST_net_12515) );
na02s01 g64833_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__Q), .b(FE_OFN633_n_4454), .o(g64833_db) );
na02m02 TIMEBOOST_cell_38520 ( .a(TIMEBOOST_net_11498), .b(g59798_sb), .o(TIMEBOOST_net_585) );
in01s01 g64834_u0 ( .a(FE_OFN1809_n_4454), .o(g64834_sb) );
na02m02 TIMEBOOST_cell_17894 ( .a(g53892_sb), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__Q), .o(TIMEBOOST_net_4204) );
na02s01 g64834_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__Q), .b(FE_OFN1809_n_4454), .o(g64834_db) );
na02m02 TIMEBOOST_cell_17895 ( .a(FE_OFN1148_n_13249), .b(TIMEBOOST_net_4204), .o(TIMEBOOST_net_505) );
in01s01 g64835_u0 ( .a(FE_OFN1809_n_4454), .o(g64835_sb) );
na02s02 TIMEBOOST_cell_45168 ( .a(TIMEBOOST_net_14822), .b(FE_OFN1284_n_4097), .o(TIMEBOOST_net_13258) );
na02s02 TIMEBOOST_cell_43328 ( .a(TIMEBOOST_net_13902), .b(g62516_sb), .o(n_6546) );
na02f02 TIMEBOOST_cell_40080 ( .a(TIMEBOOST_net_12278), .b(g57141_sb), .o(n_11607) );
in01s01 g64836_u0 ( .a(FE_OFN629_n_4454), .o(g64836_sb) );
na02s01 TIMEBOOST_cell_36646 ( .a(TIMEBOOST_net_10561), .b(g65813_db), .o(n_2595) );
na02s01 g64836_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__Q), .b(FE_OFN629_n_4454), .o(g64836_db) );
na03f02 TIMEBOOST_cell_44457 ( .a(n_3290), .b(pciu_bar0_in_377), .c(n_3058), .o(TIMEBOOST_net_14467) );
in01s01 g64837_u0 ( .a(FE_OFN631_n_4454), .o(g64837_sb) );
na02m02 TIMEBOOST_cell_44617 ( .a(n_9649), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__Q), .o(TIMEBOOST_net_14547) );
na02s01 g64837_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__Q), .b(FE_OFN631_n_4454), .o(g64837_db) );
na03s02 TIMEBOOST_cell_40557 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__Q), .b(n_1871), .c(FE_OFN1215_n_4151), .o(TIMEBOOST_net_12517) );
in01s01 g64838_u0 ( .a(FE_OFN631_n_4454), .o(g64838_sb) );
na02f02 TIMEBOOST_cell_40082 ( .a(TIMEBOOST_net_12279), .b(g57124_sb), .o(n_11622) );
na02s01 g64838_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__28__Q), .b(FE_OFN631_n_4454), .o(g64838_db) );
na02s01 TIMEBOOST_cell_16390 ( .a(g58042_sb), .b(g58042_db), .o(TIMEBOOST_net_3452) );
in01s01 g64839_u0 ( .a(FE_OFN634_n_4454), .o(g64839_sb) );
na02s01 TIMEBOOST_cell_42093 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__20__Q), .b(n_3753), .o(TIMEBOOST_net_13285) );
na02s01 g64839_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__Q), .b(FE_OFN634_n_4454), .o(g64839_db) );
na02s01 TIMEBOOST_cell_16391 ( .a(TIMEBOOST_net_3452), .b(FE_OFN209_n_9126), .o(n_9095) );
in01s01 g64840_u0 ( .a(FE_OFN628_n_4454), .o(g64840_sb) );
na02m02 TIMEBOOST_cell_37967 ( .a(g53893_db), .b(wishbone_slave_unit_pcim_if_wbw_cbe_in_417), .o(TIMEBOOST_net_11222) );
na02s01 g64840_u2 ( .a(n_75), .b(FE_OFN628_n_4454), .o(g64840_db) );
na02f02 TIMEBOOST_cell_37966 ( .a(TIMEBOOST_net_11221), .b(TIMEBOOST_net_495), .o(n_13461) );
in01s01 g64841_u0 ( .a(FE_OFN630_n_4454), .o(g64841_sb) );
na02s01 TIMEBOOST_cell_9295 ( .a(TIMEBOOST_net_1214), .b(g65750_db), .o(n_1605) );
na02s01 g64841_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__8__Q), .b(FE_OFN630_n_4454), .o(g64841_db) );
na02s01 TIMEBOOST_cell_9297 ( .a(TIMEBOOST_net_1215), .b(g65755_db), .o(n_1604) );
in01s01 g64842_u0 ( .a(FE_OFN689_n_4438), .o(g64842_sb) );
na02s01 TIMEBOOST_cell_16392 ( .a(pci_target_unit_pcit_if_strd_addr_in_688), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_52), .o(TIMEBOOST_net_3453) );
na02s01 g64842_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__Q), .b(FE_OFN689_n_4438), .o(g64842_db) );
na02f02 TIMEBOOST_cell_44458 ( .a(TIMEBOOST_net_14467), .b(n_2855), .o(n_4644) );
in01s01 g64843_u0 ( .a(FE_OFN1625_n_4438), .o(g64843_sb) );
na02s01 TIMEBOOST_cell_42614 ( .a(TIMEBOOST_net_13545), .b(g57984_db), .o(n_9814) );
na02m02 TIMEBOOST_cell_44097 ( .a(n_9490), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__Q), .o(TIMEBOOST_net_14287) );
na02s01 TIMEBOOST_cell_43139 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__Q), .b(n_3743), .o(TIMEBOOST_net_13808) );
in01s01 g64844_u0 ( .a(FE_OFN1624_n_4438), .o(g64844_sb) );
na02s01 TIMEBOOST_cell_40546 ( .a(TIMEBOOST_net_12511), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_11553) );
na02s01 g64844_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__Q), .b(FE_OFN1624_n_4438), .o(g64844_db) );
na02f02 TIMEBOOST_cell_44459 ( .a(FE_OFN1398_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_), .o(TIMEBOOST_net_14468) );
in01s01 g64845_u0 ( .a(FE_OFN1625_n_4438), .o(g64845_sb) );
na02s01 TIMEBOOST_cell_36648 ( .a(TIMEBOOST_net_10562), .b(g65858_sb), .o(n_2594) );
na02s01 g64845_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__Q), .b(FE_OFN1625_n_4438), .o(g64845_db) );
na02s01 TIMEBOOST_cell_44984 ( .a(TIMEBOOST_net_14730), .b(g63599_db), .o(TIMEBOOST_net_13153) );
in01s01 g64846_u0 ( .a(FE_OFN1624_n_4438), .o(g64846_sb) );
na02s01 TIMEBOOST_cell_36651 ( .a(parchk_pci_ad_reg_in_1224), .b(g65813_sb), .o(TIMEBOOST_net_10564) );
na02s01 g64846_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__14__Q), .b(FE_OFN1624_n_4438), .o(g64846_db) );
na02f02 TIMEBOOST_cell_40084 ( .a(TIMEBOOST_net_12280), .b(g57089_sb), .o(n_11652) );
in01s01 g64847_u0 ( .a(FE_OFN1625_n_4438), .o(g64847_sb) );
na02s02 TIMEBOOST_cell_43604 ( .a(TIMEBOOST_net_14040), .b(FE_OFN1317_n_6624), .o(TIMEBOOST_net_12236) );
na02s01 g64847_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__Q), .b(FE_OFN1625_n_4438), .o(g64847_db) );
na02m02 TIMEBOOST_cell_43761 ( .a(n_9845), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__Q), .o(TIMEBOOST_net_14119) );
in01s01 g64848_u0 ( .a(FE_OFN1625_n_4438), .o(g64848_sb) );
na02s01 TIMEBOOST_cell_41775 ( .a(FE_OFN247_n_9112), .b(g58194_sb), .o(TIMEBOOST_net_13126) );
na02s01 g64848_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__Q), .b(FE_OFN1625_n_4438), .o(g64848_db) );
na02s01 TIMEBOOST_cell_44885 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__Q), .b(FE_OFN1678_n_4655), .o(TIMEBOOST_net_14681) );
in01s01 g64849_u0 ( .a(FE_OFN1626_n_4438), .o(g64849_sb) );
na02m02 TIMEBOOST_cell_44327 ( .a(n_9461), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__Q), .o(TIMEBOOST_net_14402) );
na02s01 g64849_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__Q), .b(FE_OFN1626_n_4438), .o(g64849_db) );
na02f02 TIMEBOOST_cell_44328 ( .a(TIMEBOOST_net_14402), .b(FE_OFN1401_n_8567), .o(TIMEBOOST_net_12726) );
in01s01 g64850_u0 ( .a(FE_OFN1628_n_4438), .o(g64850_sb) );
na02s01 TIMEBOOST_cell_42626 ( .a(TIMEBOOST_net_13551), .b(FE_OFN217_n_9889), .o(TIMEBOOST_net_3793) );
na02m02 TIMEBOOST_cell_44395 ( .a(n_9771), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__Q), .o(TIMEBOOST_net_14436) );
na02f02 TIMEBOOST_cell_43800 ( .a(TIMEBOOST_net_14138), .b(FE_OFN1392_n_8567), .o(TIMEBOOST_net_13375) );
in01s01 g64851_u0 ( .a(FE_OFN1624_n_4438), .o(g64851_sb) );
na02m08 TIMEBOOST_cell_36282 ( .a(TIMEBOOST_net_10379), .b(n_783), .o(n_11877) );
na02s01 g64851_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__Q), .b(FE_OFN1624_n_4438), .o(g64851_db) );
na02s01 TIMEBOOST_cell_16769 ( .a(TIMEBOOST_net_3641), .b(g65931_db), .o(n_1849) );
in01s01 g64852_u0 ( .a(FE_OFN1625_n_4438), .o(g64852_sb) );
na02s01 TIMEBOOST_cell_36650 ( .a(TIMEBOOST_net_10563), .b(g65892_sb), .o(n_2569) );
na02f02 TIMEBOOST_cell_41514 ( .a(TIMEBOOST_net_12995), .b(g57260_sb), .o(n_11493) );
na02s02 TIMEBOOST_cell_45037 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__Q), .b(n_1613), .o(TIMEBOOST_net_14757) );
in01s01 g64853_u0 ( .a(FE_OFN1626_n_4438), .o(g64853_sb) );
na02s02 TIMEBOOST_cell_42094 ( .a(TIMEBOOST_net_13285), .b(FE_OFN1230_n_6391), .o(TIMEBOOST_net_11573) );
na02s01 g64853_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__Q), .b(FE_OFN1626_n_4438), .o(g64853_db) );
na02s02 TIMEBOOST_cell_45109 ( .a(g63196_db), .b(TIMEBOOST_net_9826), .o(TIMEBOOST_net_14793) );
in01s01 g64854_u0 ( .a(FE_OFN1626_n_4438), .o(g64854_sb) );
na02s01 TIMEBOOST_cell_36652 ( .a(TIMEBOOST_net_10564), .b(g65963_db), .o(n_2571) );
na02f02 TIMEBOOST_cell_44098 ( .a(TIMEBOOST_net_14287), .b(FE_OFN1388_n_8567), .o(TIMEBOOST_net_12927) );
na02f02 TIMEBOOST_cell_40086 ( .a(TIMEBOOST_net_12281), .b(g57264_sb), .o(n_11489) );
in01s01 g64855_u0 ( .a(FE_OFN1626_n_4438), .o(g64855_sb) );
na02m02 TIMEBOOST_cell_44329 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q), .b(n_9481), .o(TIMEBOOST_net_14403) );
na02s01 g64855_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__Q), .b(FE_OFN1626_n_4438), .o(g64855_db) );
na02f02 TIMEBOOST_cell_44330 ( .a(TIMEBOOST_net_14403), .b(FE_OFN1373_n_8567), .o(TIMEBOOST_net_12712) );
in01s01 g64856_u0 ( .a(FE_OFN689_n_4438), .o(g64856_sb) );
na02m02 TIMEBOOST_cell_44331 ( .a(n_9197), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__Q), .o(TIMEBOOST_net_14404) );
na02f02 TIMEBOOST_cell_44460 ( .a(TIMEBOOST_net_14468), .b(n_9341), .o(n_9342) );
na02f02 TIMEBOOST_cell_44332 ( .a(TIMEBOOST_net_14404), .b(FE_OFN1416_n_8567), .o(TIMEBOOST_net_12742) );
in01s01 g64857_u0 ( .a(FE_OFN1623_n_4438), .o(g64857_sb) );
na03f04 TIMEBOOST_cell_34445 ( .a(FE_OCPN1823_n_16560), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q), .c(n_16521), .o(n_16442) );
na02s02 g64857_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__Q), .b(FE_OFN1623_n_4438), .o(g64857_db) );
na02s01 TIMEBOOST_cell_42758 ( .a(TIMEBOOST_net_13617), .b(g58169_db), .o(n_9622) );
in01s01 g64858_u0 ( .a(FE_OFN615_n_4501), .o(g64858_sb) );
na02s01 TIMEBOOST_cell_31188 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__Q), .b(pci_target_unit_fifos_pcir_data_in_176), .o(TIMEBOOST_net_9505) );
na02s01 g64858_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__Q), .b(FE_OFN615_n_4501), .o(g64858_db) );
na02s01 TIMEBOOST_cell_42900 ( .a(TIMEBOOST_net_13688), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_11191) );
in01s01 g64859_u0 ( .a(FE_OFN612_n_4501), .o(g64859_sb) );
na02s02 TIMEBOOST_cell_16770 ( .a(n_3770), .b(g64753_sb), .o(TIMEBOOST_net_3642) );
na02s01 g64859_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__Q), .b(FE_OFN612_n_4501), .o(g64859_db) );
na02s01 TIMEBOOST_cell_16771 ( .a(TIMEBOOST_net_3642), .b(g64753_db), .o(n_3790) );
in01s01 g64860_u0 ( .a(FE_OFN647_n_4497), .o(g64860_sb) );
na02s01 g64860_u2 ( .a(n_4429), .b(FE_OFN647_n_4497), .o(g64860_db) );
na02s01 TIMEBOOST_cell_40750 ( .a(TIMEBOOST_net_12613), .b(g63144_sb), .o(n_5852) );
in01s01 g64861_u0 ( .a(FE_OFN1663_n_4490), .o(g64861_sb) );
na02m02 TIMEBOOST_cell_44099 ( .a(n_9541), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__Q), .o(TIMEBOOST_net_14288) );
na02s01 g64861_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__Q), .b(FE_OFN1663_n_4490), .o(g64861_db) );
na02s01 TIMEBOOST_cell_31186 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__Q), .b(pci_target_unit_fifos_pcir_data_in_177), .o(TIMEBOOST_net_9504) );
in01s01 g64862_u0 ( .a(FE_OFN615_n_4501), .o(g64862_sb) );
na02s01 TIMEBOOST_cell_42901 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__Q), .b(FE_OFN554_n_9864), .o(TIMEBOOST_net_13689) );
na02s01 g64862_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__15__Q), .b(FE_OFN615_n_4501), .o(g64862_db) );
na03s02 TIMEBOOST_cell_41887 ( .a(g64089_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__Q), .c(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_13182) );
in01s01 g64863_u0 ( .a(FE_OFN615_n_4501), .o(g64863_sb) );
na02f02 TIMEBOOST_cell_31183 ( .a(n_2022), .b(TIMEBOOST_net_9502), .o(TIMEBOOST_net_6242) );
na02s01 g64863_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__Q), .b(FE_OFN615_n_4501), .o(g64863_db) );
na02m02 TIMEBOOST_cell_31182 ( .a(g57779_da), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_9502) );
in01s01 g64864_u0 ( .a(FE_OFN1807_n_4501), .o(g64864_sb) );
na02s01 TIMEBOOST_cell_17980 ( .a(pci_target_unit_fifos_pciw_addr_data_in_146), .b(g64221_sb), .o(TIMEBOOST_net_4247) );
na02s01 g64864_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__Q), .b(FE_OFN1807_n_4501), .o(g64864_db) );
na02s02 TIMEBOOST_cell_44863 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__Q), .b(FE_OFN1643_n_4671), .o(TIMEBOOST_net_14670) );
in01s01 g64865_u0 ( .a(FE_OFN615_n_4501), .o(g64865_sb) );
na02f02 TIMEBOOST_cell_41862 ( .a(TIMEBOOST_net_13169), .b(TIMEBOOST_net_496), .o(n_13446) );
na02s01 g64865_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__Q), .b(FE_OFN615_n_4501), .o(g64865_db) );
na02s02 TIMEBOOST_cell_41863 ( .a(TIMEBOOST_net_332), .b(g61899_sb), .o(TIMEBOOST_net_13170) );
in01s01 g64866_u0 ( .a(FE_OFN612_n_4501), .o(g64866_sb) );
na02s01 g64866_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__Q), .b(FE_OFN612_n_4501), .o(g64866_db) );
na02f04 TIMEBOOST_cell_44871 ( .a(n_4675), .b(n_4874), .o(TIMEBOOST_net_14674) );
in01s01 g64867_u0 ( .a(FE_OFN1807_n_4501), .o(g64867_sb) );
na02s01 TIMEBOOST_cell_17982 ( .a(pci_target_unit_fifos_pciw_addr_data_in_145), .b(g64222_sb), .o(TIMEBOOST_net_4248) );
na02s01 g64867_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__Q), .b(FE_OFN1807_n_4501), .o(g64867_db) );
na02m02 TIMEBOOST_cell_38937 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_15__Q), .o(TIMEBOOST_net_11707) );
in01s01 g64868_u0 ( .a(FE_OFN615_n_4501), .o(g64868_sb) );
na02s01 TIMEBOOST_cell_41864 ( .a(TIMEBOOST_net_13170), .b(g61899_db), .o(n_8027) );
na02f02 TIMEBOOST_cell_44100 ( .a(TIMEBOOST_net_14288), .b(FE_OFN1382_n_8567), .o(TIMEBOOST_net_13382) );
na02s01 TIMEBOOST_cell_42870 ( .a(TIMEBOOST_net_13673), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_11210) );
in01s01 g64869_u0 ( .a(FE_OFN1806_n_4501), .o(g64869_sb) );
na02f02 TIMEBOOST_cell_42255 ( .a(n_9655), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__Q), .o(TIMEBOOST_net_13366) );
na02s02 g64869_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q), .b(FE_OFN1806_n_4501), .o(g64869_db) );
na02s02 TIMEBOOST_cell_36785 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__Q), .b(n_4004), .o(TIMEBOOST_net_10631) );
in01s01 g64870_u0 ( .a(FE_OFN1807_n_4501), .o(g64870_sb) );
na02s01 TIMEBOOST_cell_39277 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q), .b(g64301_sb), .o(TIMEBOOST_net_11877) );
na02s01 g64870_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__Q), .b(FE_OFN1807_n_4501), .o(g64870_db) );
na02s01 TIMEBOOST_cell_39278 ( .a(TIMEBOOST_net_11877), .b(g64301_db), .o(n_3874) );
in01s01 g64871_u0 ( .a(FE_OFN612_n_4501), .o(g64871_sb) );
na02s01 TIMEBOOST_cell_42871 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__Q), .b(FE_OFN587_n_9692), .o(TIMEBOOST_net_13674) );
na02s01 g64871_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__Q), .b(FE_OFN612_n_4501), .o(g64871_db) );
na02s02 TIMEBOOST_cell_31175 ( .a(TIMEBOOST_net_9498), .b(g64881_sb), .o(n_3706) );
in01s01 g64872_u0 ( .a(FE_OFN615_n_4501), .o(g64872_sb) );
na02s01 TIMEBOOST_cell_45127 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__Q), .b(n_3971), .o(TIMEBOOST_net_14802) );
na02s01 g64872_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__Q), .b(FE_OFN615_n_4501), .o(g64872_db) );
na02f02 TIMEBOOST_cell_40088 ( .a(TIMEBOOST_net_12282), .b(g57568_sb), .o(n_11184) );
in01s01 g64873_u0 ( .a(FE_OFN1807_n_4501), .o(g64873_sb) );
na02s01 TIMEBOOST_cell_17988 ( .a(pci_target_unit_fifos_pciw_addr_data_in_141), .b(g64084_sb), .o(TIMEBOOST_net_4251) );
na02s01 g64873_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__Q), .b(FE_OFN614_n_4501), .o(g64873_db) );
na03s02 TIMEBOOST_cell_38333 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__Q), .b(FE_OFN1137_g64577_p), .c(n_3870), .o(TIMEBOOST_net_11405) );
in01s01 g64874_u0 ( .a(FE_OFN614_n_4501), .o(g64874_sb) );
na02m02 TIMEBOOST_cell_44101 ( .a(n_9056), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__Q), .o(TIMEBOOST_net_14289) );
na02s01 g64874_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__Q), .b(FE_OFN614_n_4501), .o(g64874_db) );
na02s01 TIMEBOOST_cell_31173 ( .a(TIMEBOOST_net_9497), .b(g64859_db), .o(n_3717) );
in01s01 g64875_u0 ( .a(FE_OFN664_n_4495), .o(g64875_sb) );
na03s02 TIMEBOOST_cell_42095 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__Q), .b(n_4258), .c(FE_OFN1236_n_6391), .o(TIMEBOOST_net_13286) );
na02s01 g64875_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__Q), .b(FE_OFN664_n_4495), .o(g64875_db) );
na03s02 TIMEBOOST_cell_45525 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__Q), .b(FE_OFN1094_g64577_p), .c(n_4595), .o(TIMEBOOST_net_15001) );
in01s01 g64876_u0 ( .a(FE_OFN612_n_4501), .o(g64876_sb) );
na02f06 TIMEBOOST_cell_41704 ( .a(TIMEBOOST_net_13090), .b(n_16424), .o(n_16425) );
na02s01 g64876_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__Q), .b(FE_OFN612_n_4501), .o(g64876_db) );
na02s02 TIMEBOOST_cell_17285 ( .a(TIMEBOOST_net_3899), .b(FE_OFN254_n_9825), .o(n_9432) );
in01s01 g64877_u0 ( .a(FE_OFN612_n_4501), .o(g64877_sb) );
na02f04 TIMEBOOST_cell_39046 ( .a(TIMEBOOST_net_11761), .b(FE_OFN2243_g52675_p), .o(TIMEBOOST_net_10739) );
na02s02 TIMEBOOST_cell_15938 ( .a(n_2756), .b(n_2305), .o(TIMEBOOST_net_3226) );
na02f04 TIMEBOOST_cell_39048 ( .a(TIMEBOOST_net_11762), .b(FE_OFN2243_g52675_p), .o(TIMEBOOST_net_10747) );
in01s01 g64878_u0 ( .a(FE_OFN665_n_4495), .o(g64878_sb) );
na02m02 TIMEBOOST_cell_44203 ( .a(n_9459), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__Q), .o(TIMEBOOST_net_14340) );
na02f02 TIMEBOOST_cell_43762 ( .a(TIMEBOOST_net_14119), .b(FE_OFN1392_n_8567), .o(TIMEBOOST_net_12946) );
na02s01 TIMEBOOST_cell_16122 ( .a(parchk_pci_ad_reg_in_1226), .b(pci_target_unit_del_sync_addr_in_225), .o(TIMEBOOST_net_3318) );
in01s01 g64879_u0 ( .a(FE_OFN686_n_4417), .o(g64879_sb) );
na02s02 TIMEBOOST_cell_37436 ( .a(TIMEBOOST_net_10956), .b(FE_OFN227_n_9841), .o(n_9735) );
na02f02 TIMEBOOST_cell_44102 ( .a(TIMEBOOST_net_14289), .b(FE_OFN1380_n_8567), .o(TIMEBOOST_net_12913) );
na02s01 TIMEBOOST_cell_36654 ( .a(TIMEBOOST_net_10565), .b(g65892_sb), .o(n_2572) );
in01s01 g64880_u0 ( .a(FE_OFN686_n_4417), .o(g64880_sb) );
na02s01 TIMEBOOST_cell_37439 ( .a(TIMEBOOST_net_3459), .b(g52647_sb), .o(TIMEBOOST_net_10958) );
na02m02 TIMEBOOST_cell_44103 ( .a(n_9498), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__Q), .o(TIMEBOOST_net_14290) );
na02s02 TIMEBOOST_cell_37438 ( .a(TIMEBOOST_net_10957), .b(n_3453), .o(n_5723) );
in01s01 g64881_u0 ( .a(FE_OFN685_n_4417), .o(g64881_sb) );
na02m02 TIMEBOOST_cell_44461 ( .a(n_9218), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__Q), .o(TIMEBOOST_net_14469) );
na02s02 TIMEBOOST_cell_43445 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__20__Q), .b(n_3540), .o(TIMEBOOST_net_13961) );
na02f02 TIMEBOOST_cell_40090 ( .a(TIMEBOOST_net_12283), .b(g57287_sb), .o(n_11466) );
in01s01 g64882_u0 ( .a(FE_OFN685_n_4417), .o(g64882_sb) );
na02f02 TIMEBOOST_cell_40092 ( .a(TIMEBOOST_net_12284), .b(g57490_sb), .o(n_11246) );
na02s01 g64882_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__14__Q), .b(FE_OFN685_n_4417), .o(g64882_db) );
na02s01 TIMEBOOST_cell_42096 ( .a(TIMEBOOST_net_13286), .b(g62981_sb), .o(n_5920) );
in01s01 g64883_u0 ( .a(FE_OFN686_n_4417), .o(g64883_sb) );
na02f02 TIMEBOOST_cell_44462 ( .a(TIMEBOOST_net_14469), .b(FE_OFN2175_n_8567), .o(TIMEBOOST_net_13018) );
na02s01 g64883_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__Q), .b(FE_OFN686_n_4417), .o(g64883_db) );
na02s01 TIMEBOOST_cell_36656 ( .a(TIMEBOOST_net_10566), .b(g65892_sb), .o(n_2573) );
in01s01 g64884_u0 ( .a(FE_OFN686_n_4417), .o(g64884_sb) );
na02f02 TIMEBOOST_cell_44104 ( .a(TIMEBOOST_net_14290), .b(FE_OFN1408_n_8567), .o(TIMEBOOST_net_12914) );
na02s01 g64884_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__Q), .b(FE_OFN686_n_4417), .o(g64884_db) );
na02s02 TIMEBOOST_cell_43446 ( .a(TIMEBOOST_net_13961), .b(FE_OFN1230_n_6391), .o(TIMEBOOST_net_12622) );
in01s01 g64885_u0 ( .a(FE_OFN686_n_4417), .o(g64885_sb) );
na02f02 TIMEBOOST_cell_40094 ( .a(TIMEBOOST_net_12285), .b(g57071_sb), .o(n_11670) );
na02s01 g64885_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__Q), .b(FE_OFN686_n_4417), .o(g64885_db) );
na02s01 TIMEBOOST_cell_31369 ( .a(TIMEBOOST_net_9595), .b(g65331_da), .o(n_4265) );
in01s01 g64886_u0 ( .a(FE_OFN686_n_4417), .o(g64886_sb) );
na02f02 TIMEBOOST_cell_40096 ( .a(TIMEBOOST_net_12286), .b(g57576_sb), .o(n_11175) );
na02s01 g64886_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__Q), .b(FE_OFN686_n_4417), .o(g64886_db) );
na02s01 TIMEBOOST_cell_36266 ( .a(TIMEBOOST_net_10371), .b(wbu_addr_in_273), .o(n_9841) );
in01s01 g64887_u0 ( .a(FE_OFN687_n_4417), .o(g64887_sb) );
na02m02 TIMEBOOST_cell_44105 ( .a(n_9742), .b(n_15569), .o(TIMEBOOST_net_14291) );
na02f02 TIMEBOOST_cell_44106 ( .a(TIMEBOOST_net_14291), .b(FE_OFN1387_n_8567), .o(TIMEBOOST_net_12990) );
na02m02 TIMEBOOST_cell_44107 ( .a(n_9842), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__Q), .o(TIMEBOOST_net_14292) );
in01s01 g64888_u0 ( .a(FE_OFN685_n_4417), .o(g64888_sb) );
na02s02 TIMEBOOST_cell_39555 ( .a(wbm_adr_o_28_), .b(FE_OFN1698_n_5751), .o(TIMEBOOST_net_12016) );
na02s01 g64888_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__Q), .b(FE_OFN685_n_4417), .o(g64888_db) );
na02s01 TIMEBOOST_cell_40548 ( .a(TIMEBOOST_net_12512), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_11557) );
in01s01 g64889_u0 ( .a(FE_OFN685_n_4417), .o(g64889_sb) );
na02s01 TIMEBOOST_cell_40261 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__Q), .b(n_2161), .o(TIMEBOOST_net_12369) );
na02s01 g64889_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__Q), .b(FE_OFN685_n_4417), .o(g64889_db) );
na02f02 TIMEBOOST_cell_40098 ( .a(TIMEBOOST_net_12287), .b(g57349_sb), .o(n_11401) );
in01s01 g64890_u0 ( .a(FE_OFN686_n_4417), .o(g64890_sb) );
na02m02 TIMEBOOST_cell_44463 ( .a(n_9539), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__Q), .o(TIMEBOOST_net_14470) );
na02s01 g64890_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__Q), .b(FE_OFN686_n_4417), .o(g64890_db) );
na02f02 TIMEBOOST_cell_40100 ( .a(TIMEBOOST_net_12288), .b(g57328_sb), .o(n_11421) );
in01s01 g64891_u0 ( .a(FE_OFN687_n_4417), .o(g64891_sb) );
na02s01 TIMEBOOST_cell_16404 ( .a(pci_target_unit_pcit_if_strd_addr_in_690), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_54), .o(TIMEBOOST_net_3459) );
na02s01 g64891_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__Q), .b(FE_OFN687_n_4417), .o(g64891_db) );
na02f02 TIMEBOOST_cell_44464 ( .a(TIMEBOOST_net_14470), .b(FE_OFN2173_n_8567), .o(TIMEBOOST_net_13433) );
in01s01 g64892_u0 ( .a(FE_OFN687_n_4417), .o(g64892_sb) );
na02s01 TIMEBOOST_cell_45075 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__Q), .b(FE_OFN518_n_9697), .o(TIMEBOOST_net_14776) );
na02s01 g64892_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__Q), .b(FE_OFN687_n_4417), .o(g64892_db) );
na02s01 TIMEBOOST_cell_31368 ( .a(n_4473), .b(FE_OFN654_n_4508), .o(TIMEBOOST_net_9595) );
in01s01 g64893_u0 ( .a(FE_OFN686_n_4417), .o(g64893_sb) );
na02f02 TIMEBOOST_cell_44465 ( .a(n_9506), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__Q), .o(TIMEBOOST_net_14471) );
na02f02 TIMEBOOST_cell_44108 ( .a(TIMEBOOST_net_14292), .b(FE_OFN1422_n_8567), .o(TIMEBOOST_net_12860) );
na02f02 TIMEBOOST_cell_44466 ( .a(TIMEBOOST_net_14471), .b(FE_OFN2173_n_8567), .o(TIMEBOOST_net_13434) );
in01s01 g64894_u0 ( .a(FE_OFN687_n_4417), .o(g64894_sb) );
na02m02 TIMEBOOST_cell_44109 ( .a(n_9689), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__Q), .o(TIMEBOOST_net_14293) );
na02s02 TIMEBOOST_cell_40678 ( .a(TIMEBOOST_net_12577), .b(g62661_sb), .o(n_6221) );
in01s01 g64895_u0 ( .a(FE_OFN687_n_4417), .o(g64895_sb) );
na02m02 TIMEBOOST_cell_43729 ( .a(n_9820), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__Q), .o(TIMEBOOST_net_14103) );
na02s01 g64895_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__Q), .b(FE_OFN687_n_4417), .o(g64895_db) );
na02s02 TIMEBOOST_cell_43378 ( .a(TIMEBOOST_net_13927), .b(n_6319), .o(TIMEBOOST_net_12158) );
in01s01 g64896_u0 ( .a(n_4417), .o(g64896_sb) );
na02m02 TIMEBOOST_cell_10159 ( .a(FE_OFN1151_n_13249), .b(TIMEBOOST_net_1646), .o(TIMEBOOST_net_493) );
na02s01 g64896_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__Q), .b(n_4417), .o(g64896_db) );
na02f02 TIMEBOOST_cell_10161 ( .a(TIMEBOOST_net_1647), .b(FE_OFN1149_n_13249), .o(TIMEBOOST_net_494) );
in01s01 g64897_u0 ( .a(FE_OFN684_n_4417), .o(g64897_sb) );
na02f02 TIMEBOOST_cell_43730 ( .a(TIMEBOOST_net_14103), .b(FE_OFN1423_n_8567), .o(TIMEBOOST_net_12694) );
na02s01 g64897_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__Q), .b(FE_OFN684_n_4417), .o(g64897_db) );
na02f02 TIMEBOOST_cell_40102 ( .a(TIMEBOOST_net_12289), .b(g57526_sb), .o(n_11215) );
in01s01 g64898_u0 ( .a(FE_OFN684_n_4417), .o(g64898_sb) );
na02m02 TIMEBOOST_cell_44467 ( .a(n_9872), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__Q), .o(TIMEBOOST_net_14472) );
na02s01 g64898_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__Q), .b(FE_OFN684_n_4417), .o(g64898_db) );
na02f02 TIMEBOOST_cell_44396 ( .a(TIMEBOOST_net_14436), .b(FE_OFN1421_n_8567), .o(TIMEBOOST_net_12727) );
in01s01 g64899_u0 ( .a(FE_OFN624_n_4409), .o(g64899_sb) );
na02s02 TIMEBOOST_cell_15939 ( .a(TIMEBOOST_net_3226), .b(n_2753), .o(TIMEBOOST_net_214) );
na02s01 g64899_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__Q), .b(FE_OFN624_n_4409), .o(g64899_db) );
na02s01 TIMEBOOST_cell_15940 ( .a(pci_target_unit_fifos_pcir_data_in_178), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__Q), .o(TIMEBOOST_net_3227) );
in01s01 g64900_u0 ( .a(FE_OFN624_n_4409), .o(g64900_sb) );
na02s02 TIMEBOOST_cell_38599 ( .a(TIMEBOOST_net_9933), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_11538) );
na02s01 g64900_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__Q), .b(FE_OFN624_n_4409), .o(g64900_db) );
in01s01 g64901_u0 ( .a(FE_OFN625_n_4409), .o(g64901_sb) );
na02f02 TIMEBOOST_cell_40104 ( .a(TIMEBOOST_net_12290), .b(g57454_sb), .o(n_11280) );
na02s01 g64901_u2 ( .a(n_4410), .b(FE_OFN625_n_4409), .o(g64901_db) );
na02f02 TIMEBOOST_cell_44468 ( .a(TIMEBOOST_net_14472), .b(FE_OFN2174_n_8567), .o(TIMEBOOST_net_13435) );
in01s01 g64902_u0 ( .a(FE_OFN625_n_4409), .o(g64902_sb) );
na02f02 TIMEBOOST_cell_40106 ( .a(TIMEBOOST_net_12291), .b(g57296_sb), .o(n_11456) );
na02s01 g64902_u2 ( .a(n_0), .b(FE_OFN625_n_4409), .o(g64902_db) );
na02s01 TIMEBOOST_cell_16412 ( .a(n_3764), .b(g64808_sb), .o(TIMEBOOST_net_3463) );
in01s01 g64903_u0 ( .a(FE_OFN623_n_4409), .o(g64903_sb) );
na02s02 TIMEBOOST_cell_38598 ( .a(TIMEBOOST_net_11537), .b(g60627_sb), .o(n_5710) );
na02s01 g64903_u2 ( .a(n_3691), .b(FE_OFN623_n_4409), .o(g64903_db) );
na02s01 TIMEBOOST_cell_15942 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__Q), .o(TIMEBOOST_net_3228) );
in01s01 g64904_u0 ( .a(FE_OFN623_n_4409), .o(g64904_sb) );
na02s01 TIMEBOOST_cell_42972 ( .a(TIMEBOOST_net_13724), .b(n_4743), .o(TIMEBOOST_net_509) );
na02s01 TIMEBOOST_cell_44985 ( .a(g61962_sb), .b(g61986_db), .o(TIMEBOOST_net_14731) );
na02m02 TIMEBOOST_cell_38933 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_12__Q), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__Q), .o(TIMEBOOST_net_11705) );
in01s01 g64905_u0 ( .a(FE_OFN624_n_4409), .o(g64905_sb) );
na02s01 TIMEBOOST_cell_16413 ( .a(TIMEBOOST_net_3463), .b(g64808_db), .o(n_3751) );
na02s01 g64905_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__Q), .b(FE_OFN624_n_4409), .o(g64905_db) );
na02s02 TIMEBOOST_cell_16414 ( .a(n_3739), .b(g64966_sb), .o(TIMEBOOST_net_3464) );
in01s01 g64906_u0 ( .a(FE_OFN624_n_4409), .o(g64906_sb) );
na02s01 TIMEBOOST_cell_15944 ( .a(pci_target_unit_fifos_pcir_data_in_173), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__Q), .o(TIMEBOOST_net_3229) );
na02s01 g64906_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__20__Q), .b(FE_OFN624_n_4409), .o(g64906_db) );
in01s01 g64907_u0 ( .a(FE_OFN624_n_4409), .o(g64907_sb) );
na02f02 TIMEBOOST_cell_40904 ( .a(TIMEBOOST_net_12690), .b(g57515_sb), .o(n_11226) );
na02s01 g64907_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__22__Q), .b(FE_OFN624_n_4409), .o(g64907_db) );
no02f06 TIMEBOOST_cell_15947 ( .a(TIMEBOOST_net_3230), .b(n_832), .o(g65808_p) );
in01s01 g64908_u0 ( .a(FE_OFN625_n_4409), .o(g64908_sb) );
na02s01 TIMEBOOST_cell_16415 ( .a(TIMEBOOST_net_3464), .b(g64966_db), .o(n_3654) );
na02s01 g64908_u2 ( .a(n_156), .b(FE_OFN625_n_4409), .o(g64908_db) );
na02s01 TIMEBOOST_cell_16416 ( .a(n_3747), .b(g65091_sb), .o(TIMEBOOST_net_3465) );
in01s01 g64909_u0 ( .a(FE_OFN625_n_4409), .o(g64909_sb) );
na02s01 TIMEBOOST_cell_16417 ( .a(TIMEBOOST_net_3465), .b(g65091_db), .o(n_3597) );
na02s01 g64909_u2 ( .a(n_4403), .b(FE_OFN625_n_4409), .o(g64909_db) );
na02s01 TIMEBOOST_cell_36658 ( .a(TIMEBOOST_net_10567), .b(g65892_sb), .o(n_2582) );
in01s01 g64910_u0 ( .a(FE_OFN625_n_4409), .o(g64910_sb) );
na02m02 TIMEBOOST_cell_44469 ( .a(n_9485), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q), .o(TIMEBOOST_net_14473) );
na02s01 g64910_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__Q), .b(FE_OFN625_n_4409), .o(g64910_db) );
na02f02 TIMEBOOST_cell_40108 ( .a(TIMEBOOST_net_12292), .b(g57517_sb), .o(n_11223) );
in01s01 g64911_u0 ( .a(FE_OFN622_n_4409), .o(g64911_sb) );
na02s01 TIMEBOOST_cell_16420 ( .a(n_3741), .b(g64998_sb), .o(TIMEBOOST_net_3467) );
na02s01 g64911_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__Q), .b(FE_OFN622_n_4409), .o(g64911_db) );
na02s02 TIMEBOOST_cell_16421 ( .a(TIMEBOOST_net_3467), .b(g64998_db), .o(n_3643) );
in01s01 g64912_u0 ( .a(FE_OFN623_n_4409), .o(g64912_sb) );
na02s01 TIMEBOOST_cell_45076 ( .a(TIMEBOOST_net_14776), .b(FE_OFN270_n_9836), .o(TIMEBOOST_net_11941) );
na02s01 g64912_u2 ( .a(n_4399), .b(FE_OFN623_n_4409), .o(g64912_db) );
na02f02 TIMEBOOST_cell_40110 ( .a(TIMEBOOST_net_12293), .b(g57254_sb), .o(n_11500) );
in01s01 g64913_u0 ( .a(FE_OFN625_n_4409), .o(g64913_sb) );
na02s01 TIMEBOOST_cell_16424 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__Q), .b(g64327_sb), .o(TIMEBOOST_net_3469) );
na02s01 g64913_u2 ( .a(n_50), .b(FE_OFN625_n_4409), .o(g64913_db) );
na02s02 TIMEBOOST_cell_45169 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__Q), .b(n_3542), .o(TIMEBOOST_net_14823) );
in01s01 g64914_u0 ( .a(FE_OFN622_n_4409), .o(g64914_sb) );
na02s02 TIMEBOOST_cell_31365 ( .a(TIMEBOOST_net_9593), .b(FE_OFN254_n_9825), .o(n_9702) );
na02s01 g64914_u2 ( .a(n_4396), .b(FE_OFN622_n_4409), .o(g64914_db) );
na02s01 TIMEBOOST_cell_16426 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__Q), .b(g64333_sb), .o(TIMEBOOST_net_3470) );
in01s01 g64915_u0 ( .a(FE_OFN624_n_4409), .o(g64915_sb) );
na02f02 TIMEBOOST_cell_38572 ( .a(TIMEBOOST_net_11524), .b(TIMEBOOST_net_869), .o(g54039_da) );
na02s01 g64915_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__Q), .b(FE_OFN624_n_4409), .o(g64915_db) );
na02s01 TIMEBOOST_cell_15948 ( .a(pci_target_unit_fifos_pcir_data_in_172), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__Q), .o(TIMEBOOST_net_3231) );
in01s01 g64916_u0 ( .a(FE_OFN622_n_4409), .o(g64916_sb) );
na02s01 TIMEBOOST_cell_15949 ( .a(TIMEBOOST_net_3231), .b(FE_OFN946_n_2248), .o(TIMEBOOST_net_1172) );
na02s02 TIMEBOOST_cell_45192 ( .a(TIMEBOOST_net_14834), .b(FE_OFN1253_n_4143), .o(TIMEBOOST_net_12074) );
in01s01 g64917_u0 ( .a(FE_OFN1663_n_4490), .o(g64917_sb) );
na02s01 TIMEBOOST_cell_31172 ( .a(n_3777), .b(g64859_sb), .o(TIMEBOOST_net_9497) );
na02s01 g64917_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__15__Q), .b(FE_OFN1663_n_4490), .o(g64917_db) );
na02s01 TIMEBOOST_cell_31171 ( .a(TIMEBOOST_net_9496), .b(g64851_db), .o(n_3722) );
in01s01 g64918_u0 ( .a(FE_OFN662_n_4392), .o(g64918_sb) );
na02s02 TIMEBOOST_cell_43379 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q), .b(n_3576), .o(TIMEBOOST_net_13928) );
na02f02 TIMEBOOST_cell_44110 ( .a(TIMEBOOST_net_14293), .b(FE_OFN1420_n_8567), .o(TIMEBOOST_net_12915) );
na02s02 TIMEBOOST_cell_43380 ( .a(TIMEBOOST_net_13928), .b(n_6287), .o(TIMEBOOST_net_12171) );
in01s01 g64919_u0 ( .a(FE_OFN1810_n_4454), .o(g64919_sb) );
na02f02 TIMEBOOST_cell_44470 ( .a(TIMEBOOST_net_14473), .b(FE_OFN2167_n_8567), .o(TIMEBOOST_net_13436) );
na02s01 g64919_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__Q), .b(FE_OFN1810_n_4454), .o(g64919_db) );
na02f02 TIMEBOOST_cell_40112 ( .a(TIMEBOOST_net_12294), .b(g57560_sb), .o(n_10298) );
in01s01 g64920_u0 ( .a(FE_OFN618_n_4490), .o(g64920_sb) );
na02m02 TIMEBOOST_cell_38483 ( .a(TIMEBOOST_net_2048), .b(TIMEBOOST_net_9981), .o(TIMEBOOST_net_11480) );
na02f02 TIMEBOOST_cell_39539 ( .a(n_2918), .b(n_2846), .o(TIMEBOOST_net_12008) );
na03s02 TIMEBOOST_cell_38153 ( .a(TIMEBOOST_net_3552), .b(g64362_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__Q), .o(TIMEBOOST_net_11315) );
in01s01 g64921_u0 ( .a(FE_OFN660_n_4392), .o(g64921_sb) );
na02f02 TIMEBOOST_cell_44618 ( .a(TIMEBOOST_net_14547), .b(FE_OFN2185_n_8567), .o(TIMEBOOST_net_13005) );
na02s01 g64921_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__Q), .b(FE_OFN660_n_4392), .o(g64921_db) );
na02s01 TIMEBOOST_cell_16695 ( .a(TIMEBOOST_net_3604), .b(g64917_db), .o(n_3686) );
in01s01 g64922_u0 ( .a(FE_OFN660_n_4392), .o(g64922_sb) );
na02s01 TIMEBOOST_cell_45077 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__Q), .b(FE_OFN881_g64577_p), .o(TIMEBOOST_net_14777) );
na02s01 g64922_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__Q), .b(FE_OFN660_n_4392), .o(g64922_db) );
na02s01 TIMEBOOST_cell_16428 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__Q), .b(g64334_sb), .o(TIMEBOOST_net_3471) );
in01s01 g64923_u0 ( .a(FE_OFN661_n_4392), .o(g64923_sb) );
na02s02 TIMEBOOST_cell_45170 ( .a(TIMEBOOST_net_14823), .b(FE_OFN1285_n_4097), .o(TIMEBOOST_net_12022) );
na02m02 TIMEBOOST_cell_44111 ( .a(n_9483), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q), .o(TIMEBOOST_net_14294) );
na02s02 TIMEBOOST_cell_43447 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__Q), .b(n_4401), .o(TIMEBOOST_net_13962) );
in01s01 g64924_u0 ( .a(FE_OFN660_n_4392), .o(g64924_sb) );
na03s02 TIMEBOOST_cell_38109 ( .a(TIMEBOOST_net_4241), .b(g64212_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__28__Q), .o(TIMEBOOST_net_11293) );
na02s02 TIMEBOOST_cell_40752 ( .a(TIMEBOOST_net_12614), .b(g62338_sb), .o(n_6922) );
na03s02 TIMEBOOST_cell_38421 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__Q), .b(FE_OFN1124_g64577_p), .c(n_3213), .o(TIMEBOOST_net_11449) );
in01s01 g64925_u0 ( .a(FE_OFN619_n_4490), .o(g64925_sb) );
na02s01 TIMEBOOST_cell_31170 ( .a(n_3785), .b(g64851_sb), .o(TIMEBOOST_net_9496) );
na02s01 g64925_u2 ( .a(n_38), .b(FE_OFN619_n_4490), .o(g64925_db) );
na04m02 TIMEBOOST_cell_34480 ( .a(n_3485), .b(g52397_sb), .c(g52397_db), .d(TIMEBOOST_net_588), .o(n_14824) );
in01s01 g64926_u0 ( .a(FE_OFN662_n_4392), .o(g64926_sb) );
na02s01 TIMEBOOST_cell_16430 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__Q), .b(g64335_sb), .o(TIMEBOOST_net_3472) );
na02s02 g64926_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__Q), .b(FE_OFN662_n_4392), .o(g64926_db) );
na02s02 TIMEBOOST_cell_45171 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__Q), .b(n_4455), .o(TIMEBOOST_net_14824) );
in01s01 g64927_u0 ( .a(FE_OFN662_n_4392), .o(g64927_sb) );
na02s02 TIMEBOOST_cell_45710 ( .a(TIMEBOOST_net_15093), .b(FE_OFN1218_n_6886), .o(TIMEBOOST_net_12541) );
na02s01 g64927_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__Q), .b(FE_OFN662_n_4392), .o(g64927_db) );
na02m02 TIMEBOOST_cell_44619 ( .a(n_9711), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__Q), .o(TIMEBOOST_net_14548) );
in01s01 g64928_u0 ( .a(FE_OFN661_n_4392), .o(g64928_sb) );
na02m02 TIMEBOOST_cell_44471 ( .a(n_9874), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__Q), .o(TIMEBOOST_net_14474) );
na02s01 g64928_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__Q), .b(FE_OFN661_n_4392), .o(g64928_db) );
na02s02 TIMEBOOST_cell_43381 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__14__Q), .b(n_4240), .o(TIMEBOOST_net_13929) );
in01s01 g64929_u0 ( .a(FE_OFN661_n_4392), .o(g64929_sb) );
na02m02 TIMEBOOST_cell_41592 ( .a(FE_OFN1439_n_9372), .b(TIMEBOOST_net_13034), .o(TIMEBOOST_net_11667) );
na02s01 g64929_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__Q), .b(FE_OFN661_n_4392), .o(g64929_db) );
na02s01 TIMEBOOST_cell_31363 ( .a(TIMEBOOST_net_9592), .b(FE_OFN241_n_9830), .o(n_9729) );
in01s01 g64930_u0 ( .a(FE_OFN660_n_4392), .o(g64930_sb) );
na02s02 TIMEBOOST_cell_43382 ( .a(TIMEBOOST_net_13929), .b(n_6232), .o(TIMEBOOST_net_12170) );
na02s01 g64930_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__Q), .b(FE_OFN660_n_4392), .o(g64930_db) );
na02s02 TIMEBOOST_cell_42098 ( .a(TIMEBOOST_net_13287), .b(g62982_sb), .o(n_5918) );
in01s01 g64931_u0 ( .a(FE_OFN659_n_4392), .o(g64931_sb) );
na02s01 TIMEBOOST_cell_36660 ( .a(TIMEBOOST_net_10568), .b(g65892_sb), .o(n_2587) );
na02s01 g64931_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__Q), .b(FE_OFN659_n_4392), .o(g64931_db) );
na02f02 TIMEBOOST_cell_40114 ( .a(TIMEBOOST_net_12295), .b(g57159_sb), .o(n_11590) );
in01s01 g64932_u0 ( .a(FE_OFN660_n_4392), .o(g64932_sb) );
na02f02 TIMEBOOST_cell_44472 ( .a(TIMEBOOST_net_14474), .b(FE_OFN2179_n_8567), .o(TIMEBOOST_net_13437) );
na02s01 g64932_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__26__Q), .b(FE_OFN660_n_4392), .o(g64932_db) );
na02f02 TIMEBOOST_cell_40116 ( .a(TIMEBOOST_net_12296), .b(g57277_sb), .o(n_11477) );
in01s01 g64933_u0 ( .a(FE_OFN664_n_4495), .o(g64933_sb) );
na02m02 TIMEBOOST_cell_44473 ( .a(n_9411), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__Q), .o(TIMEBOOST_net_14475) );
na02s01 g64933_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__Q), .b(FE_OFN664_n_4495), .o(g64933_db) );
na02f02 TIMEBOOST_cell_40118 ( .a(TIMEBOOST_net_12297), .b(g57176_sb), .o(n_11579) );
in01s01 g64934_u0 ( .a(FE_OFN660_n_4392), .o(g64934_sb) );
na02f02 TIMEBOOST_cell_44474 ( .a(TIMEBOOST_net_14475), .b(FE_OFN2184_n_8567), .o(TIMEBOOST_net_13438) );
na02s01 g64934_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__Q), .b(FE_OFN660_n_4392), .o(g64934_db) );
na02f02 TIMEBOOST_cell_40120 ( .a(TIMEBOOST_net_12298), .b(g57246_sb), .o(n_11510) );
in01s01 g64935_u0 ( .a(FE_OFN661_n_4392), .o(g64935_sb) );
na02s02 TIMEBOOST_cell_36663 ( .a(TIMEBOOST_net_9562), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_10570) );
na02s01 g64935_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__Q), .b(FE_OFN661_n_4392), .o(g64935_db) );
na02m02 TIMEBOOST_cell_44475 ( .a(n_9572), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__Q), .o(TIMEBOOST_net_14476) );
in01s01 g64936_u0 ( .a(FE_OFN661_n_4392), .o(g64936_sb) );
na02s01 TIMEBOOST_cell_36662 ( .a(TIMEBOOST_net_10569), .b(g65892_sb), .o(n_2592) );
na02f02 TIMEBOOST_cell_44112 ( .a(TIMEBOOST_net_14294), .b(FE_OFN1409_n_8567), .o(TIMEBOOST_net_12753) );
na02s02 TIMEBOOST_cell_31357 ( .a(TIMEBOOST_net_9589), .b(g65329_da), .o(n_4266) );
in01s01 g64937_u0 ( .a(FE_OFN659_n_4392), .o(g64937_sb) );
na02f02 TIMEBOOST_cell_40122 ( .a(TIMEBOOST_net_12299), .b(g57269_sb), .o(n_11483) );
na02s01 g64937_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__Q), .b(FE_OFN659_n_4392), .o(g64937_db) );
na02f02 TIMEBOOST_cell_44476 ( .a(TIMEBOOST_net_14476), .b(FE_OFN2190_n_8567), .o(TIMEBOOST_net_13439) );
in01s01 g64938_u0 ( .a(FE_OFN659_n_4392), .o(g64938_sb) );
na02s02 TIMEBOOST_cell_31356 ( .a(n_4476), .b(FE_OFN653_n_4508), .o(TIMEBOOST_net_9589) );
na02s01 g64938_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__Q), .b(FE_OFN659_n_4392), .o(g64938_db) );
na02s01 TIMEBOOST_cell_31355 ( .a(TIMEBOOST_net_9588), .b(g65271_da), .o(n_4293) );
in01s01 g64939_u0 ( .a(FE_OFN659_n_4392), .o(g64939_sb) );
na02f02 TIMEBOOST_cell_40124 ( .a(TIMEBOOST_net_12300), .b(g57062_sb), .o(n_11677) );
na02s01 TIMEBOOST_cell_31354 ( .a(n_4465), .b(FE_OFN652_n_4508), .o(TIMEBOOST_net_9588) );
in01s01 g64940_u0 ( .a(FE_OFN659_n_4392), .o(g64940_sb) );
na02s01 TIMEBOOST_cell_16444 ( .a(n_3752), .b(g64849_sb), .o(TIMEBOOST_net_3479) );
na02s01 g64940_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__Q), .b(FE_OFN660_n_4392), .o(g64940_db) );
na02s01 TIMEBOOST_cell_16445 ( .a(TIMEBOOST_net_3479), .b(g64849_db), .o(n_3723) );
in01s01 g64941_u0 ( .a(FE_OFN649_n_4497), .o(g64941_sb) );
na02s02 TIMEBOOST_cell_45172 ( .a(TIMEBOOST_net_14824), .b(FE_OFN1208_n_6356), .o(TIMEBOOST_net_12211) );
na02s01 g64941_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__Q), .b(FE_OFN649_n_4497), .o(g64941_db) );
na02f02 TIMEBOOST_cell_40126 ( .a(TIMEBOOST_net_12301), .b(g57495_sb), .o(n_11242) );
in01s01 g64942_u0 ( .a(FE_OFN646_n_4497), .o(g64942_sb) );
na02s01 TIMEBOOST_cell_40323 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__Q), .b(g58453_sb), .o(TIMEBOOST_net_12400) );
na02s01 g64942_u2 ( .a(n_3672), .b(FE_OFN646_n_4497), .o(g64942_db) );
na02f02 TIMEBOOST_cell_40128 ( .a(TIMEBOOST_net_12302), .b(g57358_sb), .o(n_11390) );
in01s01 g64943_u0 ( .a(FE_OFN648_n_4497), .o(g64943_sb) );
na02s01 TIMEBOOST_cell_17082 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__Q), .b(g65967_sb), .o(TIMEBOOST_net_3798) );
na02s01 TIMEBOOST_cell_42771 ( .a(FE_OFN215_n_9856), .b(g57983_sb), .o(TIMEBOOST_net_13624) );
na02f02 TIMEBOOST_cell_44652 ( .a(TIMEBOOST_net_14564), .b(FE_OFN2180_n_8567), .o(TIMEBOOST_net_13486) );
in01s01 g64944_u0 ( .a(FE_OFN649_n_4497), .o(g64944_sb) );
na02m02 TIMEBOOST_cell_44477 ( .a(n_9686), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__Q), .o(TIMEBOOST_net_14477) );
na02s01 g64944_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__Q), .b(FE_OFN649_n_4497), .o(g64944_db) );
na02f02 TIMEBOOST_cell_40130 ( .a(TIMEBOOST_net_12303), .b(g58574_sb), .o(n_9194) );
in01s01 g64945_u0 ( .a(FE_OFN649_n_4497), .o(g64945_sb) );
na02s01 TIMEBOOST_cell_9018 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__Q), .o(TIMEBOOST_net_1076) );
na02s01 g64945_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__Q), .b(FE_OFN649_n_4497), .o(g64945_db) );
na02s01 TIMEBOOST_cell_9019 ( .a(TIMEBOOST_net_1076), .b(n_2299), .o(TIMEBOOST_net_117) );
in01s01 g64946_u0 ( .a(FE_OFN649_n_4497), .o(g64946_sb) );
na02s01 TIMEBOOST_cell_9020 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__Q), .o(TIMEBOOST_net_1077) );
na02s01 g64946_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__1__Q), .b(FE_OFN649_n_4497), .o(g64946_db) );
na02s01 TIMEBOOST_cell_9021 ( .a(TIMEBOOST_net_1077), .b(n_2299), .o(TIMEBOOST_net_118) );
in01s01 g64947_u0 ( .a(FE_OFN649_n_4497), .o(g64947_sb) );
na02s01 TIMEBOOST_cell_9022 ( .a(pci_target_unit_fifos_pcir_data_in_165), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q), .o(TIMEBOOST_net_1078) );
na02s01 g64947_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__Q), .b(FE_OFN649_n_4497), .o(g64947_db) );
na02s01 TIMEBOOST_cell_9023 ( .a(TIMEBOOST_net_1078), .b(n_2299), .o(TIMEBOOST_net_119) );
in01s01 g64948_u0 ( .a(FE_OFN649_n_4497), .o(g64948_sb) );
na02s01 g64948_u1 ( .a(n_3749), .b(g64948_sb), .o(g64948_da) );
na02s01 g64948_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__Q), .b(FE_OFN649_n_4497), .o(g64948_db) );
na02s01 g64948_u3 ( .a(g64948_da), .b(g64948_db), .o(n_3668) );
in01s01 g64949_u0 ( .a(FE_OFN647_n_4497), .o(g64949_sb) );
na02s01 TIMEBOOST_cell_9024 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__Q), .o(TIMEBOOST_net_1079) );
na02s01 g64949_u2 ( .a(n_65), .b(FE_OFN647_n_4497), .o(g64949_db) );
na02m02 TIMEBOOST_cell_45110 ( .a(TIMEBOOST_net_14793), .b(TIMEBOOST_net_9670), .o(TIMEBOOST_net_4766) );
in01s01 g64950_u0 ( .a(FE_OFN647_n_4497), .o(g64950_sb) );
na02s01 TIMEBOOST_cell_44986 ( .a(TIMEBOOST_net_14731), .b(g63614_db), .o(TIMEBOOST_net_13154) );
na02s01 g64950_u2 ( .a(n_3665), .b(FE_OFN647_n_4497), .o(g64950_db) );
na02f02 TIMEBOOST_cell_40132 ( .a(TIMEBOOST_net_12304), .b(g57238_sb), .o(n_10430) );
in01s01 g64951_u0 ( .a(FE_OFN649_n_4497), .o(g64951_sb) );
na02s01 TIMEBOOST_cell_16926 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__Q), .b(g65339_sb), .o(TIMEBOOST_net_3720) );
na02s01 g64951_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__Q), .b(FE_OFN649_n_4497), .o(g64951_db) );
na02s01 TIMEBOOST_cell_16927 ( .a(TIMEBOOST_net_3720), .b(g65339_db), .o(n_3549) );
in01s01 g64952_u0 ( .a(FE_OFN646_n_4497), .o(g64952_sb) );
na02m02 TIMEBOOST_cell_9030 ( .a(n_15924), .b(n_2078), .o(TIMEBOOST_net_1082) );
na02s01 g64952_u2 ( .a(n_74), .b(FE_OFN646_n_4497), .o(g64952_db) );
na02f02 TIMEBOOST_cell_9031 ( .a(TIMEBOOST_net_1082), .b(n_15923), .o(TIMEBOOST_net_121) );
in01s01 g64953_u0 ( .a(n_4460), .o(g64953_sb) );
na03s02 TIMEBOOST_cell_33148 ( .a(wbu_addr_in_277), .b(g58787_sb), .c(TIMEBOOST_net_3649), .o(n_9836) );
na02s01 g64953_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__Q), .b(n_4460), .o(g64953_db) );
na02s02 TIMEBOOST_cell_43068 ( .a(TIMEBOOST_net_13772), .b(FE_OFN1216_n_4151), .o(TIMEBOOST_net_12027) );
in01s01 g64954_u0 ( .a(FE_OFN649_n_4497), .o(g64954_sb) );
na02s01 TIMEBOOST_cell_17006 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(g65727_sb), .o(TIMEBOOST_net_3760) );
na02s01 g64954_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__Q), .b(FE_OFN649_n_4497), .o(g64954_db) );
na02s02 TIMEBOOST_cell_36722 ( .a(TIMEBOOST_net_10599), .b(g63616_sb), .o(TIMEBOOST_net_9823) );
in01s01 g64955_u0 ( .a(FE_OFN648_n_4497), .o(g64955_sb) );
na02f02 TIMEBOOST_cell_44478 ( .a(TIMEBOOST_net_14477), .b(FE_OFN2179_n_8567), .o(TIMEBOOST_net_13440) );
na02s02 TIMEBOOST_cell_43448 ( .a(TIMEBOOST_net_13962), .b(FE_OFN1233_n_6391), .o(TIMEBOOST_net_12151) );
na02f02 TIMEBOOST_cell_40134 ( .a(TIMEBOOST_net_12305), .b(g57206_sb), .o(n_11551) );
in01s01 g64956_u0 ( .a(FE_OFN648_n_4497), .o(g64956_sb) );
na02s01 TIMEBOOST_cell_39279 ( .a(pci_target_unit_fifos_pcir_data_in_174), .b(g65791_sb), .o(TIMEBOOST_net_11878) );
na02s01 g64956_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__Q), .b(FE_OFN648_n_4497), .o(g64956_db) );
na02s01 TIMEBOOST_cell_39280 ( .a(TIMEBOOST_net_11878), .b(g65791_db), .o(n_1595) );
in01s01 g64957_u0 ( .a(FE_OFN646_n_4497), .o(g64957_sb) );
na02s01 TIMEBOOST_cell_39281 ( .a(pci_target_unit_fifos_pcir_data_in_173), .b(g65793_sb), .o(TIMEBOOST_net_11879) );
na02s01 g64957_u2 ( .a(n_40), .b(FE_OFN646_n_4497), .o(g64957_db) );
na02s01 TIMEBOOST_cell_39282 ( .a(TIMEBOOST_net_11879), .b(g65793_db), .o(n_1593) );
in01s01 g64958_u0 ( .a(FE_OFN646_n_4497), .o(g64958_sb) );
na03f02 TIMEBOOST_cell_35325 ( .a(TIMEBOOST_net_10050), .b(FE_OFN1369_n_8567), .c(g58617_sb), .o(n_9185) );
na02s01 g64958_u2 ( .a(n_119), .b(FE_OFN646_n_4497), .o(g64958_db) );
na02f02 TIMEBOOST_cell_44113 ( .a(n_9132), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__Q), .o(TIMEBOOST_net_14295) );
in01s01 g64959_u0 ( .a(FE_OFN612_n_4501), .o(g64959_sb) );
na02s01 TIMEBOOST_cell_31169 ( .a(TIMEBOOST_net_9495), .b(g64837_db), .o(n_3728) );
na02s01 g64959_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__Q), .b(FE_OFN612_n_4501), .o(g64959_db) );
na02s02 TIMEBOOST_cell_31168 ( .a(n_3785), .b(g64837_sb), .o(TIMEBOOST_net_9495) );
in01s01 g64960_u0 ( .a(FE_OFN612_n_4501), .o(g64960_sb) );
na02s01 g64960_u1 ( .a(n_3783), .b(g64960_sb), .o(g64960_da) );
na02s01 g64960_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__Q), .b(FE_OFN612_n_4501), .o(g64960_db) );
na02s01 g64960_u3 ( .a(g64960_da), .b(g64960_db), .o(n_3658) );
in01s01 g64961_u0 ( .a(FE_OFN614_n_4501), .o(g64961_sb) );
na02s02 TIMEBOOST_cell_31167 ( .a(TIMEBOOST_net_9494), .b(g64811_sb), .o(n_3746) );
na02s01 g64961_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__Q), .b(FE_OFN614_n_4501), .o(g64961_db) );
na02f02 TIMEBOOST_cell_44114 ( .a(TIMEBOOST_net_14295), .b(FE_OFN1397_n_8567), .o(TIMEBOOST_net_12705) );
in01s01 g64962_u0 ( .a(FE_OFN615_n_4501), .o(g64962_sb) );
na02f04 TIMEBOOST_cell_39050 ( .a(TIMEBOOST_net_11763), .b(FE_OFN2242_g52675_p), .o(TIMEBOOST_net_10752) );
na02f02 TIMEBOOST_cell_39052 ( .a(TIMEBOOST_net_11764), .b(g52600_db), .o(n_11871) );
in01s01 g64963_u0 ( .a(FE_OFN618_n_4490), .o(g64963_sb) );
na02s01 TIMEBOOST_cell_31165 ( .a(TIMEBOOST_net_9493), .b(g65302_db), .o(n_3574) );
na02s01 g64963_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__Q), .b(FE_OFN618_n_4490), .o(g64963_db) );
na02s01 TIMEBOOST_cell_31164 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__Q), .b(g65302_sb), .o(TIMEBOOST_net_9493) );
na02m02 TIMEBOOST_cell_44479 ( .a(n_9086), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__Q), .o(TIMEBOOST_net_14478) );
na02s01 g64964_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__Q), .b(FE_OFN679_n_4460), .o(g64964_db) );
na02f02 TIMEBOOST_cell_40136 ( .a(TIMEBOOST_net_12306), .b(g57240_sb), .o(n_10426) );
in01s01 g64965_u0 ( .a(FE_OFN1807_n_4501), .o(g64965_sb) );
na02s02 TIMEBOOST_cell_17990 ( .a(pci_target_unit_fifos_pciw_addr_data_in_130), .b(g64086_sb), .o(TIMEBOOST_net_4252) );
na02s01 TIMEBOOST_cell_36472 ( .a(TIMEBOOST_net_10474), .b(g65770_db), .o(n_1913) );
na02f01 TIMEBOOST_cell_38467 ( .a(TIMEBOOST_net_828), .b(n_16452), .o(TIMEBOOST_net_11472) );
in01s01 g64966_u0 ( .a(FE_OFN665_n_4495), .o(g64966_sb) );
na02s01 TIMEBOOST_cell_16123 ( .a(TIMEBOOST_net_3318), .b(FE_OFN2095_n_2520), .o(TIMEBOOST_net_1303) );
na02s01 g64966_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__Q), .b(FE_OFN665_n_4495), .o(g64966_db) );
na02s01 TIMEBOOST_cell_16124 ( .a(parchk_pci_ad_reg_in_1218), .b(pci_target_unit_del_sync_addr_in_217), .o(TIMEBOOST_net_3319) );
in01s01 g64967_u0 ( .a(FE_OFN619_n_4490), .o(g64967_sb) );
na02s01 TIMEBOOST_cell_31163 ( .a(TIMEBOOST_net_9492), .b(g65098_db), .o(n_3595) );
na02s01 g64967_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__Q), .b(FE_OFN619_n_4490), .o(g64967_db) );
na02s01 TIMEBOOST_cell_31162 ( .a(n_3739), .b(g65098_sb), .o(TIMEBOOST_net_9492) );
in01s01 g64968_u0 ( .a(FE_OFN618_n_4490), .o(g64968_sb) );
na02s01 TIMEBOOST_cell_31161 ( .a(TIMEBOOST_net_9491), .b(g64780_db), .o(n_3771) );
na02s01 g64968_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q), .b(FE_OFN1663_n_4490), .o(g64968_db) );
na02s01 TIMEBOOST_cell_31160 ( .a(n_3770), .b(g64780_sb), .o(TIMEBOOST_net_9491) );
in01s01 g64969_u0 ( .a(FE_OFN615_n_4501), .o(g64969_sb) );
na02s01 TIMEBOOST_cell_31159 ( .a(TIMEBOOST_net_9490), .b(g64777_db), .o(n_3772) );
na02s01 g64969_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__Q), .b(FE_OFN615_n_4501), .o(g64969_db) );
na02s01 TIMEBOOST_cell_31158 ( .a(n_3785), .b(g64777_sb), .o(TIMEBOOST_net_9490) );
in01s01 g64970_u0 ( .a(FE_OFN667_n_4495), .o(g64970_sb) );
na02f02 TIMEBOOST_cell_44480 ( .a(TIMEBOOST_net_14478), .b(FE_OFN2168_n_8567), .o(TIMEBOOST_net_13441) );
na02s01 g64970_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__Q), .b(FE_OFN667_n_4495), .o(g64970_db) );
na02f02 TIMEBOOST_cell_40138 ( .a(TIMEBOOST_net_12307), .b(g57041_sb), .o(n_11693) );
in01s01 g64971_u0 ( .a(FE_OFN615_n_4501), .o(g64971_sb) );
na02s02 TIMEBOOST_cell_31157 ( .a(TIMEBOOST_net_9489), .b(g65074_sb), .o(n_3605) );
na02s01 g64971_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q), .b(FE_OFN615_n_4501), .o(g64971_db) );
na02s01 TIMEBOOST_cell_43449 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__Q), .b(n_3708), .o(TIMEBOOST_net_13963) );
in01s01 g64972_u0 ( .a(FE_OFN1807_n_4501), .o(g64972_sb) );
na02s02 TIMEBOOST_cell_17992 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(g64115_sb), .o(TIMEBOOST_net_4253) );
na02s01 TIMEBOOST_cell_39283 ( .a(pci_target_unit_fifos_pcir_data_in_178), .b(g65724_sb), .o(TIMEBOOST_net_11880) );
in01s01 TIMEBOOST_cell_45936 ( .a(TIMEBOOST_net_15242), .o(TIMEBOOST_net_15243) );
in01s01 g64973_u0 ( .a(FE_OFN1807_n_4501), .o(g64973_sb) );
na02s02 TIMEBOOST_cell_17994 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(g64140_sb), .o(TIMEBOOST_net_4254) );
na02s01 TIMEBOOST_cell_36474 ( .a(TIMEBOOST_net_10475), .b(g65715_sb), .o(n_1918) );
na03s02 TIMEBOOST_cell_38325 ( .a(n_3876), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q), .c(FE_OFN1119_g64577_p), .o(TIMEBOOST_net_11401) );
in01s01 g64974_u0 ( .a(FE_OFN647_n_4497), .o(g64974_sb) );
na02s01 g64974_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__31__Q), .b(FE_OFN647_n_4497), .o(g64974_db) );
na02s02 TIMEBOOST_cell_40754 ( .a(TIMEBOOST_net_12615), .b(g62355_sb), .o(n_6889) );
in01s01 g64975_u0 ( .a(FE_OFN622_n_4409), .o(g64975_sb) );
na02s02 TIMEBOOST_cell_16448 ( .a(n_3783), .b(g64857_sb), .o(TIMEBOOST_net_3481) );
na02s01 g64975_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__Q), .b(FE_OFN622_n_4409), .o(g64975_db) );
na02s02 TIMEBOOST_cell_16449 ( .a(TIMEBOOST_net_3481), .b(g64857_db), .o(n_3719) );
in01s01 g64976_u0 ( .a(FE_OFN615_n_4501), .o(g64976_sb) );
na02f02 TIMEBOOST_cell_44278 ( .a(TIMEBOOST_net_14377), .b(FE_OFN1417_n_8567), .o(TIMEBOOST_net_12691) );
na02s01 g64976_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__Q), .b(FE_OFN615_n_4501), .o(g64976_db) );
na02s02 TIMEBOOST_cell_43450 ( .a(TIMEBOOST_net_13963), .b(FE_OFN1232_n_6391), .o(TIMEBOOST_net_12179) );
in01s01 g64977_u0 ( .a(FE_OFN1623_n_4438), .o(g64977_sb) );
na02s01 TIMEBOOST_cell_31353 ( .a(TIMEBOOST_net_9587), .b(g65370_da), .o(n_4519) );
na02s01 g64977_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__Q), .b(FE_OFN1623_n_4438), .o(g64977_db) );
na02s02 TIMEBOOST_cell_16450 ( .a(n_3741), .b(g64888_sb), .o(TIMEBOOST_net_3482) );
in01s01 g64978_u0 ( .a(FE_OFN665_n_4495), .o(g64978_sb) );
na02s02 TIMEBOOST_cell_16451 ( .a(TIMEBOOST_net_3482), .b(g64888_db), .o(n_3702) );
na02s01 g64978_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__Q), .b(FE_OFN665_n_4495), .o(g64978_db) );
na02s01 TIMEBOOST_cell_16452 ( .a(n_3755), .b(g64895_sb), .o(TIMEBOOST_net_3483) );
in01s01 g64979_u0 ( .a(FE_OFN619_n_4490), .o(g64979_sb) );
na02s02 TIMEBOOST_cell_43451 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__Q), .b(n_4229), .o(TIMEBOOST_net_13964) );
na02s01 g64979_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__Q), .b(FE_OFN619_n_4490), .o(g64979_db) );
na02m02 TIMEBOOST_cell_44115 ( .a(n_9637), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__Q), .o(TIMEBOOST_net_14296) );
in01s01 g64980_u0 ( .a(FE_OFN685_n_4417), .o(g64980_sb) );
na02s01 TIMEBOOST_cell_16453 ( .a(TIMEBOOST_net_3483), .b(g64895_db), .o(n_3698) );
na02s01 g64980_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q), .b(FE_OFN685_n_4417), .o(g64980_db) );
na02s01 TIMEBOOST_cell_16454 ( .a(FE_OFN223_n_9844), .b(g57927_sb), .o(TIMEBOOST_net_3484) );
na02s01 TIMEBOOST_cell_9305 ( .a(TIMEBOOST_net_1219), .b(g65790_db), .o(n_1596) );
na02s01 g64981_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__0__Q), .b(n_4501), .o(g64981_db) );
na02m02 TIMEBOOST_cell_40550 ( .a(TIMEBOOST_net_12513), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_11554) );
in01s01 g64982_u0 ( .a(FE_OFN1624_n_4438), .o(g64982_sb) );
na02s01 TIMEBOOST_cell_16455 ( .a(TIMEBOOST_net_3484), .b(g57927_db), .o(n_9882) );
na02s01 g64982_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__8__Q), .b(FE_OFN1624_n_4438), .o(g64982_db) );
na02s02 TIMEBOOST_cell_45526 ( .a(TIMEBOOST_net_15001), .b(g61958_sb), .o(n_6956) );
in01s01 g64983_u0 ( .a(FE_OFN647_n_4497), .o(g64983_sb) );
na02m02 TIMEBOOST_cell_44481 ( .a(n_9565), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__Q), .o(TIMEBOOST_net_14479) );
na02s01 g64983_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__Q), .b(FE_OFN647_n_4497), .o(g64983_db) );
na02f02 TIMEBOOST_cell_40140 ( .a(TIMEBOOST_net_12308), .b(g57360_sb), .o(n_11386) );
in01s01 g64984_u0 ( .a(FE_OFN649_n_4497), .o(g64984_sb) );
na02s01 g64984_u1 ( .a(n_3761), .b(g64984_sb), .o(g64984_da) );
na02s01 g64984_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__Q), .b(FE_OFN649_n_4497), .o(g64984_db) );
na02s01 TIMEBOOST_cell_39259 ( .a(pci_target_unit_fifos_pciw_cbe_in), .b(g64186_sb), .o(TIMEBOOST_net_11868) );
in01s01 g64985_u0 ( .a(FE_OFN1628_n_4438), .o(g64985_sb) );
na02s02 TIMEBOOST_cell_36774 ( .a(TIMEBOOST_net_10625), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_1997) );
na02s01 g64985_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__Q), .b(FE_OFN1628_n_4438), .o(g64985_db) );
na02s01 TIMEBOOST_cell_17819 ( .a(TIMEBOOST_net_4166), .b(g61816_sb), .o(n_8159) );
in01s01 g64986_u0 ( .a(FE_OFN667_n_4495), .o(g64986_sb) );
na02s01 TIMEBOOST_cell_16125 ( .a(TIMEBOOST_net_3319), .b(FE_OFN2095_n_2520), .o(TIMEBOOST_net_1308) );
na02s01 g64986_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__Q), .b(FE_OFN667_n_4495), .o(g64986_db) );
na02s01 TIMEBOOST_cell_16126 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__Q), .b(pci_target_unit_fifos_pcir_data_in_164), .o(TIMEBOOST_net_3320) );
in01s01 g64987_u0 ( .a(FE_OFN689_n_4438), .o(g64987_sb) );
na02f02 TIMEBOOST_cell_40142 ( .a(TIMEBOOST_net_12309), .b(g57531_sb), .o(n_11211) );
na02s01 g64987_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__Q), .b(FE_OFN689_n_4438), .o(g64987_db) );
na02f02 TIMEBOOST_cell_44482 ( .a(TIMEBOOST_net_14479), .b(FE_OFN2170_n_8567), .o(TIMEBOOST_net_13442) );
in01s01 g64988_u0 ( .a(FE_OFN646_n_4497), .o(g64988_sb) );
na02m02 TIMEBOOST_cell_44397 ( .a(n_9800), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__Q), .o(TIMEBOOST_net_14437) );
na02s01 g64988_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__Q), .b(FE_OFN646_n_4497), .o(g64988_db) );
na02s01 TIMEBOOST_cell_40552 ( .a(TIMEBOOST_net_12514), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_11556) );
in01s01 g64989_u0 ( .a(FE_OFN684_n_4417), .o(g64989_sb) );
na02f02 TIMEBOOST_cell_40144 ( .a(TIMEBOOST_net_12310), .b(g57428_sb), .o(n_11306) );
na02s01 g64989_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__Q), .b(FE_OFN684_n_4417), .o(g64989_db) );
na02m02 TIMEBOOST_cell_44483 ( .a(n_9209), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__Q), .o(TIMEBOOST_net_14480) );
in01s01 g64990_u0 ( .a(FE_OFN1625_n_4438), .o(g64990_sb) );
na02f02 TIMEBOOST_cell_44484 ( .a(TIMEBOOST_net_14480), .b(FE_OFN2177_n_8567), .o(TIMEBOOST_net_13443) );
na02s01 g64990_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__Q), .b(FE_OFN1625_n_4438), .o(g64990_db) );
na02f02 TIMEBOOST_cell_40146 ( .a(TIMEBOOST_net_12311), .b(g57351_sb), .o(n_11398) );
in01s01 g64991_u0 ( .a(FE_OFN1628_n_4438), .o(g64991_sb) );
in01s01 TIMEBOOST_cell_45885 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_), .o(TIMEBOOST_net_15192) );
na02s01 g64991_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__Q), .b(FE_OFN1628_n_4438), .o(g64991_db) );
na03f02 TIMEBOOST_cell_36137 ( .a(n_16234), .b(n_16237), .c(n_16239), .o(n_16240) );
in01s01 g64992_u0 ( .a(FE_OFN659_n_4392), .o(g64992_sb) );
na02f02 TIMEBOOST_cell_40148 ( .a(TIMEBOOST_net_12312), .b(g57347_sb), .o(n_11403) );
na02s01 g64992_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__Q), .b(FE_OFN659_n_4392), .o(g64992_db) );
na02s01 TIMEBOOST_cell_31352 ( .a(n_4498), .b(FE_OFN1644_n_4671), .o(TIMEBOOST_net_9587) );
in01s01 g64993_u0 ( .a(FE_OFN1624_n_4438), .o(g64993_sb) );
na02s01 TIMEBOOST_cell_16462 ( .a(n_3752), .b(g64928_sb), .o(TIMEBOOST_net_3488) );
na02s01 g64993_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q), .b(FE_OFN1624_n_4438), .o(g64993_db) );
na02s01 TIMEBOOST_cell_16463 ( .a(TIMEBOOST_net_3488), .b(g64928_db), .o(n_3680) );
in01s01 g64994_u0 ( .a(FE_OFN661_n_4392), .o(g64994_sb) );
na02s01 TIMEBOOST_cell_31351 ( .a(TIMEBOOST_net_9586), .b(g65379_da), .o(n_4246) );
na02s01 g64994_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__Q), .b(FE_OFN661_n_4392), .o(g64994_db) );
na02m02 TIMEBOOST_cell_44485 ( .a(n_9648), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__Q), .o(TIMEBOOST_net_14481) );
in01s01 g64995_u0 ( .a(FE_OFN664_n_4495), .o(g64995_sb) );
na02f02 TIMEBOOST_cell_40150 ( .a(TIMEBOOST_net_12313), .b(g57482_sb), .o(n_11254) );
na02s01 g64995_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__Q), .b(FE_OFN664_n_4495), .o(g64995_db) );
na02f02 TIMEBOOST_cell_44486 ( .a(TIMEBOOST_net_14481), .b(FE_OFN2188_n_8567), .o(TIMEBOOST_net_13444) );
in01s01 g64996_u0 ( .a(FE_OFN1624_n_4438), .o(g64996_sb) );
na02f02 TIMEBOOST_cell_40152 ( .a(TIMEBOOST_net_12314), .b(g57309_sb), .o(n_11441) );
na02s01 g64996_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__26__Q), .b(FE_OFN1624_n_4438), .o(g64996_db) );
na02m02 TIMEBOOST_cell_44487 ( .a(n_9556), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q), .o(TIMEBOOST_net_14482) );
in01s01 g64997_u0 ( .a(FE_OFN689_n_4438), .o(g64997_sb) );
na02f02 TIMEBOOST_cell_40154 ( .a(TIMEBOOST_net_12315), .b(g57448_sb), .o(n_11285) );
na02s01 g64997_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__Q), .b(FE_OFN689_n_4438), .o(g64997_db) );
na02f02 TIMEBOOST_cell_44488 ( .a(TIMEBOOST_net_14482), .b(FE_OFN2185_n_8567), .o(TIMEBOOST_net_13445) );
in01s01 g64998_u0 ( .a(FE_OFN1624_n_4438), .o(g64998_sb) );
na02s01 TIMEBOOST_cell_31350 ( .a(n_4498), .b(FE_OFN652_n_4508), .o(TIMEBOOST_net_9586) );
na02s01 g64998_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__Q), .b(FE_OFN1624_n_4438), .o(g64998_db) );
na02s01 TIMEBOOST_cell_31349 ( .a(TIMEBOOST_net_9585), .b(g65421_da), .o(n_4226) );
in01s01 g64999_u0 ( .a(FE_OFN667_n_4495), .o(g64999_sb) );
na02m02 TIMEBOOST_cell_44489 ( .a(n_9025), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__Q), .o(TIMEBOOST_net_14483) );
na02s01 g64999_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__Q), .b(FE_OFN667_n_4495), .o(g64999_db) );
na02f02 TIMEBOOST_cell_40156 ( .a(TIMEBOOST_net_12316), .b(g57524_sb), .o(n_11217) );
ao22f02 g64_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__Q), .b(FE_OFN1529_n_10853), .c(FE_OFN1453_n_10588), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__Q), .o(n_15528) );
in01s01 g65000_u0 ( .a(FE_OFN1628_n_4438), .o(g65000_sb) );
na02f02 TIMEBOOST_cell_44286 ( .a(TIMEBOOST_net_14381), .b(FE_OFN1406_n_8567), .o(TIMEBOOST_net_12787) );
na02s01 g65000_u2 ( .a(n_27), .b(FE_OFN1628_n_4438), .o(g65000_db) );
na02s01 TIMEBOOST_cell_17525 ( .a(TIMEBOOST_net_4019), .b(g65936_sb), .o(n_1564) );
in01s01 g65001_u0 ( .a(FE_OFN662_n_4392), .o(g65001_sb) );
na02f02 TIMEBOOST_cell_44490 ( .a(TIMEBOOST_net_14483), .b(FE_OFN2168_n_8567), .o(TIMEBOOST_net_13446) );
na02s01 g65001_u2 ( .a(n_84), .b(FE_OFN662_n_4392), .o(g65001_db) );
na02f02 TIMEBOOST_cell_40158 ( .a(TIMEBOOST_net_12317), .b(g57350_sb), .o(n_11399) );
in01s01 g65002_u0 ( .a(FE_OFN647_n_4497), .o(g65002_sb) );
na02s01 TIMEBOOST_cell_45111 ( .a(FE_OFN237_n_9118), .b(g57994_sb), .o(TIMEBOOST_net_14794) );
na02s01 g65002_u2 ( .a(n_139), .b(FE_OFN647_n_4497), .o(g65002_db) );
na02s02 TIMEBOOST_cell_45078 ( .a(TIMEBOOST_net_14777), .b(g63165_sb), .o(TIMEBOOST_net_11236) );
in01s01 g65003_u0 ( .a(FE_OFN685_n_4417), .o(g65003_sb) );
na02f02 TIMEBOOST_cell_40160 ( .a(TIMEBOOST_net_12318), .b(g57523_sb), .o(n_11218) );
na02s01 g65003_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__Q), .b(FE_OFN685_n_4417), .o(g65003_db) );
na03m04 TIMEBOOST_cell_45527 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_6__Q), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__Q), .c(FE_OFN2157_n_16439), .o(TIMEBOOST_net_15002) );
in01s01 g65004_u0 ( .a(FE_OFN666_n_4495), .o(g65004_sb) );
na02s01 TIMEBOOST_cell_40545 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_0__Q), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_0__Q), .o(TIMEBOOST_net_12511) );
na02m02 TIMEBOOST_cell_42211 ( .a(n_9747), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__Q), .o(TIMEBOOST_net_13344) );
na02s01 TIMEBOOST_cell_16128 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__Q), .b(pci_target_unit_fifos_pcir_data_in_177), .o(TIMEBOOST_net_3321) );
in01s01 g65005_u0 ( .a(FE_OFN661_n_4392), .o(g65005_sb) );
na02f02 TIMEBOOST_cell_40162 ( .a(TIMEBOOST_net_12319), .b(g57227_sb), .o(n_11530) );
na02s01 g65005_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__Q), .b(FE_OFN661_n_4392), .o(g65005_db) );
na02m02 TIMEBOOST_cell_44491 ( .a(n_9046), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__Q), .o(TIMEBOOST_net_14484) );
in01s01 g65006_u0 ( .a(FE_OFN661_n_4392), .o(g65006_sb) );
na02s01 TIMEBOOST_cell_31348 ( .a(n_4442), .b(FE_OFN653_n_4508), .o(TIMEBOOST_net_9585) );
na02s01 g65006_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__Q), .b(FE_OFN659_n_4392), .o(g65006_db) );
na02f02 TIMEBOOST_cell_40164 ( .a(TIMEBOOST_net_12320), .b(g57342_sb), .o(n_11408) );
in01s01 g65007_u0 ( .a(FE_OFN1625_n_4438), .o(g65007_sb) );
na02m02 TIMEBOOST_cell_41621 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_19__Q), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_13049) );
na02s01 g65007_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__Q), .b(FE_OFN1625_n_4438), .o(g65007_db) );
na02s01 TIMEBOOST_cell_16707 ( .a(TIMEBOOST_net_3610), .b(g58401_sb), .o(n_9004) );
in01s01 g65008_u0 ( .a(FE_OFN1625_n_4438), .o(g65008_sb) );
na02f02 TIMEBOOST_cell_44492 ( .a(TIMEBOOST_net_14484), .b(FE_OFN2169_n_8567), .o(TIMEBOOST_net_13447) );
na02s01 g65008_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__Q), .b(FE_OFN1625_n_4438), .o(g65008_db) );
na02f02 TIMEBOOST_cell_40166 ( .a(TIMEBOOST_net_12321), .b(g57373_sb), .o(n_11375) );
in01s01 g65009_u0 ( .a(FE_OFN648_n_4497), .o(g65009_sb) );
na02s01 TIMEBOOST_cell_9050 ( .a(pci_ad_i_5_), .b(parchk_pci_ad_reg_in_1209), .o(TIMEBOOST_net_1092) );
na02s01 g65009_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__Q), .b(FE_OFN648_n_4497), .o(g65009_db) );
na02s01 TIMEBOOST_cell_9051 ( .a(TIMEBOOST_net_1092), .b(FE_OFN989_n_574), .o(TIMEBOOST_net_767) );
in01s01 g65010_u0 ( .a(FE_OFN622_n_4409), .o(g65010_sb) );
na02s02 TIMEBOOST_cell_32122 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_), .b(n_655), .o(TIMEBOOST_net_9972) );
na02s01 g65010_u2 ( .a(n_3636), .b(FE_OFN622_n_4409), .o(g65010_db) );
na02s02 TIMEBOOST_cell_40756 ( .a(TIMEBOOST_net_12616), .b(g62977_sb), .o(n_5928) );
in01s01 g65011_u0 ( .a(FE_OFN1625_n_4438), .o(g65011_sb) );
na02s02 TIMEBOOST_cell_45173 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__Q), .b(n_1958), .o(TIMEBOOST_net_14825) );
na02s01 g65011_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__Q), .b(FE_OFN1625_n_4438), .o(g65011_db) );
na02f02 TIMEBOOST_cell_40168 ( .a(TIMEBOOST_net_12322), .b(g57365_sb), .o(n_11382) );
in01s01 g65012_u0 ( .a(FE_OFN661_n_4392), .o(g65012_sb) );
na02m02 TIMEBOOST_cell_44493 ( .a(n_9548), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__Q), .o(TIMEBOOST_net_14485) );
na02s01 g65012_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__Q), .b(FE_OFN661_n_4392), .o(g65012_db) );
na02f02 TIMEBOOST_cell_40170 ( .a(TIMEBOOST_net_12323), .b(g57255_sb), .o(n_11499) );
in01s01 g65013_u0 ( .a(FE_OFN625_n_4409), .o(g65013_sb) );
na02s01 TIMEBOOST_cell_16480 ( .a(FE_OFN243_n_9116), .b(g57940_sb), .o(TIMEBOOST_net_3497) );
na02s01 g65013_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__Q), .b(FE_OFN622_n_4409), .o(g65013_db) );
na02s02 TIMEBOOST_cell_36665 ( .a(n_4450), .b(g64864_sb), .o(TIMEBOOST_net_10571) );
in01s01 g65014_u0 ( .a(FE_OFN647_n_4497), .o(g65014_sb) );
na02f02 TIMEBOOST_cell_42156 ( .a(TIMEBOOST_net_13316), .b(FE_OFN1386_n_8567), .o(TIMEBOOST_net_12302) );
na02s01 g65014_u2 ( .a(n_4343), .b(FE_OFN647_n_4497), .o(g65014_db) );
na02s01 TIMEBOOST_cell_42894 ( .a(TIMEBOOST_net_13685), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_11192) );
in01s01 g65015_u0 ( .a(FE_OFN1628_n_4438), .o(g65015_sb) );
na02m02 TIMEBOOST_cell_44269 ( .a(n_9117), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__Q), .o(TIMEBOOST_net_14373) );
na02s02 g65015_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__Q), .b(FE_OFN1628_n_4438), .o(g65015_db) );
na02s01 TIMEBOOST_cell_17527 ( .a(TIMEBOOST_net_4020), .b(g65848_sb), .o(n_1587) );
in01s01 g65016_u0 ( .a(FE_OFN622_n_4409), .o(g65016_sb) );
na02s01 TIMEBOOST_cell_45112 ( .a(TIMEBOOST_net_14794), .b(g57998_db), .o(n_9107) );
na02s01 g65016_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__Q), .b(FE_OFN622_n_4409), .o(g65016_db) );
na02f02 TIMEBOOST_cell_38574 ( .a(g60691_sb), .b(TIMEBOOST_net_11525), .o(n_4199) );
in01s01 g65017_u0 ( .a(FE_OFN646_n_4497), .o(g65017_sb) );
na02s01 TIMEBOOST_cell_9054 ( .a(n_2742), .b(n_3503), .o(TIMEBOOST_net_1094) );
na02s01 g65017_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__Q), .b(FE_OFN646_n_4497), .o(g65017_db) );
na02s01 TIMEBOOST_cell_9055 ( .a(TIMEBOOST_net_1094), .b(n_2125), .o(TIMEBOOST_net_137) );
in01s01 g65018_u0 ( .a(FE_OFN1625_n_4438), .o(g65018_sb) );
na02s01 TIMEBOOST_cell_16481 ( .a(TIMEBOOST_net_3497), .b(g57940_db), .o(n_9130) );
na02s01 g65018_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__Q), .b(FE_OFN1625_n_4438), .o(g65018_db) );
na02f02 TIMEBOOST_cell_44494 ( .a(TIMEBOOST_net_14485), .b(FE_OFN2191_n_8567), .o(TIMEBOOST_net_13019) );
in01s01 g65019_u0 ( .a(FE_OFN687_n_4417), .o(g65019_sb) );
na02f02 TIMEBOOST_cell_40172 ( .a(TIMEBOOST_net_12324), .b(g57084_sb), .o(n_11659) );
na02s01 g65019_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__Q), .b(FE_OFN687_n_4417), .o(g65019_db) );
na02m02 TIMEBOOST_cell_44495 ( .a(n_9898), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__8__Q), .o(TIMEBOOST_net_14486) );
in01s01 g65020_u0 ( .a(FE_OFN670_n_4505), .o(g65020_sb) );
na02s01 TIMEBOOST_cell_9311 ( .a(TIMEBOOST_net_1222), .b(g65805_db), .o(n_1668) );
na02s01 g65020_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__Q), .b(FE_OFN670_n_4505), .o(g65020_db) );
na02s01 TIMEBOOST_cell_40554 ( .a(TIMEBOOST_net_12515), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_11559) );
in01s01 g65021_u0 ( .a(FE_OFN630_n_4454), .o(g65021_sb) );
na02s02 TIMEBOOST_cell_40758 ( .a(TIMEBOOST_net_12617), .b(g62550_sb), .o(n_6465) );
na02s01 g65021_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__Q), .b(FE_OFN630_n_4454), .o(g65021_db) );
na02s02 TIMEBOOST_cell_32120 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_), .o(TIMEBOOST_net_9971) );
in01s01 g65022_u0 ( .a(FE_OFN687_n_4417), .o(g65022_sb) );
na02f02 TIMEBOOST_cell_40174 ( .a(TIMEBOOST_net_12325), .b(g57278_sb), .o(n_11476) );
na02s01 g65022_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__Q), .b(FE_OFN687_n_4417), .o(g65022_db) );
na02s02 TIMEBOOST_cell_36664 ( .a(TIMEBOOST_net_10570), .b(g52638_sb), .o(n_14750) );
in01s01 g65023_u0 ( .a(FE_OFN667_n_4495), .o(g65023_sb) );
na02m04 TIMEBOOST_cell_39021 ( .a(wbs_wbb3_2_wbb2_dat_o_i_127), .b(wbs_dat_o_28_), .o(TIMEBOOST_net_11749) );
na02s01 g65023_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__Q), .b(FE_OFN667_n_4495), .o(g65023_db) );
na02s02 TIMEBOOST_cell_39198 ( .a(TIMEBOOST_net_11837), .b(wbu_addr_in_267), .o(n_9851) );
in01s01 g65024_u0 ( .a(FE_OFN630_n_4454), .o(g65024_sb) );
na02s01 TIMEBOOST_cell_38576 ( .a(TIMEBOOST_net_11526), .b(n_7136), .o(n_7393) );
na02s01 g65024_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__Q), .b(FE_OFN630_n_4454), .o(g65024_db) );
na02s02 TIMEBOOST_cell_32118 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_), .b(n_669), .o(TIMEBOOST_net_9970) );
in01s01 g65025_u0 ( .a(FE_OFN624_n_4409), .o(g65025_sb) );
na02s01 TIMEBOOST_cell_16708 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(g64146_sb), .o(TIMEBOOST_net_3611) );
na02s01 g65025_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q), .b(FE_OFN624_n_4409), .o(g65025_db) );
na02s01 TIMEBOOST_cell_16709 ( .a(TIMEBOOST_net_3611), .b(g64146_db), .o(n_4019) );
in01s01 g65026_u0 ( .a(FE_OFN634_n_4454), .o(g65026_sb) );
na02s02 TIMEBOOST_cell_45113 ( .a(n_3984), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__Q), .o(TIMEBOOST_net_14795) );
na02s01 TIMEBOOST_cell_42751 ( .a(FE_OFN247_n_9112), .b(g58256_sb), .o(TIMEBOOST_net_13614) );
na02s02 TIMEBOOST_cell_38578 ( .a(TIMEBOOST_net_11527), .b(g59384_sb), .o(n_7539) );
in01s01 g65027_u0 ( .a(FE_OFN630_n_4454), .o(g65027_sb) );
na02s01 TIMEBOOST_cell_9351 ( .a(TIMEBOOST_net_1242), .b(g65757_db), .o(n_3212) );
na02s02 TIMEBOOST_cell_32116 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_), .b(n_741), .o(TIMEBOOST_net_9969) );
na02s01 TIMEBOOST_cell_17201 ( .a(TIMEBOOST_net_3857), .b(g65348_db), .o(n_3543) );
in01s01 g65028_u0 ( .a(FE_OFN665_n_4495), .o(g65028_sb) );
na02f02 TIMEBOOST_cell_40176 ( .a(TIMEBOOST_net_12326), .b(g57286_sb), .o(n_11467) );
na02s01 g65028_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__Q), .b(FE_OFN665_n_4495), .o(g65028_db) );
na02f02 TIMEBOOST_cell_44538 ( .a(TIMEBOOST_net_14507), .b(FE_OFN1428_n_8567), .o(TIMEBOOST_net_13460) );
in01s01 g65029_u0 ( .a(FE_OFN685_n_4417), .o(g65029_sb) );
na02f02 TIMEBOOST_cell_40178 ( .a(TIMEBOOST_net_12327), .b(FE_OFN2179_n_8567), .o(n_11546) );
na02s01 g65029_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__Q), .b(FE_OFN685_n_4417), .o(g65029_db) );
na02m02 TIMEBOOST_cell_44539 ( .a(n_9750), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q), .o(TIMEBOOST_net_14508) );
in01s01 g65030_u0 ( .a(FE_OFN634_n_4454), .o(g65030_sb) );
na02s02 TIMEBOOST_cell_40760 ( .a(TIMEBOOST_net_12618), .b(g62346_sb), .o(n_6908) );
na02s01 g65030_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__Q), .b(FE_OFN634_n_4454), .o(g65030_db) );
in01s01 g65031_u0 ( .a(FE_OFN685_n_4417), .o(g65031_sb) );
na02m02 TIMEBOOST_cell_36667 ( .a(pci_target_unit_pcit_if_strd_addr_in_715), .b(g52645_sb), .o(TIMEBOOST_net_10572) );
na02s01 g65031_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__26__Q), .b(FE_OFN685_n_4417), .o(g65031_db) );
na02f02 TIMEBOOST_cell_40180 ( .a(TIMEBOOST_net_12328), .b(FE_OFN2180_n_8567), .o(n_11566) );
in01s01 g65032_u0 ( .a(FE_OFN660_n_4392), .o(g65032_sb) );
na02f02 TIMEBOOST_cell_44620 ( .a(TIMEBOOST_net_14548), .b(FE_OFN2189_n_8567), .o(TIMEBOOST_net_13492) );
na02s01 g65032_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__Q), .b(FE_OFN660_n_4392), .o(g65032_db) );
na02m02 TIMEBOOST_cell_44621 ( .a(n_9855), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__Q), .o(TIMEBOOST_net_14549) );
in01s01 g65033_u0 ( .a(FE_OFN629_n_4454), .o(g65033_sb) );
na02f02 TIMEBOOST_cell_44540 ( .a(TIMEBOOST_net_14508), .b(FE_OFN1428_n_8567), .o(TIMEBOOST_net_13461) );
na02f02 TIMEBOOST_cell_40182 ( .a(TIMEBOOST_net_12329), .b(FE_OFN2179_n_8567), .o(n_11205) );
in01s01 g65034_u0 ( .a(FE_OFN633_n_4454), .o(g65034_sb) );
na02m02 TIMEBOOST_cell_44541 ( .a(n_9431), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__Q), .o(TIMEBOOST_net_14509) );
na02s01 g65034_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__Q), .b(FE_OFN633_n_4454), .o(g65034_db) );
na02f02 TIMEBOOST_cell_40184 ( .a(TIMEBOOST_net_12330), .b(FE_OFN2179_n_8567), .o(n_11287) );
in01s01 g65035_u0 ( .a(FE_OFN1810_n_4454), .o(g65035_sb) );
na02f02 TIMEBOOST_cell_44496 ( .a(TIMEBOOST_net_14486), .b(FE_OFN2173_n_8567), .o(TIMEBOOST_net_13448) );
na02s01 g65035_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__Q), .b(FE_OFN1810_n_4454), .o(g65035_db) );
na02f02 TIMEBOOST_cell_40186 ( .a(TIMEBOOST_net_12331), .b(FE_OFN2177_n_8567), .o(n_11682) );
in01s01 g65036_u0 ( .a(FE_OFN618_n_4490), .o(g65036_sb) );
na02s01 TIMEBOOST_cell_31153 ( .a(TIMEBOOST_net_9487), .b(g64921_db), .o(n_3683) );
na02s01 g65036_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__Q), .b(FE_OFN618_n_4490), .o(g65036_db) );
na02s02 TIMEBOOST_cell_41820 ( .a(TIMEBOOST_net_13148), .b(g58406_db), .o(n_9001) );
in01s01 g65037_u0 ( .a(FE_OFN684_n_4417), .o(g65037_sb) );
na02f02 TIMEBOOST_cell_44542 ( .a(TIMEBOOST_net_14509), .b(FE_OFN2168_n_8567), .o(TIMEBOOST_net_13462) );
na02s01 g65037_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__Q), .b(FE_OFN684_n_4417), .o(g65037_db) );
na02f02 TIMEBOOST_cell_40188 ( .a(TIMEBOOST_net_12332), .b(g57323_sb), .o(n_11427) );
in01s01 g65038_u0 ( .a(FE_OFN633_n_4454), .o(g65038_sb) );
na02s01 TIMEBOOST_cell_36666 ( .a(TIMEBOOST_net_10571), .b(g64864_db), .o(n_4427) );
na02s01 TIMEBOOST_cell_42752 ( .a(TIMEBOOST_net_13614), .b(g58256_db), .o(n_9040) );
na02f02 TIMEBOOST_cell_44558 ( .a(TIMEBOOST_net_14517), .b(FE_OFN2175_n_8567), .o(TIMEBOOST_net_13468) );
in01s01 g65039_u0 ( .a(FE_OFN623_n_4409), .o(g65039_sb) );
na02f02 TIMEBOOST_cell_40190 ( .a(TIMEBOOST_net_12333), .b(g57510_sb), .o(n_10323) );
na02s01 g65039_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__Q), .b(FE_OFN623_n_4409), .o(g65039_db) );
na02s02 TIMEBOOST_cell_45688 ( .a(TIMEBOOST_net_15082), .b(FE_OFN1248_n_4093), .o(TIMEBOOST_net_13304) );
in01s01 g65040_u0 ( .a(FE_OFN1809_n_4454), .o(g65040_sb) );
na02s01 TIMEBOOST_cell_9750 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__Q), .b(g65877_sb), .o(TIMEBOOST_net_1442) );
na02s01 g65040_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__Q), .b(FE_OFN1809_n_4454), .o(g65040_db) );
na02s01 TIMEBOOST_cell_9751 ( .a(TIMEBOOST_net_1442), .b(g65877_db), .o(n_1867) );
in01s01 g65041_u0 ( .a(FE_OFN625_n_4409), .o(g65041_sb) );
na02f02 TIMEBOOST_cell_44622 ( .a(TIMEBOOST_net_14549), .b(FE_OFN2182_n_8567), .o(TIMEBOOST_net_13479) );
na02s01 g65041_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__Q), .b(FE_OFN625_n_4409), .o(g65041_db) );
na02m02 TIMEBOOST_cell_44623 ( .a(n_9054), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__Q), .o(TIMEBOOST_net_14550) );
in01s01 g65042_u0 ( .a(FE_OFN649_n_4497), .o(g65042_sb) );
na02s01 TIMEBOOST_cell_9056 ( .a(n_245), .b(n_193), .o(TIMEBOOST_net_1095) );
na02s01 g65042_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__Q), .b(FE_OFN649_n_4497), .o(g65042_db) );
na02s02 TIMEBOOST_cell_9057 ( .a(TIMEBOOST_net_1095), .b(n_785), .o(TIMEBOOST_net_166) );
in01s01 g65043_u0 ( .a(FE_OFN647_n_4497), .o(g65043_sb) );
na02s01 TIMEBOOST_cell_39199 ( .a(TIMEBOOST_net_3320), .b(FE_OFN1003_n_2047), .o(TIMEBOOST_net_11838) );
na02s01 g65043_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__Q), .b(FE_OFN647_n_4497), .o(g65043_db) );
na02f02 TIMEBOOST_cell_39054 ( .a(TIMEBOOST_net_11765), .b(g54337_sb), .o(n_13482) );
in01s01 g65044_u0 ( .a(FE_OFN625_n_4409), .o(g65044_sb) );
na02s02 TIMEBOOST_cell_40762 ( .a(TIMEBOOST_net_12619), .b(g62367_sb), .o(n_6868) );
na02s01 g65044_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__Q), .b(FE_OFN625_n_4409), .o(g65044_db) );
in01s01 g65045_u0 ( .a(FE_OFN1810_n_4454), .o(g65045_sb) );
na02s01 TIMEBOOST_cell_9752 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__Q), .b(g65976_sb), .o(TIMEBOOST_net_1443) );
na02s01 g65045_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__Q), .b(FE_OFN1810_n_4454), .o(g65045_db) );
na02s01 TIMEBOOST_cell_9753 ( .a(TIMEBOOST_net_1443), .b(g65976_db), .o(n_1838) );
in01s01 g65046_u0 ( .a(FE_OFN624_n_4409), .o(g65046_sb) );
na02f02 TIMEBOOST_cell_40192 ( .a(TIMEBOOST_net_12334), .b(g57067_sb), .o(n_11675) );
na02s01 g65046_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__Q), .b(FE_OFN624_n_4409), .o(g65046_db) );
na02s01 TIMEBOOST_cell_31343 ( .a(TIMEBOOST_net_9582), .b(g65326_da), .o(n_4267) );
in01s01 g65047_u0 ( .a(FE_OFN631_n_4454), .o(g65047_sb) );
na02s02 TIMEBOOST_cell_40698 ( .a(TIMEBOOST_net_12587), .b(g62494_sb), .o(n_6596) );
na02s01 g65047_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__Q), .b(FE_OFN631_n_4454), .o(g65047_db) );
na03s02 TIMEBOOST_cell_40699 ( .a(n_4403), .b(n_4404), .c(FE_OFN1218_n_6886), .o(TIMEBOOST_net_12588) );
in01s01 g65048_u0 ( .a(FE_OFN646_n_4497), .o(g65048_sb) );
na02s02 TIMEBOOST_cell_45751 ( .a(n_4331), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__Q), .o(TIMEBOOST_net_15114) );
na02s01 g65048_u2 ( .a(n_4323), .b(FE_OFN646_n_4497), .o(g65048_db) );
na02f04 TIMEBOOST_cell_9059 ( .a(TIMEBOOST_net_1096), .b(n_3123), .o(FE_RN_273_0) );
in01s01 g65049_u0 ( .a(FE_OFN687_n_4417), .o(g65049_sb) );
na02m02 TIMEBOOST_cell_44497 ( .a(n_9726), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__8__Q), .o(TIMEBOOST_net_14487) );
na02s01 g65049_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__Q), .b(FE_OFN687_n_4417), .o(g65049_db) );
na02f02 TIMEBOOST_cell_40194 ( .a(TIMEBOOST_net_12335), .b(g57163_sb), .o(n_11587) );
in01s01 g65050_u0 ( .a(FE_OFN687_n_4417), .o(g65050_sb) );
na02s01 TIMEBOOST_cell_16502 ( .a(pci_target_unit_fifos_pcir_data_in_185), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__Q), .o(TIMEBOOST_net_3508) );
na02s01 g65050_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__Q), .b(FE_OFN686_n_4417), .o(g65050_db) );
na02f02 TIMEBOOST_cell_44630 ( .a(TIMEBOOST_net_14553), .b(FE_OFN2177_n_8567), .o(TIMEBOOST_net_13025) );
in01s01 g65051_u0 ( .a(FE_OFN648_n_4497), .o(g65051_sb) );
na02s01 g65051_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__Q), .b(FE_OFN646_n_4497), .o(g65051_db) );
na02s02 TIMEBOOST_cell_40764 ( .a(TIMEBOOST_net_12620), .b(g62627_sb), .o(n_6301) );
in01s01 g65052_u0 ( .a(FE_OFN666_n_4495), .o(g65052_sb) );
na02s01 g65052_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__Q), .b(FE_OFN666_n_4495), .o(g65052_db) );
na02m02 TIMEBOOST_cell_40196 ( .a(TIMEBOOST_net_12336), .b(g58842_sb), .o(n_8672) );
in01s01 g65053_u0 ( .a(FE_OFN620_n_4490), .o(g65053_sb) );
na02m04 TIMEBOOST_cell_45528 ( .a(TIMEBOOST_net_15002), .b(g58833_sb), .o(n_8604) );
na02s01 g65053_u2 ( .a(n_17), .b(FE_OFN620_n_4490), .o(g65053_db) );
na02f02 TIMEBOOST_cell_40198 ( .a(TIMEBOOST_net_12337), .b(FE_OFN1471_g52675_p), .o(TIMEBOOST_net_11747) );
in01s01 g65054_u0 ( .a(FE_OFN618_n_4490), .o(g65054_sb) );
na02s01 TIMEBOOST_cell_31152 ( .a(n_3777), .b(g64921_sb), .o(TIMEBOOST_net_9487) );
na02s01 g65054_u2 ( .a(n_3616), .b(FE_OFN618_n_4490), .o(g65054_db) );
na02s02 TIMEBOOST_cell_31151 ( .a(TIMEBOOST_net_9486), .b(g64893_sb), .o(n_3700) );
in01s01 g65055_u0 ( .a(FE_OFN620_n_4490), .o(g65055_sb) );
na02f02 TIMEBOOST_cell_39056 ( .a(TIMEBOOST_net_11766), .b(FE_OFN1774_n_13800), .o(g53171_p) );
na02s02 TIMEBOOST_cell_40694 ( .a(TIMEBOOST_net_12585), .b(g62428_sb), .o(n_6743) );
na02f02 TIMEBOOST_cell_39058 ( .a(TIMEBOOST_net_11767), .b(FE_OFN1774_n_13800), .o(g53214_p) );
in01s01 g65056_u0 ( .a(FE_OFN624_n_4409), .o(g65056_sb) );
na02m02 TIMEBOOST_cell_40199 ( .a(wbs_wbb3_2_wbb2_dat_o_i_106), .b(wbs_dat_o_7_), .o(TIMEBOOST_net_12338) );
na02s01 g65056_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__Q), .b(FE_OFN624_n_4409), .o(g65056_db) );
na02s01 TIMEBOOST_cell_42646 ( .a(TIMEBOOST_net_13561), .b(g57941_db), .o(n_9129) );
in01s01 g65057_u0 ( .a(n_4460), .o(g65057_sb) );
na02s01 TIMEBOOST_cell_18645 ( .a(TIMEBOOST_net_4579), .b(g63132_sb), .o(n_4986) );
na02s01 g65057_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__Q), .b(n_4460), .o(g65057_db) );
na03s02 TIMEBOOST_cell_38213 ( .a(TIMEBOOST_net_4008), .b(g64137_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__Q), .o(TIMEBOOST_net_11345) );
in01s01 g65058_u0 ( .a(FE_OFN619_n_4490), .o(g65058_sb) );
na02s02 TIMEBOOST_cell_41821 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__Q), .b(g58346_sb), .o(TIMEBOOST_net_13149) );
na02s01 g65058_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__Q), .b(FE_OFN619_n_4490), .o(g65058_db) );
na02s02 TIMEBOOST_cell_43452 ( .a(TIMEBOOST_net_13964), .b(FE_OFN1233_n_6391), .o(TIMEBOOST_net_12162) );
in01s01 g65059_u0 ( .a(FE_OFN1663_n_4490), .o(g65059_sb) );
na02s01 TIMEBOOST_cell_31149 ( .a(TIMEBOOST_net_9485), .b(g64886_db), .o(n_3704) );
na02s01 g65059_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__Q), .b(FE_OFN1663_n_4490), .o(g65059_db) );
na02s01 TIMEBOOST_cell_31105 ( .a(TIMEBOOST_net_9463), .b(g64821_db), .o(n_3737) );
in01s01 g65060_u0 ( .a(FE_OFN667_n_4495), .o(g65060_sb) );
na02s01 TIMEBOOST_cell_16129 ( .a(TIMEBOOST_net_3321), .b(FE_OFN1003_n_2047), .o(TIMEBOOST_net_1267) );
na02s01 g65060_u2 ( .a(n_83), .b(FE_OFN667_n_4495), .o(g65060_db) );
na02s01 TIMEBOOST_cell_16130 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__Q), .b(pci_target_unit_fifos_pcir_data_in_175), .o(TIMEBOOST_net_3322) );
in01s01 g65061_u0 ( .a(FE_OFN1663_n_4490), .o(g65061_sb) );
na02s01 TIMEBOOST_cell_16578 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__Q), .b(g64344_sb), .o(TIMEBOOST_net_3546) );
na02s01 g65061_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__Q), .b(FE_OFN1663_n_4490), .o(g65061_db) );
na02s01 TIMEBOOST_cell_44987 ( .a(g61962_sb), .b(g61988_db), .o(TIMEBOOST_net_14732) );
in01s01 g65062_u0 ( .a(FE_OFN1663_n_4490), .o(g65062_sb) );
na02s02 TIMEBOOST_cell_16580 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q), .b(g64353_sb), .o(TIMEBOOST_net_3547) );
na02s01 g65062_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__Q), .b(FE_OFN1663_n_4490), .o(g65062_db) );
na02s01 TIMEBOOST_cell_45079 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__Q), .b(FE_OFN576_n_9902), .o(TIMEBOOST_net_14778) );
in01s01 g65063_u0 ( .a(FE_OFN681_n_4460), .o(g65063_sb) );
na02s01 TIMEBOOST_cell_31342 ( .a(n_4465), .b(FE_OFN1644_n_4671), .o(TIMEBOOST_net_9582) );
na02s01 g65063_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__Q), .b(FE_OFN681_n_4460), .o(g65063_db) );
na02s02 TIMEBOOST_cell_45198 ( .a(TIMEBOOST_net_14837), .b(FE_OFN1260_n_4143), .o(TIMEBOOST_net_12097) );
in01s01 g65064_u0 ( .a(FE_OFN1810_n_4454), .o(g65064_sb) );
na02s01 TIMEBOOST_cell_9754 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__Q), .b(g65977_sb), .o(TIMEBOOST_net_1444) );
na02s01 g65064_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__Q), .b(FE_OFN1810_n_4454), .o(g65064_db) );
na02s01 TIMEBOOST_cell_9755 ( .a(TIMEBOOST_net_1444), .b(g65977_db), .o(n_1837) );
in01s01 g65065_u0 ( .a(FE_OFN662_n_4392), .o(g65065_sb) );
na02f02 TIMEBOOST_cell_40200 ( .a(TIMEBOOST_net_12338), .b(FE_OFN1471_g52675_p), .o(TIMEBOOST_net_11742) );
na02s01 g65065_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__Q), .b(FE_OFN662_n_4392), .o(g65065_db) );
na02s02 TIMEBOOST_cell_31341 ( .a(TIMEBOOST_net_9581), .b(g65416_da), .o(n_4229) );
in01s01 g65066_u0 ( .a(FE_OFN620_n_4490), .o(g65066_sb) );
na02s01 TIMEBOOST_cell_16582 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__Q), .b(g64357_sb), .o(TIMEBOOST_net_3548) );
na02s01 g65066_u2 ( .a(n_3608), .b(FE_OFN620_n_4490), .o(g65066_db) );
na02s02 TIMEBOOST_cell_45114 ( .a(TIMEBOOST_net_14795), .b(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_11447) );
in01s01 g65067_u0 ( .a(FE_OFN1663_n_4490), .o(g65067_sb) );
na02m02 TIMEBOOST_cell_40201 ( .a(wbs_wbb3_2_wbb2_dat_o_i_105), .b(wbs_dat_o_6_), .o(TIMEBOOST_net_12339) );
na02s01 g65067_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__Q), .b(FE_OFN1663_n_4490), .o(g65067_db) );
na02f02 TIMEBOOST_cell_40202 ( .a(TIMEBOOST_net_12339), .b(FE_OFN1471_g52675_p), .o(TIMEBOOST_net_11741) );
in01s01 g65068_u0 ( .a(FE_OFN618_n_4490), .o(g65068_sb) );
na02s01 TIMEBOOST_cell_17411 ( .a(TIMEBOOST_net_3962), .b(g64263_db), .o(n_3910) );
na02s02 TIMEBOOST_cell_38580 ( .a(TIMEBOOST_net_11528), .b(g60622_sb), .o(n_4832) );
na02f04 TIMEBOOST_cell_37112 ( .a(TIMEBOOST_net_10794), .b(n_12589), .o(n_12851) );
in01s01 g65069_u0 ( .a(n_4460), .o(g65069_sb) );
na02s01 TIMEBOOST_cell_22292 ( .a(g52474_da), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_6403) );
na02s01 g65069_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__Q), .b(n_4460), .o(g65069_db) );
na02m02 TIMEBOOST_cell_10163 ( .a(FE_OFN1151_n_13249), .b(TIMEBOOST_net_1648), .o(TIMEBOOST_net_492) );
in01s01 g65070_u0 ( .a(FE_OFN665_n_4495), .o(g65070_sb) );
na02f02 TIMEBOOST_cell_42212 ( .a(TIMEBOOST_net_13344), .b(FE_OFN1408_n_8567), .o(TIMEBOOST_net_12297) );
na02s01 TIMEBOOST_cell_16132 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__Q), .b(pci_target_unit_fifos_pcir_data_in_165), .o(TIMEBOOST_net_3323) );
in01s01 g65071_u0 ( .a(FE_OFN631_n_4454), .o(g65071_sb) );
na02m02 TIMEBOOST_cell_40203 ( .a(wbs_wbb3_2_wbb2_dat_o_i), .b(wbs_dat_o_0_), .o(TIMEBOOST_net_12340) );
na02s01 g65071_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__Q), .b(FE_OFN631_n_4454), .o(g65071_db) );
na02s02 TIMEBOOST_cell_31340 ( .a(n_4479), .b(FE_OFN1640_n_4671), .o(TIMEBOOST_net_9581) );
in01s01 g65072_u0 ( .a(FE_OFN681_n_4460), .o(g65072_sb) );
na02s01 TIMEBOOST_cell_31339 ( .a(TIMEBOOST_net_9580), .b(g65430_da), .o(n_4222) );
na02s01 g65072_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q), .b(FE_OFN681_n_4460), .o(g65072_db) );
na02f02 TIMEBOOST_cell_40204 ( .a(TIMEBOOST_net_12340), .b(FE_OFN1471_g52675_p), .o(TIMEBOOST_net_11746) );
in01s01 g65073_u0 ( .a(FE_OFN660_n_4392), .o(g65073_sb) );
na02s01 TIMEBOOST_cell_31338 ( .a(n_4645), .b(FE_OFN653_n_4508), .o(TIMEBOOST_net_9580) );
na02s01 g65073_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__Q), .b(FE_OFN660_n_4392), .o(g65073_db) );
na02s02 TIMEBOOST_cell_31337 ( .a(TIMEBOOST_net_9579), .b(g65429_da), .o(n_4223) );
in01s01 g65074_u0 ( .a(FE_OFN681_n_4460), .o(g65074_sb) );
na02f02 TIMEBOOST_cell_40206 ( .a(TIMEBOOST_net_12341), .b(FE_OFN1471_g52675_p), .o(TIMEBOOST_net_11744) );
na02m02 TIMEBOOST_cell_44543 ( .a(n_9891), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__Q), .o(TIMEBOOST_net_14510) );
na02m02 TIMEBOOST_cell_40207 ( .a(wbs_wbb3_2_wbb2_dat_o_i_123), .b(wbs_dat_o_24_), .o(TIMEBOOST_net_12342) );
in01s01 g65075_u0 ( .a(FE_OFN666_n_4495), .o(g65075_sb) );
na02f02 TIMEBOOST_cell_40208 ( .a(TIMEBOOST_net_12342), .b(FE_OFN1471_g52675_p), .o(TIMEBOOST_net_11743) );
na02s01 g65075_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__Q), .b(FE_OFN666_n_4495), .o(g65075_db) );
na02s01 TIMEBOOST_cell_42872 ( .a(TIMEBOOST_net_13674), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_11209) );
in01s01 g65076_u0 ( .a(FE_OFN662_n_4392), .o(g65076_sb) );
na02s02 TIMEBOOST_cell_31336 ( .a(n_4447), .b(FE_OFN654_n_4508), .o(TIMEBOOST_net_9579) );
na02m02 TIMEBOOST_cell_39557 ( .a(TIMEBOOST_net_4079), .b(n_8750), .o(TIMEBOOST_net_12017) );
na02s01 TIMEBOOST_cell_36476 ( .a(TIMEBOOST_net_10476), .b(g65691_sb), .o(n_1916) );
in01s01 g65077_u0 ( .a(n_4460), .o(g65077_sb) );
na02f02 TIMEBOOST_cell_10165 ( .a(TIMEBOOST_net_1649), .b(FE_OFN1147_n_13249), .o(TIMEBOOST_net_556) );
na02s01 g65077_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__Q), .b(n_4460), .o(g65077_db) );
na02m02 TIMEBOOST_cell_10167 ( .a(TIMEBOOST_net_1650), .b(FE_OFN1149_n_13249), .o(TIMEBOOST_net_495) );
in01s01 g65078_u0 ( .a(FE_OFN681_n_4460), .o(g65078_sb) );
na02s01 TIMEBOOST_cell_16510 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__Q), .b(g64227_sb), .o(TIMEBOOST_net_3512) );
na02s01 g65078_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q), .b(FE_OFN681_n_4460), .o(g65078_db) );
na02s01 TIMEBOOST_cell_44988 ( .a(TIMEBOOST_net_14732), .b(g63613_db), .o(TIMEBOOST_net_13151) );
in01s01 g65079_u0 ( .a(FE_OFN631_n_4454), .o(g65079_sb) );
na02s01 TIMEBOOST_cell_42873 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__Q), .b(FE_OFN540_n_9690), .o(TIMEBOOST_net_13675) );
na02s01 g65079_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__Q), .b(FE_OFN631_n_4454), .o(g65079_db) );
na02s01 TIMEBOOST_cell_42874 ( .a(TIMEBOOST_net_13675), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_11214) );
in01s01 g65080_u0 ( .a(FE_OFN682_n_4460), .o(g65080_sb) );
na02s01 TIMEBOOST_cell_31334 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__Q), .o(TIMEBOOST_net_9578) );
na02s02 g65080_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__Q), .b(FE_OFN682_n_4460), .o(g65080_db) );
na02s01 TIMEBOOST_cell_16512 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__Q), .b(g64254_sb), .o(TIMEBOOST_net_3513) );
in01s01 g65081_u0 ( .a(FE_OFN624_n_4409), .o(g65081_sb) );
na02s02 TIMEBOOST_cell_32114 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_), .b(n_599), .o(TIMEBOOST_net_9968) );
na02s01 g65081_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__Q), .b(FE_OFN624_n_4409), .o(g65081_db) );
na02m02 TIMEBOOST_cell_32113 ( .a(TIMEBOOST_net_9967), .b(TIMEBOOST_net_2307), .o(n_3456) );
in01s01 g65082_u0 ( .a(FE_OFN678_n_4460), .o(g65082_sb) );
na02s02 TIMEBOOST_cell_45174 ( .a(TIMEBOOST_net_14825), .b(FE_OFN1265_n_4095), .o(TIMEBOOST_net_12055) );
na02s01 g65082_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__Q), .b(FE_OFN678_n_4460), .o(g65082_db) );
na02m02 TIMEBOOST_cell_40205 ( .a(wbs_wbb3_2_wbb2_dat_o_i_111), .b(wbs_dat_o_12_), .o(TIMEBOOST_net_12341) );
in01s01 g65083_u0 ( .a(FE_OFN624_n_4409), .o(g65083_sb) );
na02m02 TIMEBOOST_cell_32112 ( .a(wbm_adr_o_11_), .b(g63204_sb), .o(TIMEBOOST_net_9967) );
na02s01 g65083_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__Q), .b(FE_OFN624_n_4409), .o(g65083_db) );
in01s01 g65084_u0 ( .a(FE_OFN682_n_4460), .o(g65084_sb) );
na02f02 TIMEBOOST_cell_40210 ( .a(TIMEBOOST_net_12343), .b(FE_OFN1471_g52675_p), .o(TIMEBOOST_net_11740) );
na02s01 g65084_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__Q), .b(FE_OFN682_n_4460), .o(g65084_db) );
na02s01 TIMEBOOST_cell_16516 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(g65676_sb), .o(TIMEBOOST_net_3515) );
in01s01 g65085_u0 ( .a(FE_OFN662_n_4392), .o(g65085_sb) );
na02s01 g65085_u1 ( .a(n_4473), .b(g65085_sb), .o(g65085_da) );
na02s01 g65085_u2 ( .a(n_26), .b(FE_OFN662_n_4392), .o(g65085_db) );
na02s01 g65085_u3 ( .a(g65085_da), .b(g65085_db), .o(n_4303) );
in01s01 g65086_u0 ( .a(FE_OFN682_n_4460), .o(g65086_sb) );
na02s01 TIMEBOOST_cell_36479 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__Q), .b(FE_OFN527_n_9899), .o(TIMEBOOST_net_10478) );
na02f02 TIMEBOOST_cell_44116 ( .a(TIMEBOOST_net_14296), .b(FE_OFN1424_n_8567), .o(TIMEBOOST_net_13383) );
na02s01 TIMEBOOST_cell_36478 ( .a(TIMEBOOST_net_10477), .b(g65769_db), .o(n_1914) );
in01s01 g65087_u0 ( .a(FE_OFN662_n_4392), .o(g65087_sb) );
na02s01 TIMEBOOST_cell_16517 ( .a(TIMEBOOST_net_3515), .b(g65676_db), .o(n_1957) );
na02m02 TIMEBOOST_cell_44117 ( .a(n_9487), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__Q), .o(TIMEBOOST_net_14297) );
na02m02 TIMEBOOST_cell_40211 ( .a(wbs_wbb3_2_wbb2_dat_o_i_108), .b(wbs_dat_o_9_), .o(TIMEBOOST_net_12344) );
in01s01 g65088_u0 ( .a(FE_OFN659_n_4392), .o(g65088_sb) );
na02f02 TIMEBOOST_cell_40212 ( .a(TIMEBOOST_net_12344), .b(FE_OFN1471_g52675_p), .o(TIMEBOOST_net_11745) );
na02s01 g65088_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__Q), .b(FE_OFN659_n_4392), .o(g65088_db) );
na02s01 TIMEBOOST_cell_16520 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(g65708_sb), .o(TIMEBOOST_net_3517) );
in01s01 g65089_u0 ( .a(FE_OFN669_n_4505), .o(g65089_sb) );
na02s01 TIMEBOOST_cell_16521 ( .a(TIMEBOOST_net_3517), .b(g65708_db), .o(n_1947) );
na02s01 g65089_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__Q), .b(FE_OFN669_n_4505), .o(g65089_db) );
na02s01 TIMEBOOST_cell_31331 ( .a(TIMEBOOST_net_9576), .b(g65395_db), .o(n_4156) );
in01s01 g65090_u0 ( .a(FE_OFN666_n_4495), .o(g65090_sb) );
na02s01 TIMEBOOST_cell_16522 ( .a(pci_target_unit_fifos_pcir_data_in_164), .b(g65722_sb), .o(TIMEBOOST_net_3518) );
na02s01 g65090_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__28__Q), .b(FE_OFN666_n_4495), .o(g65090_db) );
na02s01 TIMEBOOST_cell_16523 ( .a(TIMEBOOST_net_3518), .b(g65722_db), .o(n_1940) );
in01s01 g65091_u0 ( .a(FE_OFN667_n_4495), .o(g65091_sb) );
na02s01 TIMEBOOST_cell_16133 ( .a(TIMEBOOST_net_3323), .b(FE_OFN1003_n_2047), .o(TIMEBOOST_net_1294) );
na02s01 g65091_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__Q), .b(FE_OFN667_n_4495), .o(g65091_db) );
na02s01 TIMEBOOST_cell_40497 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__Q), .b(wishbone_slave_unit_pcim_sm_data_in_660), .o(TIMEBOOST_net_12487) );
in01s01 g65092_u0 ( .a(FE_OFN618_n_4490), .o(g65092_sb) );
na02m02 TIMEBOOST_cell_38820 ( .a(TIMEBOOST_net_11648), .b(g58476_sb), .o(n_9363) );
na02s02 TIMEBOOST_cell_37969 ( .a(TIMEBOOST_net_1682), .b(g61887_sb), .o(TIMEBOOST_net_11223) );
na02s01 TIMEBOOST_cell_9141 ( .a(TIMEBOOST_net_1137), .b(n_4730), .o(TIMEBOOST_net_170) );
in01s01 g65093_u0 ( .a(FE_OFN686_n_4417), .o(g65093_sb) );
na02f02 TIMEBOOST_cell_39055 ( .a(TIMEBOOST_net_10144), .b(FE_OFN1770_n_14054), .o(TIMEBOOST_net_11766) );
na02s01 g65093_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__Q), .b(FE_OFN686_n_4417), .o(g65093_db) );
na02f02 TIMEBOOST_cell_39060 ( .a(TIMEBOOST_net_11768), .b(FE_OFN1774_n_13800), .o(g53203_p) );
in01s01 g65094_u0 ( .a(FE_OFN625_n_4409), .o(g65094_sb) );
na02s01 TIMEBOOST_cell_42875 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__Q), .b(FE_OFN517_n_9697), .o(TIMEBOOST_net_13676) );
na02s01 g65094_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__Q), .b(FE_OFN625_n_4409), .o(g65094_db) );
na02s01 TIMEBOOST_cell_44989 ( .a(g61943_sb), .b(g61966_db), .o(TIMEBOOST_net_14733) );
in01s01 g65095_u0 ( .a(FE_OFN679_n_4460), .o(g65095_sb) );
na02s01 TIMEBOOST_cell_16524 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(g65723_sb), .o(TIMEBOOST_net_3519) );
na02s01 g65095_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__Q), .b(FE_OFN679_n_4460), .o(g65095_db) );
na02s01 TIMEBOOST_cell_31330 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__Q), .b(g65395_sb), .o(TIMEBOOST_net_9576) );
in01s01 g65096_u0 ( .a(n_4417), .o(g65096_sb) );
na02s02 TIMEBOOST_cell_45175 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__26__Q), .b(n_4387), .o(TIMEBOOST_net_14826) );
na03s02 TIMEBOOST_cell_43329 ( .a(n_3740), .b(FE_OFN1222_n_6391), .c(n_3738), .o(TIMEBOOST_net_13903) );
na02s01 TIMEBOOST_cell_40556 ( .a(TIMEBOOST_net_12516), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_11555) );
in01s01 g65097_u0 ( .a(FE_OFN679_n_4460), .o(g65097_sb) );
na02s01 TIMEBOOST_cell_16525 ( .a(TIMEBOOST_net_3519), .b(g65723_db), .o(n_1748) );
na02s01 g65097_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__Q), .b(FE_OFN679_n_4460), .o(g65097_db) );
no02f02 TIMEBOOST_cell_40213 ( .a(n_15769), .b(n_2416), .o(TIMEBOOST_net_12345) );
in01s01 g65098_u0 ( .a(FE_OFN1660_n_4490), .o(g65098_sb) );
na02s01 TIMEBOOST_cell_16586 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__Q), .b(g64360_sb), .o(TIMEBOOST_net_3550) );
na02s01 g65098_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__Q), .b(FE_OFN1660_n_4490), .o(g65098_db) );
na02f02 TIMEBOOST_cell_42213 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__Q), .b(n_9685), .o(TIMEBOOST_net_13345) );
in01s01 g65099_u0 ( .a(FE_OFN669_n_4505), .o(g65099_sb) );
na02m02 TIMEBOOST_cell_37968 ( .a(g54164_sb), .b(TIMEBOOST_net_11222), .o(TIMEBOOST_net_4342) );
na02s01 g65099_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__Q), .b(FE_OFN669_n_4505), .o(g65099_db) );
na02f02 TIMEBOOST_cell_21906 ( .a(FE_RN_739_0), .b(n_2927), .o(TIMEBOOST_net_6210) );
ao22f02 g65101_u0 ( .a(configuration_wb_err_addr_547), .b(n_15444), .c(n_16000), .d(n_2831), .o(n_3072) );
in01f02 g65102_u0 ( .a(n_2871), .o(n_3071) );
ao22f02 g65103_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_517), .c(configuration_wb_err_data_586), .d(FE_OFN1069_n_15729), .o(n_2871) );
ao22f02 g65104_u0 ( .a(n_14919), .b(n_16810), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_525), .o(n_3070) );
ao22f02 g65105_u0 ( .a(configuration_wb_err_data_587), .b(FE_OFN1069_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2869), .o(n_2870) );
ao22f02 g65106_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_365), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_526), .o(n_3068) );
ao22f02 g65107_u0 ( .a(configuration_wb_err_addr_549), .b(n_15444), .c(n_16000), .d(n_2869), .o(n_3066) );
ao22f02 g65109_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_519), .c(n_14921), .d(n_16810), .o(n_2868) );
ao22f02 g65110_u0 ( .a(configuration_wb_err_data_588), .b(FE_OFN1069_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2866), .o(n_2867) );
ao22f02 g65111_u0 ( .a(configuration_wb_err_addr_550), .b(n_15444), .c(n_16000), .d(n_2866), .o(n_3064) );
ao22f02 g65112_u0 ( .a(configuration_wb_err_data_592), .b(FE_OFN1068_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2864), .o(n_2865) );
ao22f02 g65115_u0 ( .a(FE_OFN1066_n_15808), .b(configuration_pci_err_data_502), .c(n_3371), .d(wbu_pref_en_in_136), .o(n_3374) );
ao22f01 g65116_u0 ( .a(configuration_isr_bit_2975), .b(n_3246), .c(n_3248), .d(configuration_sync_command_bit1), .o(n_3245) );
ao22f02 g65117_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_521), .c(n_14923), .d(n_16810), .o(n_2775) );
ao22f02 g65118_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_368), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_529), .o(n_3062) );
ao22f02 g65119_u0 ( .a(configuration_wb_err_addr_552), .b(n_15444), .c(n_16000), .d(n_2835), .o(n_3061) );
ao22f02 g65120_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_522), .c(n_14924), .d(n_16810), .o(n_2860) );
ao22f01 g65121_u0 ( .a(n_3231), .b(pciu_bar0_in_370), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_531), .o(n_3060) );
ao22f01 g65122_u0 ( .a(configuration_wb_err_addr_554), .b(n_15444), .c(n_16000), .d(n_2864), .o(n_3059) );
ao22f02 g65125_u0 ( .a(FE_OFN1065_n_15808), .b(configuration_pci_err_data_523), .c(n_14925), .d(n_16810), .o(n_2859) );
ao22f02 g65126_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_518), .c(n_14920), .d(n_16810), .o(n_2858) );
ao22f02 g65127_u0 ( .a(configuration_wb_err_data_596), .b(FE_OFN1070_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2856), .o(n_2857) );
ao22f02 g65128_u0 ( .a(configuration_status_bit_435), .b(n_3248), .c(n_16000), .d(n_2841), .o(n_17048) );
ao22f02 g65129_u0 ( .a(FE_OFN1066_n_15808), .b(configuration_pci_err_data_529), .c(configuration_wb_err_cs_bit_567), .d(n_16543), .o(n_3241) );
ao22f02 g65130_u0 ( .a(configuration_status_bit_379), .b(n_3248), .c(n_16000), .d(n_2854), .o(n_17039) );
ao22f02 g65131_u0 ( .a(FE_OFN1066_n_15808), .b(configuration_pci_err_data_530), .c(configuration_wb_err_cs_bit_568), .d(n_16543), .o(n_17027) );
ao22f02 g65132_u0 ( .a(n_14932), .b(n_16810), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_538), .o(n_3058) );
ao22f02 g65133_u0 ( .a(configuration_wb_err_data_599), .b(FE_OFN1070_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2854), .o(n_2855) );
ao22f02 g65134_u0 ( .a(configuration_wb_err_data_573), .b(FE_OFN1071_n_15729), .c(configuration_wb_err_addr_535), .d(n_15445), .o(n_2853) );
ao22f02 g65135_u0 ( .a(n_3372), .b(n_14906), .c(n_3371), .d(n_14907), .o(n_3373) );
ao22f02 g65136_u0 ( .a(configuration_status_bit_351), .b(n_3248), .c(n_16000), .d(n_2851), .o(n_3238) );
ao22f02 g65137_u0 ( .a(FE_OFN1066_n_15808), .b(configuration_pci_err_data_531), .c(configuration_wb_err_cs_bit_569), .d(n_16543), .o(n_3237) );
ao22f02 g65138_u0 ( .a(n_14933), .b(n_16810), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_539), .o(n_3057) );
ao22f02 g65139_u0 ( .a(configuration_wb_err_data_600), .b(FE_OFN1070_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2851), .o(n_2852) );
ao22m02 g65141_u0 ( .a(configuration_wb_err_data_574), .b(FE_OFN1071_n_15729), .c(configuration_wb_err_addr_536), .d(n_15445), .o(n_2849) );
ao22f02 g65142_u0 ( .a(configuration_interrupt_line_40), .b(n_3295), .c(FE_OFN1695_n_3368), .d(wbu_cache_line_size_in_208), .o(n_3370) );
ao22f02 g65143_u0 ( .a(configuration_wb_err_data_575), .b(FE_OFN1071_n_15729), .c(configuration_wb_err_addr_537), .d(n_15445), .o(n_2848) );
ao22f02 g65144_u0 ( .a(configuration_wb_err_cs_bit_564), .b(n_16543), .c(n_3231), .d(pciu_bar0_in_373), .o(n_3236) );
ao22f02 g65145_u0 ( .a(configuration_wb_err_data_576), .b(FE_OFN1071_n_15729), .c(n_3248), .d(configuration_sync_command_bit6), .o(n_3235) );
ao22f02 g65146_u0 ( .a(FE_OFN1066_n_15808), .b(configuration_pci_err_data_507), .c(configuration_wb_err_addr_538), .d(n_15445), .o(n_2847) );
ao22f02 g65147_u0 ( .a(configuration_wb_err_data_577), .b(FE_OFN1071_n_15729), .c(configuration_wb_err_addr_539), .d(n_15445), .o(n_2846) );
ao22f02 g65148_u0 ( .a(configuration_interrupt_line_43), .b(n_3295), .c(FE_OFN1695_n_3368), .d(wbu_cache_line_size_in_211), .o(n_3367) );
ao22m02 g65151_u0 ( .a(configuration_wb_err_addr_546), .b(n_15444), .c(n_16000), .d(n_2809), .o(n_3055) );
ao22f02 g65152_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_366), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_527), .o(n_3054) );
ao22f02 g65153_u0 ( .a(configuration_status_bit_407), .b(n_3248), .c(n_16000), .d(n_2825), .o(n_3233) );
na02s02 TIMEBOOST_cell_17655 ( .a(TIMEBOOST_net_4084), .b(g65364_db), .o(n_4507) );
ao22f02 g65155_u0 ( .a(FE_OFN1065_n_15808), .b(configuration_pci_err_data_526), .c(n_16791), .d(pciu_bar0_in_373), .o(n_2843) );
ao22f02 g65156_u0 ( .a(configuration_wb_err_data_597), .b(FE_OFN1070_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2841), .o(n_2842) );
ao22f02 g65157_u0 ( .a(configuration_wb_err_cs_bit_565), .b(n_16543), .c(n_3231), .d(pciu_bar0_in_374), .o(n_3232) );
ao22f02 g65158_u0 ( .a(configuration_status_bit_322), .b(n_3504), .c(n_16000), .d(n_3592), .o(n_3593) );
ao22f02 g65159_u0 ( .a(FE_OFN1066_n_15808), .b(configuration_pci_err_data_528), .c(configuration_wb_err_cs_bit_566), .d(n_16543), .o(n_17034) );
ao22f02 g65160_u0 ( .a(FE_OFN1065_n_15808), .b(configuration_pci_err_data_527), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_535), .o(n_3053) );
ao22f02 g65161_u0 ( .a(configuration_wb_err_data_601), .b(FE_OFN1070_n_15729), .c(n_16810), .d(n_14934), .o(n_2840) );
ao22f02 g65162_u0 ( .a(n_3231), .b(pciu_bar0_in_379), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_540), .o(n_3052) );
ao22m02 g65163_u0 ( .a(n_16000), .b(n_2838), .c(n_15444), .d(configuration_wb_err_addr_541), .o(n_3051) );
ao22f02 g65164_u0 ( .a(n_14930), .b(n_16810), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_536), .o(n_3050) );
ao22f02 g65165_u0 ( .a(n_15808), .b(configuration_pci_err_data_532), .c(configuration_wb_err_cs_bit_570), .d(n_16543), .o(n_3229) );
ao22f02 g65166_u0 ( .a(FE_OCPN1845_n_16427), .b(n_2838), .c(FE_OFN1068_n_15729), .d(configuration_wb_err_data_579), .o(n_2839) );
ao22f02 g65168_u0 ( .a(n_3252), .b(configuration_pci_err_cs_bit9), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_243), .o(n_2969) );
ao22f02 g65169_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_363), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_524), .o(n_3049) );
ao22f02 g65170_u0 ( .a(configuration_wb_err_data_590), .b(FE_OFN1069_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2835), .o(n_2836) );
ao22f02 g65171_u0 ( .a(configuration_wb_err_data_595), .b(FE_OFN1070_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2833), .o(n_2834) );
ao22f02 g65173_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_369), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_530), .o(n_3048) );
ao22f02 g65174_u0 ( .a(n_14929), .b(n_16810), .c(n_16791), .d(pciu_bar0_in_374), .o(n_2830) );
ao22f02 g65175_u0 ( .a(configuration_wb_err_data_591), .b(FE_OFN1069_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2828), .o(n_2829) );
ao22f04 g65177_u0 ( .a(n_1724), .b(parchk_pci_trdy_en_in), .c(n_2804), .d(conf_wb_err_bc_in), .o(n_3047) );
ao22f02 g65178_u0 ( .a(configuration_wb_err_data_598), .b(FE_OFN1070_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2825), .o(n_2826) );
ao22f02 g65179_u0 ( .a(n_3371), .b(wbu_mrl_en_in_141), .c(FE_OCPN1845_n_16427), .d(pciu_am1_in_540), .o(n_3366) );
ao22f02 g65180_u0 ( .a(configuration_wb_err_cs_bit0), .b(n_16543), .c(n_3372), .d(wbu_mrl_en_in_142), .o(n_3228) );
ao22m02 g65181_u0 ( .a(configuration_cache_line_size_reg), .b(FE_OFN1695_n_3368), .c(n_16000), .d(pciu_am1_in_540), .o(n_3046) );
ao22m01 g65182_u0 ( .a(n_3252), .b(configuration_pci_err_cs_bit0), .c(configuration_interrupt_line), .d(n_3295), .o(n_3365) );
ao22f02 g65183_u0 ( .a(configuration_wb_err_addr_553), .b(n_15445), .c(n_16000), .d(n_2828), .o(n_3045) );
ao22f02 g65184_u0 ( .a(n_3252), .b(configuration_pci_err_cs_bit10), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_244), .o(n_2824) );
ao22f02 g65185_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_511), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_519), .o(n_3044) );
ao22f02 g65186_u0 ( .a(configuration_wb_err_data_580), .b(FE_OFN1068_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2822), .o(n_2823) );
ao22f02 g65187_u0 ( .a(configuration_wb_err_addr_542), .b(n_15445), .c(n_16000), .d(n_2822), .o(n_3043) );
in01s01 TIMEBOOST_cell_45871 ( .a(n_11857), .o(TIMEBOOST_net_15178) );
in01f02 g65189_u0 ( .a(n_2821), .o(n_3042) );
ao22f02 g65190_u0 ( .a(FE_OFN1065_n_15808), .b(configuration_pci_err_data_524), .c(configuration_wb_err_data_593), .d(FE_OFN1068_n_15729), .o(n_2821) );
ao22f02 g65191_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_512), .c(n_14914), .d(n_16810), .o(n_2820) );
ao22f02 g65192_u0 ( .a(configuration_wb_err_data_581), .b(FE_OFN1068_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2818), .o(n_2819) );
in01f02 g65193_u0 ( .a(n_3041), .o(n_3227) );
ao22f02 g65194_u0 ( .a(configuration_wb_err_addr_543), .b(n_15445), .c(n_16000), .d(n_2818), .o(n_3041) );
ao22f02 g65195_u0 ( .a(n_14931), .b(n_16810), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_537), .o(n_3040) );
ao22f01 g65196_u0 ( .a(n_14926), .b(n_16810), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_532), .o(n_3039) );
na02m02 TIMEBOOST_cell_41695 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__Q), .b(n_13447), .o(TIMEBOOST_net_13086) );
ao22f01 g65201_u0 ( .a(n_14915), .b(n_16810), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_521), .o(n_3037) );
ao22m01 g65202_u0 ( .a(configuration_wb_err_addr_544), .b(n_15445), .c(n_16000), .d(n_16428), .o(n_3036) );
ao22f02 g65203_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_514), .c(n_14916), .d(n_16810), .o(n_2814) );
ao22f02 g65204_u0 ( .a(configuration_wb_err_data_583), .b(FE_OFN1069_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2812), .o(n_2813) );
ao22f02 g65205_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_361), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_522), .o(n_3034) );
ao22f01 g65206_u0 ( .a(configuration_wb_err_addr_545), .b(n_15445), .c(n_16000), .d(n_2812), .o(n_3033) );
ao22f02 g65209_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_362), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_523), .o(n_3032) );
in01s01 g65210_u0 ( .a(FE_OFN785_n_2678), .o(g65210_sb) );
na02s01 TIMEBOOST_cell_17042 ( .a(n_3764), .b(g64957_sb), .o(TIMEBOOST_net_3778) );
na02s01 TIMEBOOST_cell_9247 ( .a(TIMEBOOST_net_1190), .b(g65687_db), .o(n_2293) );
na02s01 TIMEBOOST_cell_40558 ( .a(TIMEBOOST_net_12517), .b(g63180_sb), .o(n_5790) );
in01s01 g65211_u0 ( .a(FE_OFN786_n_2678), .o(g65211_sb) );
na02m04 TIMEBOOST_cell_39033 ( .a(wbs_wbb3_2_wbb2_dat_o_i_116), .b(wbs_dat_o_17_), .o(TIMEBOOST_net_11755) );
na02s01 g65211_u2 ( .a(pci_target_unit_pcit_if_strd_bc_in_719), .b(FE_OFN786_n_2678), .o(g65211_db) );
na02f06 TIMEBOOST_cell_41703 ( .a(n_15757), .b(n_15474), .o(TIMEBOOST_net_13090) );
na02s02 TIMEBOOST_cell_42113 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__Q), .b(n_3638), .o(TIMEBOOST_net_13295) );
na02s01 g65212_u2 ( .a(pci_target_unit_wbm_sm_pci_tar_burst_ok), .b(n_2678), .o(g65212_db) );
na02s01 TIMEBOOST_cell_42729 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__Q), .b(n_1700), .o(TIMEBOOST_net_13603) );
in01s01 g65213_u0 ( .a(FE_OFN789_n_2678), .o(g65213_sb) );
na02s01 TIMEBOOST_cell_9299 ( .a(TIMEBOOST_net_1216), .b(g65756_db), .o(n_1700) );
na02s02 g65213_u2 ( .a(pci_target_unit_pcit_if_strd_addr_in_713), .b(FE_OFN789_n_2678), .o(g65213_db) );
na02f02 TIMEBOOST_cell_42492 ( .a(TIMEBOOST_net_13484), .b(g57060_sb), .o(n_10847) );
in01s01 g65214_u0 ( .a(FE_OFN785_n_2678), .o(g65214_sb) );
na03s02 TIMEBOOST_cell_449 ( .a(n_1646), .b(g61810_sb), .c(g61810_db), .o(n_8173) );
na02s02 TIMEBOOST_cell_40560 ( .a(TIMEBOOST_net_12518), .b(g62462_sb), .o(n_6672) );
na02f02 TIMEBOOST_cell_44118 ( .a(TIMEBOOST_net_14297), .b(FE_OFN1376_n_8567), .o(TIMEBOOST_net_13384) );
in01s02 g65215_u0 ( .a(FE_OFN787_n_2678), .o(g65215_sb) );
na02m02 TIMEBOOST_cell_44119 ( .a(n_9026), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__Q), .o(TIMEBOOST_net_14298) );
na02f02 TIMEBOOST_cell_39061 ( .a(TIMEBOOST_net_10136), .b(FE_OFN1770_n_14054), .o(TIMEBOOST_net_11769) );
na02m02 TIMEBOOST_cell_43763 ( .a(n_9141), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__Q), .o(TIMEBOOST_net_14120) );
in01s01 g65216_u0 ( .a(FE_OFN786_n_2678), .o(g65216_sb) );
na02m02 TIMEBOOST_cell_39541 ( .a(FE_OFN1085_n_13221), .b(TIMEBOOST_net_1840), .o(TIMEBOOST_net_12009) );
na02s01 g65216_u2 ( .a(pci_target_unit_del_sync_be_out_reg_0__Q), .b(FE_OFN786_n_2678), .o(g65216_db) );
no02f02 TIMEBOOST_cell_40214 ( .a(TIMEBOOST_net_12345), .b(FE_OFN1506_n_15768), .o(n_11448) );
in01s01 g65217_u0 ( .a(FE_OFN785_n_2678), .o(g65217_sb) );
na02s01 TIMEBOOST_cell_40562 ( .a(TIMEBOOST_net_12519), .b(g63166_sb), .o(n_5806) );
na02s02 TIMEBOOST_cell_40564 ( .a(TIMEBOOST_net_12520), .b(g62681_sb), .o(n_6177) );
in01s01 g65218_u0 ( .a(FE_OFN785_n_2678), .o(g65218_sb) );
na02s01 TIMEBOOST_cell_39200 ( .a(TIMEBOOST_net_11838), .b(g65710_sb), .o(n_1945) );
na02s02 TIMEBOOST_cell_40706 ( .a(TIMEBOOST_net_12591), .b(g62341_sb), .o(n_6917) );
na02s01 TIMEBOOST_cell_16812 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__Q), .b(g65313_sb), .o(TIMEBOOST_net_3663) );
in01s01 g65219_u0 ( .a(FE_OFN785_n_2678), .o(g65219_sb) );
na02m02 TIMEBOOST_cell_41797 ( .a(g52471_da), .b(FE_OFN1023_n_11877), .o(TIMEBOOST_net_13137) );
na02s02 TIMEBOOST_cell_43631 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__Q), .b(n_3788), .o(TIMEBOOST_net_14054) );
na02s01 TIMEBOOST_cell_42601 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__Q), .b(FE_OFN527_n_9899), .o(TIMEBOOST_net_13539) );
in01s01 g65220_u0 ( .a(FE_OFN784_n_2678), .o(g65220_sb) );
na02s02 TIMEBOOST_cell_41790 ( .a(TIMEBOOST_net_13133), .b(g64991_sb), .o(n_4358) );
na02s01 TIMEBOOST_cell_42578 ( .a(TIMEBOOST_net_13527), .b(g60689_sb), .o(n_7215) );
na02s02 TIMEBOOST_cell_41791 ( .a(pci_target_unit_fifos_pciw_addr_data_in_142), .b(g64213_sb), .o(TIMEBOOST_net_13134) );
in01s01 g65221_u0 ( .a(FE_OFN789_n_2678), .o(g65221_sb) );
in01s01 TIMEBOOST_cell_45912 ( .a(TIMEBOOST_net_15218), .o(TIMEBOOST_net_15219) );
na02s01 TIMEBOOST_cell_16140 ( .a(parchk_pci_ad_reg_in_1220), .b(pci_target_unit_del_sync_addr_in_219), .o(TIMEBOOST_net_3327) );
in01s01 g65222_u0 ( .a(FE_OFN784_n_2678), .o(g65222_sb) );
na02f02 TIMEBOOST_cell_42338 ( .a(TIMEBOOST_net_13407), .b(g57479_sb), .o(n_11258) );
na02s01 TIMEBOOST_cell_16141 ( .a(TIMEBOOST_net_3327), .b(FE_OFN2096_n_2520), .o(TIMEBOOST_net_1295) );
na03m04 TIMEBOOST_cell_45529 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_2__Q), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__Q), .c(FE_OFN2157_n_16439), .o(TIMEBOOST_net_15003) );
in01s01 g65223_u0 ( .a(FE_OFN785_n_2678), .o(g65223_sb) );
na02s02 TIMEBOOST_cell_43266 ( .a(TIMEBOOST_net_13871), .b(FE_OFN1247_n_4093), .o(TIMEBOOST_net_12107) );
na02s01 TIMEBOOST_cell_16142 ( .a(parchk_pci_ad_reg_in_1230), .b(pci_target_unit_del_sync_addr_in_229), .o(TIMEBOOST_net_3328) );
na02m04 TIMEBOOST_cell_45530 ( .a(TIMEBOOST_net_15003), .b(g58823_sb), .o(n_8618) );
in01s01 g65224_u0 ( .a(FE_OFN784_n_2678), .o(g65224_sb) );
na02f02 TIMEBOOST_cell_42340 ( .a(TIMEBOOST_net_13408), .b(g57577_sb), .o(n_11174) );
na02s01 TIMEBOOST_cell_16143 ( .a(TIMEBOOST_net_3328), .b(FE_OFN2095_n_2520), .o(TIMEBOOST_net_1297) );
na02m02 TIMEBOOST_cell_42341 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__Q), .b(n_9722), .o(TIMEBOOST_net_13409) );
in01s01 g65225_u0 ( .a(FE_OFN786_n_2678), .o(g65225_sb) );
na02f02 TIMEBOOST_cell_42342 ( .a(TIMEBOOST_net_13409), .b(g57210_sb), .o(TIMEBOOST_net_12327) );
na02s01 g65225_u2 ( .a(pci_target_unit_pcit_if_strd_bc_in_718), .b(FE_OFN786_n_2678), .o(g65225_db) );
na02m02 TIMEBOOST_cell_42343 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__Q), .b(n_9738), .o(TIMEBOOST_net_13410) );
in01s01 g65226_u0 ( .a(FE_OFN785_n_2678), .o(g65226_sb) );
na04m02 TIMEBOOST_cell_34477 ( .a(g52396_db), .b(g52396_sb), .c(n_3137), .d(TIMEBOOST_net_592), .o(n_14825) );
na02s01 TIMEBOOST_cell_16144 ( .a(parchk_pci_ad_reg_in_1223), .b(pci_target_unit_del_sync_addr_in_222), .o(TIMEBOOST_net_3329) );
na03s02 TIMEBOOST_cell_470 ( .a(n_1925), .b(g61752_sb), .c(g61752_db), .o(n_8311) );
in01s01 g65227_u0 ( .a(FE_OFN785_n_2678), .o(g65227_sb) );
na02s01 TIMEBOOST_cell_9259 ( .a(TIMEBOOST_net_1196), .b(g65686_db), .o(n_2209) );
na02s01 TIMEBOOST_cell_16145 ( .a(TIMEBOOST_net_3329), .b(FE_OFN2096_n_2520), .o(TIMEBOOST_net_1300) );
na02s01 TIMEBOOST_cell_9261 ( .a(TIMEBOOST_net_1197), .b(g65689_db), .o(n_2207) );
in01s01 g65228_u0 ( .a(FE_OFN785_n_2678), .o(g65228_sb) );
na02f02 TIMEBOOST_cell_39062 ( .a(TIMEBOOST_net_11769), .b(FE_OFN1774_n_13800), .o(g53167_p) );
na02s01 TIMEBOOST_cell_16146 ( .a(parchk_pci_ad_reg_in_1215), .b(pci_target_unit_del_sync_addr_in_214), .o(TIMEBOOST_net_3330) );
na02f02 TIMEBOOST_cell_39064 ( .a(TIMEBOOST_net_11770), .b(FE_OFN1774_n_13800), .o(g53183_p) );
in01s01 g65229_u0 ( .a(FE_OFN785_n_2678), .o(g65229_sb) );
na02f02 TIMEBOOST_cell_39066 ( .a(TIMEBOOST_net_11771), .b(FE_OFN1774_n_13800), .o(g53210_p) );
na02s01 TIMEBOOST_cell_16147 ( .a(TIMEBOOST_net_3330), .b(FE_OFN2095_n_2520), .o(TIMEBOOST_net_1302) );
na03s01 TIMEBOOST_cell_33965 ( .a(n_1601), .b(g61809_sb), .c(g61809_db), .o(n_8175) );
in01s01 g65230_u0 ( .a(FE_OFN786_n_2678), .o(g65230_sb) );
na02f02 TIMEBOOST_cell_37114 ( .a(TIMEBOOST_net_10795), .b(n_13926), .o(n_16256) );
na02s01 g65230_u2 ( .a(FE_OFN787_n_2678), .b(pci_target_unit_pcit_if_strd_bc_in_717), .o(g65230_db) );
na02f02 TIMEBOOST_cell_37116 ( .a(TIMEBOOST_net_10796), .b(FE_OFN1601_n_13995), .o(g53310_p) );
in01s01 g65231_u0 ( .a(FE_OFN784_n_2678), .o(g65231_sb) );
na03s01 TIMEBOOST_cell_37397 ( .a(n_1584), .b(n_8272), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__Q), .o(TIMEBOOST_net_10937) );
na02s01 TIMEBOOST_cell_16148 ( .a(parchk_pci_ad_reg_in_1235), .b(pci_target_unit_del_sync_addr_in_234), .o(TIMEBOOST_net_3331) );
na02f02 TIMEBOOST_cell_37118 ( .a(TIMEBOOST_net_10797), .b(FE_OFN1600_n_13995), .o(g53163_p) );
in01s01 g65232_u0 ( .a(FE_OFN789_n_2678), .o(g65232_sb) );
na02s02 TIMEBOOST_cell_18573 ( .a(TIMEBOOST_net_4543), .b(g62849_sb), .o(n_5272) );
na02s01 TIMEBOOST_cell_16149 ( .a(TIMEBOOST_net_3331), .b(FE_OFN795_n_2520), .o(TIMEBOOST_net_1307) );
na02f02 TIMEBOOST_cell_37120 ( .a(TIMEBOOST_net_10798), .b(FE_OFN1602_n_13995), .o(g53298_p) );
in01s01 g65233_u0 ( .a(FE_OFN784_n_2678), .o(g65233_sb) );
na02s02 TIMEBOOST_cell_16817 ( .a(TIMEBOOST_net_3665), .b(g65315_db), .o(n_3566) );
na02s01 TIMEBOOST_cell_16150 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__Q), .b(pci_target_unit_fifos_pcir_data_in_179), .o(TIMEBOOST_net_3332) );
na02m02 TIMEBOOST_cell_45531 ( .a(n_2269), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q), .o(TIMEBOOST_net_15004) );
na02s01 TIMEBOOST_cell_8892 ( .a(pci_ad_i_13_), .b(parchk_pci_ad_reg_in_1217), .o(TIMEBOOST_net_1013) );
na02s02 TIMEBOOST_cell_44414 ( .a(TIMEBOOST_net_14445), .b(FE_OFN1305_n_13124), .o(TIMEBOOST_net_13418) );
na02s01 TIMEBOOST_cell_8893 ( .a(TIMEBOOST_net_1013), .b(n_2373), .o(TIMEBOOST_net_742) );
in01s01 g65235_u0 ( .a(FE_OFN786_n_2678), .o(g65235_sb) );
no02f02 TIMEBOOST_cell_40215 ( .a(n_4145), .b(n_12595), .o(TIMEBOOST_net_12346) );
na02s01 g65235_u2 ( .a(pci_target_unit_del_sync_be_out_reg_1__Q), .b(FE_OFN786_n_2678), .o(g65235_db) );
no02f02 TIMEBOOST_cell_40216 ( .a(TIMEBOOST_net_12346), .b(n_4807), .o(g60339_p) );
in01s01 g65236_u0 ( .a(FE_OFN786_n_2678), .o(g65236_sb) );
na02f02 TIMEBOOST_cell_40217 ( .a(n_16836), .b(n_16837), .o(TIMEBOOST_net_12347) );
na02s01 g65236_u2 ( .a(pci_target_unit_del_sync_be_out_reg_2__Q), .b(FE_OFN786_n_2678), .o(g65236_db) );
na02f02 TIMEBOOST_cell_40218 ( .a(TIMEBOOST_net_12347), .b(n_10547), .o(TIMEBOOST_net_683) );
in01s01 g65237_u0 ( .a(FE_OFN785_n_2678), .o(g65237_sb) );
na02m02 TIMEBOOST_cell_30786 ( .a(n_2435), .b(n_2428), .o(TIMEBOOST_net_9304) );
na02f02 TIMEBOOST_cell_45532 ( .a(TIMEBOOST_net_15004), .b(n_13617), .o(TIMEBOOST_net_14588) );
in01s01 g65238_u0 ( .a(FE_OFN789_n_2678), .o(g65238_sb) );
na03f02 TIMEBOOST_cell_45533 ( .a(wbu_addr_in_262), .b(g52597_sb), .c(TIMEBOOST_net_3028), .o(TIMEBOOST_net_15005) );
na02s01 TIMEBOOST_cell_16152 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__Q), .b(pci_target_unit_fifos_pcir_data_in_173), .o(TIMEBOOST_net_3333) );
na02s01 TIMEBOOST_cell_42647 ( .a(FE_OFN250_n_9789), .b(g58257_sb), .o(TIMEBOOST_net_13562) );
na02s01 TIMEBOOST_cell_8894 ( .a(pci_ad_i_22_), .b(parchk_pci_ad_reg_in_1226), .o(TIMEBOOST_net_1014) );
na02s01 g65239_u2 ( .a(FE_OFN787_n_2678), .b(pci_target_unit_pcit_if_strd_bc_in), .o(g65239_db) );
na02s01 TIMEBOOST_cell_8895 ( .a(TIMEBOOST_net_1014), .b(n_2373), .o(TIMEBOOST_net_736) );
in01s01 g65240_u0 ( .a(FE_OFN786_n_2678), .o(g65240_sb) );
na03f02 TIMEBOOST_cell_40219 ( .a(n_9285), .b(n_10093), .c(n_9284), .o(TIMEBOOST_net_12348) );
na02s01 g65240_u2 ( .a(pci_target_unit_del_sync_be_out_reg_3__Q), .b(FE_OFN786_n_2678), .o(g65240_db) );
na02f02 TIMEBOOST_cell_40220 ( .a(TIMEBOOST_net_12348), .b(n_10090), .o(n_12151) );
in01s01 g65241_u0 ( .a(FE_OFN789_n_2678), .o(g65241_sb) );
na02f02 TIMEBOOST_cell_45534 ( .a(TIMEBOOST_net_15005), .b(g52597_db), .o(n_11874) );
na02s01 TIMEBOOST_cell_40499 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__Q), .b(wishbone_slave_unit_pcim_sm_data_in_640), .o(TIMEBOOST_net_12488) );
na02s01 TIMEBOOST_cell_22296 ( .a(g52460_da), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_6405) );
in01s01 g65242_u0 ( .a(FE_OFN789_n_2678), .o(g65242_sb) );
na02f02 TIMEBOOST_cell_32553 ( .a(n_12313), .b(TIMEBOOST_net_10187), .o(TIMEBOOST_net_6559) );
na03s02 TIMEBOOST_cell_37623 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__Q), .b(FE_OFN710_n_8232), .c(n_1940), .o(TIMEBOOST_net_11050) );
na02m02 TIMEBOOST_cell_43731 ( .a(n_9870), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__Q), .o(TIMEBOOST_net_14104) );
in01s01 g65243_u0 ( .a(FE_OFN784_n_2678), .o(g65243_sb) );
na03s02 TIMEBOOST_cell_33371 ( .a(n_4442), .b(g64838_sb), .c(g64838_db), .o(n_4443) );
na02s01 TIMEBOOST_cell_16154 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__Q), .b(pci_target_unit_fifos_pcir_data_in_178), .o(TIMEBOOST_net_3334) );
na02s01 TIMEBOOST_cell_15831 ( .a(TIMEBOOST_net_3172), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_403), .o(TIMEBOOST_net_63) );
in01s01 g65244_u0 ( .a(FE_OFN785_n_2678), .o(g65244_sb) );
na02s02 TIMEBOOST_cell_18693 ( .a(TIMEBOOST_net_4603), .b(g62832_sb), .o(n_5311) );
na02s01 TIMEBOOST_cell_40501 ( .a(wishbone_slave_unit_pcim_sm_data_in_651), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__Q), .o(TIMEBOOST_net_12489) );
na02f02 TIMEBOOST_cell_39068 ( .a(TIMEBOOST_net_11772), .b(FE_OFN1774_n_13800), .o(g53314_p) );
in01s01 g65245_u0 ( .a(FE_OFN789_n_2678), .o(g65245_sb) );
na02f02 TIMEBOOST_cell_39070 ( .a(TIMEBOOST_net_11773), .b(FE_OFN1768_n_14054), .o(n_14507) );
na02s01 TIMEBOOST_cell_16156 ( .a(n_3752), .b(g65077_sb), .o(TIMEBOOST_net_3335) );
na02s01 TIMEBOOST_cell_38522 ( .a(TIMEBOOST_net_11499), .b(g62049_sb), .o(n_7761) );
in01s01 g65246_u0 ( .a(FE_OFN785_n_2678), .o(g65246_sb) );
na02s02 TIMEBOOST_cell_18701 ( .a(TIMEBOOST_net_4607), .b(g62726_sb), .o(n_5528) );
na02s01 TIMEBOOST_cell_16157 ( .a(TIMEBOOST_net_3335), .b(g65077_db), .o(n_3602) );
na02s01 TIMEBOOST_cell_18703 ( .a(TIMEBOOST_net_4608), .b(g62769_sb), .o(n_5456) );
in01s01 g65247_u0 ( .a(FE_OFN785_n_2678), .o(g65247_sb) );
na02s01 TIMEBOOST_cell_38524 ( .a(TIMEBOOST_net_11500), .b(g62065_sb), .o(n_7744) );
na02f02 TIMEBOOST_cell_45535 ( .a(TIMEBOOST_net_10156), .b(FE_OCPN1877_n_13903), .o(TIMEBOOST_net_15006) );
na02s02 TIMEBOOST_cell_18707 ( .a(TIMEBOOST_net_4610), .b(g63065_sb), .o(n_5120) );
in01s01 g65248_u0 ( .a(FE_OFN785_n_2678), .o(g65248_sb) );
na02s01 TIMEBOOST_cell_39202 ( .a(TIMEBOOST_net_11839), .b(n_1586), .o(TIMEBOOST_net_11455) );
na02s02 TIMEBOOST_cell_42648 ( .a(TIMEBOOST_net_13562), .b(g58257_db), .o(n_9540) );
na02s01 TIMEBOOST_cell_18491 ( .a(TIMEBOOST_net_4502), .b(g62745_sb), .o(n_5491) );
in01s01 g65249_u0 ( .a(FE_OFN784_n_2678), .o(g65249_sb) );
na02s02 TIMEBOOST_cell_18717 ( .a(TIMEBOOST_net_4615), .b(g63104_sb), .o(n_5046) );
na02s01 TIMEBOOST_cell_40541 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_3__Q), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_3__Q), .o(TIMEBOOST_net_12509) );
na02s02 TIMEBOOST_cell_18493 ( .a(TIMEBOOST_net_4503), .b(g62748_sb), .o(n_5483) );
in01s01 g65250_u0 ( .a(FE_OFN784_n_2678), .o(g65250_sb) );
na02s02 TIMEBOOST_cell_18719 ( .a(TIMEBOOST_net_4616), .b(g62750_sb), .o(n_5481) );
na02s02 TIMEBOOST_cell_40566 ( .a(TIMEBOOST_net_12521), .b(g62393_sb), .o(n_6812) );
na02s02 TIMEBOOST_cell_18721 ( .a(TIMEBOOST_net_4617), .b(g62751_sb), .o(n_5478) );
in01s01 g65251_u0 ( .a(FE_OFN923_n_4740), .o(g65251_sb) );
na02f02 TIMEBOOST_cell_40222 ( .a(FE_OFN1757_n_12681), .b(TIMEBOOST_net_12349), .o(TIMEBOOST_net_11810) );
na02s01 g65251_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__Q), .b(FE_OFN923_n_4740), .o(g65251_db) );
na02s02 TIMEBOOST_cell_18607 ( .a(TIMEBOOST_net_4560), .b(g62840_sb), .o(n_5293) );
in01s01 g65252_u0 ( .a(FE_OFN1046_n_16657), .o(g65252_sb) );
na02s01 g65252_u1 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(g65252_sb), .o(g65252_da) );
na02s01 g65252_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__Q), .b(FE_OFN1046_n_16657), .o(g65252_db) );
na02m02 TIMEBOOST_cell_45014 ( .a(TIMEBOOST_net_14745), .b(g52646_db), .o(n_14743) );
ao12s01 g65253_u0 ( .a(n_2469), .b(n_2468), .c(pci_target_unit_wbm_sm_pci_tar_read_request), .o(n_2979) );
no02s01 g65254_u0 ( .a(n_568), .b(conf_wb_err_addr_in_945), .o(g65254_p) );
ao12s01 g65254_u1 ( .a(g65254_p), .b(conf_wb_err_addr_in_945), .c(n_568), .o(n_1673) );
no02m02 g65255_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q), .b(n_1224), .o(g65255_p) );
ao12m02 g65255_u1 ( .a(g65255_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q), .c(n_1224), .o(n_2269) );
na03s02 TIMEBOOST_cell_37971 ( .a(TIMEBOOST_net_4174), .b(g65815_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__Q), .o(TIMEBOOST_net_11224) );
na03s02 TIMEBOOST_cell_39461 ( .a(TIMEBOOST_net_3969), .b(g64238_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__18__Q), .o(TIMEBOOST_net_11969) );
na02s01 TIMEBOOST_cell_37970 ( .a(TIMEBOOST_net_11223), .b(g61887_db), .o(n_8056) );
no02s01 g65257_u0 ( .a(n_1674), .b(wbm_adr_o_4_), .o(g65257_p) );
ao12s01 g65257_u1 ( .a(g65257_p), .b(wbm_adr_o_4_), .c(n_1674), .o(n_1675) );
no02s01 g65258_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_), .b(n_1418), .o(g65258_p) );
ao12s01 g65258_u1 ( .a(g65258_p), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_), .c(n_1418), .o(n_1678) );
no02s01 g65259_u0 ( .a(wbu_addr_in_256), .b(n_2225), .o(g65259_p) );
ao12s01 g65259_u1 ( .a(g65259_p), .b(wbu_addr_in_256), .c(n_2225), .o(n_2226) );
no02s01 g65260_u0 ( .a(wbu_addr_in_253), .b(n_1679), .o(g65260_p) );
ao12s01 g65260_u1 ( .a(g65260_p), .b(wbu_addr_in_253), .c(n_1679), .o(n_1680) );
no02s01 g65261_u0 ( .a(n_1985), .b(wbm_adr_o_7_), .o(g65261_p) );
ao12s01 g65261_u1 ( .a(g65261_p), .b(wbm_adr_o_7_), .c(n_1985), .o(n_2224) );
in01s01 g65262_u0 ( .a(FE_OFN1012_n_4734), .o(g65262_sb) );
na02s01 g65262_u1 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(g65262_sb), .o(g65262_da) );
na02s01 g65262_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__Q), .b(FE_OFN1012_n_4734), .o(g65262_db) );
na02s01 g65262_u3 ( .a(g65262_da), .b(g65262_db), .o(n_3588) );
no02s01 g65263_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_2_), .b(n_733), .o(g65263_p) );
ao12s01 g65263_u1 ( .a(g65263_p), .b(pci_target_unit_del_sync_comp_cycle_count_2_), .c(n_733), .o(n_1424) );
no02s01 g65264_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_), .b(n_554), .o(g65264_p) );
ao12s01 g65264_u1 ( .a(g65264_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_), .c(n_554), .o(n_1423) );
no02s02 g65265_u0 ( .a(conf_wb_err_addr_in_948), .b(n_1561), .o(g65265_p) );
ao12s02 g65265_u1 ( .a(g65265_p), .b(conf_wb_err_addr_in_948), .c(n_1561), .o(n_2395) );
no02s01 g65266_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_2_), .b(n_566), .o(g65266_p) );
ao12s01 g65266_u1 ( .a(g65266_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_2_), .c(n_566), .o(n_1422) );
no02s01 g65267_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_), .b(n_1215), .o(g65267_p) );
ao12s01 g65267_u1 ( .a(g65267_p), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_), .c(n_1215), .o(n_1421) );
in01s01 g65268_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .o(g65268_sb) );
na02s01 g65268_u1 ( .a(n_1109), .b(g65268_sb), .o(g65268_da) );
na02s02 TIMEBOOST_cell_43383 ( .a(n_3616), .b(n_3617), .o(TIMEBOOST_net_13930) );
na03f02 TIMEBOOST_cell_36217 ( .a(FE_OCP_RBN1974_n_12381), .b(TIMEBOOST_net_10301), .c(FE_OFN1755_n_12681), .o(n_12767) );
in01s01 g65269_u0 ( .a(FE_OCPN1839_n_1238), .o(g65269_sb) );
na02s01 TIMEBOOST_cell_17222 ( .a(n_4645), .b(FE_OFN1640_n_4671), .o(TIMEBOOST_net_3868) );
na02m02 TIMEBOOST_cell_41696 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_399), .b(TIMEBOOST_net_13086), .o(TIMEBOOST_net_9630) );
na02m02 TIMEBOOST_cell_41593 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_17__Q), .b(FE_OFN219_n_9853), .o(TIMEBOOST_net_13035) );
in01s01 g65270_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .o(g65270_sb) );
na02s01 TIMEBOOST_cell_41937 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__Q), .b(g58439_sb), .o(TIMEBOOST_net_13207) );
in01s01 TIMEBOOST_cell_45884 ( .a(TIMEBOOST_net_15190), .o(TIMEBOOST_net_15191) );
na03f20 TIMEBOOST_cell_42 ( .a(n_15317), .b(n_16818), .c(n_15314), .o(n_15414) );
in01s01 g65271_u0 ( .a(FE_OFN652_n_4508), .o(g65271_sb) );
na02s01 g65271_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__Q), .b(g65271_sb), .o(g65271_da) );
na02f04 TIMEBOOST_cell_40224 ( .a(FE_OFN1755_n_12681), .b(TIMEBOOST_net_12350), .o(TIMEBOOST_net_11811) );
na02f02 TIMEBOOST_cell_40225 ( .a(FE_OFN1739_n_11019), .b(TIMEBOOST_net_10289), .o(TIMEBOOST_net_12351) );
in01s01 g65272_u0 ( .a(n_4677), .o(g65272_sb) );
na02s01 g65272_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__Q), .b(g65272_sb), .o(g65272_da) );
na03f02 TIMEBOOST_cell_36113 ( .a(FE_RN_471_0), .b(n_10676), .c(n_12578), .o(n_12840) );
na02f02 TIMEBOOST_cell_37122 ( .a(TIMEBOOST_net_10799), .b(FE_OFN1599_n_13995), .o(g53231_p) );
in01s01 g65273_u0 ( .a(FE_OFN643_n_4677), .o(g65273_sb) );
na02s01 g65273_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__Q), .b(g65273_sb), .o(g65273_da) );
na02s02 TIMEBOOST_cell_31329 ( .a(TIMEBOOST_net_9575), .b(g65362_db), .o(n_3536) );
na02f02 TIMEBOOST_cell_40226 ( .a(TIMEBOOST_net_12351), .b(FE_OFN1734_n_16317), .o(n_12501) );
in01s01 g65274_u0 ( .a(FE_OFN1642_n_4671), .o(g65274_sb) );
na02s02 TIMEBOOST_cell_44427 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_766), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_1__Q), .o(TIMEBOOST_net_14452) );
na02f02 TIMEBOOST_cell_40227 ( .a(FE_OFN1759_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__Q), .o(TIMEBOOST_net_12352) );
na02f02 TIMEBOOST_cell_40228 ( .a(TIMEBOOST_net_963), .b(TIMEBOOST_net_12352), .o(n_12516) );
in01s01 g65275_u0 ( .a(FE_OFN643_n_4677), .o(g65275_sb) );
na02s01 g65275_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__Q), .b(g65275_sb), .o(g65275_da) );
na02f02 TIMEBOOST_cell_44498 ( .a(TIMEBOOST_net_14487), .b(FE_OFN1427_n_8567), .o(TIMEBOOST_net_13449) );
na02f02 TIMEBOOST_cell_40230 ( .a(n_12312), .b(TIMEBOOST_net_12353), .o(n_12747) );
in01s01 g65276_u0 ( .a(FE_OFN643_n_4677), .o(g65276_sb) );
na02s01 TIMEBOOST_cell_8896 ( .a(pci_ad_i_17_), .b(parchk_pci_ad_reg_in_1221), .o(TIMEBOOST_net_1015) );
na02s01 g65276_u2 ( .a(n_3747), .b(FE_OFN643_n_4677), .o(g65276_db) );
na02s01 TIMEBOOST_cell_8897 ( .a(TIMEBOOST_net_1015), .b(n_2373), .o(TIMEBOOST_net_737) );
in01s01 g65277_u0 ( .a(FE_OFN642_n_4677), .o(g65277_sb) );
na02s01 TIMEBOOST_cell_8898 ( .a(pci_ad_i_7_), .b(parchk_pci_ad_reg_in_1211), .o(TIMEBOOST_net_1016) );
na02s01 g65277_u2 ( .a(n_3777), .b(FE_OFN642_n_4677), .o(g65277_db) );
na02s01 TIMEBOOST_cell_8899 ( .a(TIMEBOOST_net_1016), .b(n_2373), .o(TIMEBOOST_net_738) );
in01s01 g65278_u0 ( .a(FE_OFN642_n_4677), .o(g65278_sb) );
na02s01 TIMEBOOST_cell_8900 ( .a(pci_ad_i_0_), .b(parchk_pci_ad_reg_in), .o(TIMEBOOST_net_1017) );
na02s01 g65278_u2 ( .a(n_4476), .b(FE_OFN642_n_4677), .o(g65278_db) );
na02s01 TIMEBOOST_cell_8901 ( .a(TIMEBOOST_net_1017), .b(n_2373), .o(TIMEBOOST_net_739) );
in01s01 g65279_u0 ( .a(FE_OFN643_n_4677), .o(g65279_sb) );
na02s01 TIMEBOOST_cell_8902 ( .a(pci_ad_i_4_), .b(parchk_pci_ad_reg_in_1208), .o(TIMEBOOST_net_1018) );
na02s01 g65279_u2 ( .a(n_3744), .b(FE_OFN643_n_4677), .o(g65279_db) );
na02s01 TIMEBOOST_cell_8903 ( .a(TIMEBOOST_net_1018), .b(n_2373), .o(TIMEBOOST_net_740) );
in01s01 g65280_u0 ( .a(FE_OFN643_n_4677), .o(g65280_sb) );
na02s01 g65280_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__Q), .b(g65280_sb), .o(g65280_da) );
na02s02 TIMEBOOST_cell_40568 ( .a(TIMEBOOST_net_12522), .b(g62994_sb), .o(n_5894) );
na02s01 TIMEBOOST_cell_44990 ( .a(TIMEBOOST_net_14733), .b(g63611_db), .o(TIMEBOOST_net_13155) );
in01s01 g65281_u0 ( .a(FE_OFN643_n_4677), .o(g65281_sb) );
na02s01 g65281_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__Q), .b(g65281_sb), .o(g65281_da) );
na02f02 TIMEBOOST_cell_40232 ( .a(n_12433), .b(TIMEBOOST_net_12354), .o(n_12733) );
na02s01 TIMEBOOST_cell_42649 ( .a(g64102_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__Q), .o(TIMEBOOST_net_13563) );
in01s01 g65282_u0 ( .a(FE_OFN644_n_4677), .o(g65282_sb) );
na02s01 TIMEBOOST_cell_8904 ( .a(n_1412), .b(n_1674), .o(TIMEBOOST_net_1019) );
na02s01 g65282_u2 ( .a(n_4470), .b(FE_OFN644_n_4677), .o(g65282_db) );
na02s01 TIMEBOOST_cell_8905 ( .a(TIMEBOOST_net_1019), .b(n_2235), .o(TIMEBOOST_net_102) );
in01s01 g65283_u0 ( .a(FE_OFN642_n_4677), .o(g65283_sb) );
na02f02 TIMEBOOST_cell_44398 ( .a(TIMEBOOST_net_14437), .b(FE_OFN1383_n_8567), .o(TIMEBOOST_net_12688) );
na02s01 g65283_u2 ( .a(n_3741), .b(FE_OFN642_n_4677), .o(g65283_db) );
na02f02 TIMEBOOST_cell_43732 ( .a(TIMEBOOST_net_14104), .b(FE_OFN1397_n_8567), .o(TIMEBOOST_net_12699) );
in01s01 g65284_u0 ( .a(FE_OFN642_n_4677), .o(g65284_sb) );
na02s01 TIMEBOOST_cell_8908 ( .a(pci_target_unit_del_sync_comp_cycle_count_10_), .b(pci_target_unit_del_sync_comp_cycle_count_11_), .o(TIMEBOOST_net_1021) );
na02s01 g65284_u2 ( .a(n_3785), .b(FE_OFN642_n_4677), .o(g65284_db) );
na02s01 TIMEBOOST_cell_8909 ( .a(TIMEBOOST_net_1021), .b(n_523), .o(TIMEBOOST_net_164) );
in01s01 g65285_u0 ( .a(FE_OFN644_n_4677), .o(g65285_sb) );
na02s01 g65285_u2 ( .a(n_4482), .b(FE_OFN644_n_4677), .o(g65285_db) );
na02f02 TIMEBOOST_cell_44438 ( .a(TIMEBOOST_net_14457), .b(g57875_sb), .o(n_8921) );
in01s01 g65286_u0 ( .a(n_4677), .o(g65286_sb) );
in01s01 TIMEBOOST_cell_45913 ( .a(wbm_dat_i_16_), .o(TIMEBOOST_net_15220) );
na02m02 TIMEBOOST_cell_38822 ( .a(TIMEBOOST_net_11649), .b(g58459_sb), .o(n_9396) );
na02f02 TIMEBOOST_cell_44410 ( .a(TIMEBOOST_net_14443), .b(FE_OFN1404_n_8567), .o(n_10400) );
in01s01 g65287_u0 ( .a(FE_OFN643_n_4677), .o(g65287_sb) );
na02s01 g65287_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__Q), .b(g65287_sb), .o(g65287_da) );
na02f02 TIMEBOOST_cell_40233 ( .a(FE_OFN1554_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__Q), .o(TIMEBOOST_net_12355) );
na02f02 TIMEBOOST_cell_40234 ( .a(n_12113), .b(TIMEBOOST_net_12355), .o(n_12624) );
in01s01 g65288_u0 ( .a(FE_OFN644_n_4677), .o(g65288_sb) );
na02s01 TIMEBOOST_cell_8912 ( .a(TIMEBOOST_net_718), .b(wishbone_slave_unit_wishbone_slave_pref_en_reg_Q), .o(TIMEBOOST_net_1023) );
na02s01 g65288_u2 ( .a(n_3739), .b(FE_OFN644_n_4677), .o(g65288_db) );
na02s01 TIMEBOOST_cell_8913 ( .a(TIMEBOOST_net_1023), .b(wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q), .o(n_1721) );
in01s01 g65289_u0 ( .a(FE_OFN644_n_4677), .o(g65289_sb) );
na02s01 TIMEBOOST_cell_8914 ( .a(pci_target_unit_del_sync_comp_cycle_count_9_), .b(pci_target_unit_del_sync_comp_cycle_count_10_), .o(TIMEBOOST_net_1024) );
na02s01 g65289_u2 ( .a(n_3755), .b(FE_OFN644_n_4677), .o(g65289_db) );
na02s01 TIMEBOOST_cell_8915 ( .a(TIMEBOOST_net_1024), .b(n_1989), .o(TIMEBOOST_net_96) );
na02s01 g65290_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__Q), .b(g65272_sb), .o(g65290_da) );
na02f02 TIMEBOOST_cell_41106 ( .a(TIMEBOOST_net_12791), .b(g57378_sb), .o(n_11370) );
na02s01 TIMEBOOST_cell_15829 ( .a(TIMEBOOST_net_3171), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_400), .o(TIMEBOOST_net_61) );
in01s01 g65291_u0 ( .a(n_4677), .o(g65291_sb) );
na02s01 g65291_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__Q), .b(g65291_sb), .o(g65291_da) );
na02f02 TIMEBOOST_cell_10169 ( .a(TIMEBOOST_net_1651), .b(FE_OFN1147_n_13249), .o(TIMEBOOST_net_487) );
na03s02 TIMEBOOST_cell_318 ( .a(FE_OFN2079_n_8069), .b(pci_target_unit_fifos_pcir_whole_waddr_94), .c(n_8503), .o(n_8505) );
in01s01 g65292_u0 ( .a(FE_OFN642_n_4677), .o(g65292_sb) );
na02s01 g65292_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__26__Q), .b(g65292_sb), .o(g65292_da) );
na02s01 TIMEBOOST_cell_16532 ( .a(pci_target_unit_fifos_pcir_data_in_188), .b(g65739_sb), .o(TIMEBOOST_net_3523) );
na02s01 TIMEBOOST_cell_16533 ( .a(TIMEBOOST_net_3523), .b(g65739_db), .o(n_1932) );
in01s01 g65293_u0 ( .a(FE_OFN644_n_4677), .o(g65293_sb) );
na02s02 g65293_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__Q), .b(g65293_sb), .o(g65293_da) );
na02s01 TIMEBOOST_cell_16534 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(g65740_sb), .o(TIMEBOOST_net_3524) );
na02s02 TIMEBOOST_cell_31328 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__Q), .b(g65362_sb), .o(TIMEBOOST_net_9575) );
in01s01 g65294_u0 ( .a(FE_OFN636_n_4669), .o(g65294_sb) );
na02s02 TIMEBOOST_cell_45176 ( .a(TIMEBOOST_net_14826), .b(FE_OFN1241_n_4092), .o(TIMEBOOST_net_12550) );
na02s01 g65294_u2 ( .a(n_4488), .b(FE_OFN636_n_4669), .o(g65294_db) );
na02s01 TIMEBOOST_cell_16588 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__Q), .b(g64361_sb), .o(TIMEBOOST_net_3551) );
in01s01 g65295_u0 ( .a(FE_OFN640_n_4669), .o(g65295_sb) );
na02s02 TIMEBOOST_cell_45115 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__Q), .b(n_3985), .o(TIMEBOOST_net_14796) );
na02m02 TIMEBOOST_cell_40221 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__Q), .o(TIMEBOOST_net_12349) );
na02s01 TIMEBOOST_cell_16590 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__Q), .b(g64362_sb), .o(TIMEBOOST_net_3552) );
in01s01 g65296_u0 ( .a(FE_OFN639_n_4669), .o(g65296_sb) );
na02s02 TIMEBOOST_cell_45116 ( .a(TIMEBOOST_net_14796), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_11418) );
na02s01 g65296_u2 ( .a(n_3777), .b(FE_OFN639_n_4669), .o(g65296_db) );
na02s01 TIMEBOOST_cell_16592 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__Q), .b(g64363_sb), .o(TIMEBOOST_net_3553) );
in01s01 g65297_u0 ( .a(FE_OFN639_n_4669), .o(g65297_sb) );
na02s02 TIMEBOOST_cell_45193 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__Q), .b(n_3751), .o(TIMEBOOST_net_14835) );
na02s02 g65297_u2 ( .a(n_4476), .b(FE_OFN639_n_4669), .o(g65297_db) );
na02s01 TIMEBOOST_cell_44991 ( .a(g61943_sb), .b(g61970_db), .o(TIMEBOOST_net_14734) );
in01s01 g65298_u0 ( .a(FE_OFN640_n_4669), .o(g65298_sb) );
na02f02 TIMEBOOST_cell_40236 ( .a(n_11927), .b(TIMEBOOST_net_12356), .o(n_12493) );
na02s01 TIMEBOOST_cell_17650 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__Q), .b(g65389_sb), .o(TIMEBOOST_net_4082) );
na02f02 TIMEBOOST_cell_40237 ( .a(FE_OFN1558_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__Q), .o(TIMEBOOST_net_12357) );
in01s01 g65299_u0 ( .a(FE_OFN640_n_4669), .o(g65299_sb) );
na02f02 TIMEBOOST_cell_40238 ( .a(n_12227), .b(TIMEBOOST_net_12357), .o(n_12656) );
na02s01 TIMEBOOST_cell_17658 ( .a(n_4273), .b(g65306_sb), .o(TIMEBOOST_net_4086) );
na02s01 TIMEBOOST_cell_16598 ( .a(n_3739), .b(g64822_sb), .o(TIMEBOOST_net_3556) );
in01s01 g65300_u0 ( .a(FE_OFN640_n_4669), .o(g65300_sb) );
na02s01 TIMEBOOST_cell_16599 ( .a(TIMEBOOST_net_3556), .b(g64822_db), .o(n_3736) );
na02s01 TIMEBOOST_cell_16600 ( .a(n_3755), .b(g64823_sb), .o(TIMEBOOST_net_3557) );
in01s01 g65301_u0 ( .a(FE_OFN640_n_4669), .o(g65301_sb) );
na02s01 TIMEBOOST_cell_16601 ( .a(TIMEBOOST_net_3557), .b(g64823_db), .o(n_3735) );
na02s01 TIMEBOOST_cell_38772 ( .a(TIMEBOOST_net_11624), .b(g53900_sb), .o(n_13543) );
na02s02 TIMEBOOST_cell_16602 ( .a(n_3783), .b(g64825_sb), .o(TIMEBOOST_net_3558) );
in01s01 g65302_u0 ( .a(FE_OFN639_n_4669), .o(g65302_sb) );
na02s02 TIMEBOOST_cell_16603 ( .a(TIMEBOOST_net_3558), .b(g64825_db), .o(n_3733) );
na02s01 g65302_u2 ( .a(n_3741), .b(FE_OFN639_n_4669), .o(g65302_db) );
na02s02 TIMEBOOST_cell_43543 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__Q), .b(n_3683), .o(TIMEBOOST_net_14010) );
in01s01 g65303_u0 ( .a(FE_OFN642_n_4677), .o(g65303_sb) );
na02s01 TIMEBOOST_cell_16928 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__Q), .b(g65283_sb), .o(TIMEBOOST_net_3721) );
na02s01 g65303_u2 ( .a(n_4465), .b(FE_OFN642_n_4677), .o(g65303_db) );
na02s01 TIMEBOOST_cell_16929 ( .a(TIMEBOOST_net_3721), .b(g65283_db), .o(n_3583) );
in01s01 g65304_u0 ( .a(FE_OFN639_n_4669), .o(g65304_sb) );
na02s03 TIMEBOOST_cell_40240 ( .a(TIMEBOOST_net_12358), .b(n_928), .o(TIMEBOOST_net_244) );
na02s01 g65304_u2 ( .a(n_3785), .b(FE_OFN639_n_4669), .o(g65304_db) );
na02s02 TIMEBOOST_cell_40570 ( .a(TIMEBOOST_net_12523), .b(g62502_sb), .o(n_6578) );
in01s01 g65305_u0 ( .a(FE_OFN640_n_4669), .o(g65305_sb) );
na02s01 TIMEBOOST_cell_16607 ( .a(TIMEBOOST_net_3560), .b(n_4488), .o(n_4261) );
na02s01 g65305_u2 ( .a(n_4482), .b(FE_OFN640_n_4669), .o(g65305_db) );
na02s01 TIMEBOOST_cell_40241 ( .a(g58783_sb), .b(n_8831), .o(TIMEBOOST_net_12359) );
in01s01 g65306_u0 ( .a(FE_OFN636_n_4669), .o(g65306_sb) );
na02s01 TIMEBOOST_cell_40242 ( .a(TIMEBOOST_net_12359), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_24__Q), .o(TIMEBOOST_net_10371) );
na02s01 g65306_u2 ( .a(n_4479), .b(FE_OFN636_n_4669), .o(g65306_db) );
na02s01 TIMEBOOST_cell_16610 ( .a(n_4479), .b(g64891_sb), .o(TIMEBOOST_net_3562) );
in01s01 g65307_u0 ( .a(FE_OFN640_n_4669), .o(g65307_sb) );
na02s01 TIMEBOOST_cell_40359 ( .a(n_4473), .b(g65042_sb), .o(TIMEBOOST_net_12418) );
na02s01 g65307_u2 ( .a(n_3770), .b(FE_OFN640_n_4669), .o(g65307_db) );
na02s03 TIMEBOOST_cell_40239 ( .a(n_245), .b(n_193), .o(TIMEBOOST_net_12358) );
in01s01 g65308_u0 ( .a(FE_OFN636_n_4669), .o(g65308_sb) );
na02m02 TIMEBOOST_cell_40244 ( .a(g58793_db), .b(TIMEBOOST_net_12360), .o(n_9116) );
na02s01 g65308_u2 ( .a(n_4498), .b(FE_OFN636_n_4669), .o(g65308_db) );
na02f02 TIMEBOOST_cell_45536 ( .a(TIMEBOOST_net_15006), .b(FE_OCP_RBN1962_FE_OFN1591_n_13741), .o(n_14298) );
in01s01 g65309_u0 ( .a(n_4669), .o(g65309_sb) );
na02s01 g65309_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__Q), .b(g65309_sb), .o(g65309_da) );
na02s01 g65309_u2 ( .a(n_3739), .b(n_4669), .o(g65309_db) );
na02s01 g65309_u3 ( .a(g65309_da), .b(g65309_db), .o(n_3571) );
in01s01 g65310_u0 ( .a(n_4669), .o(g65310_sb) );
na02s01 g65310_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__Q), .b(g65310_sb), .o(g65310_da) );
na02s01 g65310_u2 ( .a(n_3755), .b(n_4669), .o(g65310_db) );
na02s01 g65310_u3 ( .a(g65310_da), .b(g65310_db), .o(n_3570) );
in01s01 g65311_u0 ( .a(FE_OFN636_n_4669), .o(g65311_sb) );
no02f02 TIMEBOOST_cell_40246 ( .a(TIMEBOOST_net_12361), .b(FE_RN_330_0), .o(FE_RN_333_0) );
na02s01 g65311_u2 ( .a(n_3764), .b(FE_OFN636_n_4669), .o(g65311_db) );
no02f02 TIMEBOOST_cell_40245 ( .a(FE_RN_328_0), .b(FE_RN_332_0), .o(TIMEBOOST_net_12361) );
in01s01 g65312_u0 ( .a(FE_OFN636_n_4669), .o(g65312_sb) );
na02s01 TIMEBOOST_cell_17852 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__Q), .b(g65349_sb), .o(TIMEBOOST_net_4183) );
na02f02 TIMEBOOST_cell_21907 ( .a(TIMEBOOST_net_6210), .b(n_4654), .o(n_5724) );
na02s02 TIMEBOOST_cell_40626 ( .a(TIMEBOOST_net_12551), .b(g62335_sb), .o(n_6929) );
in01s01 g65313_u0 ( .a(FE_OFN1642_n_4671), .o(g65313_sb) );
na02s02 TIMEBOOST_cell_40248 ( .a(TIMEBOOST_net_12362), .b(n_2426), .o(TIMEBOOST_net_145) );
na02s01 g65313_u2 ( .a(n_3761), .b(FE_OFN1642_n_4671), .o(g65313_db) );
na02s02 TIMEBOOST_cell_40766 ( .a(TIMEBOOST_net_12621), .b(g63003_sb), .o(n_5876) );
in01s01 g65314_u0 ( .a(FE_OFN1643_n_4671), .o(g65314_sb) );
na02s01 TIMEBOOST_cell_16619 ( .a(TIMEBOOST_net_3566), .b(g64816_sb), .o(n_4458) );
na02s01 g65314_u2 ( .a(n_3777), .b(FE_OFN1643_n_4671), .o(g65314_db) );
na02m02 TIMEBOOST_cell_40209 ( .a(wbs_wbb3_2_wbb2_dat_o_i_107), .b(wbs_dat_o_8_), .o(TIMEBOOST_net_12343) );
in01s01 g65315_u0 ( .a(FE_OFN1642_n_4671), .o(g65315_sb) );
na02m02 TIMEBOOST_cell_40250 ( .a(n_14070), .b(TIMEBOOST_net_12363), .o(TIMEBOOST_net_703) );
na02s01 g65315_u2 ( .a(n_3744), .b(FE_OFN1642_n_4671), .o(g65315_db) );
na02s01 TIMEBOOST_cell_40251 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__Q), .b(FE_OFN607_n_9904), .o(TIMEBOOST_net_12364) );
in01s01 g65316_u0 ( .a(FE_OFN1642_n_4671), .o(g65316_sb) );
na02s02 g65316_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__Q), .b(g65316_sb), .o(g65316_da) );
na02f02 TIMEBOOST_cell_36964 ( .a(TIMEBOOST_net_10720), .b(g58832_sb), .o(n_8605) );
na02s02 TIMEBOOST_cell_42858 ( .a(TIMEBOOST_net_13667), .b(FE_OFN2212_n_8407), .o(TIMEBOOST_net_11146) );
in01s01 g65317_u0 ( .a(FE_OFN1642_n_4671), .o(g65317_sb) );
na02s01 TIMEBOOST_cell_40252 ( .a(TIMEBOOST_net_12364), .b(g58051_sb), .o(TIMEBOOST_net_9340) );
na02s01 g65317_u2 ( .a(n_3774), .b(FE_OFN1642_n_4671), .o(g65317_db) );
na02f02 TIMEBOOST_cell_40253 ( .a(FE_RN_593_0), .b(FE_RN_602_0), .o(TIMEBOOST_net_12365) );
in01s01 g65318_u0 ( .a(FE_OFN1642_n_4671), .o(g65318_sb) );
na02f02 TIMEBOOST_cell_40254 ( .a(TIMEBOOST_net_12365), .b(FE_RN_606_0), .o(TIMEBOOST_net_459) );
na02s01 g65318_u2 ( .a(n_3752), .b(FE_OFN1642_n_4671), .o(g65318_db) );
na02s01 TIMEBOOST_cell_16626 ( .a(n_3755), .b(g64800_sb), .o(TIMEBOOST_net_3570) );
in01s01 g65319_u0 ( .a(FE_OFN1643_n_4671), .o(g65319_sb) );
na02s01 TIMEBOOST_cell_16627 ( .a(TIMEBOOST_net_3570), .b(g64800_db), .o(n_3756) );
na02s01 g65319_u2 ( .a(n_3741), .b(FE_OFN1643_n_4671), .o(g65319_db) );
na02s01 TIMEBOOST_cell_16628 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__Q), .b(g65417_sb), .o(TIMEBOOST_net_3571) );
in01s01 g65320_u0 ( .a(FE_OFN1644_n_4671), .o(g65320_sb) );
na02s01 g65320_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__Q), .b(g65320_sb), .o(g65320_da) );
na02s01 TIMEBOOST_cell_16535 ( .a(TIMEBOOST_net_3524), .b(g65740_db), .o(n_1931) );
na02s01 TIMEBOOST_cell_16536 ( .a(pci_target_unit_fifos_pcir_data_in_187), .b(g65742_sb), .o(TIMEBOOST_net_3525) );
in01s01 g65321_u0 ( .a(FE_OFN1642_n_4671), .o(g65321_sb) );
na02s02 TIMEBOOST_cell_16631 ( .a(TIMEBOOST_net_3572), .b(g65330_db), .o(n_3554) );
na02s01 g65321_u2 ( .a(n_3770), .b(FE_OFN1642_n_4671), .o(g65321_db) );
na02s02 TIMEBOOST_cell_31077 ( .a(TIMEBOOST_net_9449), .b(g65013_db), .o(n_4345) );
in01s01 g65322_u0 ( .a(FE_OFN1640_n_4671), .o(g65322_sb) );
na02s01 g65322_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__Q), .b(g65322_sb), .o(g65322_da) );
na02s01 TIMEBOOST_cell_16537 ( .a(TIMEBOOST_net_3525), .b(g65742_db), .o(n_1929) );
na02s01 TIMEBOOST_cell_16538 ( .a(pci_target_unit_fifos_pcir_data_in_174), .b(g65743_sb), .o(TIMEBOOST_net_3526) );
in01s01 g65323_u0 ( .a(FE_OFN1640_n_4671), .o(g65323_sb) );
na02s02 TIMEBOOST_cell_31076 ( .a(n_4465), .b(g65013_sb), .o(TIMEBOOST_net_9449) );
na02s01 g65323_u2 ( .a(n_3739), .b(FE_OFN1640_n_4671), .o(g65323_db) );
na02s02 TIMEBOOST_cell_45689 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__Q), .b(n_4287), .o(TIMEBOOST_net_15083) );
in01s01 g65324_u0 ( .a(FE_OFN1645_n_4671), .o(g65324_sb) );
na02s01 TIMEBOOST_cell_16636 ( .a(n_3755), .b(g64971_sb), .o(TIMEBOOST_net_3575) );
na02s01 g65324_u2 ( .a(n_3780), .b(FE_OFN1645_n_4671), .o(g65324_db) );
na03s02 TIMEBOOST_cell_45117 ( .a(TIMEBOOST_net_443), .b(FE_OFN1138_g64577_p), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__Q), .o(TIMEBOOST_net_14797) );
in01s01 g65325_u0 ( .a(n_4671), .o(g65325_sb) );
na02s01 g65325_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__Q), .b(g65325_sb), .o(g65325_da) );
na03s02 TIMEBOOST_cell_319 ( .a(FE_OFN2079_n_8069), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_), .c(n_8503), .o(n_8504) );
na02f02 TIMEBOOST_cell_45537 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q), .b(n_13903), .o(TIMEBOOST_net_15007) );
in01s01 g65326_u0 ( .a(FE_OFN1644_n_4671), .o(g65326_sb) );
na02s01 g65326_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__Q), .b(g65326_sb), .o(g65326_da) );
na02s01 TIMEBOOST_cell_16539 ( .a(TIMEBOOST_net_3526), .b(g65743_db), .o(n_1928) );
na02s01 TIMEBOOST_cell_31327 ( .a(TIMEBOOST_net_9574), .b(g65353_db), .o(n_3540) );
in01s01 g65327_u0 ( .a(FE_OFN654_n_4508), .o(g65327_sb) );
na02s01 TIMEBOOST_cell_31074 ( .a(n_4482), .b(g65012_sb), .o(TIMEBOOST_net_9448) );
na02s01 g65327_u2 ( .a(n_3747), .b(FE_OFN654_n_4508), .o(g65327_db) );
na02s01 TIMEBOOST_cell_40255 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__Q), .b(n_2300), .o(TIMEBOOST_net_12366) );
in01s01 g65328_u0 ( .a(FE_OFN652_n_4508), .o(g65328_sb) );
na02s02 TIMEBOOST_cell_40680 ( .a(TIMEBOOST_net_12578), .b(g62474_sb), .o(n_6641) );
na02s01 g65328_u2 ( .a(n_3777), .b(FE_OFN652_n_4508), .o(g65328_db) );
na02s01 TIMEBOOST_cell_36354 ( .a(TIMEBOOST_net_10415), .b(g65268_da), .o(n_2005) );
in01s01 g65329_u0 ( .a(FE_OFN653_n_4508), .o(g65329_sb) );
na02s01 g65329_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__Q), .b(g65329_sb), .o(g65329_da) );
na02f02 TIMEBOOST_cell_40229 ( .a(FE_OFN1762_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__Q), .o(TIMEBOOST_net_12353) );
na02s01 TIMEBOOST_cell_31326 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__20__Q), .b(g65353_sb), .o(TIMEBOOST_net_9574) );
in01s01 g65330_u0 ( .a(FE_OFN654_n_4508), .o(g65330_sb) );
na02s01 TIMEBOOST_cell_40256 ( .a(TIMEBOOST_net_12366), .b(n_8232), .o(TIMEBOOST_net_11954) );
na02s01 g65330_u2 ( .a(n_3744), .b(FE_OFN654_n_4508), .o(g65330_db) );
na02s02 TIMEBOOST_cell_16672 ( .a(n_3744), .b(g64863_sb), .o(TIMEBOOST_net_3593) );
in01s01 g65331_u0 ( .a(FE_OFN654_n_4508), .o(g65331_sb) );
na02s01 g65331_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__Q), .b(g65331_sb), .o(g65331_da) );
na02s01 TIMEBOOST_cell_45118 ( .a(TIMEBOOST_net_14797), .b(FE_OFN1135_g64577_p), .o(n_5373) );
na02s02 TIMEBOOST_cell_40768 ( .a(TIMEBOOST_net_12622), .b(g62985_sb), .o(n_5912) );
in01s01 g65332_u0 ( .a(FE_OFN654_n_4508), .o(g65332_sb) );
na02s02 TIMEBOOST_cell_16673 ( .a(TIMEBOOST_net_3593), .b(g64863_db), .o(n_3715) );
na02s01 g65332_u2 ( .a(n_3774), .b(FE_OFN654_n_4508), .o(g65332_db) );
na02s01 TIMEBOOST_cell_16674 ( .a(n_3764), .b(g64959_sb), .o(TIMEBOOST_net_3594) );
in01s01 g65333_u0 ( .a(FE_OFN651_n_4508), .o(g65333_sb) );
na02s01 g65333_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__Q), .b(g65333_sb), .o(g65333_da) );
na02s01 TIMEBOOST_cell_40258 ( .a(TIMEBOOST_net_12367), .b(n_2166), .o(TIMEBOOST_net_11950) );
na02s01 TIMEBOOST_cell_16542 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(g65758_sb), .o(TIMEBOOST_net_3528) );
in01s01 g65334_u0 ( .a(FE_OFN653_n_4508), .o(g65334_sb) );
na02f02 TIMEBOOST_cell_44624 ( .a(TIMEBOOST_net_14550), .b(FE_OFN2180_n_8567), .o(TIMEBOOST_net_13480) );
na02s01 g65334_u2 ( .a(n_3741), .b(FE_OFN653_n_4508), .o(g65334_db) );
na02s01 TIMEBOOST_cell_31019 ( .a(TIMEBOOST_net_9420), .b(g64836_db), .o(n_4445) );
in01s01 g65335_u0 ( .a(FE_OFN653_n_4508), .o(g65335_sb) );
na02s01 TIMEBOOST_cell_16675 ( .a(TIMEBOOST_net_3594), .b(g64959_db), .o(n_3659) );
na02s01 g65335_u2 ( .a(n_3785), .b(FE_OFN653_n_4508), .o(g65335_db) );
na02s01 TIMEBOOST_cell_16676 ( .a(n_3761), .b(g64858_sb), .o(TIMEBOOST_net_3595) );
in01s01 g65336_u0 ( .a(FE_OFN654_n_4508), .o(g65336_sb) );
na02s01 g65336_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__Q), .b(g65336_sb), .o(g65336_da) );
na02s02 TIMEBOOST_cell_31325 ( .a(TIMEBOOST_net_9573), .b(g65397_db), .o(n_3521) );
na02s02 TIMEBOOST_cell_31324 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q), .b(g65397_sb), .o(TIMEBOOST_net_9573) );
in01s01 g65337_u0 ( .a(FE_OFN652_n_4508), .o(g65337_sb) );
na02s01 TIMEBOOST_cell_17854 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__1__Q), .b(g65352_sb), .o(TIMEBOOST_net_4184) );
na02s01 TIMEBOOST_cell_36481 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(g65691_db), .o(TIMEBOOST_net_10479) );
na02s01 TIMEBOOST_cell_36480 ( .a(TIMEBOOST_net_10478), .b(g58017_sb), .o(TIMEBOOST_net_4323) );
in01s01 g65338_u0 ( .a(FE_OFN654_n_4508), .o(g65338_sb) );
na02s01 TIMEBOOST_cell_40260 ( .a(TIMEBOOST_net_12368), .b(n_2183), .o(TIMEBOOST_net_11956) );
na02s01 g65338_u2 ( .a(n_3770), .b(FE_OFN654_n_4508), .o(g65338_db) );
na02s01 TIMEBOOST_cell_38644 ( .a(TIMEBOOST_net_11560), .b(g59111_sb), .o(n_8697) );
in01s01 g65339_u0 ( .a(FE_OFN644_n_4677), .o(g65339_sb) );
na02s03 TIMEBOOST_cell_8918 ( .a(pci_target_unit_del_sync_comp_cycle_count_4_), .b(pci_target_unit_del_sync_comp_cycle_count_7_), .o(TIMEBOOST_net_1026) );
na02s01 g65339_u2 ( .a(n_3792), .b(FE_OFN644_n_4677), .o(g65339_db) );
na02s03 TIMEBOOST_cell_8919 ( .a(TIMEBOOST_net_1026), .b(n_1690), .o(TIMEBOOST_net_182) );
in01s01 g65340_u0 ( .a(FE_OFN651_n_4508), .o(g65340_sb) );
na02s01 TIMEBOOST_cell_42876 ( .a(TIMEBOOST_net_13676), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_11215) );
na02s01 TIMEBOOST_cell_45119 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__Q), .b(n_3524), .o(TIMEBOOST_net_14798) );
na02s02 TIMEBOOST_cell_40770 ( .a(TIMEBOOST_net_12623), .b(g62378_sb), .o(n_6847) );
in01s01 g65341_u0 ( .a(FE_OFN651_n_4508), .o(g65341_sb) );
na02s01 g65341_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__Q), .b(g65341_sb), .o(g65341_da) );
na02s01 TIMEBOOST_cell_45120 ( .a(TIMEBOOST_net_14798), .b(FE_OFN1128_g64577_p), .o(TIMEBOOST_net_11394) );
na02s02 TIMEBOOST_cell_40772 ( .a(TIMEBOOST_net_12624), .b(g62688_sb), .o(n_6166) );
in01s01 g65342_u0 ( .a(FE_OFN652_n_4508), .o(g65342_sb) );
na02s01 TIMEBOOST_cell_16677 ( .a(TIMEBOOST_net_3595), .b(g64858_db), .o(n_3718) );
na02s01 g65342_u2 ( .a(n_3764), .b(FE_OFN652_n_4508), .o(g65342_db) );
na03s02 TIMEBOOST_cell_40681 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__Q), .b(n_4359), .c(FE_OFN1208_n_6356), .o(TIMEBOOST_net_12579) );
in01s01 g65343_u0 ( .a(FE_OFN652_n_4508), .o(g65343_sb) );
na02s01 TIMEBOOST_cell_16644 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(g64162_sb), .o(TIMEBOOST_net_3579) );
na02s01 g65343_u2 ( .a(n_3783), .b(FE_OFN652_n_4508), .o(g65343_db) );
na02s01 TIMEBOOST_cell_16645 ( .a(TIMEBOOST_net_3579), .b(g64162_db), .o(n_4003) );
na02s01 TIMEBOOST_cell_40507 ( .a(wishbone_slave_unit_pcim_sm_data_in_643), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__Q), .o(TIMEBOOST_net_12492) );
na02f02 TIMEBOOST_cell_42344 ( .a(TIMEBOOST_net_13410), .b(g57186_sb), .o(TIMEBOOST_net_12328) );
na02f02 TIMEBOOST_cell_44654 ( .a(TIMEBOOST_net_14565), .b(FE_OFN2167_n_8567), .o(TIMEBOOST_net_13487) );
in01s01 g65345_u0 ( .a(FE_OFN1643_n_4671), .o(g65345_sb) );
na02s01 TIMEBOOST_cell_16647 ( .a(TIMEBOOST_net_3580), .b(g64163_db), .o(n_4002) );
na02s01 g65345_u2 ( .a(n_3785), .b(FE_OFN1643_n_4671), .o(g65345_db) );
na02s02 TIMEBOOST_cell_16648 ( .a(n_3780), .b(g64961_sb), .o(TIMEBOOST_net_3581) );
in01s01 g65346_u0 ( .a(FE_OFN640_n_4669), .o(g65346_sb) );
na02s02 TIMEBOOST_cell_16649 ( .a(TIMEBOOST_net_3581), .b(g64961_db), .o(n_3657) );
na02s01 TIMEBOOST_cell_39204 ( .a(TIMEBOOST_net_11840), .b(n_1657), .o(TIMEBOOST_net_11457) );
na02s01 TIMEBOOST_cell_40262 ( .a(TIMEBOOST_net_12369), .b(n_8232), .o(TIMEBOOST_net_11953) );
in01s01 g65347_u0 ( .a(FE_OFN1676_n_4655), .o(g65347_sb) );
na02s01 g65347_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__Q), .b(g65347_sb), .o(g65347_da) );
na02f02 TIMEBOOST_cell_45538 ( .a(TIMEBOOST_net_15007), .b(n_14060), .o(n_16243) );
na02m02 TIMEBOOST_cell_44559 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__15__Q), .b(n_9424), .o(TIMEBOOST_net_14518) );
in01s01 g65348_u0 ( .a(FE_OFN1677_n_4655), .o(g65348_sb) );
na02s01 TIMEBOOST_cell_17452 ( .a(n_4452), .b(FE_OFN642_n_4677), .o(TIMEBOOST_net_3983) );
na02s01 g65348_u2 ( .a(n_3747), .b(FE_OFN1677_n_4655), .o(g65348_db) );
na02s02 TIMEBOOST_cell_17453 ( .a(TIMEBOOST_net_3983), .b(g65407_da), .o(n_4232) );
in01s01 g65349_u0 ( .a(FE_OFN1679_n_4655), .o(g65349_sb) );
na02s01 TIMEBOOST_cell_17454 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(g64079_sb), .o(TIMEBOOST_net_3984) );
na02s01 g65349_u2 ( .a(n_3777), .b(FE_OFN1679_n_4655), .o(g65349_db) );
na02s01 TIMEBOOST_cell_44992 ( .a(TIMEBOOST_net_14734), .b(g63602_db), .o(TIMEBOOST_net_13156) );
in01s01 g65350_u0 ( .a(FE_OFN1680_n_4655), .o(g65350_sb) );
na02s01 g65350_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__Q), .b(g65350_sb), .o(g65350_da) );
na02f02 TIMEBOOST_cell_40231 ( .a(FE_OFN1554_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__22__Q), .o(TIMEBOOST_net_12354) );
na02s01 TIMEBOOST_cell_40264 ( .a(TIMEBOOST_net_12370), .b(n_2163), .o(TIMEBOOST_net_11952) );
in01s01 g65351_u0 ( .a(FE_OFN1677_n_4655), .o(g65351_sb) );
na02s01 TIMEBOOST_cell_16930 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__Q), .b(g65276_sb), .o(TIMEBOOST_net_3722) );
na02s01 g65351_u2 ( .a(n_4473), .b(FE_OFN1677_n_4655), .o(g65351_db) );
na02s01 TIMEBOOST_cell_16931 ( .a(TIMEBOOST_net_3722), .b(g65276_db), .o(n_3587) );
in01s01 g65352_u0 ( .a(FE_OFN1677_n_4655), .o(g65352_sb) );
na02s01 TIMEBOOST_cell_16932 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__Q), .b(g65368_sb), .o(TIMEBOOST_net_3723) );
na02s01 g65352_u2 ( .a(n_3774), .b(FE_OFN1677_n_4655), .o(g65352_db) );
na02s01 TIMEBOOST_cell_16933 ( .a(TIMEBOOST_net_3723), .b(g65368_db), .o(n_3533) );
in01s01 g65353_u0 ( .a(FE_OFN1677_n_4655), .o(g65353_sb) );
na02s01 TIMEBOOST_cell_17456 ( .a(pci_target_unit_fifos_pciw_addr_data_in_128), .b(g64090_sb), .o(TIMEBOOST_net_3985) );
na02s01 g65353_u2 ( .a(n_3752), .b(FE_OFN1677_n_4655), .o(g65353_db) );
na03s02 TIMEBOOST_cell_38603 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__Q), .b(n_4237), .c(FE_OFN1212_n_4151), .o(TIMEBOOST_net_11540) );
in01s01 g65354_u0 ( .a(FE_OFN1679_n_4655), .o(g65354_sb) );
na02s01 TIMEBOOST_cell_17458 ( .a(n_3774), .b(FE_OFN643_n_4677), .o(TIMEBOOST_net_3986) );
na02s01 g65354_u2 ( .a(n_3741), .b(FE_OFN1679_n_4655), .o(g65354_db) );
na02s01 TIMEBOOST_cell_17459 ( .a(TIMEBOOST_net_3986), .b(g65281_da), .o(n_3584) );
in01s01 g65355_u0 ( .a(FE_OFN1676_n_4655), .o(g65355_sb) );
na02s01 TIMEBOOST_cell_17460 ( .a(n_4645), .b(FE_OFN644_n_4677), .o(TIMEBOOST_net_3987) );
na02s01 g65355_u2 ( .a(n_4444), .b(FE_OFN1676_n_4655), .o(g65355_db) );
na02s02 TIMEBOOST_cell_17461 ( .a(TIMEBOOST_net_3987), .b(g65293_da), .o(n_4282) );
in01s01 g65356_u0 ( .a(FE_OFN1680_n_4655), .o(g65356_sb) );
na02s02 TIMEBOOST_cell_17462 ( .a(n_4442), .b(FE_OFN642_n_4677), .o(TIMEBOOST_net_3988) );
na02s01 g65356_u2 ( .a(n_3785), .b(FE_OFN1680_n_4655), .o(g65356_db) );
na02s02 TIMEBOOST_cell_17463 ( .a(TIMEBOOST_net_3988), .b(g65372_da), .o(n_4250) );
in01s01 g65357_u0 ( .a(FE_OFN1678_n_4655), .o(g65357_sb) );
na02s01 TIMEBOOST_cell_17464 ( .a(n_4447), .b(FE_OFN643_n_4677), .o(TIMEBOOST_net_3989) );
na02s01 TIMEBOOST_cell_17896 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__Q), .b(g61943_sb), .o(TIMEBOOST_net_4205) );
na02s01 TIMEBOOST_cell_17465 ( .a(TIMEBOOST_net_3989), .b(g65273_da), .o(n_4291) );
in01s01 g65358_u0 ( .a(FE_OFN1680_n_4655), .o(g65358_sb) );
na02s02 g65358_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__Q), .b(g65358_sb), .o(g65358_da) );
na02s01 TIMEBOOST_cell_40266 ( .a(TIMEBOOST_net_12371), .b(n_8069), .o(TIMEBOOST_net_11955) );
na02m02 TIMEBOOST_cell_40268 ( .a(TIMEBOOST_net_12372), .b(wbu_addr_in_272), .o(n_9880) );
in01s01 g65359_u0 ( .a(FE_OFN1676_n_4655), .o(g65359_sb) );
na03s02 TIMEBOOST_cell_38365 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__Q), .b(FE_OFN1134_g64577_p), .c(n_3871), .o(TIMEBOOST_net_11421) );
na02s01 TIMEBOOST_cell_16894 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__Q), .b(g64317_sb), .o(TIMEBOOST_net_3704) );
na02m02 TIMEBOOST_cell_36668 ( .a(TIMEBOOST_net_10572), .b(g52645_db), .o(n_14744) );
in01s01 g65360_u0 ( .a(FE_OFN1678_n_4655), .o(g65360_sb) );
na02m02 TIMEBOOST_cell_38774 ( .a(TIMEBOOST_net_11625), .b(g53906_sb), .o(n_13535) );
na02s01 g65360_u2 ( .a(n_3739), .b(FE_OFN1678_n_4655), .o(g65360_db) );
na02s01 TIMEBOOST_cell_40270 ( .a(TIMEBOOST_net_12373), .b(n_1708), .o(TIMEBOOST_net_11992) );
in01s01 g65361_u0 ( .a(FE_OFN1676_n_4655), .o(g65361_sb) );
na02s01 TIMEBOOST_cell_40265 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__Q), .b(n_2168), .o(TIMEBOOST_net_12371) );
na02s01 g65361_u2 ( .a(n_4498), .b(FE_OFN1676_n_4655), .o(g65361_db) );
na02s01 TIMEBOOST_cell_39530 ( .a(TIMEBOOST_net_12003), .b(g61715_sb), .o(n_8395) );
in01s01 g65362_u0 ( .a(FE_OFN1677_n_4655), .o(g65362_sb) );
na02s02 TIMEBOOST_cell_43512 ( .a(TIMEBOOST_net_13994), .b(FE_OFN1231_n_6391), .o(TIMEBOOST_net_12629) );
na02s01 g65362_u2 ( .a(n_3755), .b(FE_OFN1677_n_4655), .o(g65362_db) );
na02s01 TIMEBOOST_cell_42591 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__Q), .b(FE_OFN597_n_9694), .o(TIMEBOOST_net_13534) );
in01s01 g65363_u0 ( .a(FE_OFN1676_n_4655), .o(g65363_sb) );
na02m02 TIMEBOOST_cell_39513 ( .a(g54178_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_398), .o(TIMEBOOST_net_11995) );
na02s01 g65363_u2 ( .a(n_3764), .b(FE_OFN1676_n_4655), .o(g65363_db) );
na02m02 TIMEBOOST_cell_39514 ( .a(TIMEBOOST_net_11995), .b(g54178_db), .o(n_13214) );
in01s01 g65364_u0 ( .a(FE_OFN1676_n_4655), .o(g65364_sb) );
na02s01 TIMEBOOST_cell_39515 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__Q), .b(g58419_sb), .o(TIMEBOOST_net_11996) );
na02s01 g65364_u2 ( .a(n_4465), .b(FE_OFN1676_n_4655), .o(g65364_db) );
na02s01 TIMEBOOST_cell_39516 ( .a(TIMEBOOST_net_11996), .b(g58419_db), .o(n_9430) );
in01s01 g65365_u0 ( .a(FE_OFN1676_n_4655), .o(g65365_sb) );
na02s01 TIMEBOOST_cell_39517 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__8__Q), .b(g58452_sb), .o(TIMEBOOST_net_11997) );
na02s01 g65365_u2 ( .a(n_3783), .b(FE_OFN1676_n_4655), .o(g65365_db) );
na02s01 TIMEBOOST_cell_39500 ( .a(TIMEBOOST_net_11988), .b(g62803_sb), .o(n_5376) );
in01s01 g65366_u0 ( .a(FE_OFN1643_n_4671), .o(g65366_sb) );
na02s01 TIMEBOOST_cell_40263 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__Q), .b(n_8119), .o(TIMEBOOST_net_12370) );
na02s01 g65366_u2 ( .a(n_4452), .b(FE_OFN1643_n_4671), .o(g65366_db) );
na02s02 TIMEBOOST_cell_40272 ( .a(TIMEBOOST_net_12374), .b(g65047_sb), .o(n_3621) );
in01s01 g65367_u0 ( .a(FE_OFN1642_n_4671), .o(g65367_sb) );
na02m02 TIMEBOOST_cell_44625 ( .a(n_9426), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__Q), .o(TIMEBOOST_net_14551) );
na02s01 g65367_u2 ( .a(n_4473), .b(FE_OFN1642_n_4671), .o(g65367_db) );
na02m02 TIMEBOOST_cell_44153 ( .a(n_9096), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__Q), .o(TIMEBOOST_net_14315) );
in01s01 g65368_u0 ( .a(FE_OFN644_n_4677), .o(g65368_sb) );
na02s01 TIMEBOOST_cell_16934 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__Q), .b(g65871_sb), .o(TIMEBOOST_net_3724) );
na02s01 g65368_u2 ( .a(n_3749), .b(FE_OFN644_n_4677), .o(g65368_db) );
na02s01 TIMEBOOST_cell_16935 ( .a(TIMEBOOST_net_3724), .b(g65871_db), .o(n_1871) );
in01s01 g65369_u0 ( .a(FE_OFN1640_n_4671), .o(g65369_sb) );
na02s01 g65369_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__Q), .b(g65369_sb), .o(g65369_da) );
na02s02 TIMEBOOST_cell_40774 ( .a(TIMEBOOST_net_12625), .b(g62495_sb), .o(n_6594) );
in01s01 g65370_u0 ( .a(FE_OFN1644_n_4671), .o(g65370_sb) );
na02s01 g65370_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__Q), .b(g65370_sb), .o(g65370_da) );
na02s02 TIMEBOOST_cell_31321 ( .a(TIMEBOOST_net_9571), .b(g65385_db), .o(n_3525) );
na02s02 TIMEBOOST_cell_31320 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__22__Q), .b(g65385_sb), .o(TIMEBOOST_net_9571) );
na02s01 g65371_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__Q), .b(g65325_sb), .o(g65371_da) );
na02s02 TIMEBOOST_cell_17717 ( .a(TIMEBOOST_net_4115), .b(g62058_sb), .o(n_7836) );
na03s01 TIMEBOOST_cell_5987 ( .a(n_1943), .b(g61732_sb), .c(g61732_db), .o(n_8355) );
in01s01 g65372_u0 ( .a(FE_OFN642_n_4677), .o(g65372_sb) );
na02s02 g65372_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__Q), .b(g65372_sb), .o(g65372_da) );
na02s01 TIMEBOOST_cell_16543 ( .a(TIMEBOOST_net_3528), .b(g65758_db), .o(n_2045) );
na02s01 TIMEBOOST_cell_16544 ( .a(pci_target_unit_fifos_pcir_data_in_175), .b(g65759_sb), .o(TIMEBOOST_net_3529) );
in01s01 g65373_u0 ( .a(n_4669), .o(g65373_sb) );
na02s01 TIMEBOOST_cell_40851 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__Q), .b(n_13544), .o(TIMEBOOST_net_12664) );
na02s01 g65373_u2 ( .a(n_3749), .b(n_4669), .o(g65373_db) );
na02s02 TIMEBOOST_cell_39468 ( .a(TIMEBOOST_net_11972), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_4629) );
in01s01 g65374_u0 ( .a(FE_OFN640_n_4669), .o(g65374_sb) );
na02f02 TIMEBOOST_cell_44154 ( .a(TIMEBOOST_net_14315), .b(FE_OFN1413_n_8567), .o(TIMEBOOST_net_12866) );
na02s01 TIMEBOOST_cell_17652 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__Q), .b(g65361_sb), .o(TIMEBOOST_net_4083) );
na02s01 TIMEBOOST_cell_40273 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__Q), .b(FE_OFN631_n_4454), .o(TIMEBOOST_net_12375) );
in01s01 g65375_u0 ( .a(FE_OFN653_n_4508), .o(g65375_sb) );
na02s01 g65375_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__Q), .b(g65375_sb), .o(g65375_da) );
na02s01 TIMEBOOST_cell_16545 ( .a(TIMEBOOST_net_3529), .b(g65759_db), .o(n_1920) );
na02s01 TIMEBOOST_cell_42868 ( .a(TIMEBOOST_net_13672), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_11211) );
in01s01 g65376_u0 ( .a(FE_OFN1059_n_4727), .o(g65376_sb) );
na02s01 g65376_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__Q), .b(g65376_sb), .o(g65376_da) );
na02s01 g65376_u2 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(FE_OFN1059_n_4727), .o(g65376_db) );
na02s01 TIMEBOOST_cell_45121 ( .a(n_4007), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q), .o(TIMEBOOST_net_14799) );
in01s01 g65377_u0 ( .a(n_4669), .o(g65377_sb) );
na02s01 g65377_u1 ( .a(n_14), .b(g65377_sb), .o(g65377_da) );
na02s01 g65377_u2 ( .a(n_4672), .b(n_4669), .o(g65377_db) );
na02s02 TIMEBOOST_cell_37844 ( .a(TIMEBOOST_net_11160), .b(g57971_sb), .o(n_9829) );
in01s01 g65378_u0 ( .a(FE_OFN652_n_4508), .o(g65378_sb) );
na02s01 g65378_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__Q), .b(g65378_sb), .o(g65378_da) );
na02s01 TIMEBOOST_cell_40259 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__Q), .b(n_8069), .o(TIMEBOOST_net_12368) );
na02s02 TIMEBOOST_cell_40274 ( .a(TIMEBOOST_net_12375), .b(g64830_sb), .o(TIMEBOOST_net_306) );
in01s01 g65379_u0 ( .a(FE_OFN652_n_4508), .o(g65379_sb) );
na02s01 g65379_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__Q), .b(g65379_sb), .o(g65379_da) );
na02s02 TIMEBOOST_cell_41865 ( .a(TIMEBOOST_net_334), .b(g61918_sb), .o(TIMEBOOST_net_13171) );
na02s01 TIMEBOOST_cell_40275 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__Q), .b(n_8232), .o(TIMEBOOST_net_12376) );
in01s01 g65380_u0 ( .a(FE_OFN1642_n_4671), .o(g65380_sb) );
na02s01 g65380_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__Q), .b(g65380_sb), .o(g65380_da) );
na02s01 TIMEBOOST_cell_45122 ( .a(TIMEBOOST_net_14799), .b(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_11409) );
na02s02 TIMEBOOST_cell_40776 ( .a(TIMEBOOST_net_12626), .b(g62987_sb), .o(n_5908) );
in01s01 g65381_u0 ( .a(FE_OFN1680_n_4655), .o(g65381_sb) );
na02s01 g65381_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__31__Q), .b(g65381_sb), .o(g65381_da) );
na03m02 TIMEBOOST_cell_40267 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_23__Q), .b(n_8884), .c(g58782_sb), .o(TIMEBOOST_net_12372) );
na02s02 TIMEBOOST_cell_45177 ( .a(n_4905), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__Q), .o(TIMEBOOST_net_14827) );
in01s01 g65382_u0 ( .a(FE_OFN1677_n_4655), .o(g65382_sb) );
na02s02 TIMEBOOST_cell_39501 ( .a(n_1284), .b(g63378_db), .o(TIMEBOOST_net_11989) );
na02s01 g65382_u2 ( .a(n_3770), .b(FE_OFN1677_n_4655), .o(g65382_db) );
na02s02 TIMEBOOST_cell_39502 ( .a(TIMEBOOST_net_11989), .b(g63378_sb), .o(n_4138) );
in01s01 g65383_u0 ( .a(FE_OFN1678_n_4655), .o(g65383_sb) );
na02s01 TIMEBOOST_cell_18222 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_402), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_4368) );
na02s01 TIMEBOOST_cell_40276 ( .a(TIMEBOOST_net_12376), .b(n_1573), .o(TIMEBOOST_net_12005) );
na02s01 TIMEBOOST_cell_40277 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__Q), .b(n_8176), .o(TIMEBOOST_net_12377) );
in01s01 g65384_u0 ( .a(FE_OFN1680_n_4655), .o(g65384_sb) );
na02s01 g65384_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__Q), .b(g65384_sb), .o(g65384_da) );
na02s01 TIMEBOOST_cell_40278 ( .a(TIMEBOOST_net_12377), .b(n_2066), .o(TIMEBOOST_net_11999) );
na02s01 TIMEBOOST_cell_16862 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__Q), .b(g64268_sb), .o(TIMEBOOST_net_3688) );
in01s01 g65385_u0 ( .a(FE_OFN1677_n_4655), .o(g65385_sb) );
na03s02 TIMEBOOST_cell_39503 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__Q), .b(FE_OFN1125_g64577_p), .c(n_4521), .o(TIMEBOOST_net_11990) );
na02s01 g65385_u2 ( .a(n_3749), .b(FE_OFN1677_n_4655), .o(g65385_db) );
na02s01 TIMEBOOST_cell_39504 ( .a(TIMEBOOST_net_11990), .b(g62820_sb), .o(n_6115) );
na03f02 TIMEBOOST_cell_5988 ( .a(g63530_db), .b(g63530_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q), .o(n_3429) );
na02s02 TIMEBOOST_cell_42364 ( .a(TIMEBOOST_net_13420), .b(g54365_sb), .o(n_13077) );
na02s02 TIMEBOOST_cell_42114 ( .a(TIMEBOOST_net_13295), .b(FE_OFN1313_n_6624), .o(TIMEBOOST_net_11600) );
in01s01 g65387_u0 ( .a(FE_OFN1677_n_4655), .o(g65387_sb) );
na02s01 g65387_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__Q), .b(g65387_sb), .o(g65387_da) );
na02m02 TIMEBOOST_cell_36670 ( .a(TIMEBOOST_net_10573), .b(FE_OFN1147_n_13249), .o(TIMEBOOST_net_4339) );
na02f02 TIMEBOOST_cell_16864 ( .a(configuration_cache_line_size_reg_2996), .b(FE_OFN1695_n_3368), .o(TIMEBOOST_net_3689) );
in01s01 g65388_u0 ( .a(FE_OFN639_n_4669), .o(g65388_sb) );
na02s04 TIMEBOOST_cell_45811 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_25__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_790), .o(TIMEBOOST_net_15144) );
na03s02 TIMEBOOST_cell_39505 ( .a(n_3851), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__Q), .c(FE_OFN1119_g64577_p), .o(TIMEBOOST_net_11991) );
na02s01 TIMEBOOST_cell_16651 ( .a(TIMEBOOST_net_3582), .b(g64963_db), .o(n_3656) );
in01s01 g65389_u0 ( .a(FE_OFN1677_n_4655), .o(g65389_sb) );
na03s02 TIMEBOOST_cell_39495 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__Q), .b(FE_OFN1125_g64577_p), .c(n_3212), .o(TIMEBOOST_net_11986) );
na02s01 g65389_u2 ( .a(n_4470), .b(FE_OFN1677_n_4655), .o(g65389_db) );
na02s01 TIMEBOOST_cell_39506 ( .a(TIMEBOOST_net_11991), .b(g63120_sb), .o(n_5016) );
in01s01 g65390_u0 ( .a(n_2629), .o(g65390_sb) );
na02s01 g65390_u1 ( .a(n_2675), .b(g65390_sb), .o(g65390_da) );
na02s01 g65390_u2 ( .a(n_16307), .b(n_2629), .o(g65390_db) );
na02s01 g65390_u3 ( .a(g65390_da), .b(g65390_db), .o(n_2630) );
in01s01 g65391_u0 ( .a(FE_OFN642_n_4677), .o(g65391_sb) );
na02s01 TIMEBOOST_cell_36331 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__Q), .b(g65907_db), .o(TIMEBOOST_net_10404) );
na02s01 g65391_u2 ( .a(n_4444), .b(n_4677), .o(g65391_db) );
na02s01 TIMEBOOST_cell_36356 ( .a(TIMEBOOST_net_10416), .b(g66399_sb), .o(n_2522) );
in01s01 g65392_u0 ( .a(FE_OFN1680_n_4655), .o(g65392_sb) );
na02s01 g65392_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__14__Q), .b(g65392_sb), .o(g65392_da) );
na02m02 TIMEBOOST_cell_44207 ( .a(n_9720), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__Q), .o(TIMEBOOST_net_14342) );
na02s01 TIMEBOOST_cell_40279 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__Q), .b(n_8232), .o(TIMEBOOST_net_12378) );
in01s01 g65393_u0 ( .a(FE_OFN640_n_4669), .o(g65393_sb) );
na02s01 TIMEBOOST_cell_16652 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(g64156_sb), .o(TIMEBOOST_net_3583) );
na02s01 g65393_u2 ( .a(n_3752), .b(FE_OFN640_n_4669), .o(g65393_db) );
na02s01 TIMEBOOST_cell_16653 ( .a(TIMEBOOST_net_3583), .b(g64156_db), .o(n_4009) );
in01s01 g65394_u0 ( .a(FE_OFN1677_n_4655), .o(g65394_sb) );
na02s02 TIMEBOOST_cell_43502 ( .a(TIMEBOOST_net_13989), .b(FE_OFN1236_n_6391), .o(TIMEBOOST_net_12620) );
na02s01 g65394_u2 ( .a(n_3744), .b(FE_OFN1677_n_4655), .o(g65394_db) );
na02s01 TIMEBOOST_cell_39508 ( .a(TIMEBOOST_net_11992), .b(g61924_sb), .o(n_7975) );
in01s01 g65395_u0 ( .a(FE_OFN1678_n_4655), .o(g65395_sb) );
na02f02 TIMEBOOST_cell_42214 ( .a(TIMEBOOST_net_13345), .b(FE_OFN1408_n_8567), .o(TIMEBOOST_net_12298) );
na02s01 g65395_u2 ( .a(n_3792), .b(FE_OFN1678_n_4655), .o(g65395_db) );
na02s01 TIMEBOOST_cell_17529 ( .a(TIMEBOOST_net_4021), .b(g65859_sb), .o(n_1580) );
in01s01 g65396_u0 ( .a(FE_OFN1680_n_4655), .o(g65396_sb) );
na02s01 g65396_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__Q), .b(g65396_sb), .o(g65396_da) );
na02s01 TIMEBOOST_cell_40280 ( .a(TIMEBOOST_net_12378), .b(n_2195), .o(TIMEBOOST_net_12003) );
na02s01 TIMEBOOST_cell_42911 ( .a(g58049_sb), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_13694) );
in01s01 g65397_u0 ( .a(FE_OFN1677_n_4655), .o(g65397_sb) );
na02s02 TIMEBOOST_cell_43048 ( .a(TIMEBOOST_net_13762), .b(n_1967), .o(n_8591) );
na02s01 g65397_u2 ( .a(n_3761), .b(FE_OFN1677_n_4655), .o(g65397_db) );
na02s01 TIMEBOOST_cell_38727 ( .a(n_1854), .b(g61870_sb), .o(TIMEBOOST_net_11602) );
in01s01 g65398_u0 ( .a(FE_OFN644_n_4677), .o(g65398_sb) );
na02s01 TIMEBOOST_cell_40282 ( .a(TIMEBOOST_net_12379), .b(n_2202), .o(TIMEBOOST_net_12001) );
na02s01 g65398_u2 ( .a(n_3752), .b(FE_OFN644_n_4677), .o(g65398_db) );
na02s02 TIMEBOOST_cell_8925 ( .a(TIMEBOOST_net_1029), .b(n_236), .o(n_13544) );
in01s01 g65399_u0 ( .a(FE_OFN1643_n_4671), .o(g65399_sb) );
na02s02 TIMEBOOST_cell_17856 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__Q), .b(g65356_sb), .o(TIMEBOOST_net_4185) );
na02s02 TIMEBOOST_cell_31317 ( .a(TIMEBOOST_net_9569), .b(FE_OFN2079_n_8069), .o(TIMEBOOST_net_4150) );
na02s01 TIMEBOOST_cell_31316 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_), .b(n_1117), .o(TIMEBOOST_net_9569) );
in01s01 g65400_u0 ( .a(FE_OFN639_n_4669), .o(g65400_sb) );
na02s02 TIMEBOOST_cell_16654 ( .a(n_3747), .b(g64976_sb), .o(TIMEBOOST_net_3584) );
na02s01 g65400_u2 ( .a(n_4450), .b(FE_OFN639_n_4669), .o(g65400_db) );
na02s01 TIMEBOOST_cell_16662 ( .a(pci_target_unit_fifos_pciw_addr_data_in_124), .b(g64144_sb), .o(TIMEBOOST_net_3588) );
in01s01 g65401_u0 ( .a(FE_OFN1676_n_4655), .o(g65401_sb) );
na02f02 TIMEBOOST_cell_44270 ( .a(TIMEBOOST_net_14373), .b(FE_OFN1403_n_8567), .o(TIMEBOOST_net_12836) );
na02s01 g65401_u2 ( .a(n_3780), .b(FE_OFN1676_n_4655), .o(g65401_db) );
na02s01 TIMEBOOST_cell_41913 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__Q), .b(g58302_sb), .o(TIMEBOOST_net_13195) );
in01s01 g65402_u0 ( .a(FE_OFN1643_n_4671), .o(g65402_sb) );
na02s01 g65402_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__Q), .b(g65402_sb), .o(g65402_da) );
na02s02 TIMEBOOST_cell_31315 ( .a(TIMEBOOST_net_9568), .b(n_8892), .o(n_9435) );
na02m02 TIMEBOOST_cell_41651 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_24__Q), .b(FE_OFN227_n_9841), .o(TIMEBOOST_net_13064) );
in01s01 g65403_u0 ( .a(FE_OFN1642_n_4671), .o(g65403_sb) );
na02s02 g65403_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__Q), .b(g65403_sb), .o(g65403_da) );
na02s01 TIMEBOOST_cell_40284 ( .a(TIMEBOOST_net_12380), .b(n_2191), .o(TIMEBOOST_net_12002) );
na02f08 TIMEBOOST_cell_36268 ( .a(TIMEBOOST_net_10372), .b(n_16936), .o(n_2687) );
in01s01 g65404_u0 ( .a(FE_OFN636_n_4669), .o(g65404_sb) );
na02s02 TIMEBOOST_cell_16655 ( .a(TIMEBOOST_net_3584), .b(g64976_db), .o(n_3651) );
na02s01 g65404_u2 ( .a(n_4465), .b(FE_OFN636_n_4669), .o(g65404_db) );
na02s01 TIMEBOOST_cell_16663 ( .a(TIMEBOOST_net_3588), .b(g64144_db), .o(n_4020) );
in01s01 g65405_u0 ( .a(FE_OFN636_n_4669), .o(g65405_sb) );
na02s01 TIMEBOOST_cell_40295 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__Q), .b(FE_OFN562_n_9895), .o(TIMEBOOST_net_12386) );
na02s02 TIMEBOOST_cell_17654 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__Q), .b(g65364_sb), .o(TIMEBOOST_net_4084) );
na02s01 TIMEBOOST_cell_40286 ( .a(TIMEBOOST_net_12381), .b(n_2058), .o(TIMEBOOST_net_12006) );
in01s01 g65406_u0 ( .a(FE_OFN1643_n_4671), .o(g65406_sb) );
na02s01 TIMEBOOST_cell_38651 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__Q), .b(n_8119), .o(TIMEBOOST_net_11564) );
na02m02 TIMEBOOST_cell_31312 ( .a(configuration_pci_err_data_515), .b(n_2809), .o(TIMEBOOST_net_9567) );
na04f04 TIMEBOOST_cell_36236 ( .a(n_12863), .b(n_13117), .c(n_12778), .d(n_12864), .o(n_13318) );
in01s01 g65407_u0 ( .a(FE_OFN642_n_4677), .o(g65407_sb) );
na02s01 g65407_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__Q), .b(g65407_sb), .o(g65407_da) );
na02s01 TIMEBOOST_cell_31310 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__Q), .b(FE_OFN205_n_9140), .o(TIMEBOOST_net_9566) );
na02s02 TIMEBOOST_cell_43453 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__Q), .b(n_3760), .o(TIMEBOOST_net_13965) );
in01s01 g65408_u0 ( .a(FE_OFN651_n_4508), .o(g65408_sb) );
na02s01 g65408_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__Q), .b(g65408_sb), .o(g65408_da) );
na02s02 TIMEBOOST_cell_37922 ( .a(TIMEBOOST_net_11199), .b(g58046_sb), .o(n_9728) );
in01s01 g65409_u0 ( .a(FE_OFN1642_n_4671), .o(g65409_sb) );
na02s01 TIMEBOOST_cell_40363 ( .a(n_1956), .b(g61735_sb), .o(TIMEBOOST_net_12420) );
na02s02 TIMEBOOST_cell_43454 ( .a(TIMEBOOST_net_13965), .b(FE_OFN1234_n_6391), .o(TIMEBOOST_net_12192) );
na02s01 TIMEBOOST_cell_36238 ( .a(TIMEBOOST_net_10357), .b(pci_target_unit_del_sync_comp_cycle_count_2_), .o(TIMEBOOST_net_34) );
in01s01 g65410_u0 ( .a(FE_OFN643_n_4677), .o(g65410_sb) );
na02s01 TIMEBOOST_cell_40288 ( .a(TIMEBOOST_net_12382), .b(n_2188), .o(TIMEBOOST_net_12000) );
na02s01 g65410_u2 ( .a(n_3761), .b(FE_OFN643_n_4677), .o(g65410_db) );
na02s02 TIMEBOOST_cell_8927 ( .a(TIMEBOOST_net_1030), .b(n_398), .o(n_13541) );
na02s01 g65411_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__Q), .b(g65286_sb), .o(g65411_da) );
na02m02 TIMEBOOST_cell_42345 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__Q), .b(n_9438), .o(TIMEBOOST_net_13411) );
na02s01 TIMEBOOST_cell_40290 ( .a(TIMEBOOST_net_12383), .b(n_2208), .o(TIMEBOOST_net_12004) );
in01s01 g65412_u0 ( .a(FE_OFN639_n_4669), .o(g65412_sb) );
na02s01 TIMEBOOST_cell_40287 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__Q), .b(n_8407), .o(TIMEBOOST_net_12382) );
na02s01 g65412_u2 ( .a(n_4645), .b(FE_OFN639_n_4669), .o(g65412_db) );
na02s01 TIMEBOOST_cell_40292 ( .a(TIMEBOOST_net_12384), .b(n_2197), .o(TIMEBOOST_net_12007) );
in01s01 g65413_u0 ( .a(FE_OFN1640_n_4671), .o(g65413_sb) );
na02s02 TIMEBOOST_cell_40294 ( .a(TIMEBOOST_net_12385), .b(g64994_sb), .o(n_3644) );
na02s01 g65413_u2 ( .a(n_3792), .b(FE_OFN1640_n_4671), .o(g65413_db) );
na02s01 TIMEBOOST_cell_40293 ( .a(n_3755), .b(g64994_db), .o(TIMEBOOST_net_12385) );
in01s01 g65414_u0 ( .a(FE_OFN651_n_4508), .o(g65414_sb) );
na02s01 g65414_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__Q), .b(g65414_sb), .o(g65414_da) );
na02s01 g65414_u2 ( .a(n_4672), .b(FE_OFN651_n_4508), .o(g65414_db) );
na03s02 TIMEBOOST_cell_38055 ( .a(g64193_da), .b(g64193_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__15__Q), .o(TIMEBOOST_net_11266) );
in01s01 g65415_u0 ( .a(FE_OFN1640_n_4671), .o(g65415_sb) );
na02s01 TIMEBOOST_cell_40296 ( .a(TIMEBOOST_net_12386), .b(g57924_sb), .o(TIMEBOOST_net_352) );
na02s01 g65415_u2 ( .a(n_3749), .b(FE_OFN1640_n_4671), .o(g65415_db) );
na02s01 TIMEBOOST_cell_16686 ( .a(pci_target_unit_fifos_pciw_addr_data_in_130), .b(g64178_sb), .o(TIMEBOOST_net_3600) );
in01s01 g65416_u0 ( .a(FE_OFN1640_n_4671), .o(g65416_sb) );
na02s01 g65416_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__Q), .b(g65416_sb), .o(g65416_da) );
na02s01 TIMEBOOST_cell_31306 ( .a(pci_target_unit_del_sync_addr_in_221), .b(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(TIMEBOOST_net_9564) );
na02f02 TIMEBOOST_cell_44120 ( .a(TIMEBOOST_net_14298), .b(FE_OFN1370_n_8567), .o(TIMEBOOST_net_13385) );
in01s01 g65417_u0 ( .a(FE_OFN654_n_4508), .o(g65417_sb) );
na02s01 TIMEBOOST_cell_16687 ( .a(TIMEBOOST_net_3600), .b(g64178_db), .o(n_3988) );
na02s01 g65417_u2 ( .a(n_3761), .b(FE_OFN654_n_4508), .o(g65417_db) );
na02s01 TIMEBOOST_cell_16688 ( .a(pci_target_unit_fifos_pciw_addr_data_in_139), .b(g64180_sb), .o(TIMEBOOST_net_3601) );
in01s01 g65418_u0 ( .a(FE_OFN638_n_4669), .o(g65418_sb) );
na02s01 TIMEBOOST_cell_16689 ( .a(TIMEBOOST_net_3601), .b(g64180_db), .o(n_3986) );
na02s01 TIMEBOOST_cell_39191 ( .a(TIMEBOOST_net_3333), .b(FE_OFN1003_n_2047), .o(TIMEBOOST_net_11834) );
na02s01 TIMEBOOST_cell_16690 ( .a(pci_target_unit_fifos_pciw_addr_data_in_151), .b(g64181_sb), .o(TIMEBOOST_net_3602) );
na02s01 g65419_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__Q), .b(g65272_sb), .o(g65419_da) );
na02s01 TIMEBOOST_cell_45080 ( .a(TIMEBOOST_net_14778), .b(FE_OFN270_n_9836), .o(TIMEBOOST_net_11172) );
na02s01 TIMEBOOST_cell_22260 ( .a(FE_OFN8_n_11877), .b(g52482_da), .o(TIMEBOOST_net_6387) );
na02s01 g65420_u1 ( .a(n_12), .b(g65377_sb), .o(g65420_da) );
na02s01 g65420_u2 ( .a(n_3792), .b(n_4669), .o(g65420_db) );
na02m02 TIMEBOOST_cell_44499 ( .a(n_9663), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__Q), .o(TIMEBOOST_net_14488) );
in01s01 g65421_u0 ( .a(FE_OFN653_n_4508), .o(g65421_sb) );
na02s01 g65421_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__Q), .b(g65421_sb), .o(g65421_da) );
na02s02 TIMEBOOST_cell_43455 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__Q), .b(n_1860), .o(TIMEBOOST_net_13966) );
na03f02 TIMEBOOST_cell_36214 ( .a(FE_OCP_RBN1973_n_12381), .b(TIMEBOOST_net_10304), .c(FE_OFN1755_n_12681), .o(n_12713) );
in01s01 g65422_u0 ( .a(FE_OFN653_n_4508), .o(g65422_sb) );
na02s01 TIMEBOOST_cell_39257 ( .a(pci_target_unit_fifos_pciw_addr_data_in_150), .b(g64130_sb), .o(TIMEBOOST_net_11867) );
na02s02 TIMEBOOST_cell_31302 ( .a(pci_target_unit_pcit_if_strd_addr_in_711), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_75), .o(TIMEBOOST_net_9562) );
na02f02 TIMEBOOST_cell_44212 ( .a(TIMEBOOST_net_14344), .b(FE_OFN1411_n_8567), .o(TIMEBOOST_net_12991) );
in01s01 g65423_u0 ( .a(FE_OFN644_n_4677), .o(g65423_sb) );
na02s02 TIMEBOOST_cell_43513 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q), .b(n_3521), .o(TIMEBOOST_net_13995) );
na02s01 TIMEBOOST_cell_31300 ( .a(configuration_wb_err_data_593), .b(parchk_pci_ad_out_in_1190), .o(TIMEBOOST_net_9561) );
na02s01 TIMEBOOST_cell_40285 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__Q), .b(n_8069), .o(TIMEBOOST_net_12381) );
in01s01 g65424_u0 ( .a(FE_OFN652_n_4508), .o(g65424_sb) );
na02s01 g65424_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__Q), .b(g65424_sb), .o(g65424_da) );
na03s02 TIMEBOOST_cell_34474 ( .a(wbm_adr_o_23_), .b(FE_OFN1699_n_5751), .c(g62030_sb), .o(TIMEBOOST_net_594) );
in01s01 g65425_u0 ( .a(n_4725), .o(g65425_sb) );
na03s02 TIMEBOOST_cell_39469 ( .a(TIMEBOOST_net_3959), .b(g64342_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__Q), .o(TIMEBOOST_net_11973) );
na02s01 g65425_u2 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(n_4725), .o(g65425_db) );
na02s02 TIMEBOOST_cell_39470 ( .a(TIMEBOOST_net_11973), .b(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_4648) );
in01s01 g65426_u0 ( .a(FE_OFN651_n_4508), .o(g65426_sb) );
na02s01 TIMEBOOST_cell_16691 ( .a(TIMEBOOST_net_3602), .b(g64181_db), .o(n_3985) );
na02s01 g65426_u2 ( .a(n_3749), .b(FE_OFN651_n_4508), .o(g65426_db) );
na02s01 TIMEBOOST_cell_40297 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__Q), .b(FE_OFN554_n_9864), .o(TIMEBOOST_net_12387) );
in01s01 g65427_u0 ( .a(FE_OFN651_n_4508), .o(g65427_sb) );
na02s01 g65427_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__Q), .b(g65427_sb), .o(g65427_da) );
na02s02 TIMEBOOST_cell_40778 ( .a(TIMEBOOST_net_12627), .b(g62339_sb), .o(n_6920) );
in01s01 g65428_u0 ( .a(FE_OFN652_n_4508), .o(g65428_sb) );
na02s01 g65428_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__Q), .b(g65428_sb), .o(g65428_da) );
na02s01 TIMEBOOST_cell_36483 ( .a(TIMEBOOST_net_3322), .b(FE_OFN1003_n_2047), .o(TIMEBOOST_net_10480) );
na02s01 TIMEBOOST_cell_36482 ( .a(TIMEBOOST_net_10479), .b(g65691_sb), .o(n_2048) );
in01s01 g65429_u0 ( .a(FE_OFN654_n_4508), .o(g65429_sb) );
na02s01 g65429_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__Q), .b(g65429_sb), .o(g65429_da) );
na02s01 TIMEBOOST_cell_31298 ( .a(configuration_wb_err_data_572), .b(parchk_pci_ad_out_in_1169), .o(TIMEBOOST_net_9560) );
in01s01 g65430_u0 ( .a(FE_OFN653_n_4508), .o(g65430_sb) );
na02s01 g65430_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__31__Q), .b(g65430_sb), .o(g65430_da) );
na02s01 TIMEBOOST_cell_31296 ( .a(configuration_wb_err_addr_562), .b(conf_wb_err_addr_in_971), .o(TIMEBOOST_net_9559) );
na02s02 TIMEBOOST_cell_43480 ( .a(TIMEBOOST_net_13978), .b(FE_OFN1233_n_6391), .o(TIMEBOOST_net_12188) );
in01s01 g65431_u0 ( .a(FE_OFN1036_n_4732), .o(g65431_sb) );
na02s01 g65431_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__Q), .b(g65431_sb), .o(g65431_da) );
na02s01 g65431_u2 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(FE_OFN1036_n_4732), .o(g65431_db) );
na02s02 TIMEBOOST_cell_38515 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__Q), .b(g58374_sb), .o(TIMEBOOST_net_11496) );
in01s01 g65432_u0 ( .a(FE_OFN1640_n_4671), .o(g65432_sb) );
na02s01 TIMEBOOST_cell_16660 ( .a(pci_target_unit_fifos_pciw_addr_data_in_140), .b(g64198_sb), .o(TIMEBOOST_net_3587) );
na02s01 g65432_u2 ( .a(n_4672), .b(FE_OFN1640_n_4671), .o(g65432_db) );
na02s01 TIMEBOOST_cell_40298 ( .a(TIMEBOOST_net_12387), .b(g57956_sb), .o(TIMEBOOST_net_444) );
in01s01 g65433_u0 ( .a(FE_OFN653_n_4508), .o(g65433_sb) );
na02s01 TIMEBOOST_cell_31050 ( .a(n_4498), .b(g65095_sb), .o(TIMEBOOST_net_9436) );
na02s02 TIMEBOOST_cell_38505 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__Q), .b(g58358_sb), .o(TIMEBOOST_net_11491) );
na02s01 TIMEBOOST_cell_32018 ( .a(configuration_pci_err_data_502), .b(wbm_dat_o_1_), .o(TIMEBOOST_net_9920) );
in01s01 g65434_u0 ( .a(FE_OFN639_n_4669), .o(g65434_sb) );
na02m02 TIMEBOOST_cell_44155 ( .a(n_9567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__Q), .o(TIMEBOOST_net_14316) );
na02s02 TIMEBOOST_cell_36724 ( .a(TIMEBOOST_net_10600), .b(g63596_sb), .o(n_4772) );
na02f02 TIMEBOOST_cell_44156 ( .a(TIMEBOOST_net_14316), .b(FE_OFN1392_n_8567), .o(TIMEBOOST_net_12709) );
in01s01 g65435_u0 ( .a(FE_OFN636_n_4669), .o(g65435_sb) );
na02f02 TIMEBOOST_cell_44626 ( .a(TIMEBOOST_net_14551), .b(FE_OFN2188_n_8567), .o(TIMEBOOST_net_13006) );
na02s01 TIMEBOOST_cell_39509 ( .a(g64354_da), .b(g64354_db), .o(TIMEBOOST_net_11993) );
na02s01 TIMEBOOST_cell_45719 ( .a(TIMEBOOST_net_4795), .b(FE_OFN1200_n_4090), .o(TIMEBOOST_net_15098) );
no02s01 g65436_u0 ( .a(pci_target_unit_wishbone_master_read_count_reg_2__Q), .b(n_987), .o(g65436_p) );
ao12s01 g65436_u1 ( .a(g65436_p), .b(pci_target_unit_wishbone_master_read_count_reg_2__Q), .c(n_987), .o(n_1180) );
no02s01 g65437_u0 ( .a(pci_target_unit_wishbone_master_read_count_0_), .b(n_1999), .o(g65437_p) );
ao12s01 g65437_u1 ( .a(g65437_p), .b(pci_target_unit_wishbone_master_read_count_0_), .c(n_1999), .o(n_3226) );
ao22s01 g65438_u0 ( .a(n_1281), .b(wbm_rty_i), .c(pci_target_unit_wishbone_master_rty_counter_1_), .d(n_705), .o(n_2223) );
no02f04 g65439_u0 ( .a(n_582), .b(n_588), .o(g65439_p) );
ao12f04 g65439_u1 ( .a(g65439_p), .b(n_582), .c(n_588), .o(n_1461) );
in01s01 g65440_u0 ( .a(pci_target_unit_fifos_pciw_control_in), .o(n_3806) );
no02s02 g65484_u0 ( .a(n_2747), .b(pci_target_unit_del_sync_comp_cycle_count_reg_16__Q), .o(n_3795) );
na03s02 TIMEBOOST_cell_38235 ( .a(g64203_da), .b(g64203_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__Q), .o(TIMEBOOST_net_11356) );
na02s01 g65486_u0 ( .a(n_1696), .b(wishbone_slave_unit_pcim_if_del_req_in), .o(g65486_p) );
in01s01 g65486_u1 ( .a(g65486_p), .o(n_1697) );
no02f03 g65487_u0 ( .a(n_1554), .b(n_978), .o(n_13820) );
na02f08 g65488_u0 ( .a(n_1679), .b(wbu_addr_in_253), .o(g65488_p) );
in01f06 g65488_u1 ( .a(g65488_p), .o(n_2013) );
na02m02 g65489_u0 ( .a(n_1331), .b(wbu_am1_in), .o(g65489_p) );
in01m02 g65489_u1 ( .a(g65489_p), .o(n_2699) );
na02m08 g65490_u0 ( .a(n_1413), .b(conf_wb_err_addr_in_945), .o(g65490_p) );
in01m04 g65490_u1 ( .a(g65490_p), .o(n_1669) );
no02f04 g65491_u0 ( .a(n_1371), .b(n_602), .o(g65491_p) );
in01f04 g65491_u1 ( .a(g65491_p), .o(n_2399) );
no02f04 g65492_u0 ( .a(n_1346), .b(n_668), .o(n_2409) );
no02m02 g65493_u0 ( .a(n_3023), .b(n_2803), .o(g65493_p) );
in01m02 g65493_u1 ( .a(g65493_p), .o(n_3163) );
na02m02 g65494_u0 ( .a(n_3386), .b(n_3022), .o(n_4084) );
na02s01 g65495_u0 ( .a(n_1418), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_), .o(g65495_p) );
in01s01 g65495_u1 ( .a(g65495_p), .o(n_1419) );
na02m06 g65497_u0 ( .a(n_1674), .b(wbm_adr_o_4_), .o(g65497_p) );
in01m04 g65497_u1 ( .a(g65497_p), .o(n_2012) );
no02s01 g65498_u0 ( .a(n_1215), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_), .o(g65498_p) );
in01s02 g65498_u1 ( .a(g65498_p), .o(n_1216) );
na02m02 g65499_u0 ( .a(n_15445), .b(configuration_wb_err_addr_558), .o(n_2626) );
na02f02 g65505_u0 ( .a(configuration_wb_err_addr_557), .b(n_15445), .o(n_2625) );
no02s02 g65506_u0 ( .a(wishbone_slave_unit_pci_initiator_if_read_count_2_), .b(n_660), .o(n_1659) );
na02s01 g65507_u0 ( .a(n_3250), .b(pci_target_unit_wishbone_master_read_bound), .o(n_2807) );
no02s01 g65508_u0 ( .a(n_988), .b(n_3250), .o(n_2806) );
in01s01 g65509_u0 ( .a(n_1226), .o(n_1178) );
no02s03 g65510_u0 ( .a(n_1011), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_2_), .o(g65510_p) );
in01s02 g65510_u1 ( .a(g65510_p), .o(n_1226) );
na02s03 g65511_u0 ( .a(n_948), .b(pci_target_unit_del_sync_comp_cycle_count_2_), .o(g65511_p) );
in01s02 g65511_u1 ( .a(g65511_p), .o(n_1438) );
no02m02 g65512_u0 ( .a(pci_target_unit_pci_target_sm_cnf_progress), .b(n_1554), .o(n_14070) );
na02m02 g65513_u0 ( .a(n_1333), .b(wbu_am2_in), .o(g65513_p) );
in01m02 g65513_u1 ( .a(g65513_p), .o(n_2698) );
na02s06 g65514_u0 ( .a(n_947), .b(wishbone_slave_unit_del_sync_comp_cycle_count_2_), .o(g65514_p) );
in01m02 g65514_u1 ( .a(g65514_p), .o(n_1476) );
no02f04 g65515_u0 ( .a(n_1345), .b(n_596), .o(g65515_p) );
in01f02 g65515_u1 ( .a(g65515_p), .o(n_1976) );
na02f02 g65516_u0 ( .a(FE_OFN1695_n_3368), .b(wbu_cache_line_size_in_207), .o(n_2624) );
no02m08 g65517_u0 ( .a(n_3123), .b(parchk_pci_frame_reg_in), .o(g65517_p) );
in01m04 g65517_u1 ( .a(g65517_p), .o(n_2623) );
na02m02 g65518_u0 ( .a(n_2347), .b(n_2556), .o(g65518_p) );
in01s02 g65518_u1 ( .a(g65518_p), .o(n_3027) );
no02f04 g65519_u0 ( .a(n_3026), .b(n_3295), .o(n_4880) );
no02f04 g65520_u0 ( .a(n_3231), .b(n_16791), .o(g65520_p) );
in01f04 g65520_u1 ( .a(g65520_p), .o(n_3290) );
na03s02 TIMEBOOST_cell_39497 ( .a(n_3878), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__12__Q), .c(FE_OFN2106_g64577_p), .o(TIMEBOOST_net_11987) );
no02s01 g65522_u0 ( .a(n_1011), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_3_), .o(g65522_p1) );
no02s01 g65522_u1 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_4_), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_2_), .o(g65522_p2) );
na02s02 g65522_u2 ( .a(g65522_p1), .b(g65522_p2), .o(n_1015) );
na02m04 g65523_u0 ( .a(n_1985), .b(n_1374), .o(g65523_p) );
in01m02 g65523_u1 ( .a(g65523_p), .o(n_2419) );
na02f02 g65524_u0 ( .a(n_16791), .b(pciu_bar0_in_379), .o(n_2621) );
na02f10 g65525_u0 ( .a(n_1027), .b(pci_target_unit_wishbone_master_rty_counter_4_), .o(n_1177) );
no02s02 g65526_u0 ( .a(n_1477), .b(n_1974), .o(n_1975) );
na02s01 g65528_u0 ( .a(n_1999), .b(n_3164), .o(n_3166) );
na02f02 g65529_u0 ( .a(FE_OFN1695_n_3368), .b(wbu_cache_line_size_in_209), .o(n_2620) );
no02s01 g65530_u0 ( .a(n_3223), .b(n_1999), .o(g65530_p) );
in01s01 g65530_u1 ( .a(FE_OFN147_g65530_p), .o(n_3224) );
na02f02 g65531_u0 ( .a(FE_OFN1061_n_16720), .b(pciu_am1_in_518), .o(n_2984) );
no02m02 g65532_u0 ( .a(n_1548), .b(n_1972), .o(n_1973) );
na02f02 g65533_u0 ( .a(n_1391), .b(n_1971), .o(g65533_p) );
in01f02 g65533_u1 ( .a(g65533_p), .o(n_2461) );
no02f02 g65534_u0 ( .a(n_3504), .b(n_3295), .o(n_3505) );
in01s04 g65536_u0 ( .a(n_2218), .o(n_2219) );
na02m02 TIMEBOOST_cell_42215 ( .a(n_9662), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__Q), .o(TIMEBOOST_net_13346) );
na02f01 g65538_u0 ( .a(n_2804), .b(n_2803), .o(n_2805) );
no02m04 g65539_u0 ( .a(n_2750), .b(n_1639), .o(n_2457) );
na02f02 g65540_u0 ( .a(FE_OFN2129_n_16720), .b(pciu_am1_in_534), .o(n_2802) );
na02s02 TIMEBOOST_cell_42967 ( .a(TIMEBOOST_net_9832), .b(g54198_sb), .o(TIMEBOOST_net_13722) );
na02f02 g65543_u0 ( .a(n_1415), .b(n_1679), .o(g65543_p) );
in01f02 g65543_u1 ( .a(g65543_p), .o(n_2256) );
na02f04 g65549_u0 ( .a(n_2225), .b(n_1478), .o(g65549_p) );
in01f04 g65549_u1 ( .a(g65549_p), .o(n_2694) );
na02m02 g65550_u0 ( .a(n_1969), .b(n_1968), .o(g65550_p) );
in01m02 g65550_u1 ( .a(g65550_p), .o(n_1970) );
in01s02 g65551_u0 ( .a(n_2049), .o(n_2406) );
ao12s02 g65552_u0 ( .a(n_692), .b(n_527), .c(n_1624), .o(n_2049) );
no02f02 g65555_u0 ( .a(n_15762), .b(n_3023), .o(g65555_p) );
in01f02 g65555_u1 ( .a(g65555_p), .o(n_3378) );
na02f06 g65556_u0 ( .a(n_1363), .b(n_1369), .o(n_2708) );
no02s02 g65557_u0 ( .a(n_1805), .b(pci_gnt_i), .o(g65557_p) );
in01s02 g65557_u1 ( .a(g65557_p), .o(n_3810) );
na02s02 g65558_u0 ( .a(n_3222), .b(n_3221), .o(n_3798) );
no02s01 g65559_u0 ( .a(n_3123), .b(output_backup_devsel_out_reg_Q), .o(g65559_p) );
in01s01 g65559_u1 ( .a(g65559_p), .o(n_2619) );
na02f02 TIMEBOOST_cell_42216 ( .a(TIMEBOOST_net_13346), .b(FE_OFN1399_n_8567), .o(TIMEBOOST_net_12299) );
no02m02 g65561_u0 ( .a(n_3023), .b(n_3022), .o(n_4086) );
na02s02 g65562_u0 ( .a(n_1175), .b(n_1416), .o(g65562_p) );
in01s01 g65562_u1 ( .a(g65562_p), .o(n_1176) );
na02s01 g65563_u0 ( .a(n_1337), .b(n_1038), .o(n_2051) );
na02s01 g65564_u0 ( .a(n_1338), .b(n_1093), .o(n_1967) );
na02f01 g65565_u0 ( .a(FE_OFN1695_n_3368), .b(wbu_cache_line_size_in_206), .o(n_2615) );
no02s02 g65566_u0 ( .a(n_2468), .b(pci_target_unit_del_sync_sync_comp_req_pending), .o(n_2469) );
na02m02 g65567_u0 ( .a(n_1414), .b(n_1413), .o(g65567_p) );
in01m02 g65567_u1 ( .a(g65567_p), .o(n_2260) );
na02m04 g65568_u0 ( .a(n_1965), .b(n_1966), .o(g65568_p) );
in01m04 g65568_u1 ( .a(g65568_p), .o(n_2691) );
na02f02 g65569_u0 ( .a(n_2214), .b(n_2390), .o(g65569_p) );
in01f02 g65569_u1 ( .a(g65569_p), .o(n_4675) );
na02s01 g65570_u0 ( .a(n_15762), .b(n_1471), .o(g65570_p) );
in01s01 g65570_u1 ( .a(g65570_p), .o(n_2065) );
na02f02 g65571_u0 ( .a(n_1412), .b(n_1674), .o(g65571_p) );
in01f02 g65571_u1 ( .a(g65571_p), .o(n_2258) );
no02f08 g65572_u0 ( .a(n_1016), .b(n_861), .o(g65572_p1) );
no02f08 g65572_u1 ( .a(n_845), .b(n_872), .o(g65572_p2) );
na02f08 g65572_u2 ( .a(g65572_p1), .b(g65572_p2), .o(n_4686) );
no02f04 TIMEBOOST_cell_44766 ( .a(TIMEBOOST_net_14621), .b(n_300), .o(TIMEBOOST_net_13519) );
in01s01 g65573_u1 ( .a(g65573_p), .o(n_2801) );
no02s01 g65574_u0 ( .a(n_3123), .b(n_205), .o(n_2799) );
in01f06 g65576_u0 ( .a(FE_OFN2121_n_2687), .o(n_1964) );
na02s01 TIMEBOOST_cell_31294 ( .a(configuration_wb_err_addr_535), .b(conf_wb_err_addr_in_944), .o(TIMEBOOST_net_9558) );
na02s01 TIMEBOOST_cell_39327 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__Q), .b(g58332_sb), .o(TIMEBOOST_net_11902) );
na02m01 g65579_u0 ( .a(n_2001), .b(pci_target_unit_wishbone_master_rty_counter_6_), .o(n_2002) );
na02s02 g65580_u0 ( .a(n_1985), .b(n_1986), .o(n_1987) );
na02m02 TIMEBOOST_cell_44319 ( .a(n_9710), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__Q), .o(TIMEBOOST_net_14398) );
no02f04 g65582_u0 ( .a(n_1819), .b(n_15210), .o(n_3115) );
na02m01 g65583_u0 ( .a(n_15407), .b(pci_target_unit_pci_target_sm_rd_progress), .o(g65583_p) );
in01s02 g65583_u1 ( .a(g65583_p), .o(n_13745) );
na02m02 TIMEBOOST_cell_42217 ( .a(n_9871), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__Q), .o(TIMEBOOST_net_13347) );
no02s01 g65585_u0 ( .a(n_3020), .b(n_1133), .o(n_3021) );
na02f02 g65586_u0 ( .a(n_16810), .b(n_14913), .o(n_2614) );
na02f02 g65587_u0 ( .a(FE_OFN1061_n_16720), .b(pciu_am1_in_520), .o(n_2797) );
na02f04 g65588_u0 ( .a(n_3018), .b(n_3019), .o(g65588_p) );
in01f04 g65588_u1 ( .a(g65588_p), .o(n_5230) );
no02s01 g65589_u0 ( .a(n_1696), .b(wishbone_slave_unit_del_sync_sync_comp_req_pending), .o(n_1635) );
na02m02 g65590_u0 ( .a(n_2392), .b(n_3107), .o(g65590_p) );
in01m02 g65590_u1 ( .a(g65590_p), .o(n_7110) );
in01s06 g65592_u0 ( .a(n_4512), .o(n_4904) );
no02s02 g65595_u0 ( .a(n_3001), .b(n_2685), .o(g65595_p) );
in01s04 g65595_u1 ( .a(g65595_p), .o(n_4512) );
na02s01 TIMEBOOST_cell_40300 ( .a(TIMEBOOST_net_12388), .b(g64296_db), .o(n_3878) );
na02s01 g65597_u0 ( .a(n_1329), .b(n_1283), .o(n_2057) );
in01s01 g65598_u0 ( .a(n_1632), .o(n_1633) );
no02s02 g65599_u0 ( .a(n_1425), .b(n_878), .o(n_1632) );
in01s01 g65600_u0 ( .a(n_1630), .o(n_1631) );
no02s02 g65601_u0 ( .a(n_1426), .b(n_883), .o(n_1630) );
na02s01 TIMEBOOST_cell_42650 ( .a(TIMEBOOST_net_13563), .b(g64102_da), .o(TIMEBOOST_net_11276) );
ao12s02 g65603_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_reg_16__Q), .b(n_1126), .c(pci_target_unit_pci_target_if_same_read_reg), .o(n_1961) );
na02s02 TIMEBOOST_cell_45699 ( .a(n_4371), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__Q), .o(TIMEBOOST_net_15088) );
oa12s01 g65605_u0 ( .a(n_2779), .b(pci_target_unit_del_sync_addr_in_204), .c(n_2301), .o(n_2794) );
oa12s01 g65606_u0 ( .a(g74689_p), .b(n_1698), .c(FE_OFN2214_n_15366), .o(n_2793) );
na04f04 TIMEBOOST_cell_36221 ( .a(n_16617), .b(n_16616), .c(n_13923), .d(n_13846), .o(n_14577) );
na02s01 TIMEBOOST_cell_38526 ( .a(TIMEBOOST_net_11501), .b(g62048_sb), .o(n_7762) );
oa12s01 g65609_u0 ( .a(n_2612), .b(pci_target_unit_del_sync_addr_in_212), .c(n_2301), .o(n_2613) );
na02f02 TIMEBOOST_cell_21979 ( .a(TIMEBOOST_net_6246), .b(n_13901), .o(TIMEBOOST_net_3017) );
oa12s01 g65611_u0 ( .a(n_2610), .b(pci_target_unit_del_sync_addr_in_211), .c(n_2301), .o(n_2611) );
oa12s01 g65612_u0 ( .a(n_2790), .b(pci_target_unit_del_sync_addr_in_205), .c(n_2301), .o(n_2792) );
oa12s01 g65613_u0 ( .a(n_2788), .b(pci_target_unit_del_sync_addr_in_206), .c(n_2301), .o(n_2789) );
na02m02 g65614_u0 ( .a(n_3107), .b(n_2609), .o(g65614_p) );
in01m02 g65614_u1 ( .a(g65614_p), .o(n_3089) );
oa12s01 g65615_u0 ( .a(n_2783), .b(pci_target_unit_del_sync_addr_in_209), .c(n_2301), .o(n_2787) );
oa12s01 g65616_u0 ( .a(n_2790), .b(n_2742), .c(n_2301), .o(n_4214) );
na02s02 g65617_u0 ( .a(n_3108), .b(n_3107), .o(g65617_p) );
in01s02 g65617_u1 ( .a(g65617_p), .o(n_7108) );
na02s01 g65618_u0 ( .a(n_2361), .b(n_3217), .o(n_3220) );
na02s01 g65619_u0 ( .a(n_2356), .b(n_2610), .o(n_2786) );
na02s01 g65620_u0 ( .a(n_2366), .b(n_2612), .o(n_2785) );
na02s01 g65621_u0 ( .a(n_2363), .b(n_2783), .o(n_2784) );
na02s01 g65622_u0 ( .a(n_2362), .b(n_2604), .o(n_2782) );
na02s01 g65623_u0 ( .a(n_2364), .b(n_2732), .o(n_2781) );
no02f04 g65626_u0 ( .a(n_2345), .b(n_15805), .o(g65626_p) );
in01f04 g65626_u1 ( .a(g65626_p), .o(n_3314) );
oa12s01 g65627_u0 ( .a(n_2779), .b(n_16027), .c(n_2301), .o(n_2780) );
na02s01 g65628_u0 ( .a(n_2349), .b(n_2606), .o(n_2745) );
oa12s01 g65629_u0 ( .a(n_3217), .b(n_1724), .c(FE_OFN2093_n_2301), .o(n_3219) );
ao12s01 g65630_u0 ( .a(wbs_bte_i_0_), .b(n_1666), .c(wbs_bte_i_1_), .o(n_1667) );
oa12s01 g65631_u0 ( .a(n_2606), .b(pci_target_unit_del_sync_addr_in_210), .c(n_2301), .o(n_2608) );
na02s01 g65632_u0 ( .a(n_2767), .b(n_2788), .o(n_3216) );
ao12m02 g65633_u0 ( .a(n_1134), .b(n_1628), .c(pci_target_unit_pci_target_sm_n_3), .o(n_1629) );
oa12s01 g65634_u0 ( .a(n_2604), .b(pci_target_unit_del_sync_addr_in_208), .c(n_2301), .o(n_2605) );
no02s01 g65635_u0 ( .a(n_249), .b(pci_target_unit_del_sync_req_rty_exp_clr), .o(n_738) );
in01f02 g65636_u0 ( .a(n_2701), .o(n_2387) );
ao12s01 g65639_u0 ( .a(n_3386), .b(n_1322), .c(n_1686), .o(n_3361) );
ao12s01 g65641_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_transfer), .b(n_1436), .c(n_2043), .o(n_2726) );
ao12f02 g65642_u0 ( .a(n_2430), .b(wishbone_slave_unit_pcim_sm_be_in_558), .c(wishbone_slave_unit_pcim_sm_be_in_559), .o(n_1626) );
na02m06 g65643_u0 ( .a(n_2777), .b(n_2778), .o(n_3261) );
oa12s01 g65644_u0 ( .a(n_2601), .b(pci_target_unit_del_sync_addr_in), .c(n_2301), .o(n_2603) );
na03s02 TIMEBOOST_cell_5972 ( .a(n_4452), .b(g64983_sb), .c(g64983_db), .o(n_4362) );
no02s01 g65646_u0 ( .a(n_1327), .b(wishbone_slave_unit_del_sync_req_rty_exp_clr), .o(n_2386) );
oa12s01 g65647_u0 ( .a(n_2601), .b(n_16390), .c(n_2301), .o(n_2602) );
oa12s01 g65648_u0 ( .a(n_2732), .b(pci_target_unit_del_sync_addr_in_207), .c(n_2301), .o(n_2734) );
ao12s01 g65649_u0 ( .a(n_15371), .b(n_1524), .c(n_1326), .o(n_2446) );
ao12s01 g65650_u0 ( .a(n_434), .b(n_802), .c(n_1624), .o(n_1625) );
ao22f02 g65651_u0 ( .a(n_15755), .b(n_1332), .c(n_16001), .d(wbu_am2_in), .o(n_3016) );
oa12s01 g65652_u0 ( .a(n_1453), .b(n_3415), .c(n_1316), .o(n_1623) );
oa12s01 g65653_u0 ( .a(n_1265), .b(n_8876), .c(n_1174), .o(n_1621) );
in01m02 g65654_u0 ( .a(n_1443), .o(n_1619) );
na02f02 TIMEBOOST_cell_42218 ( .a(TIMEBOOST_net_13347), .b(FE_OFN1399_n_8567), .o(TIMEBOOST_net_12300) );
ao22f01 g65658_u0 ( .a(n_2560), .b(n_14908), .c(n_15065), .d(n_1330), .o(n_2972) );
in01s01 g65661_u0 ( .a(n_2730), .o(n_2776) );
ao22s01 g65662_u0 ( .a(n_2671), .b(n_2599), .c(n_2597), .d(parchk_pci_ad_reg_in), .o(n_2730) );
na02f02 TIMEBOOST_cell_44190 ( .a(TIMEBOOST_net_14333), .b(FE_OFN1413_n_8567), .o(TIMEBOOST_net_12745) );
in01s01 g65664_u0 ( .a(n_2600), .o(n_2973) );
ao22s01 g65665_u0 ( .a(n_2599), .b(n_2598), .c(n_2597), .d(parchk_pci_ad_reg_in_1205), .o(n_2600) );
na02m02 TIMEBOOST_cell_43538 ( .a(TIMEBOOST_net_14007), .b(FE_OFN1322_n_6436), .o(TIMEBOOST_net_12241) );
na02f02 TIMEBOOST_cell_44667 ( .a(n_9227), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__Q), .o(TIMEBOOST_net_14572) );
in01s01 g65668_u0 ( .a(FE_OFN672_n_4505), .o(g65668_sb) );
na02s02 TIMEBOOST_cell_40572 ( .a(TIMEBOOST_net_12524), .b(g62552_sb), .o(n_6461) );
na02s01 g65668_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__Q), .b(FE_OFN672_n_4505), .o(g65668_db) );
na02s01 TIMEBOOST_cell_44993 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__Q), .b(g64244_sb), .o(TIMEBOOST_net_14735) );
in01s01 g65669_u0 ( .a(FE_OFN1626_n_4438), .o(g65669_sb) );
na03f02 TIMEBOOST_cell_36184 ( .a(n_12084), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__Q), .c(n_11823), .o(n_12509) );
na02m02 TIMEBOOST_cell_44121 ( .a(n_9410), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__Q), .o(TIMEBOOST_net_14299) );
na02s01 TIMEBOOST_cell_31292 ( .a(configuration_wb_err_cs_bit_569), .b(parchk_pci_cbe_out_in_1203), .o(TIMEBOOST_net_9557) );
in01s01 g65670_u0 ( .a(FE_OFN648_n_4497), .o(g65670_sb) );
na02s01 TIMEBOOST_cell_40302 ( .a(TIMEBOOST_net_12389), .b(g65052_db), .o(n_4321) );
na02s01 g65670_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__Q), .b(FE_OFN648_n_4497), .o(g65670_db) );
na02m02 TIMEBOOST_cell_9063 ( .a(TIMEBOOST_net_1098), .b(n_2494), .o(TIMEBOOST_net_127) );
in01s01 g65671_u0 ( .a(FE_OFN665_n_4495), .o(g65671_sb) );
na02m02 TIMEBOOST_cell_32384 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_26__Q), .o(TIMEBOOST_net_10103) );
na02m02 TIMEBOOST_cell_42219 ( .a(n_2005), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .o(TIMEBOOST_net_13348) );
na02s01 TIMEBOOST_cell_42579 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(g64139_sb), .o(TIMEBOOST_net_13528) );
in01s01 g65672_u0 ( .a(FE_OFN687_n_4417), .o(g65672_sb) );
na03f02 TIMEBOOST_cell_36186 ( .a(n_12090), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__Q), .c(n_11823), .o(n_12515) );
na02s01 g65672_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__Q), .b(FE_OFN687_n_4417), .o(g65672_db) );
na02s01 TIMEBOOST_cell_31290 ( .a(configuration_wb_err_data_571), .b(parchk_pci_ad_out_in_1168), .o(TIMEBOOST_net_9556) );
in01s01 g65673_u0 ( .a(FE_OFN623_n_4409), .o(g65673_sb) );
na02s02 TIMEBOOST_cell_40574 ( .a(TIMEBOOST_net_12525), .b(g62707_sb), .o(n_6152) );
na02s01 g65673_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__Q), .b(FE_OFN623_n_4409), .o(g65673_db) );
na02s01 TIMEBOOST_cell_36485 ( .a(pci_target_unit_del_sync_addr_in_220), .b(g66404_db), .o(TIMEBOOST_net_10481) );
in01s01 g65674_u0 ( .a(FE_OFN938_n_2292), .o(g65674_sb) );
na02f02 TIMEBOOST_cell_42508 ( .a(TIMEBOOST_net_13492), .b(g57225_sb), .o(n_11531) );
na02s01 g65674_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__Q), .b(FE_OFN938_n_2292), .o(g65674_db) );
na03s02 TIMEBOOST_cell_34264 ( .a(TIMEBOOST_net_9791), .b(FE_OFN1168_n_5592), .c(g62100_sb), .o(n_5603) );
in01s01 g65675_u0 ( .a(FE_OFN1003_n_2047), .o(g65675_sb) );
na02s01 TIMEBOOST_cell_44994 ( .a(TIMEBOOST_net_14735), .b(g64244_db), .o(n_3928) );
na02s01 g65675_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__Q), .b(FE_OFN1003_n_2047), .o(g65675_db) );
na02s02 TIMEBOOST_cell_40576 ( .a(TIMEBOOST_net_12526), .b(g62640_sb), .o(n_6268) );
in01s01 g65676_u0 ( .a(FE_OFN952_n_2055), .o(g65676_sb) );
na02s02 TIMEBOOST_cell_45690 ( .a(TIMEBOOST_net_15083), .b(FE_OFN1249_n_4093), .o(TIMEBOOST_net_12559) );
na02s01 g65676_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__Q), .b(FE_OFN952_n_2055), .o(g65676_db) );
na02s01 TIMEBOOST_cell_42859 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__Q), .o(TIMEBOOST_net_13668) );
in01s01 g65677_u0 ( .a(FE_OFN936_n_2292), .o(g65677_sb) );
na03s01 TIMEBOOST_cell_34265 ( .a(TIMEBOOST_net_9790), .b(FE_OFN1163_n_5615), .c(g62104_sb), .o(n_5597) );
na02s01 g65677_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__Q), .b(FE_OFN936_n_2292), .o(g65677_db) );
na02s02 TIMEBOOST_cell_43596 ( .a(TIMEBOOST_net_14036), .b(FE_OFN1315_n_6624), .o(TIMEBOOST_net_12250) );
in01s01 g65678_u0 ( .a(FE_OFN936_n_2292), .o(g65678_sb) );
na02s02 TIMEBOOST_cell_37846 ( .a(TIMEBOOST_net_11161), .b(g58291_sb), .o(n_9513) );
na02s01 g65678_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__Q), .b(FE_OFN936_n_2292), .o(g65678_db) );
na02s02 TIMEBOOST_cell_32003 ( .a(TIMEBOOST_net_9912), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_4894) );
in01s01 g65679_u0 ( .a(FE_OFN1003_n_2047), .o(g65679_sb) );
na02m02 TIMEBOOST_cell_40249 ( .a(n_12179), .b(n_2315), .o(TIMEBOOST_net_12363) );
na02s01 g65679_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__Q), .b(FE_OFN941_n_2047), .o(g65679_db) );
na02s01 TIMEBOOST_cell_40304 ( .a(TIMEBOOST_net_12390), .b(g64890_sb), .o(TIMEBOOST_net_5307) );
in01s01 g65680_u0 ( .a(FE_OFN1074_n_4740), .o(g65680_sb) );
na02s01 TIMEBOOST_cell_40306 ( .a(TIMEBOOST_net_12391), .b(g65095_db), .o(n_4297) );
na02s01 g65680_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__Q), .b(FE_OFN1074_n_4740), .o(g65680_db) );
na02s02 TIMEBOOST_cell_18609 ( .a(TIMEBOOST_net_4561), .b(g62846_sb), .o(n_5279) );
in01s01 g65681_u0 ( .a(FE_OFN1046_n_16657), .o(g65681_sb) );
na02s01 g65681_u1 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(g65681_sb), .o(g65681_da) );
na02s01 g65681_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__Q), .b(FE_OFN1046_n_16657), .o(g65681_db) );
na02s01 TIMEBOOST_cell_38581 ( .a(TIMEBOOST_net_4790), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_11529) );
in01s01 g65682_u0 ( .a(FE_OFN953_n_2055), .o(g65682_sb) );
na03s02 TIMEBOOST_cell_37687 ( .a(n_2017), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__Q), .c(FE_OFN709_n_8232), .o(TIMEBOOST_net_11082) );
na02s01 g65682_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__Q), .b(FE_OFN953_n_2055), .o(g65682_db) );
na02s01 TIMEBOOST_cell_42812 ( .a(TIMEBOOST_net_13644), .b(g62028_sb), .o(n_7840) );
in01s01 g65683_u0 ( .a(FE_OFN2108_n_2047), .o(g65683_sb) );
na02s01 TIMEBOOST_cell_45081 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__Q), .b(FE_OFN579_n_9531), .o(TIMEBOOST_net_14779) );
na02s02 TIMEBOOST_cell_44995 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__Q), .b(g64246_sb), .o(TIMEBOOST_net_14736) );
na02s02 TIMEBOOST_cell_40308 ( .a(TIMEBOOST_net_12392), .b(g64905_db), .o(TIMEBOOST_net_4812) );
in01s01 g65684_u0 ( .a(FE_OFN941_n_2047), .o(g65684_sb) );
na02s01 TIMEBOOST_cell_36484 ( .a(TIMEBOOST_net_10480), .b(g65734_sb), .o(n_1934) );
na02s01 g65684_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__Q), .b(FE_OFN941_n_2047), .o(g65684_db) );
na03s02 TIMEBOOST_cell_40577 ( .a(n_4280), .b(n_4281), .c(FE_OFN1258_n_4143), .o(TIMEBOOST_net_12527) );
in01s01 g65685_u0 ( .a(FE_OFN938_n_2292), .o(g65685_sb) );
na02s01 TIMEBOOST_cell_32002 ( .a(configuration_pci_err_addr_474), .b(wbm_adr_o_4_), .o(TIMEBOOST_net_9912) );
na02s01 g65685_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN938_n_2292), .o(g65685_db) );
na02s02 TIMEBOOST_cell_32001 ( .a(TIMEBOOST_net_9911), .b(FE_OFN1181_n_3476), .o(TIMEBOOST_net_4893) );
in01s01 g65686_u0 ( .a(FE_OFN936_n_2292), .o(g65686_sb) );
na02s02 TIMEBOOST_cell_40398 ( .a(TIMEBOOST_net_12437), .b(g52633_db), .o(n_14674) );
na02s01 g65686_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__Q), .b(FE_OFN936_n_2292), .o(g65686_db) );
na02s02 TIMEBOOST_cell_38090 ( .a(TIMEBOOST_net_11283), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_4646) );
in01s01 g65687_u0 ( .a(FE_OFN936_n_2292), .o(g65687_sb) );
na02s01 TIMEBOOST_cell_15816 ( .a(pci_target_unit_del_sync_comp_cycle_count_14_), .b(pci_target_unit_del_sync_comp_cycle_count_13_), .o(TIMEBOOST_net_3165) );
na02s01 g65687_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__Q), .b(FE_OFN936_n_2292), .o(g65687_db) );
na02s01 TIMEBOOST_cell_15817 ( .a(TIMEBOOST_net_3165), .b(n_1989), .o(TIMEBOOST_net_175) );
in01s01 g65688_u0 ( .a(FE_OFN936_n_2292), .o(g65688_sb) );
na02f02 TIMEBOOST_cell_44200 ( .a(TIMEBOOST_net_14338), .b(FE_OFN1398_n_8567), .o(TIMEBOOST_net_12856) );
na02s01 g65688_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__Q), .b(FE_OFN936_n_2292), .o(g65688_db) );
na02f02 TIMEBOOST_cell_39072 ( .a(TIMEBOOST_net_11774), .b(FE_OFN1769_n_14054), .o(n_14510) );
in01s01 g65689_u0 ( .a(FE_OFN937_n_2292), .o(g65689_sb) );
na03f06 TIMEBOOST_cell_45539 ( .a(n_11792), .b(n_10791), .c(n_11791), .o(TIMEBOOST_net_15008) );
na02s01 g65689_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__Q), .b(FE_OFN937_n_2292), .o(g65689_db) );
na02f02 TIMEBOOST_cell_41236 ( .a(TIMEBOOST_net_12856), .b(g58597_sb), .o(n_9189) );
in01s01 g65690_u0 ( .a(FE_OFN2108_n_2047), .o(g65690_sb) );
na02s01 TIMEBOOST_cell_17002 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(g65783_sb), .o(TIMEBOOST_net_3758) );
na03s02 TIMEBOOST_cell_39493 ( .a(n_3916), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__Q), .c(FE_OFN1119_g64577_p), .o(TIMEBOOST_net_11985) );
na02s01 TIMEBOOST_cell_17003 ( .a(TIMEBOOST_net_3758), .b(g65783_db), .o(n_1599) );
in01s01 g65691_u0 ( .a(FE_OFN1003_n_2047), .o(g65691_sb) );
na02s01 TIMEBOOST_cell_40578 ( .a(TIMEBOOST_net_12527), .b(g62908_sb), .o(n_6061) );
na02s01 g65691_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__Q), .b(FE_OFN1003_n_2047), .o(g65691_db) );
na02s01 TIMEBOOST_cell_44996 ( .a(TIMEBOOST_net_14736), .b(g64246_db), .o(n_3926) );
in01s01 g65692_u0 ( .a(FE_OFN938_n_2292), .o(g65692_sb) );
na02m02 TIMEBOOST_cell_32522 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__Q), .o(TIMEBOOST_net_10172) );
na02s01 g65692_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__Q), .b(FE_OFN938_n_2292), .o(g65692_db) );
na02f02 TIMEBOOST_cell_41162 ( .a(TIMEBOOST_net_12819), .b(g57280_sb), .o(n_11474) );
in01s01 g65693_u0 ( .a(FE_OFN2108_n_2047), .o(g65693_sb) );
na02s01 TIMEBOOST_cell_40291 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__Q), .b(n_8232), .o(TIMEBOOST_net_12384) );
na02s01 g65693_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__Q), .b(FE_OFN2109_n_2047), .o(g65693_db) );
na02s01 TIMEBOOST_cell_40310 ( .a(TIMEBOOST_net_12393), .b(g64803_db), .o(n_4464) );
in01s01 g65694_u0 ( .a(FE_OFN950_n_2055), .o(g65694_sb) );
na02s02 TIMEBOOST_cell_37848 ( .a(TIMEBOOST_net_11162), .b(g57987_sb), .o(n_9810) );
na02s01 g65694_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__Q), .b(FE_OFN950_n_2055), .o(g65694_db) );
na02s02 TIMEBOOST_cell_43069 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__Q), .b(n_4453), .o(TIMEBOOST_net_13773) );
in01s01 g65695_u0 ( .a(FE_OFN938_n_2292), .o(g65695_sb) );
na03s02 TIMEBOOST_cell_7102 ( .a(TIMEBOOST_net_469), .b(g63124_sb), .c(g62724_db), .o(n_5534) );
na02s01 g65695_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__Q), .b(FE_OFN938_n_2292), .o(g65695_db) );
na02s01 TIMEBOOST_cell_42651 ( .a(g64126_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q), .o(TIMEBOOST_net_13564) );
in01s01 g65696_u0 ( .a(FE_OFN951_n_2055), .o(g65696_sb) );
na02m02 TIMEBOOST_cell_43565 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q), .b(n_4425), .o(TIMEBOOST_net_14021) );
na02s02 TIMEBOOST_cell_40580 ( .a(TIMEBOOST_net_12528), .b(g62648_sb), .o(n_6252) );
na02s02 TIMEBOOST_cell_43070 ( .a(TIMEBOOST_net_13773), .b(FE_OFN1212_n_4151), .o(TIMEBOOST_net_12028) );
in01s01 g65697_u0 ( .a(FE_OFN936_n_2292), .o(g65697_sb) );
na02f02 TIMEBOOST_cell_39073 ( .a(TIMEBOOST_net_10135), .b(FE_OFN1769_n_14054), .o(TIMEBOOST_net_11775) );
na02f02 TIMEBOOST_cell_39074 ( .a(TIMEBOOST_net_11775), .b(FE_OFN1773_n_13800), .o(g53289_p) );
in01s01 g65698_u0 ( .a(FE_OFN937_n_2292), .o(g65698_sb) );
na02f04 TIMEBOOST_cell_45540 ( .a(TIMEBOOST_net_15008), .b(n_11130), .o(n_12771) );
na02s01 g65698_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__Q), .b(FE_OFN937_n_2292), .o(g65698_db) );
na03f02 TIMEBOOST_cell_7105 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in), .b(g54330_sb), .c(g54330_db), .o(n_12986) );
in01s01 g65699_u0 ( .a(FE_OFN935_n_2292), .o(g65699_sb) );
na02f02 TIMEBOOST_cell_39075 ( .a(n_13903), .b(TIMEBOOST_net_10122), .o(TIMEBOOST_net_11776) );
na02s01 g65699_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__Q), .b(FE_OFN937_n_2292), .o(g65699_db) );
na02f02 TIMEBOOST_cell_39076 ( .a(TIMEBOOST_net_11776), .b(FE_OFN1596_n_13741), .o(n_14277) );
in01s01 g65700_u0 ( .a(FE_OFN935_n_2292), .o(g65700_sb) );
na02f02 TIMEBOOST_cell_39077 ( .a(FE_OFN1775_n_13800), .b(TIMEBOOST_net_10154), .o(TIMEBOOST_net_11777) );
na02s01 g65700_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__Q), .b(FE_OFN935_n_2292), .o(g65700_db) );
na02f02 TIMEBOOST_cell_39078 ( .a(TIMEBOOST_net_11777), .b(FE_OFN1769_n_14054), .o(g53259_p) );
in01s01 g65701_u0 ( .a(FE_OFN937_n_2292), .o(g65701_sb) );
na02m02 TIMEBOOST_cell_32586 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__Q), .o(TIMEBOOST_net_10204) );
na02s01 g65701_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__Q), .b(FE_OFN937_n_2292), .o(g65701_db) );
na02f02 TIMEBOOST_cell_32585 ( .a(n_12010), .b(TIMEBOOST_net_10203), .o(TIMEBOOST_net_6418) );
in01s01 g65702_u0 ( .a(FE_OFN2108_n_2047), .o(g65702_sb) );
na02s02 TIMEBOOST_cell_17090 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(g65773_sb), .o(TIMEBOOST_net_3802) );
na02s01 g65702_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__Q), .b(FE_OFN2108_n_2047), .o(g65702_db) );
na03m02 TIMEBOOST_cell_39193 ( .a(g58792_sb), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_3__Q), .c(n_8884), .o(TIMEBOOST_net_11835) );
in01s01 g65703_u0 ( .a(FE_OFN937_n_2292), .o(g65703_sb) );
na02m02 TIMEBOOST_cell_32584 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__Q), .o(TIMEBOOST_net_10203) );
na02s01 g65703_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__Q), .b(FE_OFN937_n_2292), .o(g65703_db) );
na02f02 TIMEBOOST_cell_32583 ( .a(n_12010), .b(TIMEBOOST_net_10202), .o(TIMEBOOST_net_6417) );
in01s01 g65704_u0 ( .a(FE_OFN955_n_1699), .o(g65704_sb) );
na02s01 TIMEBOOST_cell_17044 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__Q), .o(TIMEBOOST_net_3779) );
na02s01 g65704_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__Q), .b(FE_OFN955_n_1699), .o(g65704_db) );
na02s01 TIMEBOOST_cell_17045 ( .a(TIMEBOOST_net_3779), .b(FE_OFN1059_n_4727), .o(TIMEBOOST_net_317) );
in01s01 g65705_u0 ( .a(FE_OFN951_n_2055), .o(g65705_sb) );
na02s02 TIMEBOOST_cell_43384 ( .a(TIMEBOOST_net_13930), .b(n_6319), .o(TIMEBOOST_net_12148) );
na02s01 g65705_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__Q), .b(FE_OFN951_n_2055), .o(g65705_db) );
na02s02 TIMEBOOST_cell_37850 ( .a(TIMEBOOST_net_11163), .b(g57978_sb), .o(n_9822) );
in01s01 g65706_u0 ( .a(FE_OFN937_n_2292), .o(g65706_sb) );
na02m02 TIMEBOOST_cell_32582 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__Q), .o(TIMEBOOST_net_10202) );
na02s01 g65706_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__Q), .b(FE_OFN938_n_2292), .o(g65706_db) );
na02f02 TIMEBOOST_cell_32581 ( .a(n_12010), .b(TIMEBOOST_net_10201), .o(TIMEBOOST_net_6416) );
in01s01 g65707_u0 ( .a(FE_OFN938_n_2292), .o(g65707_sb) );
na02m02 TIMEBOOST_cell_32580 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__Q), .o(TIMEBOOST_net_10201) );
na02s01 g65707_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__Q), .b(FE_OFN938_n_2292), .o(g65707_db) );
na02f02 TIMEBOOST_cell_42518 ( .a(TIMEBOOST_net_13497), .b(g57249_sb), .o(n_10423) );
in01s01 g65708_u0 ( .a(FE_OFN952_n_2055), .o(g65708_sb) );
na02s02 TIMEBOOST_cell_44840 ( .a(TIMEBOOST_net_14658), .b(n_4470), .o(TIMEBOOST_net_11858) );
na02s01 g65708_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__Q), .b(FE_OFN952_n_2055), .o(g65708_db) );
na03s02 TIMEBOOST_cell_40431 ( .a(TIMEBOOST_net_4255), .b(g64149_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__Q), .o(TIMEBOOST_net_12454) );
in01s01 g65709_u0 ( .a(FE_OFN2109_n_2047), .o(g65709_sb) );
na02s02 TIMEBOOST_cell_17092 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(g65807_sb), .o(TIMEBOOST_net_3803) );
na02s01 g65709_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__Q), .b(FE_OFN2109_n_2047), .o(g65709_db) );
na02s02 TIMEBOOST_cell_39345 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q), .b(g64313_sb), .o(TIMEBOOST_net_11911) );
in01s01 g65710_u0 ( .a(FE_OFN1003_n_2047), .o(g65710_sb) );
na02s01 TIMEBOOST_cell_36487 ( .a(n_2544), .b(g66398_db), .o(TIMEBOOST_net_10482) );
na02s02 TIMEBOOST_cell_43605 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__26__Q), .b(n_4283), .o(TIMEBOOST_net_14041) );
na02f04 TIMEBOOST_cell_15990 ( .a(FE_RN_262_0), .b(n_5755), .o(TIMEBOOST_net_3252) );
in01s01 g65711_u0 ( .a(FE_OFN938_n_2292), .o(g65711_sb) );
na02f02 TIMEBOOST_cell_41200 ( .a(TIMEBOOST_net_12838), .b(g57584_sb), .o(n_11165) );
na02s01 g65711_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__Q), .b(FE_OFN938_n_2292), .o(g65711_db) );
na02m02 TIMEBOOST_cell_32578 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__Q), .o(TIMEBOOST_net_10200) );
in01s01 g65712_u0 ( .a(FE_OFN936_n_2292), .o(g65712_sb) );
na02f02 TIMEBOOST_cell_32577 ( .a(n_12010), .b(TIMEBOOST_net_10199), .o(TIMEBOOST_net_6414) );
na02s01 g65712_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__Q), .b(FE_OFN936_n_2292), .o(g65712_db) );
na02m02 TIMEBOOST_cell_32576 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__Q), .o(TIMEBOOST_net_10199) );
in01s01 g65713_u0 ( .a(FE_OFN1786_n_1699), .o(g65713_sb) );
na02s01 TIMEBOOST_cell_36486 ( .a(TIMEBOOST_net_10481), .b(g66402_sb), .o(n_2536) );
na02s01 g65713_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__Q), .b(FE_OFN1786_n_1699), .o(g65713_db) );
na02s02 TIMEBOOST_cell_32099 ( .a(TIMEBOOST_net_9960), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4878) );
in01s01 g65714_u0 ( .a(FE_OFN941_n_2047), .o(g65714_sb) );
na02s01 TIMEBOOST_cell_32098 ( .a(configuration_pci_err_data_521), .b(wbm_dat_o_20_), .o(TIMEBOOST_net_9960) );
na02s01 g65714_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__Q), .b(FE_OFN941_n_2047), .o(g65714_db) );
na02s01 TIMEBOOST_cell_9143 ( .a(TIMEBOOST_net_1138), .b(n_4730), .o(TIMEBOOST_net_171) );
in01s01 g65715_u0 ( .a(FE_OFN1003_n_2047), .o(g65715_sb) );
na02s02 TIMEBOOST_cell_40582 ( .a(TIMEBOOST_net_12529), .b(g62564_sb), .o(n_6430) );
na02s02 TIMEBOOST_cell_45206 ( .a(TIMEBOOST_net_14841), .b(FE_OFN1268_n_4095), .o(TIMEBOOST_net_12106) );
na02s01 TIMEBOOST_cell_40523 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__Q), .b(wishbone_slave_unit_pcim_sm_data_in), .o(TIMEBOOST_net_12500) );
na02m02 TIMEBOOST_cell_43801 ( .a(n_9589), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__Q), .o(TIMEBOOST_net_14139) );
na02s01 g65716_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__Q), .b(FE_OFN1003_n_2047), .o(g65716_db) );
no02f06 TIMEBOOST_cell_38776 ( .a(TIMEBOOST_net_11626), .b(n_15513), .o(n_15514) );
in01s01 g65717_u0 ( .a(FE_OFN1784_n_1699), .o(g65717_sb) );
na02s01 TIMEBOOST_cell_17442 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__Q), .b(g64248_sb), .o(TIMEBOOST_net_3978) );
na02s01 g65717_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__Q), .b(FE_OFN1784_n_1699), .o(g65717_db) );
na02f02 TIMEBOOST_cell_37124 ( .a(FE_OFN1602_n_13995), .b(TIMEBOOST_net_10800), .o(g53199_p) );
in01s01 g65718_u0 ( .a(FE_OFN935_n_2292), .o(g65718_sb) );
na02f02 TIMEBOOST_cell_39079 ( .a(FE_OFN1768_n_14054), .b(TIMEBOOST_net_10133), .o(TIMEBOOST_net_11778) );
na02s01 g65718_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__Q), .b(FE_OFN935_n_2292), .o(g65718_db) );
na02f02 TIMEBOOST_cell_39080 ( .a(TIMEBOOST_net_11778), .b(FE_OFN1773_n_13800), .o(g53155_p) );
in01s01 g65719_u0 ( .a(FE_OFN936_n_2292), .o(g65719_sb) );
na02f02 TIMEBOOST_cell_39081 ( .a(n_13873), .b(TIMEBOOST_net_10127), .o(TIMEBOOST_net_11779) );
na02s01 g65719_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__Q), .b(FE_OFN935_n_2292), .o(g65719_db) );
na02f02 TIMEBOOST_cell_39082 ( .a(FE_OFN1593_n_13741), .b(TIMEBOOST_net_11779), .o(n_14403) );
in01s01 g65720_u0 ( .a(FE_OFN2109_n_2047), .o(g65720_sb) );
na02s01 TIMEBOOST_cell_17094 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__Q), .b(g65909_sb), .o(TIMEBOOST_net_3804) );
na02s01 g65720_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__Q), .b(FE_OFN2109_n_2047), .o(g65720_db) );
na02f02 TIMEBOOST_cell_39129 ( .a(FE_OFN1605_n_13997), .b(TIMEBOOST_net_10172), .o(TIMEBOOST_net_11803) );
in01s01 g65721_u0 ( .a(FE_OFN953_n_2055), .o(g65721_sb) );
na02s01 g65721_u1 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(g65721_sb), .o(g65721_da) );
na02s01 g65721_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__Q), .b(FE_OFN953_n_2055), .o(g65721_db) );
na02s01 TIMEBOOST_cell_44997 ( .a(pci_target_unit_fifos_pciw_cbe_in), .b(g64113_sb), .o(TIMEBOOST_net_14737) );
in01s01 g65722_u0 ( .a(FE_OFN952_n_2055), .o(g65722_sb) );
na02s02 TIMEBOOST_cell_40420 ( .a(TIMEBOOST_net_12448), .b(FE_OFN268_n_9880), .o(n_9901) );
na02s01 g65722_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__Q), .b(FE_OFN952_n_2055), .o(g65722_db) );
na02s02 TIMEBOOST_cell_16220 ( .a(n_2306), .b(n_2755), .o(TIMEBOOST_net_3367) );
in01s01 g65723_u0 ( .a(FE_OFN950_n_2055), .o(g65723_sb) );
na02s02 TIMEBOOST_cell_16221 ( .a(TIMEBOOST_net_3367), .b(n_2487), .o(TIMEBOOST_net_178) );
na02s01 g65723_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__Q), .b(FE_OFN950_n_2055), .o(g65723_db) );
na02f06 TIMEBOOST_cell_16222 ( .a(n_16474), .b(n_168), .o(TIMEBOOST_net_3368) );
in01s01 g65724_u0 ( .a(FE_OFN956_n_1699), .o(g65724_sb) );
na02s01 TIMEBOOST_cell_45082 ( .a(TIMEBOOST_net_14779), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_11936) );
na02s01 g65724_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__Q), .b(FE_OFN956_n_1699), .o(g65724_db) );
na02s02 TIMEBOOST_cell_40312 ( .a(TIMEBOOST_net_12394), .b(n_4444), .o(n_4463) );
in01s01 g65725_u0 ( .a(FE_OFN950_n_2055), .o(g65725_sb) );
na02f06 TIMEBOOST_cell_16223 ( .a(n_16504), .b(TIMEBOOST_net_3368), .o(n_15117) );
na02s01 g65725_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__Q), .b(FE_OFN950_n_2055), .o(g65725_db) );
na02f02 TIMEBOOST_cell_42346 ( .a(TIMEBOOST_net_13411), .b(g57537_sb), .o(TIMEBOOST_net_12329) );
in01s01 g65726_u0 ( .a(FE_OFN953_n_2055), .o(g65726_sb) );
na02s02 TIMEBOOST_cell_32097 ( .a(TIMEBOOST_net_9959), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4877) );
na02s02 TIMEBOOST_cell_43071 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__Q), .b(n_3560), .o(TIMEBOOST_net_13774) );
in01s01 g65727_u0 ( .a(FE_OFN955_n_1699), .o(g65727_sb) );
na02s02 TIMEBOOST_cell_17048 ( .a(n_3770), .b(g64954_sb), .o(TIMEBOOST_net_3781) );
na02s01 g65727_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__Q), .b(FE_OFN955_n_1699), .o(g65727_db) );
na02s01 TIMEBOOST_cell_17049 ( .a(TIMEBOOST_net_3781), .b(g64954_db), .o(n_3664) );
in01s01 g65728_u0 ( .a(FE_OFN953_n_2055), .o(g65728_sb) );
na02s02 TIMEBOOST_cell_40780 ( .a(TIMEBOOST_net_12628), .b(g62465_sb), .o(n_6665) );
na02s01 g65728_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__Q), .b(FE_OFN953_n_2055), .o(g65728_db) );
no02s02 TIMEBOOST_cell_16225 ( .a(TIMEBOOST_net_3369), .b(n_1697), .o(TIMEBOOST_net_315) );
no02s01 g65729_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .b(n_905), .o(g65729_p) );
ao12s01 g65729_u1 ( .a(g65729_p), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .c(n_905), .o(n_1609) );
in01s01 g65730_u0 ( .a(FE_OFN951_n_2055), .o(g65730_sb) );
na02s01 g65730_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__Q), .b(FE_OFN952_n_2055), .o(g65730_db) );
na02s01 TIMEBOOST_cell_40584 ( .a(TIMEBOOST_net_12530), .b(g62371_sb), .o(n_6861) );
in01s01 g65731_u0 ( .a(FE_OFN953_n_2055), .o(g65731_sb) );
na02s01 g65731_u1 ( .a(pci_target_unit_fifos_pcir_data_in_167), .b(g65731_sb), .o(g65731_da) );
na02s01 g65731_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__Q), .b(FE_OFN953_n_2055), .o(g65731_db) );
na02s01 g65731_u3 ( .a(g65731_da), .b(g65731_db), .o(n_1936) );
in01s01 g65732_u0 ( .a(FE_OFN2109_n_2047), .o(g65732_sb) );
na02f02 TIMEBOOST_cell_44500 ( .a(TIMEBOOST_net_14488), .b(FE_OFN2170_n_8567), .o(TIMEBOOST_net_13450) );
na02s01 g65732_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__Q), .b(FE_OFN2109_n_2047), .o(g65732_db) );
na02s01 TIMEBOOST_cell_40314 ( .a(TIMEBOOST_net_12395), .b(g64901_db), .o(n_4411) );
in01s01 g65733_u0 ( .a(FE_OFN935_n_2292), .o(g65733_sb) );
na02s01 g65733_u1 ( .a(pci_target_unit_fifos_pcir_data_in_172), .b(g65733_sb), .o(g65733_da) );
na02s01 g65733_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__Q), .b(FE_OFN935_n_2292), .o(g65733_db) );
no02f02 TIMEBOOST_cell_38778 ( .a(TIMEBOOST_net_11627), .b(n_7214), .o(g59721_p) );
in01s01 g65734_u0 ( .a(FE_OFN1003_n_2047), .o(g65734_sb) );
na02s02 TIMEBOOST_cell_40586 ( .a(TIMEBOOST_net_12531), .b(g62538_sb), .o(n_6493) );
na02s02 TIMEBOOST_cell_45207 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__Q), .b(n_3730), .o(TIMEBOOST_net_14842) );
in01s01 g65735_u0 ( .a(FE_OFN956_n_1699), .o(g65735_sb) );
na02s01 TIMEBOOST_cell_17050 ( .a(pci_target_unit_fifos_pciw_cbe_in_152), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__Q), .o(TIMEBOOST_net_3782) );
na02s01 g65735_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__Q), .b(FE_OFN956_n_1699), .o(g65735_db) );
na02s01 TIMEBOOST_cell_17051 ( .a(TIMEBOOST_net_3782), .b(FE_OFN1059_n_4727), .o(TIMEBOOST_net_316) );
in01s01 g65736_u0 ( .a(FE_OFN955_n_1699), .o(g65736_sb) );
na02s02 TIMEBOOST_cell_17052 ( .a(n_3747), .b(g64941_sb), .o(TIMEBOOST_net_3783) );
na02s01 g65736_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__Q), .b(FE_OFN955_n_1699), .o(g65736_db) );
na02s02 TIMEBOOST_cell_17053 ( .a(TIMEBOOST_net_3783), .b(g64941_db), .o(n_3674) );
in01s01 g65737_u0 ( .a(FE_OFN941_n_2047), .o(g65737_sb) );
na02s02 TIMEBOOST_cell_40588 ( .a(TIMEBOOST_net_12532), .b(g62336_sb), .o(n_6926) );
na02s01 g65737_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__Q), .b(FE_OFN941_n_2047), .o(g65737_db) );
in01s01 g65738_u0 ( .a(FE_OFN953_n_2055), .o(g65738_sb) );
na02s01 g65738_u1 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(g65738_sb), .o(g65738_da) );
na02s01 g65738_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__Q), .b(FE_OFN953_n_2055), .o(g65738_db) );
na02s02 TIMEBOOST_cell_45178 ( .a(TIMEBOOST_net_14827), .b(FE_OFN1222_n_6391), .o(TIMEBOOST_net_12059) );
in01s01 g65739_u0 ( .a(FE_OFN952_n_2055), .o(g65739_sb) );
na03s02 TIMEBOOST_cell_40585 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__Q), .b(n_4424), .c(FE_OFN1279_n_4097), .o(TIMEBOOST_net_12531) );
na02s01 g65739_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__Q), .b(FE_OFN952_n_2055), .o(g65739_db) );
na02s02 TIMEBOOST_cell_40590 ( .a(TIMEBOOST_net_12533), .b(g62991_sb), .o(n_5900) );
in01s01 g65740_u0 ( .a(FE_OFN951_n_2055), .o(g65740_sb) );
na02s01 g65740_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__Q), .b(FE_OFN951_n_2055), .o(g65740_db) );
na02s01 TIMEBOOST_cell_37578 ( .a(TIMEBOOST_net_11027), .b(g65926_db), .o(n_2585) );
in01s01 g65741_u0 ( .a(FE_OFN953_n_2055), .o(g65741_sb) );
na02s02 TIMEBOOST_cell_40592 ( .a(TIMEBOOST_net_12534), .b(g62933_sb), .o(n_6015) );
na02s01 g65741_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__Q), .b(FE_OFN953_n_2055), .o(g65741_db) );
na02s01 TIMEBOOST_cell_40305 ( .a(n_4465), .b(g65095_sb), .o(TIMEBOOST_net_12391) );
in01s01 g65742_u0 ( .a(FE_OFN952_n_2055), .o(g65742_sb) );
na02s01 TIMEBOOST_cell_40316 ( .a(TIMEBOOST_net_12396), .b(g64908_db), .o(n_4405) );
na02s01 g65742_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__Q), .b(FE_OFN952_n_2055), .o(g65742_db) );
na02s02 TIMEBOOST_cell_40317 ( .a(g64926_sb), .b(g64926_db), .o(TIMEBOOST_net_12397) );
in01s01 g65743_u0 ( .a(FE_OFN951_n_2055), .o(g65743_sb) );
na02s01 TIMEBOOST_cell_40318 ( .a(TIMEBOOST_net_12397), .b(n_4447), .o(n_4389) );
na02s01 g65743_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__Q), .b(FE_OFN950_n_2055), .o(g65743_db) );
na02s01 TIMEBOOST_cell_40319 ( .a(g65008_sb), .b(g65008_db), .o(TIMEBOOST_net_12398) );
in01s01 g65744_u0 ( .a(FE_OFN951_n_2055), .o(g65744_sb) );
na02s02 TIMEBOOST_cell_40682 ( .a(TIMEBOOST_net_12579), .b(g62578_sb), .o(n_6398) );
na02s01 g65744_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__Q), .b(FE_OFN951_n_2055), .o(g65744_db) );
na02s01 TIMEBOOST_cell_40547 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_2__Q), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_2__Q), .o(TIMEBOOST_net_12512) );
in01s01 g65745_u0 ( .a(FE_OFN937_n_2292), .o(g65745_sb) );
na02f02 TIMEBOOST_cell_39083 ( .a(n_13903), .b(TIMEBOOST_net_10126), .o(TIMEBOOST_net_11780) );
na02s01 g65745_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__Q), .b(FE_OFN937_n_2292), .o(g65745_db) );
na02f02 TIMEBOOST_cell_39084 ( .a(TIMEBOOST_net_11780), .b(FE_OFN1596_n_13741), .o(n_14410) );
in01s01 g65746_u0 ( .a(FE_OFN950_n_2055), .o(g65746_sb) );
na02s01 TIMEBOOST_cell_31800 ( .a(configuration_wb_err_addr_552), .b(conf_wb_err_addr_in_961), .o(TIMEBOOST_net_9811) );
na02s01 g65746_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__Q), .b(FE_OFN950_n_2055), .o(g65746_db) );
na02s01 TIMEBOOST_cell_30808 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__Q), .b(pci_target_unit_fifos_pcir_data_in_183), .o(TIMEBOOST_net_9315) );
in01s01 g65747_u0 ( .a(FE_OFN2109_n_2047), .o(g65747_sb) );
na02s02 TIMEBOOST_cell_17098 ( .a(pci_target_unit_fifos_pcir_control_in_192), .b(g64145_sb), .o(TIMEBOOST_net_3806) );
na02s01 g65747_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__Q), .b(FE_OFN2108_n_2047), .o(g65747_db) );
na02m02 TIMEBOOST_cell_39175 ( .a(TIMEBOOST_net_1643), .b(wishbone_slave_unit_pcim_if_wbw_cbe_in_416), .o(TIMEBOOST_net_11826) );
in01s01 g65748_u0 ( .a(FE_OFN955_n_1699), .o(g65748_sb) );
na02s01 TIMEBOOST_cell_17054 ( .a(n_3780), .b(g65051_sb), .o(TIMEBOOST_net_3784) );
na02s01 g65748_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__Q), .b(FE_OFN955_n_1699), .o(g65748_db) );
na02s01 TIMEBOOST_cell_17055 ( .a(TIMEBOOST_net_3784), .b(g65051_db), .o(n_3619) );
in01s01 g65749_u0 ( .a(FE_OFN951_n_2055), .o(g65749_sb) );
na02s02 TIMEBOOST_cell_43385 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__31__Q), .b(n_4646), .o(TIMEBOOST_net_13931) );
na02s01 TIMEBOOST_cell_32096 ( .a(configuration_pci_err_data_520), .b(wbm_dat_o_19_), .o(TIMEBOOST_net_9959) );
na02s01 TIMEBOOST_cell_31790 ( .a(parchk_pci_ad_out_in_1180), .b(configuration_wb_err_data_583), .o(TIMEBOOST_net_9806) );
in01s01 g65750_u0 ( .a(FE_OFN1786_n_1699), .o(g65750_sb) );
na02s02 TIMEBOOST_cell_32095 ( .a(TIMEBOOST_net_9958), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4876) );
na02s01 g65750_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__Q), .b(FE_OFN1786_n_1699), .o(g65750_db) );
na02m02 TIMEBOOST_cell_43606 ( .a(TIMEBOOST_net_14041), .b(FE_OFN1322_n_6436), .o(TIMEBOOST_net_12222) );
in01s01 g65751_u0 ( .a(FE_OFN2108_n_2047), .o(g65751_sb) );
na02s02 TIMEBOOST_cell_17100 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(g65693_sb), .o(TIMEBOOST_net_3807) );
na02s01 g65751_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__Q), .b(FE_OFN2108_n_2047), .o(g65751_db) );
na02s01 TIMEBOOST_cell_39205 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__Q), .b(n_8140), .o(TIMEBOOST_net_11841) );
in01s01 g65752_u0 ( .a(FE_OFN1012_n_4734), .o(g65752_sb) );
na02s01 g65752_u1 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(g65752_sb), .o(g65752_da) );
na02s01 g65752_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__Q), .b(FE_OFN1012_n_4734), .o(g65752_db) );
na02s01 g65752_u3 ( .a(g65752_da), .b(g65752_db), .o(n_3213) );
in01s01 g65753_u0 ( .a(FE_OFN1003_n_2047), .o(g65753_sb) );
na02s02 TIMEBOOST_cell_45179 ( .a(n_3658), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__Q), .o(TIMEBOOST_net_14828) );
na02s01 g65753_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__Q), .b(FE_OFN1003_n_2047), .o(g65753_db) );
na02s01 TIMEBOOST_cell_40320 ( .a(TIMEBOOST_net_12398), .b(n_4447), .o(n_4349) );
in01s01 g65754_u0 ( .a(FE_OFN950_n_2055), .o(g65754_sb) );
na02s02 TIMEBOOST_cell_40594 ( .a(TIMEBOOST_net_12535), .b(g62466_sb), .o(n_6662) );
na02s01 g65754_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__Q), .b(FE_OFN950_n_2055), .o(g65754_db) );
na02s01 TIMEBOOST_cell_44998 ( .a(TIMEBOOST_net_14737), .b(g64113_db), .o(n_4739) );
in01s01 g65755_u0 ( .a(FE_OFN1785_n_1699), .o(g65755_sb) );
na02s01 TIMEBOOST_cell_32094 ( .a(configuration_pci_err_data_518), .b(wbm_dat_o_17_), .o(TIMEBOOST_net_9958) );
na02s01 g65755_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__Q), .b(FE_OFN1785_n_1699), .o(g65755_db) );
na02s02 TIMEBOOST_cell_38092 ( .a(TIMEBOOST_net_11284), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_4578) );
in01s01 g65756_u0 ( .a(FE_OFN1783_n_1699), .o(g65756_sb) );
na02s01 TIMEBOOST_cell_32092 ( .a(configuration_pci_err_data_515), .b(wbm_dat_o_14_), .o(TIMEBOOST_net_9957) );
na02s01 g65756_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__Q), .b(FE_OFN1783_n_1699), .o(g65756_db) );
na02s02 TIMEBOOST_cell_38094 ( .a(TIMEBOOST_net_11285), .b(FE_OFN1139_g64577_p), .o(TIMEBOOST_net_4503) );
na02s01 TIMEBOOST_cell_32090 ( .a(configuration_pci_err_data_513), .b(wbm_dat_o_12_), .o(TIMEBOOST_net_9956) );
na02s01 g65757_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__Q), .b(FE_OFN902_n_4736), .o(g65757_db) );
na02s02 TIMEBOOST_cell_40596 ( .a(TIMEBOOST_net_12536), .b(g62997_sb), .o(n_5888) );
in01s01 g65758_u0 ( .a(FE_OFN952_n_2055), .o(g65758_sb) );
na02s01 TIMEBOOST_cell_40598 ( .a(TIMEBOOST_net_12537), .b(g62460_sb), .o(n_6676) );
na02s01 g65758_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__Q), .b(FE_OFN952_n_2055), .o(g65758_db) );
na02s02 TIMEBOOST_cell_16242 ( .a(n_3792), .b(g64754_sb), .o(TIMEBOOST_net_3378) );
in01s01 g65759_u0 ( .a(FE_OFN951_n_2055), .o(g65759_sb) );
na02s01 TIMEBOOST_cell_16243 ( .a(TIMEBOOST_net_3378), .b(g64754_db), .o(n_3789) );
na02s01 g65759_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__Q), .b(FE_OFN951_n_2055), .o(g65759_db) );
na02s01 TIMEBOOST_cell_16244 ( .a(n_3747), .b(g64769_sb), .o(TIMEBOOST_net_3379) );
in01s01 g65760_u0 ( .a(FE_OFN1783_n_1699), .o(g65760_sb) );
no02f02 TIMEBOOST_cell_38777 ( .a(n_4144), .b(n_7552), .o(TIMEBOOST_net_11627) );
na02s01 g65760_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__Q), .b(FE_OFN1783_n_1699), .o(g65760_db) );
na02s01 TIMEBOOST_cell_39484 ( .a(TIMEBOOST_net_11980), .b(TIMEBOOST_net_9824), .o(n_7141) );
in01s01 g65761_u0 ( .a(FE_OFN1003_n_2047), .o(g65761_sb) );
na02s02 TIMEBOOST_cell_32089 ( .a(TIMEBOOST_net_9955), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_4873) );
na02s02 TIMEBOOST_cell_45208 ( .a(TIMEBOOST_net_14842), .b(FE_OFN1219_n_6886), .o(TIMEBOOST_net_12535) );
na02s01 TIMEBOOST_cell_32088 ( .a(configuration_pci_err_addr_479), .b(wbm_adr_o_9_), .o(TIMEBOOST_net_9955) );
in01s01 g65762_u0 ( .a(FE_OFN950_n_2055), .o(g65762_sb) );
na02s01 TIMEBOOST_cell_16245 ( .a(TIMEBOOST_net_3379), .b(g64769_db), .o(n_3779) );
na02s01 g65762_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__Q), .b(FE_OFN950_n_2055), .o(g65762_db) );
na02s01 TIMEBOOST_cell_37580 ( .a(TIMEBOOST_net_11028), .b(g61722_sb), .o(n_8379) );
na02f02 TIMEBOOST_cell_43764 ( .a(TIMEBOOST_net_14120), .b(FE_OFN1377_n_8567), .o(TIMEBOOST_net_12761) );
na02s01 g65763_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__Q), .b(FE_OFN1003_n_2047), .o(g65763_db) );
na02f02 TIMEBOOST_cell_43765 ( .a(n_9593), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__Q), .o(TIMEBOOST_net_14121) );
in01s01 g65764_u0 ( .a(FE_OFN941_n_2047), .o(g65764_sb) );
na02s02 TIMEBOOST_cell_32087 ( .a(TIMEBOOST_net_9954), .b(FE_OFN1180_n_3476), .o(TIMEBOOST_net_4872) );
na02s01 g65764_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__Q), .b(FE_OFN941_n_2047), .o(g65764_db) );
na02s01 TIMEBOOST_cell_16000 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__Q), .b(FE_OCPN1839_n_1238), .o(TIMEBOOST_net_3257) );
na02s01 TIMEBOOST_cell_32086 ( .a(configuration_pci_err_addr_475), .b(wbm_adr_o_5_), .o(TIMEBOOST_net_9954) );
na02f02 TIMEBOOST_cell_43766 ( .a(TIMEBOOST_net_14121), .b(FE_OFN1417_n_8567), .o(TIMEBOOST_net_12945) );
na02s01 TIMEBOOST_cell_16001 ( .a(TIMEBOOST_net_3257), .b(g65269_sb), .o(TIMEBOOST_net_165) );
in01s01 g65766_u0 ( .a(FE_OFN955_n_1699), .o(g65766_sb) );
na02s01 TIMEBOOST_cell_40313 ( .a(n_4452), .b(g64901_sb), .o(TIMEBOOST_net_12395) );
na02s01 g65766_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__Q), .b(FE_OFN955_n_1699), .o(g65766_db) );
na02s01 TIMEBOOST_cell_40322 ( .a(TIMEBOOST_net_12399), .b(g65031_db), .o(n_4335) );
in01s01 g65767_u0 ( .a(FE_OFN953_n_2055), .o(g65767_sb) );
na02s01 TIMEBOOST_cell_9343 ( .a(TIMEBOOST_net_1238), .b(g64197_db), .o(n_3972) );
na02s02 TIMEBOOST_cell_32085 ( .a(TIMEBOOST_net_9953), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_4871) );
na02s01 TIMEBOOST_cell_31788 ( .a(conf_wb_err_addr_in_960), .b(configuration_wb_err_addr_551), .o(TIMEBOOST_net_9805) );
in01s01 g65768_u0 ( .a(FE_OFN956_n_1699), .o(g65768_sb) );
na02s02 TIMEBOOST_cell_17058 ( .a(n_3744), .b(g64944_sb), .o(TIMEBOOST_net_3786) );
na02s01 TIMEBOOST_cell_39511 ( .a(g64253_da), .b(g64253_db), .o(TIMEBOOST_net_11994) );
na02s02 TIMEBOOST_cell_17059 ( .a(TIMEBOOST_net_3786), .b(g64944_db), .o(n_3670) );
in01s01 g65769_u0 ( .a(FE_OFN941_n_2047), .o(g65769_sb) );
na02s02 TIMEBOOST_cell_16002 ( .a(n_5769), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_3258) );
na02s01 g65769_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__Q), .b(FE_OFN941_n_2047), .o(g65769_db) );
na02m02 TIMEBOOST_cell_43733 ( .a(n_9010), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__Q), .o(TIMEBOOST_net_14105) );
in01s01 g65770_u0 ( .a(FE_OFN941_n_2047), .o(g65770_sb) );
na02s02 TIMEBOOST_cell_16004 ( .a(FE_OFN276_n_9941), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__Q), .o(TIMEBOOST_net_3259) );
na02s01 g65770_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__Q), .b(FE_OFN941_n_2047), .o(g65770_db) );
na02s01 TIMEBOOST_cell_32084 ( .a(configuration_pci_err_addr_473), .b(wbm_adr_o_3_), .o(TIMEBOOST_net_9953) );
in01s01 g65771_u0 ( .a(FE_OFN956_n_1699), .o(g65771_sb) );
na02s01 TIMEBOOST_cell_17060 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__Q), .b(g65965_sb), .o(TIMEBOOST_net_3787) );
na02s01 g65771_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__Q), .b(FE_OFN956_n_1699), .o(g65771_db) );
na02m02 TIMEBOOST_cell_44191 ( .a(n_9640), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__Q), .o(TIMEBOOST_net_14334) );
in01s01 g65772_u0 ( .a(FE_OFN935_n_2292), .o(g65772_sb) );
na02f02 TIMEBOOST_cell_45541 ( .a(TIMEBOOST_net_10162), .b(FE_OFN1606_n_13997), .o(TIMEBOOST_net_15009) );
na02s01 g65772_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__Q), .b(FE_OFN935_n_2292), .o(g65772_db) );
na02s01 TIMEBOOST_cell_39206 ( .a(TIMEBOOST_net_11841), .b(n_1569), .o(TIMEBOOST_net_11460) );
in01s01 g65773_u0 ( .a(FE_OFN2108_n_2047), .o(g65773_sb) );
na02s02 TIMEBOOST_cell_17102 ( .a(pci_target_unit_fifos_pcir_data_in_187), .b(g65702_sb), .o(TIMEBOOST_net_3808) );
na02s01 g65773_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__Q), .b(FE_OFN2108_n_2047), .o(g65773_db) );
na02f02 TIMEBOOST_cell_44192 ( .a(TIMEBOOST_net_14334), .b(FE_OFN1368_n_8567), .o(TIMEBOOST_net_12701) );
in01s01 g65774_u0 ( .a(FE_OFN935_n_2292), .o(g65774_sb) );
in01s01 TIMEBOOST_cell_32834 ( .a(TIMEBOOST_net_10335), .o(wbs_dat_i_16_) );
na02s01 g65774_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__Q), .b(FE_OFN935_n_2292), .o(g65774_db) );
na02f02 TIMEBOOST_cell_41246 ( .a(TIMEBOOST_net_12861), .b(g57070_sb), .o(n_11671) );
in01s01 g65775_u0 ( .a(FE_OFN937_n_2292), .o(g65775_sb) );
na02f02 TIMEBOOST_cell_45542 ( .a(TIMEBOOST_net_15009), .b(FE_OFN1599_n_13995), .o(n_14476) );
na02s01 g65775_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__Q), .b(FE_OFN937_n_2292), .o(g65775_db) );
na02s02 TIMEBOOST_cell_18825 ( .a(TIMEBOOST_net_4669), .b(g62723_sb), .o(n_5537) );
in01s01 g65776_u0 ( .a(FE_OFN936_n_2292), .o(g65776_sb) );
na02f02 TIMEBOOST_cell_39085 ( .a(TIMEBOOST_net_10132), .b(n_13901), .o(TIMEBOOST_net_11781) );
na02s01 g65776_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__Q), .b(FE_OFN936_n_2292), .o(g65776_db) );
na02f02 TIMEBOOST_cell_39086 ( .a(FE_OFN1593_n_13741), .b(TIMEBOOST_net_11781), .o(g53276_p) );
in01s01 g65777_u0 ( .a(FE_OFN1783_n_1699), .o(g65777_sb) );
na02s02 TIMEBOOST_cell_32083 ( .a(TIMEBOOST_net_9952), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_4870) );
na02s01 g65777_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__Q), .b(FE_OFN1783_n_1699), .o(g65777_db) );
na02s01 TIMEBOOST_cell_32082 ( .a(configuration_pci_err_addr_472), .b(wbm_adr_o_2_), .o(TIMEBOOST_net_9952) );
in01s01 g65778_u0 ( .a(FE_OFN1784_n_1699), .o(g65778_sb) );
na02s02 TIMEBOOST_cell_32081 ( .a(TIMEBOOST_net_9951), .b(FE_OFN1180_n_3476), .o(TIMEBOOST_net_4869) );
na02s01 g65778_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__Q), .b(FE_OFN1784_n_1699), .o(g65778_db) );
na02s01 TIMEBOOST_cell_32080 ( .a(configuration_pci_err_addr_496), .b(wbm_adr_o_26_), .o(TIMEBOOST_net_9951) );
in01s01 g65779_u0 ( .a(FE_OFN950_n_2055), .o(g65779_sb) );
na02s01 TIMEBOOST_cell_16246 ( .a(n_3744), .b(g64772_sb), .o(TIMEBOOST_net_3380) );
na02s01 g65779_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__Q), .b(FE_OFN950_n_2055), .o(g65779_db) );
na02f02 TIMEBOOST_cell_32497 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_10159), .o(TIMEBOOST_net_6330) );
in01s01 g65780_u0 ( .a(FE_OFN935_n_2292), .o(g65780_sb) );
na02s01 g65780_u1 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(g65780_sb), .o(g65780_da) );
na02s01 g65780_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__Q), .b(FE_OFN935_n_2292), .o(g65780_db) );
na02m02 TIMEBOOST_cell_42261 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__Q), .b(n_9676), .o(TIMEBOOST_net_13369) );
in01s01 g65781_u0 ( .a(FE_OFN950_n_2055), .o(g65781_sb) );
na03s02 TIMEBOOST_cell_39499 ( .a(g64200_da), .b(g64200_db), .c(g62803_db), .o(TIMEBOOST_net_11988) );
in01s01 TIMEBOOST_cell_32833 ( .a(TIMEBOOST_net_10334), .o(TIMEBOOST_net_10333) );
in01s01 g65782_u0 ( .a(FE_OFN1784_n_1699), .o(g65782_sb) );
no02f06 TIMEBOOST_cell_38775 ( .a(FE_RN_538_0), .b(FE_RN_539_0), .o(TIMEBOOST_net_11626) );
na02s01 g65782_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__Q), .b(FE_OFN1784_n_1699), .o(g65782_db) );
na02f02 TIMEBOOST_cell_38780 ( .a(TIMEBOOST_net_11628), .b(n_14618), .o(TIMEBOOST_net_10022) );
in01s01 g65783_u0 ( .a(FE_OFN956_n_1699), .o(g65783_sb) );
na02s01 TIMEBOOST_cell_17062 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__Q), .b(g65966_sb), .o(TIMEBOOST_net_3788) );
na02s01 g65783_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__Q), .b(FE_OFN956_n_1699), .o(g65783_db) );
na02f02 TIMEBOOST_cell_43802 ( .a(TIMEBOOST_net_14139), .b(FE_OFN1425_n_8567), .o(TIMEBOOST_net_12962) );
in01s01 g65784_u0 ( .a(FE_OFN941_n_2047), .o(g65784_sb) );
na02s02 TIMEBOOST_cell_32079 ( .a(TIMEBOOST_net_9950), .b(FE_OFN1180_n_3476), .o(TIMEBOOST_net_4868) );
na02s01 g65784_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__Q), .b(FE_OFN941_n_2047), .o(g65784_db) );
na02s01 TIMEBOOST_cell_32078 ( .a(configuration_pci_err_addr_494), .b(wbm_adr_o_24_), .o(TIMEBOOST_net_9950) );
na02s02 TIMEBOOST_cell_16006 ( .a(n_2705), .b(n_1096), .o(TIMEBOOST_net_3260) );
na02s02 TIMEBOOST_cell_32077 ( .a(TIMEBOOST_net_9949), .b(FE_OFN1179_n_3476), .o(TIMEBOOST_net_4937) );
in01s01 g65786_u0 ( .a(FE_OFN956_n_1699), .o(g65786_sb) );
na02s01 TIMEBOOST_cell_17064 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__Q), .b(g65969_sb), .o(TIMEBOOST_net_3789) );
na02m02 TIMEBOOST_cell_39173 ( .a(n_1083), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_11825) );
in01s01 g65787_u0 ( .a(FE_OFN941_n_2047), .o(g65787_sb) );
na02s02 TIMEBOOST_cell_16007 ( .a(TIMEBOOST_net_3260), .b(n_2243), .o(TIMEBOOST_net_307) );
na02s01 g65787_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__Q), .b(FE_OFN941_n_2047), .o(g65787_db) );
na03s02 TIMEBOOST_cell_39471 ( .a(TIMEBOOST_net_3960), .b(g64260_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__Q), .o(TIMEBOOST_net_11974) );
in01s01 g65788_u0 ( .a(FE_OFN955_n_1699), .o(g65788_sb) );
na02s02 TIMEBOOST_cell_17066 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(g65720_sb), .o(TIMEBOOST_net_3790) );
na02s01 g65788_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__Q), .b(FE_OFN955_n_1699), .o(g65788_db) );
na02s01 TIMEBOOST_cell_44841 ( .a(n_3774), .b(g64774_sb), .o(TIMEBOOST_net_14659) );
in01s01 g65789_u0 ( .a(FE_OFN938_n_2292), .o(g65789_sb) );
na02f02 TIMEBOOST_cell_41226 ( .a(TIMEBOOST_net_12851), .b(g57191_sb), .o(n_10447) );
na02s01 g65789_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__Q), .b(FE_OFN938_n_2292), .o(g65789_db) );
na03f04 TIMEBOOST_cell_45543 ( .a(n_10880), .b(n_10881), .c(n_11720), .o(TIMEBOOST_net_15010) );
in01s01 g65790_u0 ( .a(FE_OFN1785_n_1699), .o(g65790_sb) );
na02s01 TIMEBOOST_cell_32076 ( .a(configuration_pci_err_addr_492), .b(wbm_adr_o_22_), .o(TIMEBOOST_net_9949) );
na02s01 g65790_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__Q), .b(FE_OFN1785_n_1699), .o(g65790_db) );
na02s02 TIMEBOOST_cell_32075 ( .a(TIMEBOOST_net_9948), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4936) );
in01s01 g65791_u0 ( .a(FE_OFN955_n_1699), .o(g65791_sb) );
na02s02 TIMEBOOST_cell_17068 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(g65732_sb), .o(TIMEBOOST_net_3791) );
na02s01 g65791_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__Q), .b(FE_OFN955_n_1699), .o(g65791_db) );
na02m02 TIMEBOOST_cell_43803 ( .a(n_9787), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__Q), .o(TIMEBOOST_net_14140) );
in01s01 g65792_u0 ( .a(FE_OFN1786_n_1699), .o(g65792_sb) );
na02s01 TIMEBOOST_cell_32074 ( .a(configuration_pci_err_addr_487), .b(wbm_adr_o_17_), .o(TIMEBOOST_net_9948) );
na02s01 g65792_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__Q), .b(FE_OFN1786_n_1699), .o(g65792_db) );
na02s02 TIMEBOOST_cell_32073 ( .a(TIMEBOOST_net_9947), .b(FE_OFN1180_n_3476), .o(TIMEBOOST_net_4935) );
in01s01 g65793_u0 ( .a(FE_OFN955_n_1699), .o(g65793_sb) );
na02f02 TIMEBOOST_cell_41630 ( .a(FE_OFN1440_n_9372), .b(TIMEBOOST_net_13053), .o(TIMEBOOST_net_11678) );
na02s01 g65793_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__Q), .b(FE_OFN955_n_1699), .o(g65793_db) );
na02s02 TIMEBOOST_cell_17071 ( .a(TIMEBOOST_net_3792), .b(g58062_sb), .o(n_9090) );
in01s01 g65794_u0 ( .a(FE_OFN1786_n_1699), .o(g65794_sb) );
na02s01 TIMEBOOST_cell_32072 ( .a(configuration_pci_err_data_511), .b(wbm_dat_o_10_), .o(TIMEBOOST_net_9947) );
na02s01 g65794_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__Q), .b(FE_OFN1786_n_1699), .o(g65794_db) );
na02s02 TIMEBOOST_cell_40796 ( .a(TIMEBOOST_net_12636), .b(g62909_sb), .o(n_6060) );
in01s01 g65795_u0 ( .a(FE_OFN1784_n_1699), .o(g65795_sb) );
na02s02 TIMEBOOST_cell_17448 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(g64183_sb), .o(TIMEBOOST_net_3981) );
na02s01 g65795_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__Q), .b(FE_OFN1784_n_1699), .o(g65795_db) );
na02s02 TIMEBOOST_cell_44999 ( .a(pci_target_unit_fifos_pciw_addr_data_in_123), .b(g64099_sb), .o(TIMEBOOST_net_14738) );
na03f10 TIMEBOOST_cell_16010 ( .a(n_15414), .b(n_15417), .c(n_16854), .o(TIMEBOOST_net_3262) );
na02m02 TIMEBOOST_cell_43767 ( .a(n_9510), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__Q), .o(TIMEBOOST_net_14122) );
na02f10 TIMEBOOST_cell_16011 ( .a(n_16855), .b(TIMEBOOST_net_3262), .o(n_15347) );
in01s01 g65797_u0 ( .a(FE_OFN956_n_1699), .o(g65797_sb) );
na02m02 TIMEBOOST_cell_32496 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__Q), .o(TIMEBOOST_net_10159) );
na02f02 TIMEBOOST_cell_41228 ( .a(TIMEBOOST_net_12852), .b(g57372_sb), .o(n_11377) );
na02s02 TIMEBOOST_cell_45583 ( .a(n_4444), .b(g64967_sb), .o(TIMEBOOST_net_15030) );
in01s01 g65798_u0 ( .a(FE_OFN956_n_1699), .o(g65798_sb) );
na02s01 TIMEBOOST_cell_8984 ( .a(n_1415), .b(n_1679), .o(TIMEBOOST_net_1059) );
na02s01 g65798_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__Q), .b(FE_OFN956_n_1699), .o(g65798_db) );
na02m01 TIMEBOOST_cell_8985 ( .a(TIMEBOOST_net_1059), .b(n_2237), .o(TIMEBOOST_net_134) );
in01s01 g65799_u0 ( .a(FE_OFN956_n_1699), .o(g65799_sb) );
na02s01 TIMEBOOST_cell_8986 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q), .o(TIMEBOOST_net_1060) );
na02s01 g65799_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__Q), .b(FE_OFN956_n_1699), .o(g65799_db) );
na02s02 TIMEBOOST_cell_8987 ( .a(TIMEBOOST_net_1060), .b(n_1993), .o(TIMEBOOST_net_220) );
in01s01 g65800_u0 ( .a(FE_OFN951_n_2055), .o(g65800_sb) );
na02s01 TIMEBOOST_cell_16247 ( .a(TIMEBOOST_net_3380), .b(g64772_db), .o(n_3776) );
na02s01 g65800_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__Q), .b(FE_OFN951_n_2055), .o(g65800_db) );
na02s01 TIMEBOOST_cell_16248 ( .a(n_3741), .b(g64776_sb), .o(TIMEBOOST_net_3381) );
no02m02 g65801_u0 ( .a(n_908), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .o(g65801_p) );
ao12m02 g65801_u1 ( .a(g65801_p), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .c(n_908), .o(n_6136) );
in01s01 g65802_u0 ( .a(FE_OFN935_n_2292), .o(g65802_sb) );
na02f02 TIMEBOOST_cell_39087 ( .a(FE_OFN1774_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__Q), .o(TIMEBOOST_net_11782) );
na02s01 g65802_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__Q), .b(FE_OFN935_n_2292), .o(g65802_db) );
na02f02 TIMEBOOST_cell_39088 ( .a(TIMEBOOST_net_11782), .b(n_14174), .o(n_16233) );
in01s01 g65803_u0 ( .a(FE_OFN938_n_2292), .o(g65803_sb) );
na02f02 TIMEBOOST_cell_32615 ( .a(TIMEBOOST_net_10218), .b(n_14832), .o(n_14894) );
na02s01 g65803_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__Q), .b(FE_OFN938_n_2292), .o(g65803_db) );
na02f02 TIMEBOOST_cell_32614 ( .a(n_14895), .b(n_13487), .o(TIMEBOOST_net_10218) );
in01s01 g65804_u0 ( .a(FE_OFN952_n_2055), .o(g65804_sb) );
na02s01 TIMEBOOST_cell_16249 ( .a(TIMEBOOST_net_3381), .b(g64776_db), .o(n_3773) );
na02s01 g65804_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__Q), .b(FE_OFN952_n_2055), .o(g65804_db) );
na02s01 TIMEBOOST_cell_16250 ( .a(n_3739), .b(g64781_sb), .o(TIMEBOOST_net_3382) );
in01s01 g65805_u0 ( .a(FE_OFN1784_n_1699), .o(g65805_sb) );
na02s02 TIMEBOOST_cell_32071 ( .a(TIMEBOOST_net_9946), .b(FE_OFN1179_n_3476), .o(TIMEBOOST_net_4934) );
na02s01 g65805_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__Q), .b(FE_OFN1784_n_1699), .o(g65805_db) );
na02s01 TIMEBOOST_cell_32070 ( .a(configuration_pci_err_addr_477), .b(wbm_adr_o_7_), .o(TIMEBOOST_net_9946) );
in01s01 g65806_u0 ( .a(FE_OFN1785_n_1699), .o(g65806_sb) );
na02s02 TIMEBOOST_cell_32069 ( .a(TIMEBOOST_net_9945), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4933) );
na02s01 g65806_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__Q), .b(FE_OFN1785_n_1699), .o(g65806_db) );
na02s01 TIMEBOOST_cell_32068 ( .a(configuration_pci_err_addr_490), .b(wbm_adr_o_20_), .o(TIMEBOOST_net_9945) );
in01s01 g65807_u0 ( .a(FE_OFN2108_n_2047), .o(g65807_sb) );
na02s01 TIMEBOOST_cell_40315 ( .a(n_4444), .b(g64908_sb), .o(TIMEBOOST_net_12396) );
na02s01 g65807_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__Q), .b(FE_OFN2108_n_2047), .o(g65807_db) );
na02s01 TIMEBOOST_cell_40324 ( .a(TIMEBOOST_net_12400), .b(g58453_db), .o(n_9404) );
na02s01 TIMEBOOST_cell_42089 ( .a(g64985_db), .b(FE_OFN1226_n_6391), .o(TIMEBOOST_net_13283) );
na02m02 TIMEBOOST_cell_44399 ( .a(n_9658), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__Q), .o(TIMEBOOST_net_14438) );
na03s02 TIMEBOOST_cell_33592 ( .a(TIMEBOOST_net_3562), .b(g64891_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__Q), .o(TIMEBOOST_net_4811) );
in01f02 g65808_u3 ( .a(g65808_p), .o(n_1588) );
in01s01 g65809_u0 ( .a(FE_OFN1017_n_2053), .o(g65809_sb) );
na02s01 TIMEBOOST_cell_40281 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__Q), .b(n_8140), .o(TIMEBOOST_net_12379) );
na02s01 g65809_u2 ( .a(pci_target_unit_fifos_pcir_data_in_172), .b(FE_OFN1017_n_2053), .o(g65809_db) );
na02s01 TIMEBOOST_cell_40326 ( .a(TIMEBOOST_net_12401), .b(g65435_sb), .o(n_4219) );
in01s01 g65810_u0 ( .a(n_2299), .o(g65810_sb) );
na02f04 TIMEBOOST_cell_45544 ( .a(TIMEBOOST_net_15010), .b(n_12564), .o(n_12826) );
na02f02 TIMEBOOST_cell_45545 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__Q), .b(FE_OFN1740_n_11019), .o(TIMEBOOST_net_15011) );
na02f02 TIMEBOOST_cell_45546 ( .a(TIMEBOOST_net_15011), .b(n_11954), .o(n_12500) );
in01s01 g65811_u0 ( .a(FE_OFN1017_n_2053), .o(g65811_sb) );
na02s02 TIMEBOOST_cell_22249 ( .a(n_10213), .b(TIMEBOOST_net_6381), .o(n_11863) );
na02s01 g65811_u2 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(FE_OFN1017_n_2053), .o(g65811_db) );
na02f02 TIMEBOOST_cell_44400 ( .a(TIMEBOOST_net_14438), .b(FE_OFN1421_n_8567), .o(TIMEBOOST_net_12780) );
in01s01 g65812_u0 ( .a(FE_OFN1017_n_2053), .o(g65812_sb) );
na02s02 TIMEBOOST_cell_36672 ( .a(TIMEBOOST_net_10574), .b(g61798_db), .o(n_8200) );
na02s01 g65812_u2 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(FE_OFN1017_n_2053), .o(g65812_db) );
na02f02 TIMEBOOST_cell_40950 ( .a(TIMEBOOST_net_12713), .b(g57136_sb), .o(n_11614) );
in01s02 g65813_u0 ( .a(FE_OFN776_n_15366), .o(g65813_sb) );
na02s01 TIMEBOOST_cell_37778 ( .a(TIMEBOOST_net_11127), .b(FE_OFN712_n_8140), .o(TIMEBOOST_net_4344) );
na02s01 g65813_u2 ( .a(pci_target_unit_del_sync_addr_in_214), .b(FE_OFN776_n_15366), .o(g65813_db) );
na02f02 TIMEBOOST_cell_37121 ( .a(TIMEBOOST_net_10157), .b(FE_OFN1606_n_13997), .o(TIMEBOOST_net_10799) );
in01s01 g65814_u0 ( .a(FE_OFN1017_n_2053), .o(g65814_sb) );
na02s01 TIMEBOOST_cell_16856 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__Q), .b(g64285_sb), .o(TIMEBOOST_net_3685) );
na02s01 g65814_u2 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(FE_OFN1017_n_2053), .o(g65814_db) );
na02f02 TIMEBOOST_cell_45547 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__Q), .b(n_12020), .o(TIMEBOOST_net_15012) );
in01s01 g65815_u0 ( .a(FE_OFN2113_n_2053), .o(g65815_sb) );
na02s02 TIMEBOOST_cell_17996 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(g64149_sb), .o(TIMEBOOST_net_4255) );
na02s01 g65815_u2 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(FE_OFN2113_n_2053), .o(g65815_db) );
na02s01 TIMEBOOST_cell_39483 ( .a(wbs_dat_i_20_), .b(g63618_db), .o(TIMEBOOST_net_11980) );
in01s01 g65816_u0 ( .a(FE_OFN1016_n_2053), .o(g65816_sb) );
na02s01 TIMEBOOST_cell_41903 ( .a(g62738_sb), .b(g62738_db), .o(TIMEBOOST_net_13190) );
na02s01 g65816_u2 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(FE_OFN1016_n_2053), .o(g65816_db) );
na02s01 TIMEBOOST_cell_16915 ( .a(TIMEBOOST_net_3714), .b(g65398_db), .o(n_3520) );
na02s01 TIMEBOOST_cell_9145 ( .a(TIMEBOOST_net_1139), .b(n_4730), .o(TIMEBOOST_net_172) );
na02s01 TIMEBOOST_cell_9147 ( .a(TIMEBOOST_net_1140), .b(n_4730), .o(TIMEBOOST_net_173) );
in01s01 g65818_u0 ( .a(FE_OFN1016_n_2053), .o(g65818_sb) );
in01s01 TIMEBOOST_cell_8834 ( .a(conf_wb_err_addr_in_951), .o(TIMEBOOST_net_971) );
na02s01 g65818_u2 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(FE_OFN1016_n_2053), .o(g65818_db) );
in01s01 TIMEBOOST_cell_8835 ( .a(TIMEBOOST_net_971), .o(TIMEBOOST_net_972) );
in01s01 g65819_u0 ( .a(FE_OFN1016_n_2053), .o(g65819_sb) );
in01s01 TIMEBOOST_cell_8836 ( .a(conf_wb_err_addr_in_953), .o(TIMEBOOST_net_973) );
na02s01 g65819_u2 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(FE_OFN1016_n_2053), .o(g65819_db) );
in01s01 TIMEBOOST_cell_8837 ( .a(TIMEBOOST_net_973), .o(TIMEBOOST_net_974) );
in01s01 g65820_u0 ( .a(FE_OFN2113_n_2053), .o(g65820_sb) );
na02s02 TIMEBOOST_cell_17998 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(g65251_sb), .o(TIMEBOOST_net_4256) );
na02s01 TIMEBOOST_cell_18224 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_407), .b(FE_OFN2070_n_15978), .o(TIMEBOOST_net_4369) );
na03s02 TIMEBOOST_cell_38125 ( .a(g64148_da), .b(g64148_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__Q), .o(TIMEBOOST_net_11301) );
in01s01 g65821_u0 ( .a(FE_OFN1016_n_2053), .o(g65821_sb) );
in01s01 TIMEBOOST_cell_8838 ( .a(conf_wb_err_addr_in_954), .o(TIMEBOOST_net_975) );
na02s01 g65821_u2 ( .a(pci_target_unit_fifos_pcir_data_in_188), .b(FE_OFN1016_n_2053), .o(g65821_db) );
in01s01 TIMEBOOST_cell_8839 ( .a(TIMEBOOST_net_975), .o(TIMEBOOST_net_976) );
in01s01 g65822_u0 ( .a(FE_OFN1016_n_2053), .o(g65822_sb) );
na02s01 TIMEBOOST_cell_17898 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__Q), .b(g61943_sb), .o(TIMEBOOST_net_4206) );
na02s01 g65822_u2 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(FE_OFN1016_n_2053), .o(g65822_db) );
na02f02 TIMEBOOST_cell_44193 ( .a(n_9057), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__Q), .o(TIMEBOOST_net_14335) );
in01s01 g65823_u0 ( .a(FE_OFN1016_n_2053), .o(g65823_sb) );
in01s01 TIMEBOOST_cell_8840 ( .a(conf_wb_err_addr_in_958), .o(TIMEBOOST_net_977) );
na02s01 g65823_u2 ( .a(pci_target_unit_fifos_pcir_data_in_163), .b(FE_OFN1016_n_2053), .o(g65823_db) );
in01s01 TIMEBOOST_cell_8841 ( .a(TIMEBOOST_net_977), .o(TIMEBOOST_net_978) );
in01s01 g65824_u0 ( .a(FE_OFN1043_n_2037), .o(g65824_sb) );
na02s01 TIMEBOOST_cell_43330 ( .a(TIMEBOOST_net_13903), .b(g62611_sb), .o(n_6334) );
na02s02 TIMEBOOST_cell_45000 ( .a(TIMEBOOST_net_14738), .b(g64099_db), .o(n_4056) );
na02s02 TIMEBOOST_cell_40600 ( .a(TIMEBOOST_net_12538), .b(g62405_sb), .o(n_6789) );
in01s01 g65825_u0 ( .a(FE_OFN1044_n_2037), .o(g65825_sb) );
na02s01 g65825_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__Q), .b(g65825_sb), .o(g65825_da) );
na02s01 g65825_u2 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(FE_OFN1044_n_2037), .o(g65825_db) );
na02m02 TIMEBOOST_cell_44411 ( .a(n_9131), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__Q), .o(TIMEBOOST_net_14444) );
in01s01 g65826_u0 ( .a(FE_OFN1043_n_2037), .o(g65826_sb) );
na02s01 TIMEBOOST_cell_16017 ( .a(TIMEBOOST_net_3265), .b(n_2512), .o(n_2513) );
in01s01 TIMEBOOST_cell_8842 ( .a(conf_wb_err_addr_in_946), .o(TIMEBOOST_net_979) );
na02m02 TIMEBOOST_cell_43001 ( .a(n_4681), .b(n_3087), .o(TIMEBOOST_net_13739) );
in01s01 g65827_u0 ( .a(FE_OFN1043_n_2037), .o(g65827_sb) );
na02s01 g65827_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__Q), .b(g65827_sb), .o(g65827_da) );
na02s01 g65827_u2 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(FE_OFN1043_n_2037), .o(g65827_db) );
na02s01 g65827_u3 ( .a(g65827_da), .b(g65827_db), .o(n_1889) );
in01s01 g65828_u0 ( .a(FE_OFN1044_n_2037), .o(g65828_sb) );
na02s02 TIMEBOOST_cell_45001 ( .a(n_1702), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__Q), .o(TIMEBOOST_net_14739) );
na02s01 TIMEBOOST_cell_39561 ( .a(n_7078), .b(wishbone_slave_unit_pci_initiator_if_read_count_1_), .o(TIMEBOOST_net_12019) );
na02s02 TIMEBOOST_cell_40328 ( .a(TIMEBOOST_net_12402), .b(g64866_sb), .o(n_3714) );
in01s01 g65829_u0 ( .a(FE_OFN1043_n_2037), .o(g65829_sb) );
na02s01 TIMEBOOST_cell_42681 ( .a(n_3777), .b(g64770_sb), .o(TIMEBOOST_net_13579) );
in01s01 TIMEBOOST_cell_8844 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_), .o(TIMEBOOST_net_981) );
na02s01 TIMEBOOST_cell_30744 ( .a(pci_ad_i_27_), .b(parchk_pci_ad_reg_in_1231), .o(TIMEBOOST_net_9283) );
in01s01 g65830_u0 ( .a(FE_OFN1044_n_2037), .o(g65830_sb) );
na03s02 TIMEBOOST_cell_43331 ( .a(n_3710), .b(FE_OFN1274_n_4096), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__Q), .o(TIMEBOOST_net_13904) );
in01s01 TIMEBOOST_cell_8846 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_), .o(TIMEBOOST_net_983) );
na02f02 TIMEBOOST_cell_41224 ( .a(TIMEBOOST_net_12850), .b(g57272_sb), .o(n_10414) );
in01s01 g65831_u0 ( .a(FE_OFN1043_n_2037), .o(g65831_sb) );
na02s02 TIMEBOOST_cell_45038 ( .a(TIMEBOOST_net_14757), .b(FE_OFN720_n_8060), .o(TIMEBOOST_net_11247) );
in01s01 TIMEBOOST_cell_8848 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_), .o(TIMEBOOST_net_985) );
na02s01 TIMEBOOST_cell_18679 ( .a(TIMEBOOST_net_4596), .b(g62814_sb), .o(n_5349) );
in01s01 g65832_u0 ( .a(FE_OFN1044_n_2037), .o(g65832_sb) );
na02s01 TIMEBOOST_cell_43332 ( .a(TIMEBOOST_net_13904), .b(g62545_sb), .o(n_6477) );
in01s01 TIMEBOOST_cell_8850 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_), .o(TIMEBOOST_net_987) );
na02s01 TIMEBOOST_cell_18683 ( .a(TIMEBOOST_net_4598), .b(g63115_sb), .o(n_5025) );
in01s01 g65833_u0 ( .a(FE_OFN1044_n_2037), .o(g65833_sb) );
na02m02 TIMEBOOST_cell_44401 ( .a(n_9545), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__Q), .o(TIMEBOOST_net_14439) );
in01s01 TIMEBOOST_cell_8852 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_), .o(TIMEBOOST_net_989) );
na02s01 TIMEBOOST_cell_38528 ( .a(TIMEBOOST_net_11502), .b(g62041_sb), .o(n_7773) );
in01s01 g65834_u0 ( .a(FE_OFN1043_n_2037), .o(g65834_sb) );
na02f02 TIMEBOOST_cell_42220 ( .a(TIMEBOOST_net_13348), .b(FE_OFN1398_n_8567), .o(TIMEBOOST_net_12303) );
in01s01 TIMEBOOST_cell_8854 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_), .o(TIMEBOOST_net_991) );
na03s02 TIMEBOOST_cell_919 ( .a(n_7215), .b(g59381_sb), .c(g59381_db), .o(n_7677) );
in01s01 g65835_u0 ( .a(n_2299), .o(g65835_sb) );
na02s01 TIMEBOOST_cell_31264 ( .a(pci_target_unit_fifos_pcir_data_in_185), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__Q), .o(TIMEBOOST_net_9543) );
na02f02 TIMEBOOST_cell_32611 ( .a(FE_OFN1552_n_12104), .b(TIMEBOOST_net_10216), .o(TIMEBOOST_net_6493) );
na04s02 TIMEBOOST_cell_34181 ( .a(g64206_da), .b(g64206_db), .c(g62852_sb), .d(g62852_db), .o(n_5265) );
in01s01 g65836_u0 ( .a(FE_OFN1041_n_2037), .o(g65836_sb) );
na02s01 TIMEBOOST_cell_39183 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__Q), .b(g65904_sb), .o(TIMEBOOST_net_11830) );
na02s01 g65836_u2 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(FE_OFN1041_n_2037), .o(g65836_db) );
no02f04 TIMEBOOST_cell_38782 ( .a(TIMEBOOST_net_11629), .b(FE_RN_49_0), .o(TIMEBOOST_net_3038) );
in01s01 g65837_u0 ( .a(FE_OFN1043_n_2037), .o(g65837_sb) );
na02m02 TIMEBOOST_cell_42221 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__Q), .b(n_9727), .o(TIMEBOOST_net_13349) );
in01s01 TIMEBOOST_cell_8856 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_), .o(TIMEBOOST_net_993) );
na02s01 TIMEBOOST_cell_18817 ( .a(TIMEBOOST_net_4665), .b(g59371_sb), .o(n_7692) );
in01s01 g65838_u0 ( .a(FE_OFN1042_n_2037), .o(g65838_sb) );
na02s01 TIMEBOOST_cell_17540 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__Q), .b(g64326_sb), .o(TIMEBOOST_net_4027) );
na02s01 g65838_u2 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(FE_OFN1042_n_2037), .o(g65838_db) );
na03s02 TIMEBOOST_cell_38215 ( .a(TIMEBOOST_net_4009), .b(g64173_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__Q), .o(TIMEBOOST_net_11346) );
in01s01 g65839_u0 ( .a(FE_OFN1041_n_2037), .o(g65839_sb) );
na02s01 g65839_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__Q), .b(g65839_sb), .o(g65839_da) );
na02s01 g65839_u2 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(FE_OFN1041_n_2037), .o(g65839_db) );
na02f02 TIMEBOOST_cell_38909 ( .a(n_3358), .b(wbu_addr_in_263), .o(TIMEBOOST_net_11693) );
in01s01 g65840_u0 ( .a(FE_OFN1041_n_2037), .o(g65840_sb) );
na02f02 TIMEBOOST_cell_44668 ( .a(TIMEBOOST_net_14572), .b(FE_OFN1402_n_8567), .o(TIMEBOOST_net_12779) );
na02s01 g65840_u2 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(FE_OFN1041_n_2037), .o(g65840_db) );
na02f02 TIMEBOOST_cell_38804 ( .a(TIMEBOOST_net_11640), .b(g57291_sb), .o(n_11462) );
in01s01 g65841_u0 ( .a(FE_OFN1042_n_2037), .o(g65841_sb) );
na02f02 TIMEBOOST_cell_44122 ( .a(TIMEBOOST_net_14299), .b(FE_OFN1409_n_8567), .o(TIMEBOOST_net_12926) );
na02s02 TIMEBOOST_cell_45180 ( .a(TIMEBOOST_net_14828), .b(FE_OFN1224_n_6391), .o(TIMEBOOST_net_13252) );
na02s01 TIMEBOOST_cell_39208 ( .a(TIMEBOOST_net_11842), .b(n_1574), .o(TIMEBOOST_net_11454) );
in01s01 g65842_u0 ( .a(FE_OFN1041_n_2037), .o(g65842_sb) );
na02s01 g65842_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__Q), .b(g65842_sb), .o(g65842_da) );
na02s01 g65842_u2 ( .a(pci_target_unit_fifos_pcir_data_in_188), .b(FE_OFN1041_n_2037), .o(g65842_db) );
na02s02 TIMEBOOST_cell_44428 ( .a(TIMEBOOST_net_14452), .b(FE_OFN1306_n_13124), .o(TIMEBOOST_net_13427) );
in01s01 g65843_u0 ( .a(FE_OFN1042_n_2037), .o(g65843_sb) );
na02s01 TIMEBOOST_cell_17546 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__Q), .b(g64231_sb), .o(TIMEBOOST_net_4030) );
na02s01 g65843_u2 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(FE_OFN1042_n_2037), .o(g65843_db) );
na03s02 TIMEBOOST_cell_38395 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__Q), .b(FE_OFN1126_g64577_p), .c(n_3589), .o(TIMEBOOST_net_11436) );
in01s01 g65844_u0 ( .a(FE_OFN1042_n_2037), .o(g65844_sb) );
na02s01 g65844_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__Q), .b(g65844_sb), .o(g65844_da) );
na02s01 g65844_u2 ( .a(pci_target_unit_fifos_pcir_data_in_163), .b(FE_OFN1042_n_2037), .o(g65844_db) );
na02f02 TIMEBOOST_cell_37074 ( .a(TIMEBOOST_net_10775), .b(FE_OFN1586_n_13736), .o(n_14415) );
in01s01 g65845_u0 ( .a(FE_OFN1041_n_2037), .o(g65845_sb) );
na02s01 TIMEBOOST_cell_17548 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q), .b(g64235_sb), .o(TIMEBOOST_net_4031) );
na02s01 g65845_u2 ( .a(pci_target_unit_fifos_pcir_data_in_164), .b(FE_OFN1041_n_2037), .o(g65845_db) );
na03s02 TIMEBOOST_cell_38347 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__Q), .b(FE_OFN1132_g64577_p), .c(n_3823), .o(TIMEBOOST_net_11412) );
in01s01 g65846_u0 ( .a(FE_OFN1044_n_2037), .o(g65846_sb) );
na02m02 TIMEBOOST_cell_22382 ( .a(g57797_da), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_6448) );
in01s01 TIMEBOOST_cell_8858 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_), .o(TIMEBOOST_net_995) );
na02s01 TIMEBOOST_cell_38530 ( .a(TIMEBOOST_net_11503), .b(g62056_sb), .o(n_7753) );
in01s01 g65847_u0 ( .a(FE_OFN946_n_2248), .o(g65847_sb) );
na02f02 TIMEBOOST_cell_45548 ( .a(TIMEBOOST_net_15012), .b(FE_OFN1577_n_12028), .o(n_12735) );
na02s01 g65847_u2 ( .a(pci_target_unit_fifos_pcir_data_in), .b(FE_OFN946_n_2248), .o(g65847_db) );
na02m02 TIMEBOOST_cell_32610 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__Q), .o(TIMEBOOST_net_10216) );
in01s01 g65848_u0 ( .a(FE_OFN948_n_2248), .o(g65848_sb) );
na02m02 TIMEBOOST_cell_9924 ( .a(FE_OFN2069_n_15978), .b(conf_wb_err_addr_in_958), .o(TIMEBOOST_net_1529) );
na02s01 TIMEBOOST_cell_17960 ( .a(n_4493), .b(FE_OFN1680_n_4655), .o(TIMEBOOST_net_4237) );
na02m02 TIMEBOOST_cell_9925 ( .a(FE_OFN1145_n_15261), .b(TIMEBOOST_net_1529), .o(TIMEBOOST_net_584) );
in01s01 g65849_u0 ( .a(FE_OFN945_n_2248), .o(g65849_sb) );
na02f02 TIMEBOOST_cell_40400 ( .a(TIMEBOOST_net_12438), .b(n_3335), .o(TIMEBOOST_net_2408) );
na02s01 TIMEBOOST_cell_39221 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(g65744_sb), .o(TIMEBOOST_net_11849) );
na02m02 TIMEBOOST_cell_39410 ( .a(TIMEBOOST_net_11943), .b(g61831_db), .o(n_5642) );
in01s01 g65850_u0 ( .a(FE_OFN946_n_2248), .o(g65850_sb) );
na02f02 TIMEBOOST_cell_41218 ( .a(TIMEBOOST_net_12847), .b(g57208_sb), .o(n_11548) );
na02f02 TIMEBOOST_cell_43768 ( .a(TIMEBOOST_net_14122), .b(FE_OFN1417_n_8567), .o(TIMEBOOST_net_12944) );
na02m02 TIMEBOOST_cell_32608 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__Q), .o(TIMEBOOST_net_10215) );
in01s01 g65851_u0 ( .a(FE_OFN959_n_2299), .o(g65851_sb) );
na02s02 TIMEBOOST_cell_38096 ( .a(TIMEBOOST_net_11286), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_4712) );
na02s01 g65851_u2 ( .a(pci_target_unit_fifos_pcir_data_in_167), .b(FE_OFN959_n_2299), .o(g65851_db) );
na02s01 TIMEBOOST_cell_32066 ( .a(configuration_pci_err_data_516), .b(wbm_dat_o_15_), .o(TIMEBOOST_net_9944) );
in01s01 g65852_u0 ( .a(FE_OFN946_n_2248), .o(g65852_sb) );
na02f02 TIMEBOOST_cell_41016 ( .a(TIMEBOOST_net_12746), .b(g57422_sb), .o(n_10362) );
na02s01 g65852_u2 ( .a(pci_target_unit_fifos_pcir_data_in_175), .b(FE_OFN946_n_2248), .o(g65852_db) );
na02f02 TIMEBOOST_cell_32607 ( .a(FE_OFN1551_n_12104), .b(TIMEBOOST_net_10214), .o(TIMEBOOST_net_6495) );
in01s01 g65853_u0 ( .a(FE_OFN945_n_2248), .o(g65853_sb) );
na02f02 TIMEBOOST_cell_42266 ( .a(TIMEBOOST_net_13371), .b(FE_OFN1390_n_8567), .o(TIMEBOOST_net_12309) );
na02s01 g65853_u2 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(FE_OFN945_n_2248), .o(g65853_db) );
no03f08 TIMEBOOST_cell_32936 ( .a(FE_RN_428_0), .b(FE_RN_430_0), .c(FE_RN_764_0), .o(FE_RN_462_0) );
in01s01 g65854_u0 ( .a(FE_OFN2111_n_2248), .o(g65854_sb) );
na02s01 g65854_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__Q), .b(g65854_sb), .o(g65854_da) );
na02s01 g65854_u2 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(FE_OFN2111_n_2248), .o(g65854_db) );
na02s02 g65854_u3 ( .a(g65854_da), .b(g65854_db), .o(n_1702) );
in01s01 g65855_u0 ( .a(FE_OFN1017_n_2053), .o(g65855_sb) );
na02m02 TIMEBOOST_cell_44501 ( .a(n_9883), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__Q), .o(TIMEBOOST_net_14489) );
na02s01 g65855_u2 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(FE_OFN1017_n_2053), .o(g65855_db) );
na02s01 TIMEBOOST_cell_41814 ( .a(TIMEBOOST_net_13145), .b(g65335_db), .o(n_3551) );
in01s01 g65856_u0 ( .a(FE_OFN948_n_2248), .o(g65856_sb) );
na02s02 TIMEBOOST_cell_40330 ( .a(TIMEBOOST_net_12403), .b(n_4447), .o(n_4290) );
na02s02 TIMEBOOST_cell_17962 ( .a(n_4442), .b(FE_OFN1680_n_4655), .o(TIMEBOOST_net_4238) );
na02f04 TIMEBOOST_cell_9927 ( .a(TIMEBOOST_net_1530), .b(n_7040), .o(FE_RN_267_0) );
in01s01 g65857_u0 ( .a(FE_OFN945_n_2248), .o(g65857_sb) );
no02f04 TIMEBOOST_cell_10133 ( .a(TIMEBOOST_net_1633), .b(n_4744), .o(n_5722) );
na02s01 TIMEBOOST_cell_40813 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__Q), .b(n_2029), .o(TIMEBOOST_net_12645) );
na02m02 TIMEBOOST_cell_39412 ( .a(TIMEBOOST_net_11944), .b(TIMEBOOST_net_489), .o(n_13495) );
in01s01 g65858_u0 ( .a(FE_OFN776_n_15366), .o(g65858_sb) );
na02s01 TIMEBOOST_cell_36645 ( .a(parchk_pci_ad_reg_in_1215), .b(g65813_sb), .o(TIMEBOOST_net_10561) );
na02s02 TIMEBOOST_cell_43267 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__Q), .b(n_4235), .o(TIMEBOOST_net_13872) );
na02s01 TIMEBOOST_cell_36543 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(g65741_sb), .o(TIMEBOOST_net_10510) );
in01s01 g65859_u0 ( .a(FE_OFN948_n_2248), .o(g65859_sb) );
na02s01 TIMEBOOST_cell_39321 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__Q), .b(FE_OFN1794_n_9904), .o(TIMEBOOST_net_11899) );
na02s01 TIMEBOOST_cell_17964 ( .a(n_4645), .b(FE_OFN1678_n_4655), .o(TIMEBOOST_net_4239) );
na02m02 TIMEBOOST_cell_38702 ( .a(TIMEBOOST_net_11589), .b(g62635_sb), .o(n_6281) );
in01s01 g65860_u0 ( .a(FE_OFN945_n_2248), .o(g65860_sb) );
na02s01 TIMEBOOST_cell_17272 ( .a(n_3755), .b(FE_OFN1640_n_4671), .o(TIMEBOOST_net_3893) );
na02s01 g65860_u2 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(FE_OFN945_n_2248), .o(g65860_db) );
na02f02 TIMEBOOST_cell_39089 ( .a(FE_OCPN1877_n_13903), .b(TIMEBOOST_net_10155), .o(TIMEBOOST_net_11783) );
in01s01 g65861_u0 ( .a(n_2299), .o(g65861_sb) );
na02m02 TIMEBOOST_cell_32606 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__Q), .o(TIMEBOOST_net_10214) );
na02s01 g65861_u2 ( .a(pci_target_unit_fifos_pcir_data_in), .b(n_2299), .o(g65861_db) );
na02s02 TIMEBOOST_cell_22251 ( .a(n_10225), .b(TIMEBOOST_net_6382), .o(n_11864) );
in01s01 g65862_u0 ( .a(FE_OFN948_n_2248), .o(g65862_sb) );
na02s02 g65862_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__Q), .b(g65862_sb), .o(g65862_da) );
na02s02 g65862_u2 ( .a(pci_target_unit_fifos_pcir_data_in_164), .b(FE_OFN948_n_2248), .o(g65862_db) );
na02s01 TIMEBOOST_cell_37206 ( .a(TIMEBOOST_net_10841), .b(g65692_db), .o(n_2206) );
in01s01 g65863_u0 ( .a(FE_OFN945_n_2248), .o(g65863_sb) );
na02s01 TIMEBOOST_cell_39414 ( .a(TIMEBOOST_net_11945), .b(n_1756), .o(n_8024) );
na02s02 TIMEBOOST_cell_45002 ( .a(TIMEBOOST_net_14739), .b(FE_OFN709_n_8232), .o(TIMEBOOST_net_11081) );
na02s02 TIMEBOOST_cell_17813 ( .a(TIMEBOOST_net_4163), .b(g61760_sb), .o(n_8293) );
na02f02 TIMEBOOST_cell_38904 ( .a(TIMEBOOST_net_11690), .b(FE_OFN2198_n_10256), .o(TIMEBOOST_net_10697) );
na02s02 TIMEBOOST_cell_18010 ( .a(pci_target_unit_fifos_pciw_cbe_in_153), .b(g64125_sb), .o(TIMEBOOST_net_4262) );
na02s01 TIMEBOOST_cell_37780 ( .a(TIMEBOOST_net_11128), .b(FE_OFN707_n_8119), .o(TIMEBOOST_net_4347) );
in01s01 g65865_u0 ( .a(FE_OFN945_n_2248), .o(g65865_sb) );
na02m02 TIMEBOOST_cell_41609 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_10__Q), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_13043) );
na02s01 g65865_u2 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(FE_OFN945_n_2248), .o(g65865_db) );
in01s01 TIMEBOOST_cell_32853 ( .a(TIMEBOOST_net_10354), .o(TIMEBOOST_net_10353) );
in01s01 g65866_u0 ( .a(FE_OFN946_n_2248), .o(g65866_sb) );
na02s02 TIMEBOOST_cell_22247 ( .a(n_10250), .b(TIMEBOOST_net_6380), .o(n_11868) );
na02s01 g65866_u2 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(FE_OFN946_n_2248), .o(g65866_db) );
na02f02 TIMEBOOST_cell_32605 ( .a(FE_OFN1553_n_12104), .b(TIMEBOOST_net_10213), .o(TIMEBOOST_net_6494) );
in01s01 g65867_u0 ( .a(FE_OFN945_n_2248), .o(g65867_sb) );
na02s01 TIMEBOOST_cell_17274 ( .a(n_3747), .b(FE_OFN1642_n_4671), .o(TIMEBOOST_net_3894) );
na02s01 g65867_u2 ( .a(pci_target_unit_fifos_pcir_data_in_174), .b(FE_OFN945_n_2248), .o(g65867_db) );
na02s02 TIMEBOOST_cell_17275 ( .a(TIMEBOOST_net_3894), .b(g65380_da), .o(n_3527) );
in01s01 g65868_u0 ( .a(FE_OFN1016_n_2053), .o(g65868_sb) );
na02f02 TIMEBOOST_cell_21605 ( .a(TIMEBOOST_net_6059), .b(g57582_sb), .o(n_11167) );
na02s01 g65868_u2 ( .a(pci_target_unit_fifos_pcir_data_in_167), .b(FE_OFN1016_n_2053), .o(g65868_db) );
na02s01 TIMEBOOST_cell_40332 ( .a(TIMEBOOST_net_12404), .b(g65055_sb), .o(TIMEBOOST_net_237) );
in01s01 g65869_u0 ( .a(FE_OFN1041_n_2037), .o(g65869_sb) );
na02s01 g65869_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__Q), .b(g65869_sb), .o(g65869_da) );
na02s01 g65869_u2 ( .a(pci_target_unit_fifos_pcir_data_in_167), .b(FE_OFN1041_n_2037), .o(g65869_db) );
na02s02 TIMEBOOST_cell_44429 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_768), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_3__Q), .o(TIMEBOOST_net_14453) );
in01s01 g65870_u0 ( .a(n_2299), .o(g65870_sb) );
na02f02 TIMEBOOST_cell_40984 ( .a(TIMEBOOST_net_12730), .b(g57236_sb), .o(n_10432) );
na02s01 g65870_u2 ( .a(pci_target_unit_fifos_pcir_data_in_178), .b(n_2299), .o(g65870_db) );
na02s02 TIMEBOOST_cell_41764 ( .a(TIMEBOOST_net_13120), .b(g58372_db), .o(n_9457) );
in01s01 g65871_u0 ( .a(FE_OFN644_n_4677), .o(g65871_sb) );
na02f02 TIMEBOOST_cell_44680 ( .a(TIMEBOOST_net_14578), .b(g57426_sb), .o(n_11309) );
na02s01 g65871_u2 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(FE_OFN644_n_4677), .o(g65871_db) );
na02s02 TIMEBOOST_cell_17073 ( .a(TIMEBOOST_net_3793), .b(g57909_sb), .o(n_9906) );
in01s01 g65872_u0 ( .a(FE_OFN1042_n_2037), .o(g65872_sb) );
na02s01 g65872_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__Q), .b(g65872_sb), .o(g65872_da) );
na02s01 g65872_u2 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(FE_OFN1042_n_2037), .o(g65872_db) );
na02f02 TIMEBOOST_cell_37076 ( .a(TIMEBOOST_net_10776), .b(FE_OFN1587_n_13736), .o(g53288_p) );
in01s01 g65873_u0 ( .a(n_4490), .o(g65873_sb) );
na02s02 TIMEBOOST_cell_40782 ( .a(TIMEBOOST_net_12629), .b(g62529_sb), .o(n_6516) );
na02s01 g65873_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__Q), .b(n_4490), .o(g65873_db) );
na02s02 TIMEBOOST_cell_32065 ( .a(TIMEBOOST_net_9943), .b(FE_OFN1179_n_3476), .o(TIMEBOOST_net_4931) );
in01s01 g65874_u0 ( .a(FE_OFN1042_n_2037), .o(g65874_sb) );
na02f02 TIMEBOOST_cell_41680 ( .a(TIMEBOOST_net_13078), .b(n_14833), .o(n_14897) );
na02s01 g65874_u2 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(FE_OFN1042_n_2037), .o(g65874_db) );
na02s02 TIMEBOOST_cell_17551 ( .a(TIMEBOOST_net_4032), .b(g58375_sb), .o(n_9454) );
in01s01 g65875_u0 ( .a(n_2299), .o(g65875_sb) );
na02f02 TIMEBOOST_cell_45549 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__Q), .b(FE_OCPN1825_n_12030), .o(TIMEBOOST_net_15013) );
na02s01 g65875_u2 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(n_2299), .o(g65875_db) );
na02f02 TIMEBOOST_cell_40952 ( .a(TIMEBOOST_net_12714), .b(g57548_sb), .o(n_10304) );
in01s01 g65876_u0 ( .a(FE_OFN1015_n_2053), .o(g65876_sb) );
na02s01 TIMEBOOST_cell_38532 ( .a(TIMEBOOST_net_11504), .b(g62060_sb), .o(n_7750) );
na02s01 TIMEBOOST_cell_37255 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__Q), .b(n_3749), .o(TIMEBOOST_net_10866) );
na02s01 TIMEBOOST_cell_17409 ( .a(TIMEBOOST_net_3961), .b(g64256_db), .o(n_3917) );
in01s01 g65877_u0 ( .a(FE_OFN1016_n_2053), .o(g65877_sb) );
na02s01 TIMEBOOST_cell_40333 ( .a(n_3785), .b(g64756_db), .o(TIMEBOOST_net_12405) );
na02s01 g65877_u2 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(FE_OFN1015_n_2053), .o(g65877_db) );
na02s02 TIMEBOOST_cell_40334 ( .a(TIMEBOOST_net_12405), .b(g64756_sb), .o(n_3788) );
in01s01 g65878_u0 ( .a(FE_OFN959_n_2299), .o(g65878_sb) );
na02s02 TIMEBOOST_cell_44417 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_793), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_28__Q), .o(TIMEBOOST_net_14447) );
na02m02 TIMEBOOST_cell_32604 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q), .o(TIMEBOOST_net_10213) );
na02s01 TIMEBOOST_cell_9257 ( .a(TIMEBOOST_net_1195), .b(g65685_db), .o(n_2210) );
in01s01 g65879_u0 ( .a(n_4669), .o(g65879_sb) );
na02s01 g65879_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__Q), .b(g65879_sb), .o(g65879_da) );
na02s01 g65879_u2 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(n_4669), .o(g65879_db) );
na02s01 g65879_u3 ( .a(g65879_da), .b(g65879_db), .o(n_2181) );
in01s01 g65880_u0 ( .a(FE_OFN1017_n_2053), .o(g65880_sb) );
na02s01 TIMEBOOST_cell_40335 ( .a(n_3777), .b(g65075_db), .o(TIMEBOOST_net_12406) );
na02s01 g65880_u2 ( .a(pci_target_unit_fifos_pcir_data_in_165), .b(FE_OFN1017_n_2053), .o(g65880_db) );
na02s02 TIMEBOOST_cell_40336 ( .a(TIMEBOOST_net_12406), .b(g65075_sb), .o(n_3604) );
in01s01 g65881_u0 ( .a(FE_OFN1016_n_2053), .o(g65881_sb) );
na02s01 TIMEBOOST_cell_40337 ( .a(n_3785), .b(g64889_db), .o(TIMEBOOST_net_12407) );
na02s01 g65881_u2 ( .a(pci_target_unit_fifos_pcir_data_in_164), .b(FE_OFN1016_n_2053), .o(g65881_db) );
na02s02 TIMEBOOST_cell_40338 ( .a(TIMEBOOST_net_12407), .b(g64889_sb), .o(n_3701) );
in01s01 g65882_u0 ( .a(FE_OFN2113_n_2053), .o(g65882_sb) );
na02m02 TIMEBOOST_cell_10216 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__Q), .b(n_13447), .o(TIMEBOOST_net_1675) );
na02s01 TIMEBOOST_cell_18226 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_387), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_4370) );
na02m02 TIMEBOOST_cell_10217 ( .a(FE_OFN1148_n_13249), .b(TIMEBOOST_net_1675), .o(TIMEBOOST_net_496) );
in01s01 g65883_u0 ( .a(FE_OFN651_n_4508), .o(g65883_sb) );
na02s01 TIMEBOOST_cell_41866 ( .a(TIMEBOOST_net_13171), .b(g61918_db), .o(n_7985) );
na02s01 g65883_u2 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(FE_OFN651_n_4508), .o(g65883_db) );
no02f10 TIMEBOOST_cell_36270 ( .a(TIMEBOOST_net_10373), .b(n_15210), .o(n_15729) );
in01s01 g65884_u0 ( .a(FE_OFN2113_n_2053), .o(g65884_sb) );
na02s01 TIMEBOOST_cell_10218 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_4_), .b(n_6986), .o(TIMEBOOST_net_1676) );
na02s02 TIMEBOOST_cell_43632 ( .a(TIMEBOOST_net_14054), .b(FE_OFN1261_n_4143), .o(TIMEBOOST_net_12093) );
na02s01 TIMEBOOST_cell_10219 ( .a(TIMEBOOST_net_1676), .b(n_4662), .o(TIMEBOOST_net_581) );
na02m02 TIMEBOOST_cell_42347 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__10__Q), .b(n_9503), .o(TIMEBOOST_net_13412) );
na02s01 TIMEBOOST_cell_39223 ( .a(pci_target_unit_fifos_pcir_data_in_178), .b(g65800_sb), .o(TIMEBOOST_net_11850) );
na02s02 TIMEBOOST_cell_43100 ( .a(TIMEBOOST_net_13788), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_12590) );
na02s01 TIMEBOOST_cell_42708 ( .a(TIMEBOOST_net_13592), .b(g65952_db), .o(n_1845) );
na02s01 TIMEBOOST_cell_39225 ( .a(pci_target_unit_fifos_pcir_data_in_163), .b(g65730_sb), .o(TIMEBOOST_net_11851) );
na02s01 TIMEBOOST_cell_38534 ( .a(TIMEBOOST_net_11505), .b(g62054_sb), .o(n_7755) );
in01s01 g65887_u0 ( .a(FE_OFN1041_n_2037), .o(g65887_sb) );
na02s01 TIMEBOOST_cell_17552 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__Q), .b(g64297_sb), .o(TIMEBOOST_net_4033) );
na02s01 g65887_u2 ( .a(pci_target_unit_fifos_pcir_data_in_185), .b(FE_OFN1041_n_2037), .o(g65887_db) );
na02f02 TIMEBOOST_cell_44196 ( .a(TIMEBOOST_net_14336), .b(FE_OFN1420_n_8567), .o(TIMEBOOST_net_12743) );
in01s01 g65888_u0 ( .a(FE_OFN682_n_4460), .o(g65888_sb) );
na03f02 TIMEBOOST_cell_36188 ( .a(n_12088), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__Q), .c(n_11823), .o(n_12513) );
na02s01 g65888_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__Q), .b(FE_OFN682_n_4460), .o(g65888_db) );
na02s02 TIMEBOOST_cell_40340 ( .a(TIMEBOOST_net_12408), .b(g65079_sb), .o(n_3601) );
in01s01 g65889_u0 ( .a(FE_OFN634_n_4454), .o(g65889_sb) );
na02s01 TIMEBOOST_cell_32064 ( .a(configuration_pci_err_addr_489), .b(wbm_adr_o_19_), .o(TIMEBOOST_net_9943) );
na02s01 g65889_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__Q), .b(FE_OFN634_n_4454), .o(g65889_db) );
na02s02 TIMEBOOST_cell_32063 ( .a(TIMEBOOST_net_9942), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_4927) );
in01s01 g65890_u0 ( .a(FE_OFN1041_n_2037), .o(g65890_sb) );
na02s02 TIMEBOOST_cell_17554 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__Q), .b(g64300_sb), .o(TIMEBOOST_net_4034) );
na02s01 g65890_u2 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(FE_OFN1041_n_2037), .o(g65890_db) );
na02s02 TIMEBOOST_cell_17555 ( .a(TIMEBOOST_net_4034), .b(g64300_db), .o(n_3875) );
in01s01 g65891_u0 ( .a(FE_OFN946_n_2248), .o(g65891_sb) );
na02f02 TIMEBOOST_cell_41220 ( .a(TIMEBOOST_net_12848), .b(g57139_sb), .o(n_11610) );
na02s01 g65891_u2 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(FE_OFN946_n_2248), .o(g65891_db) );
na02m02 TIMEBOOST_cell_32602 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q), .o(TIMEBOOST_net_10212) );
in01s01 g65892_u0 ( .a(FE_OFN775_n_15366), .o(g65892_sb) );
na02s02 TIMEBOOST_cell_45691 ( .a(n_4260), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__Q), .o(TIMEBOOST_net_15084) );
na03f02 TIMEBOOST_cell_36216 ( .a(FE_OCPN1866_n_12377), .b(TIMEBOOST_net_10302), .c(FE_OFN1756_n_12681), .o(n_12673) );
na02s01 TIMEBOOST_cell_42892 ( .a(TIMEBOOST_net_13684), .b(FE_OFN1690_n_9528), .o(TIMEBOOST_net_11188) );
in01s02 g65893_u0 ( .a(FE_OFN775_n_15366), .o(g65893_sb) );
na02s01 TIMEBOOST_cell_36358 ( .a(TIMEBOOST_net_10417), .b(FE_OFN2094_n_2520), .o(n_2519) );
na02s01 g65893_u2 ( .a(pci_target_unit_del_sync_addr_in_225), .b(FE_OFN776_n_15366), .o(g65893_db) );
na02s01 TIMEBOOST_cell_37582 ( .a(TIMEBOOST_net_11029), .b(g61718_sb), .o(n_8389) );
in01s01 g65894_u0 ( .a(FE_OFN1041_n_2037), .o(g65894_sb) );
na02s01 TIMEBOOST_cell_39209 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__Q), .b(n_8176), .o(TIMEBOOST_net_11843) );
na02s01 g65894_u2 ( .a(pci_target_unit_fifos_pcir_data_in_187), .b(FE_OFN1041_n_2037), .o(g65894_db) );
na02m02 TIMEBOOST_cell_38784 ( .a(n_16332), .b(TIMEBOOST_net_11630), .o(g58582_p) );
na02s01 TIMEBOOST_cell_39213 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__Q), .b(n_8407), .o(TIMEBOOST_net_11845) );
na02f02 TIMEBOOST_cell_45550 ( .a(TIMEBOOST_net_15013), .b(n_11822), .o(n_12510) );
na02m02 TIMEBOOST_cell_10147 ( .a(FE_OFN1151_n_13249), .b(TIMEBOOST_net_1640), .o(TIMEBOOST_net_498) );
in01s01 g65896_u0 ( .a(FE_OFN1015_n_2053), .o(g65896_sb) );
na02s02 TIMEBOOST_cell_40339 ( .a(n_3777), .b(g65079_db), .o(TIMEBOOST_net_12408) );
na02s01 g65896_u2 ( .a(pci_target_unit_fifos_pcir_data_in_173), .b(FE_OFN1015_n_2053), .o(g65896_db) );
na02s02 TIMEBOOST_cell_40342 ( .a(TIMEBOOST_net_12409), .b(g64999_sb), .o(n_3642) );
in01s01 g65897_u0 ( .a(FE_OFN1678_n_4655), .o(g65897_sb) );
na02f02 TIMEBOOST_cell_38785 ( .a(n_9627), .b(g57300_sb), .o(TIMEBOOST_net_11631) );
na02s02 TIMEBOOST_cell_45181 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__Q), .b(n_4366), .o(TIMEBOOST_net_14829) );
na02f02 TIMEBOOST_cell_38906 ( .a(TIMEBOOST_net_11691), .b(FE_OFN2200_n_10256), .o(TIMEBOOST_net_10705) );
na02s01 TIMEBOOST_cell_37782 ( .a(TIMEBOOST_net_11129), .b(FE_OFN701_n_7845), .o(TIMEBOOST_net_4348) );
na02s02 TIMEBOOST_cell_18012 ( .a(pci_target_unit_fifos_pciw_addr_data_in_136), .b(g64112_sb), .o(TIMEBOOST_net_4263) );
na02s02 TIMEBOOST_cell_37784 ( .a(TIMEBOOST_net_11130), .b(FE_OFN699_n_7845), .o(TIMEBOOST_net_4345) );
in01s01 g65899_u0 ( .a(FE_OFN1042_n_2037), .o(g65899_sb) );
na02s01 TIMEBOOST_cell_17560 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__Q), .b(g64312_sb), .o(TIMEBOOST_net_4037) );
na02s01 TIMEBOOST_cell_37270 ( .a(TIMEBOOST_net_10873), .b(g65675_db), .o(n_2033) );
in01s01 g65900_u0 ( .a(FE_OFN948_n_2248), .o(g65900_sb) );
na03s02 TIMEBOOST_cell_43333 ( .a(n_4441), .b(FE_OFN1206_n_6356), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__Q), .o(TIMEBOOST_net_13905) );
na02s01 TIMEBOOST_cell_17966 ( .a(pci_target_unit_fifos_pciw_addr_data_in_147), .b(g64218_sb), .o(TIMEBOOST_net_4240) );
na02f02 TIMEBOOST_cell_44402 ( .a(TIMEBOOST_net_14439), .b(FE_OFN1414_n_8567), .o(TIMEBOOST_net_12778) );
in01s01 g65901_u0 ( .a(FE_OFN1044_n_2037), .o(g65901_sb) );
na02s01 g65901_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__Q), .b(g65901_sb), .o(g65901_da) );
na02s01 g65901_u2 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(FE_OFN1044_n_2037), .o(g65901_db) );
na02f02 TIMEBOOST_cell_43773 ( .a(n_9754), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__Q), .o(TIMEBOOST_net_14125) );
in01s01 g65902_u0 ( .a(FE_OFN946_n_2248), .o(g65902_sb) );
na02s01 g65902_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__Q), .b(g65902_sb), .o(g65902_da) );
na02s01 g65902_u2 ( .a(pci_target_unit_fifos_pcir_data_in_165), .b(FE_OFN946_n_2248), .o(g65902_db) );
na02f02 TIMEBOOST_cell_45551 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__Q), .b(n_12313), .o(TIMEBOOST_net_15014) );
in01s01 g65903_u0 ( .a(FE_OFN959_n_2299), .o(g65903_sb) );
na02s01 TIMEBOOST_cell_32062 ( .a(configuration_pci_err_cs_bit_464), .b(pci_target_unit_wishbone_master_bc_register_reg_1__Q), .o(TIMEBOOST_net_9942) );
na02s01 g65903_u2 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(FE_OFN959_n_2299), .o(g65903_db) );
na02s02 TIMEBOOST_cell_38098 ( .a(TIMEBOOST_net_11287), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_4707) );
in01s01 g65904_u0 ( .a(FE_OFN959_n_2299), .o(g65904_sb) );
na02s01 TIMEBOOST_cell_32060 ( .a(configuration_pci_err_data_510), .b(wbm_dat_o_9_), .o(TIMEBOOST_net_9941) );
na02s01 g65904_u2 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(FE_OFN959_n_2299), .o(g65904_db) );
na02s02 TIMEBOOST_cell_32059 ( .a(TIMEBOOST_net_9940), .b(FE_OFN1183_n_3476), .o(TIMEBOOST_net_4924) );
in01s01 g65905_u0 ( .a(FE_OFN912_n_4727), .o(g65905_sb) );
na02s01 TIMEBOOST_cell_39284 ( .a(TIMEBOOST_net_11880), .b(g65724_db), .o(n_1610) );
na02m02 TIMEBOOST_cell_30738 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_9__Q), .b(n_8831), .o(TIMEBOOST_net_9280) );
na02f02 TIMEBOOST_cell_39489 ( .a(n_17039), .b(n_2768), .o(TIMEBOOST_net_11983) );
in01s01 g65906_u0 ( .a(FE_OFN2113_n_2053), .o(g65906_sb) );
na02s02 TIMEBOOST_cell_45182 ( .a(TIMEBOOST_net_14829), .b(FE_OFN1295_n_4098), .o(TIMEBOOST_net_12591) );
na02s01 g65906_u2 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(FE_OFN2113_n_2053), .o(g65906_db) );
na02s01 TIMEBOOST_cell_40344 ( .a(TIMEBOOST_net_12410), .b(TIMEBOOST_net_3891), .o(n_3548) );
in01s01 g65907_u0 ( .a(n_2299), .o(g65907_sb) );
na02f02 TIMEBOOST_cell_40954 ( .a(TIMEBOOST_net_12715), .b(g57546_sb), .o(n_10308) );
na02s01 g65907_u2 ( .a(pci_target_unit_fifos_pcir_data_in_172), .b(n_2299), .o(g65907_db) );
na02f02 TIMEBOOST_cell_41222 ( .a(TIMEBOOST_net_12849), .b(g57273_sb), .o(n_11482) );
in01s01 g65908_u0 ( .a(FE_OFN1016_n_2053), .o(g65908_sb) );
na02s01 TIMEBOOST_cell_40343 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__Q), .b(g65340_sb), .o(TIMEBOOST_net_12410) );
na02s01 g65908_u2 ( .a(pci_target_unit_fifos_pcir_data_in_185), .b(FE_OFN1016_n_2053), .o(g65908_db) );
na02s01 TIMEBOOST_cell_40346 ( .a(TIMEBOOST_net_12411), .b(g61804_sb), .o(TIMEBOOST_net_12141) );
in01s01 g65909_u0 ( .a(FE_OFN1797_n_2299), .o(g65909_sb) );
na02m02 TIMEBOOST_cell_45801 ( .a(n_9524), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__Q), .o(TIMEBOOST_net_15139) );
na02s01 g65909_u2 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(FE_OFN1797_n_2299), .o(g65909_db) );
na02s01 TIMEBOOST_cell_40348 ( .a(TIMEBOOST_net_12412), .b(g61801_sb), .o(TIMEBOOST_net_12142) );
in01s01 g65910_u0 ( .a(FE_OFN1016_n_2053), .o(g65910_sb) );
na02s01 TIMEBOOST_cell_40347 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__Q), .b(n_8069), .o(TIMEBOOST_net_12412) );
na02s01 g65910_u2 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(FE_OFN1016_n_2053), .o(g65910_db) );
na02s01 TIMEBOOST_cell_40350 ( .a(TIMEBOOST_net_12413), .b(g61820_sb), .o(TIMEBOOST_net_12143) );
na02f02 TIMEBOOST_cell_42494 ( .a(TIMEBOOST_net_13485), .b(g57313_sb), .o(n_10401) );
na02s01 TIMEBOOST_cell_18014 ( .a(pci_target_unit_fifos_pciw_addr_data_in_144), .b(g64088_sb), .o(TIMEBOOST_net_4264) );
na02f02 TIMEBOOST_cell_37113 ( .a(FE_OFN1600_n_13995), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__Q), .o(TIMEBOOST_net_10795) );
in01s01 TIMEBOOST_cell_32852 ( .a(TIMEBOOST_net_10353), .o(TIMEBOOST_net_10334) );
na02s01 g65912_u2 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(FE_OFN945_n_2248), .o(g65912_db) );
na02s02 TIMEBOOST_cell_45692 ( .a(TIMEBOOST_net_15084), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_13305) );
in01s01 g65913_u0 ( .a(FE_OFN1015_n_2053), .o(g65913_sb) );
na02m01 TIMEBOOST_cell_8876 ( .a(n_288), .b(wbu_wb_init_complete_in), .o(TIMEBOOST_net_1005) );
na02s01 g65913_u2 ( .a(pci_target_unit_fifos_pcir_data_in_175), .b(FE_OFN1015_n_2053), .o(g65913_db) );
na02m01 TIMEBOOST_cell_8877 ( .a(TIMEBOOST_net_1005), .b(n_1432), .o(TIMEBOOST_net_256) );
in01s01 g65914_u0 ( .a(FE_OFN948_n_2248), .o(g65914_sb) );
na02s02 g65914_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__Q), .b(g65914_sb), .o(g65914_da) );
na02s02 g65914_u2 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(FE_OFN948_n_2248), .o(g65914_db) );
na02s01 TIMEBOOST_cell_37208 ( .a(TIMEBOOST_net_10842), .b(g65707_db), .o(n_2061) );
in01s01 g65915_u0 ( .a(FE_OFN1035_n_4732), .o(g65915_sb) );
na02s02 TIMEBOOST_cell_38704 ( .a(TIMEBOOST_net_11590), .b(g62486_sb), .o(n_6615) );
na02s01 g65915_u2 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(FE_OFN1035_n_4732), .o(g65915_db) );
na02s01 TIMEBOOST_cell_18175 ( .a(TIMEBOOST_net_4344), .b(g61888_sb), .o(n_8054) );
in01s01 g65916_u0 ( .a(FE_OFN1640_n_4671), .o(g65916_sb) );
na02s01 TIMEBOOST_cell_40352 ( .a(TIMEBOOST_net_12414), .b(g61808_sb), .o(TIMEBOOST_net_12140) );
na02s01 g65916_u2 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(FE_OFN1640_n_4671), .o(g65916_db) );
na02s02 TIMEBOOST_cell_40299 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__12__Q), .b(g64296_sb), .o(TIMEBOOST_net_12388) );
na02s01 TIMEBOOST_cell_39510 ( .a(TIMEBOOST_net_11993), .b(TIMEBOOST_net_9839), .o(n_4973) );
na02m02 TIMEBOOST_cell_42267 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q), .b(n_9080), .o(TIMEBOOST_net_13372) );
na02m04 TIMEBOOST_cell_45827 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_780), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_15__Q), .o(TIMEBOOST_net_15152) );
na02f02 TIMEBOOST_cell_41578 ( .a(TIMEBOOST_net_13027), .b(g57472_sb), .o(n_11262) );
na02s01 g65918_u2 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(FE_OFN945_n_2248), .o(g65918_db) );
na03s02 TIMEBOOST_cell_34252 ( .a(TIMEBOOST_net_9794), .b(FE_OFN1174_n_5592), .c(g62074_sb), .o(n_5637) );
in01s01 g65919_u0 ( .a(FE_OFN1017_n_2053), .o(g65919_sb) );
na02s01 g65919_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__Q), .b(g65919_sb), .o(g65919_da) );
na02s01 g65919_u2 ( .a(pci_target_unit_fifos_pcir_data_in_174), .b(FE_OFN1015_n_2053), .o(g65919_db) );
na02s01 g65919_u3 ( .a(g65919_da), .b(g65919_db), .o(n_1851) );
in01s01 g65920_u0 ( .a(FE_OFN948_n_2248), .o(g65920_sb) );
na02f02 TIMEBOOST_cell_44194 ( .a(TIMEBOOST_net_14335), .b(FE_OFN1416_n_8567), .o(TIMEBOOST_net_12744) );
na02s01 TIMEBOOST_cell_17968 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(g64212_sb), .o(TIMEBOOST_net_4241) );
na02s01 TIMEBOOST_cell_38536 ( .a(TIMEBOOST_net_11506), .b(g62055_sb), .o(n_7754) );
in01s01 g65921_u0 ( .a(FE_OFN661_n_4392), .o(g65921_sb) );
na02s01 TIMEBOOST_cell_31288 ( .a(configuration_wb_err_data_594), .b(parchk_pci_ad_out_in_1191), .o(TIMEBOOST_net_9555) );
na02s01 g65921_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__Q), .b(FE_OFN661_n_4392), .o(g65921_db) );
na02f02 TIMEBOOST_cell_38908 ( .a(TIMEBOOST_net_11692), .b(FE_OFN2200_n_10256), .o(TIMEBOOST_net_10699) );
na02s01 TIMEBOOST_cell_45734 ( .a(TIMEBOOST_net_15105), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_13227) );
na02s01 TIMEBOOST_cell_18177 ( .a(TIMEBOOST_net_4345), .b(g61890_sb), .o(n_8049) );
in01s01 g65923_u0 ( .a(FE_OFN946_n_2248), .o(g65923_sb) );
na02m02 TIMEBOOST_cell_32600 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__Q), .o(TIMEBOOST_net_10211) );
na02s01 g65923_u2 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(FE_OFN946_n_2248), .o(g65923_db) );
na02f02 TIMEBOOST_cell_32599 ( .a(FE_OFN1553_n_12104), .b(TIMEBOOST_net_10210), .o(TIMEBOOST_net_6492) );
in01s01 g65924_u0 ( .a(FE_OFN1043_n_2037), .o(g65924_sb) );
na02s01 g65924_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__Q), .b(g65924_sb), .o(g65924_da) );
na02s01 g65924_u2 ( .a(pci_target_unit_fifos_pcir_data_in_178), .b(FE_OFN1043_n_2037), .o(g65924_db) );
na02s01 g65924_u3 ( .a(g65924_da), .b(g65924_db), .o(n_1756) );
na02s02 TIMEBOOST_cell_44430 ( .a(TIMEBOOST_net_14453), .b(FE_OFN1306_n_13124), .o(TIMEBOOST_net_13422) );
na02s01 g65925_u2 ( .a(pci_target_unit_del_sync_addr_in_234), .b(FE_OFN775_n_15366), .o(g65925_db) );
na02s02 TIMEBOOST_cell_38712 ( .a(TIMEBOOST_net_11594), .b(g62758_sb), .o(n_6123) );
na03s02 TIMEBOOST_cell_38407 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__Q), .b(FE_OFN1132_g64577_p), .c(n_4021), .o(TIMEBOOST_net_11442) );
na02s01 g65926_u2 ( .a(pci_target_unit_del_sync_addr_in_231), .b(FE_OFN775_n_15366), .o(g65926_db) );
na02m06 TIMEBOOST_cell_18246 ( .a(n_12595), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_2__Q), .o(TIMEBOOST_net_4380) );
na02s01 g65927_u2 ( .a(pci_target_unit_del_sync_addr_in_230), .b(FE_OFN775_n_15366), .o(g65927_db) );
na02f02 TIMEBOOST_cell_38893 ( .a(n_3138), .b(wbu_addr_in_272), .o(TIMEBOOST_net_11685) );
na02s02 TIMEBOOST_cell_19949 ( .a(TIMEBOOST_net_5231), .b(g62920_sb), .o(n_6040) );
na02s01 g65928_u2 ( .a(pci_target_unit_del_sync_addr_in_229), .b(FE_OFN775_n_15366), .o(g65928_db) );
na02f02 TIMEBOOST_cell_39090 ( .a(TIMEBOOST_net_11783), .b(FE_OFN1596_n_13741), .o(n_14414) );
na02f02 TIMEBOOST_cell_39091 ( .a(wbu_addr_in_279), .b(g52614_sb), .o(TIMEBOOST_net_11784) );
na04f04 TIMEBOOST_cell_36220 ( .a(n_16170), .b(n_13938), .c(n_13937), .d(FE_RN_835_0), .o(n_16173) );
na02s01 TIMEBOOST_cell_39210 ( .a(TIMEBOOST_net_11843), .b(n_1583), .o(TIMEBOOST_net_11456) );
no03f08 TIMEBOOST_cell_709 ( .a(FE_RN_840_0), .b(FE_RN_838_0), .c(FE_RN_837_0), .o(n_16511) );
na02s01 TIMEBOOST_cell_18016 ( .a(pci_target_unit_fifos_pciw_addr_data_in_140), .b(g64089_sb), .o(TIMEBOOST_net_4265) );
na02s01 TIMEBOOST_cell_43031 ( .a(FE_OFN201_n_9230), .b(g57894_sb), .o(TIMEBOOST_net_13754) );
in01s01 g65931_u0 ( .a(FE_OFN614_n_4501), .o(g65931_sb) );
na02s02 TIMEBOOST_cell_40354 ( .a(TIMEBOOST_net_12415), .b(n_4672), .o(n_4678) );
na02s01 g65931_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__Q), .b(FE_OFN614_n_4501), .o(g65931_db) );
na02s02 TIMEBOOST_cell_40355 ( .a(n_3755), .b(g64956_db), .o(TIMEBOOST_net_12416) );
no02s01 g65932_u0 ( .a(n_2171), .b(n_2044), .o(g65932_p) );
ao12s01 g65932_u1 ( .a(g65932_p), .b(n_2171), .c(n_2044), .o(n_2172) );
na02s02 TIMEBOOST_cell_40356 ( .a(TIMEBOOST_net_12416), .b(g64956_sb), .o(n_3662) );
na02m02 TIMEBOOST_cell_45013 ( .a(pci_target_unit_pcit_if_strd_addr_in_716), .b(g52646_sb), .o(TIMEBOOST_net_14745) );
na03s02 TIMEBOOST_cell_34182 ( .a(g63572_sb), .b(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_), .c(g63572_db), .o(n_4109) );
in01s01 g65934_u0 ( .a(FE_OFN959_n_2299), .o(g65934_sb) );
na02s01 TIMEBOOST_cell_32058 ( .a(configuration_pci_err_addr), .b(wbm_adr_o_0_), .o(TIMEBOOST_net_9940) );
na02s01 g65934_u2 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(FE_OFN959_n_2299), .o(g65934_db) );
na02s02 TIMEBOOST_cell_32057 ( .a(TIMEBOOST_net_9939), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_4922) );
in01s01 g65935_u0 ( .a(FE_OFN959_n_2299), .o(g65935_sb) );
na02s01 TIMEBOOST_cell_32056 ( .a(configuration_pci_err_cs_bit_465), .b(pci_target_unit_wishbone_master_bc_register_reg_2__Q), .o(TIMEBOOST_net_9939) );
na02s01 g65935_u2 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(FE_OFN959_n_2299), .o(g65935_db) );
na02s02 TIMEBOOST_cell_45003 ( .a(pci_target_unit_fifos_pciw_addr_data_in_140), .b(g64215_sb), .o(TIMEBOOST_net_14740) );
in01s01 g65936_u0 ( .a(FE_OFN948_n_2248), .o(g65936_sb) );
na02s01 TIMEBOOST_cell_43334 ( .a(TIMEBOOST_net_13905), .b(g62476_sb), .o(n_6636) );
na02s02 TIMEBOOST_cell_17970 ( .a(pci_target_unit_fifos_pciw_addr_data_in_135), .b(g64214_sb), .o(TIMEBOOST_net_4242) );
no02f10 TIMEBOOST_cell_44759 ( .a(n_16538), .b(n_15744), .o(TIMEBOOST_net_14618) );
no02s01 g65937_u0 ( .a(n_2376), .b(FE_OCPN1854_n_2071), .o(g65937_p) );
ao12s01 g65937_u1 ( .a(g65937_p), .b(n_2376), .c(FE_OCPN1854_n_2071), .o(n_2377) );
no02s01 g65938_u0 ( .a(n_1847), .b(n_1698), .o(g65938_p) );
ao12s01 g65938_u1 ( .a(g65938_p), .b(n_1847), .c(n_1698), .o(n_1848) );
no02m01 g65939_u0 ( .a(n_2566), .b(n_1061), .o(g65939_p) );
ao12s01 g65939_u1 ( .a(g65939_p), .b(n_2566), .c(n_1061), .o(n_2580) );
in01s01 g65940_u0 ( .a(n_2301), .o(g65940_sb) );
na02s01 TIMEBOOST_cell_9732 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__8__Q), .b(g65880_sb), .o(TIMEBOOST_net_1433) );
na02s01 g65940_u2 ( .a(n_8511), .b(n_2301), .o(g65940_db) );
na02s01 TIMEBOOST_cell_9733 ( .a(TIMEBOOST_net_1433), .b(g65880_db), .o(n_1866) );
na02m02 TIMEBOOST_cell_32598 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__1__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__Q), .o(TIMEBOOST_net_10210) );
na02s01 g65941_u2 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(FE_OFN946_n_2248), .o(g65941_db) );
na02f02 TIMEBOOST_cell_32597 ( .a(FE_OFN1554_n_12104), .b(TIMEBOOST_net_10209), .o(TIMEBOOST_net_6491) );
in01s01 g65942_u0 ( .a(FE_OFN2111_n_2248), .o(g65942_sb) );
na02s01 g65942_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__Q), .b(g65942_sb), .o(g65942_da) );
na02s01 g65942_u2 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(FE_OFN2111_n_2248), .o(g65942_db) );
na02s01 TIMEBOOST_cell_36240 ( .a(TIMEBOOST_net_10358), .b(wishbone_slave_unit_del_sync_comp_cycle_count_0_), .o(TIMEBOOST_net_33) );
in01s01 g65943_u0 ( .a(FE_OFN1044_n_2037), .o(g65943_sb) );
na03m02 TIMEBOOST_cell_34903 ( .a(n_4086), .b(n_7618), .c(g59805_da), .o(n_7619) );
na02s01 TIMEBOOST_cell_8878 ( .a(n_16871), .b(n_16864), .o(TIMEBOOST_net_1006) );
na02s01 TIMEBOOST_cell_18829 ( .a(TIMEBOOST_net_4671), .b(g62736_sb), .o(n_5507) );
in01s01 TIMEBOOST_cell_32847 ( .a(TIMEBOOST_net_10348), .o(TIMEBOOST_net_10347) );
na02s02 TIMEBOOST_cell_18018 ( .a(pci_target_unit_fifos_pciw_addr_data_in_124), .b(g64092_sb), .o(TIMEBOOST_net_4266) );
na02s01 TIMEBOOST_cell_15825 ( .a(TIMEBOOST_net_3169), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_396), .o(TIMEBOOST_net_76) );
na02s02 TIMEBOOST_cell_45584 ( .a(TIMEBOOST_net_15030), .b(g64967_db), .o(n_4374) );
na02s01 g65945_u2 ( .a(pci_target_unit_del_sync_addr_in_215), .b(FE_OFN776_n_15366), .o(g65945_db) );
na02s01 TIMEBOOST_cell_41765 ( .a(TIMEBOOST_net_9521), .b(FE_OFN1678_n_4655), .o(TIMEBOOST_net_13121) );
na02s01 TIMEBOOST_cell_40345 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__Q), .b(n_8140), .o(TIMEBOOST_net_12411) );
na02s01 g65946_u2 ( .a(n_2648), .b(n_2301), .o(g65946_db) );
na02s02 TIMEBOOST_cell_40358 ( .a(TIMEBOOST_net_12417), .b(g64988_sb), .o(TIMEBOOST_net_4810) );
na02s02 TIMEBOOST_cell_45693 ( .a(n_40), .b(n_3661), .o(TIMEBOOST_net_15085) );
na02s01 g65947_u2 ( .a(pci_target_unit_del_sync_addr_in_218), .b(FE_OFN776_n_15366), .o(g65947_db) );
na02s01 TIMEBOOST_cell_41766 ( .a(TIMEBOOST_net_13121), .b(g65897_sb), .o(n_1718) );
na03s02 TIMEBOOST_cell_39211 ( .a(n_3783), .b(g65010_sb), .c(n_3636), .o(TIMEBOOST_net_11844) );
na04f04 TIMEBOOST_cell_36222 ( .a(n_14567), .b(n_13862), .c(n_14011), .d(n_14296), .o(n_14612) );
na02m02 TIMEBOOST_cell_39348 ( .a(TIMEBOOST_net_11912), .b(g52652_db), .o(n_14734) );
in01s01 g65949_u0 ( .a(FE_OFN948_n_2248), .o(g65949_sb) );
na02s02 TIMEBOOST_cell_43633 ( .a(n_4015), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__16__Q), .o(TIMEBOOST_net_14055) );
na02s02 TIMEBOOST_cell_17972 ( .a(pci_target_unit_fifos_pciw_addr_data_in_149), .b(g64209_sb), .o(TIMEBOOST_net_4243) );
na02s01 TIMEBOOST_cell_38538 ( .a(TIMEBOOST_net_11507), .b(g62063_sb), .o(n_7746) );
na02s02 TIMEBOOST_cell_42115 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__Q), .b(n_4471), .o(TIMEBOOST_net_13296) );
na02m02 TIMEBOOST_cell_32596 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__Q), .o(TIMEBOOST_net_10209) );
na02s02 TIMEBOOST_cell_30798 ( .a(g57797_sb), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_9310) );
in01s01 g65951_u0 ( .a(n_2299), .o(g65951_sb) );
na02f02 TIMEBOOST_cell_40956 ( .a(TIMEBOOST_net_12716), .b(g57056_sb), .o(n_10508) );
na02s01 g65951_u2 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(n_2299), .o(g65951_db) );
na02f02 TIMEBOOST_cell_45552 ( .a(TIMEBOOST_net_15014), .b(n_11910), .o(n_12630) );
in01s01 g65952_u0 ( .a(FE_OFN1015_n_2053), .o(g65952_sb) );
na02m02 TIMEBOOST_cell_8880 ( .a(n_565), .b(pci_target_unit_pci_target_sm_wr_to_fifo), .o(TIMEBOOST_net_1007) );
na02s01 g65952_u2 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(FE_OFN1015_n_2053), .o(g65952_db) );
na02m02 TIMEBOOST_cell_8881 ( .a(TIMEBOOST_net_1007), .b(n_5755), .o(FE_RN_268_0) );
in01s01 g65953_u0 ( .a(FE_OFN1797_n_2299), .o(g65953_sb) );
na02s01 TIMEBOOST_cell_40349 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__Q), .b(n_8140), .o(TIMEBOOST_net_12413) );
na02s02 TIMEBOOST_cell_36726 ( .a(TIMEBOOST_net_10601), .b(g63598_sb), .o(n_4770) );
na02s01 TIMEBOOST_cell_40360 ( .a(TIMEBOOST_net_12418), .b(g65042_db), .o(n_4327) );
in01s01 g65954_u0 ( .a(FE_OFN1015_n_2053), .o(g65954_sb) );
na02s02 TIMEBOOST_cell_43268 ( .a(TIMEBOOST_net_13872), .b(FE_OFN1289_n_4098), .o(TIMEBOOST_net_12087) );
na02s01 g65954_u2 ( .a(pci_target_unit_fifos_pcir_data_in_178), .b(FE_OFN1015_n_2053), .o(g65954_db) );
na02s01 TIMEBOOST_cell_8883 ( .a(TIMEBOOST_net_1008), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in), .o(n_13186) );
na02f02 TIMEBOOST_cell_40958 ( .a(TIMEBOOST_net_12717), .b(g57311_sb), .o(n_10402) );
na02s01 g65955_u2 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(n_2299), .o(g65955_db) );
na02f06 TIMEBOOST_cell_45553 ( .a(pci_target_unit_wbm_sm_pci_tar_burst_ok), .b(n_731), .o(TIMEBOOST_net_15015) );
na02m02 TIMEBOOST_cell_38706 ( .a(TIMEBOOST_net_11591), .b(g62439_sb), .o(n_6718) );
na04f04 TIMEBOOST_cell_36224 ( .a(n_14560), .b(n_13859), .c(n_14275), .d(n_13980), .o(n_14605) );
na02s01 TIMEBOOST_cell_18181 ( .a(TIMEBOOST_net_4347), .b(g61906_sb), .o(n_8009) );
in01s01 g65957_u0 ( .a(n_2299), .o(g65957_sb) );
na02s01 TIMEBOOST_cell_39227 ( .a(pci_target_unit_fifos_pcir_data_in_185), .b(g65804_sb), .o(TIMEBOOST_net_11852) );
na02s01 g65957_u2 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(n_2299), .o(g65957_db) );
na02s01 TIMEBOOST_cell_39286 ( .a(TIMEBOOST_net_11881), .b(g65799_db), .o(n_1590) );
in01s01 g65958_u0 ( .a(n_2299), .o(g65958_sb) );
na02s02 TIMEBOOST_cell_41767 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__Q), .b(g58354_sb), .o(TIMEBOOST_net_13122) );
na02s01 g65958_u2 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(n_2299), .o(g65958_db) );
na02f02 TIMEBOOST_cell_40960 ( .a(TIMEBOOST_net_12718), .b(g57181_sb), .o(n_11573) );
na02f02 TIMEBOOST_cell_40962 ( .a(TIMEBOOST_net_12719), .b(g57288_sb), .o(n_11464) );
na02s01 g65959_u2 ( .a(pci_target_unit_fifos_pcir_data_in_173), .b(n_2299), .o(g65959_db) );
na02f06 TIMEBOOST_cell_45554 ( .a(TIMEBOOST_net_15015), .b(FE_RN_209_0), .o(n_1535) );
in01s01 g65960_u0 ( .a(n_2299), .o(g65960_sb) );
na02f02 TIMEBOOST_cell_40964 ( .a(TIMEBOOST_net_12720), .b(g57463_sb), .o(n_11270) );
na02s01 g65960_u2 ( .a(pci_target_unit_fifos_pcir_data_in_174), .b(n_2299), .o(g65960_db) );
no02f04 TIMEBOOST_cell_45555 ( .a(n_2869), .b(FE_RN_627_0), .o(TIMEBOOST_net_15016) );
na02f02 TIMEBOOST_cell_40966 ( .a(TIMEBOOST_net_12721), .b(g57065_sb), .o(n_10499) );
na02s01 g65961_u2 ( .a(pci_target_unit_fifos_pcir_data_in_175), .b(n_2299), .o(g65961_db) );
no02f04 TIMEBOOST_cell_45556 ( .a(TIMEBOOST_net_15016), .b(n_287), .o(TIMEBOOST_net_14626) );
in01s01 g65962_u0 ( .a(FE_OFN959_n_2299), .o(g65962_sb) );
na02s01 g65962_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__Q), .b(g65962_sb), .o(g65962_da) );
na02s01 g65962_u2 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(FE_OFN959_n_2299), .o(g65962_db) );
na02m02 TIMEBOOST_cell_40243 ( .a(wbu_addr_in_253), .b(g58793_sb), .o(TIMEBOOST_net_12360) );
na02f02 TIMEBOOST_cell_39092 ( .a(TIMEBOOST_net_10194), .b(TIMEBOOST_net_11784), .o(n_11857) );
na02s01 g65963_u2 ( .a(pci_target_unit_del_sync_addr_in_223), .b(FE_OFN776_n_15366), .o(g65963_db) );
na02s02 TIMEBOOST_cell_18603 ( .a(TIMEBOOST_net_4558), .b(g62822_sb), .o(n_5335) );
in01s01 g65964_u0 ( .a(n_2299), .o(g65964_sb) );
na02f02 TIMEBOOST_cell_40968 ( .a(TIMEBOOST_net_12722), .b(g57135_sb), .o(n_10467) );
na02s01 g65964_u2 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(n_2299), .o(g65964_db) );
no02f06 TIMEBOOST_cell_45557 ( .a(FE_RN_37_0), .b(FE_RN_36_0), .o(TIMEBOOST_net_15017) );
in01s01 g65965_u0 ( .a(FE_OFN1797_n_2299), .o(g65965_sb) );
na03s02 TIMEBOOST_cell_43335 ( .a(n_3781), .b(FE_OFN1222_n_6391), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__Q), .o(TIMEBOOST_net_13906) );
na02s01 g65965_u2 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(FE_OFN1797_n_2299), .o(g65965_db) );
na02f02 TIMEBOOST_cell_44440 ( .a(TIMEBOOST_net_14458), .b(g57086_sb), .o(n_10491) );
in01s01 g65966_u0 ( .a(FE_OFN1797_n_2299), .o(g65966_sb) );
na02m02 TIMEBOOST_cell_44123 ( .a(n_9040), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__Q), .o(TIMEBOOST_net_14300) );
na02s01 g65966_u2 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(FE_OFN1797_n_2299), .o(g65966_db) );
na02s02 TIMEBOOST_cell_45592 ( .a(TIMEBOOST_net_15034), .b(g65233_sb), .o(n_2654) );
in01s01 g65967_u0 ( .a(FE_OFN1797_n_2299), .o(g65967_sb) );
na02f02 TIMEBOOST_cell_44544 ( .a(TIMEBOOST_net_14510), .b(FE_OFN2168_n_8567), .o(TIMEBOOST_net_13001) );
na02s01 g65967_u2 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(FE_OFN1797_n_2299), .o(g65967_db) );
na03f02 TIMEBOOST_cell_44441 ( .a(n_8555), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__Q), .c(FE_OFN1403_n_8567), .o(TIMEBOOST_net_14459) );
na02s02 TIMEBOOST_cell_41768 ( .a(TIMEBOOST_net_13122), .b(g58354_db), .o(n_9016) );
na02s01 g65968_u2 ( .a(pci_target_unit_del_sync_addr_in_220), .b(FE_OFN776_n_15366), .o(g65968_db) );
na02s02 TIMEBOOST_cell_42356 ( .a(TIMEBOOST_net_13416), .b(g54354_sb), .o(n_13087) );
in01s01 g65969_u0 ( .a(FE_OFN1797_n_2299), .o(g65969_sb) );
na02s02 TIMEBOOST_cell_45225 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__Q), .b(n_3646), .o(TIMEBOOST_net_14851) );
na02s01 g65969_u2 ( .a(pci_target_unit_fifos_pcir_data_in_187), .b(FE_OFN1797_n_2299), .o(g65969_db) );
na02f02 TIMEBOOST_cell_44442 ( .a(TIMEBOOST_net_14459), .b(g58593_sb), .o(n_8904) );
in01s01 g65970_u0 ( .a(FE_OFN1797_n_2299), .o(g65970_sb) );
na02s01 TIMEBOOST_cell_9116 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__Q), .b(g65875_sb), .o(TIMEBOOST_net_1125) );
na02s01 TIMEBOOST_cell_42772 ( .a(TIMEBOOST_net_13624), .b(g57983_db), .o(n_9816) );
na02s01 TIMEBOOST_cell_9117 ( .a(TIMEBOOST_net_1125), .b(g65875_db), .o(n_2059) );
in01s01 g65971_u0 ( .a(FE_OFN1797_n_2299), .o(g65971_sb) );
na03f02 TIMEBOOST_cell_44443 ( .a(n_8559), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__Q), .c(FE_OFN1403_n_8567), .o(TIMEBOOST_net_14460) );
na02s02 TIMEBOOST_cell_20669 ( .a(TIMEBOOST_net_5591), .b(FE_OFN2136_n_13124), .o(n_13078) );
na03f02 TIMEBOOST_cell_35250 ( .a(TIMEBOOST_net_10043), .b(n_9144), .c(g58489_sb), .o(n_8919) );
in01s01 g65972_u0 ( .a(FE_OFN1797_n_2299), .o(g65972_sb) );
na02s01 TIMEBOOST_cell_45586 ( .a(TIMEBOOST_net_15031), .b(g65036_db), .o(n_4332) );
no02f04 TIMEBOOST_cell_38781 ( .a(FE_RN_48_0), .b(FE_OFN1709_n_4868), .o(TIMEBOOST_net_11629) );
na02f02 TIMEBOOST_cell_44502 ( .a(TIMEBOOST_net_14489), .b(FE_OFN2177_n_8567), .o(TIMEBOOST_net_13494) );
na02m02 TIMEBOOST_cell_44261 ( .a(n_9047), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__Q), .o(TIMEBOOST_net_14369) );
na02f02 TIMEBOOST_cell_32595 ( .a(FE_OFN1554_n_12104), .b(TIMEBOOST_net_10208), .o(TIMEBOOST_net_6490) );
na02s02 TIMEBOOST_cell_42116 ( .a(TIMEBOOST_net_13296), .b(FE_OFN1310_n_6624), .o(TIMEBOOST_net_11595) );
na02s02 TIMEBOOST_cell_37816 ( .a(TIMEBOOST_net_11146), .b(g62014_sb), .o(n_7867) );
na02f02 TIMEBOOST_cell_40970 ( .a(TIMEBOOST_net_12723), .b(g57201_sb), .o(n_10445) );
na02s02 TIMEBOOST_cell_41883 ( .a(TIMEBOOST_net_485), .b(wishbone_slave_unit_wishbone_slave_do_del_request), .o(TIMEBOOST_net_13180) );
na02m02 TIMEBOOST_cell_38708 ( .a(TIMEBOOST_net_11592), .b(g62600_sb), .o(n_6350) );
na04f04 TIMEBOOST_cell_36226 ( .a(n_12866), .b(n_12867), .c(n_13044), .d(n_12779), .o(n_13128) );
na02s01 TIMEBOOST_cell_18183 ( .a(TIMEBOOST_net_4348), .b(g61911_sb), .o(n_7999) );
in01s01 g65976_u0 ( .a(FE_OFN1017_n_2053), .o(g65976_sb) );
na02f02 TIMEBOOST_cell_43734 ( .a(TIMEBOOST_net_14105), .b(FE_OFN1380_n_8567), .o(TIMEBOOST_net_12814) );
na02s01 g65976_u2 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(FE_OFN1017_n_2053), .o(g65976_db) );
na02s01 TIMEBOOST_cell_8885 ( .a(TIMEBOOST_net_1009), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_384), .o(n_13176) );
in01s01 g65977_u0 ( .a(FE_OFN1015_n_2053), .o(g65977_sb) );
na02m02 TIMEBOOST_cell_43735 ( .a(n_9723), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__Q), .o(TIMEBOOST_net_14106) );
na02s01 g65977_u2 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(FE_OFN1015_n_2053), .o(g65977_db) );
na02s01 TIMEBOOST_cell_8887 ( .a(TIMEBOOST_net_1010), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_409), .o(n_13325) );
in01s01 g65978_u0 ( .a(FE_OFN1015_n_2053), .o(g65978_sb) );
na02s01 TIMEBOOST_cell_8888 ( .a(g54229_db), .b(FE_OFN2114_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_1011) );
na02s01 g65978_u2 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(FE_OFN1015_n_2053), .o(g65978_db) );
na02s01 TIMEBOOST_cell_8889 ( .a(TIMEBOOST_net_1011), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_389), .o(n_13164) );
ao12f10 g65981_u0 ( .a(n_313), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_0_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_), .o(n_938) );
no02s01 g65983_u0 ( .a(pci_target_unit_fifos_wb_clk_inGreyCount_1_), .b(pci_target_unit_fifos_outGreyCount_reg_1__Q), .o(g65983_p) );
ao12s01 g65983_u1 ( .a(g65983_p), .b(pci_target_unit_fifos_wb_clk_inGreyCount_1_), .c(pci_target_unit_fifos_outGreyCount_reg_1__Q), .o(n_1834) );
no02s02 g65984_u0 ( .a(pci_target_unit_fifos_wb_clk_inGreyCount_0_), .b(n_202), .o(g65984_p) );
ao12s01 g65984_u1 ( .a(g65984_p), .b(pci_target_unit_fifos_wb_clk_inGreyCount_0_), .c(n_202), .o(n_1832) );
na02s02 TIMEBOOST_cell_41769 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__Q), .b(g58285_sb), .o(TIMEBOOST_net_13123) );
na02m02 TIMEBOOST_cell_41639 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_29__Q), .b(n_9834), .o(TIMEBOOST_net_13058) );
no02s01 g65992_u0 ( .a(n_1847), .b(n_2376), .o(g65992_p) );
ao12s02 g65992_u1 ( .a(g65992_p), .b(n_1847), .c(n_2376), .o(n_1407) );
no02s02 g65993_u0 ( .a(n_2566), .b(n_2171), .o(g65993_p) );
ao12s02 g65993_u1 ( .a(g65993_p), .b(n_2566), .c(n_2171), .o(n_1406) );
in01s01 g65994_u0 ( .a(FE_OFN992_n_2373), .o(g65994_sb) );
na02m02 TIMEBOOST_cell_32552 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__Q), .o(TIMEBOOST_net_10187) );
na02s01 g65994_u2 ( .a(n_2171), .b(FE_OFN992_n_2373), .o(g65994_db) );
na02f02 TIMEBOOST_cell_22263 ( .a(TIMEBOOST_net_6388), .b(n_8926), .o(n_9947) );
na02s01 TIMEBOOST_cell_32008 ( .a(configuration_pci_err_cs_bit31_24), .b(pci_target_unit_wishbone_master_bc_register_reg_0__Q), .o(TIMEBOOST_net_9915) );
no02f06 TIMEBOOST_cell_45558 ( .a(TIMEBOOST_net_15017), .b(n_16310), .o(n_16311) );
na02s02 TIMEBOOST_cell_32007 ( .a(TIMEBOOST_net_9914), .b(FE_OFN1179_n_3476), .o(TIMEBOOST_net_4896) );
na02m02 TIMEBOOST_cell_43769 ( .a(n_9893), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__Q), .o(TIMEBOOST_net_14123) );
na02s01 g65996_u2 ( .a(n_1551), .b(FE_OFN992_n_2373), .o(g65996_db) );
na02s02 TIMEBOOST_cell_39341 ( .a(TIMEBOOST_net_9548), .b(FE_OFN948_n_2248), .o(TIMEBOOST_net_11909) );
na02s01 TIMEBOOST_cell_40602 ( .a(TIMEBOOST_net_12539), .b(g62672_sb), .o(n_6195) );
na02s01 g65997_u2 ( .a(n_2566), .b(FE_OFN989_n_574), .o(g65997_db) );
na02s02 TIMEBOOST_cell_45559 ( .a(FE_OFN640_n_4669), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__Q), .o(TIMEBOOST_net_15018) );
na02m02 TIMEBOOST_cell_41697 ( .a(g58774_db), .b(g58774_sb), .o(TIMEBOOST_net_13087) );
na02s01 g65998_u2 ( .a(n_2376), .b(FE_OFN989_n_574), .o(g65998_db) );
na02s02 TIMEBOOST_cell_45560 ( .a(TIMEBOOST_net_15018), .b(n_4473), .o(TIMEBOOST_net_10912) );
na02s01 TIMEBOOST_cell_42753 ( .a(g64175_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__Q), .o(TIMEBOOST_net_13615) );
na02s01 g65999_u2 ( .a(n_1847), .b(FE_OFN989_n_574), .o(g65999_db) );
na02s01 TIMEBOOST_cell_42754 ( .a(TIMEBOOST_net_13615), .b(g64175_da), .o(TIMEBOOST_net_11330) );
na02s01 TIMEBOOST_cell_45561 ( .a(g58102_sb), .b(g58102_db), .o(TIMEBOOST_net_15019) );
na02s01 g66000_u2 ( .a(n_1192), .b(FE_OFN989_n_574), .o(g66000_db) );
na02s01 TIMEBOOST_cell_15836 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_98), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3175) );
na02f02 TIMEBOOST_cell_43774 ( .a(TIMEBOOST_net_14125), .b(FE_OFN1409_n_8567), .o(TIMEBOOST_net_12899) );
na02s01 TIMEBOOST_cell_38100 ( .a(TIMEBOOST_net_11288), .b(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_4589) );
na02s02 TIMEBOOST_cell_18457 ( .a(TIMEBOOST_net_4485), .b(g62772_sb), .o(n_5450) );
no02f04 g66002_u0 ( .a(n_595), .b(n_585), .o(g66002_p) );
ao12f04 g66002_u1 ( .a(g66002_p), .b(n_595), .c(n_585), .o(n_1405) );
no02f02 g66003_u0 ( .a(n_674), .b(n_598), .o(g66003_p) );
ao12f04 g66003_u1 ( .a(g66003_p), .b(n_674), .c(n_598), .o(n_1404) );
no02f04 g66004_u0 ( .a(n_672), .b(n_592), .o(g66004_p) );
ao12f04 g66004_u1 ( .a(g66004_p), .b(n_672), .c(n_592), .o(n_1403) );
no02f06 g66005_u0 ( .a(n_597), .b(n_663), .o(g66005_p) );
ao12f06 g66005_u1 ( .a(g66005_p), .b(n_597), .c(n_663), .o(n_1402) );
no02f06 g66006_u0 ( .a(n_678), .b(n_664), .o(g66006_p) );
ao12f06 g66006_u1 ( .a(g66006_p), .b(n_678), .c(n_664), .o(n_1401) );
no02f02 g66007_u0 ( .a(n_586), .b(n_584), .o(g66007_p) );
ao12f04 g66007_u1 ( .a(g66007_p), .b(n_586), .c(n_584), .o(n_1449) );
no02f04 g66008_u0 ( .a(n_603), .b(n_666), .o(g66008_p) );
ao12f04 g66008_u1 ( .a(g66008_p), .b(n_603), .c(n_666), .o(n_1400) );
no02f06 g66009_u0 ( .a(n_593), .b(n_656), .o(g66009_p) );
ao12f06 g66009_u1 ( .a(g66009_p), .b(n_593), .c(n_656), .o(n_1399) );
no02f04 g66010_u0 ( .a(n_667), .b(n_605), .o(g66010_p) );
ao12f04 g66010_u1 ( .a(g66010_p), .b(n_667), .c(n_605), .o(n_1398) );
no02f04 g66011_u0 ( .a(n_670), .b(n_652), .o(g66011_p) );
ao12f04 g66011_u1 ( .a(g66011_p), .b(n_670), .c(n_652), .o(n_1397) );
no02f04 g66012_u0 ( .a(n_650), .b(n_581), .o(g66012_p) );
ao12f04 g66012_u1 ( .a(g66012_p), .b(n_650), .c(n_581), .o(n_1396) );
no02f04 g66013_u0 ( .a(n_583), .b(n_606), .o(g66013_p) );
ao12f04 g66013_u1 ( .a(g66013_p), .b(n_606), .c(n_583), .o(n_1395) );
no02f04 g66014_u0 ( .a(n_673), .b(n_600), .o(g66014_p) );
ao12f04 g66014_u1 ( .a(g66014_p), .b(n_673), .c(n_600), .o(n_1439) );
no02f02 g66015_u0 ( .a(n_594), .b(n_677), .o(g66015_p) );
ao12f04 g66015_u1 ( .a(g66015_p), .b(n_677), .c(n_594), .o(n_1394) );
no02f02 g66016_u0 ( .a(n_675), .b(n_607), .o(g66016_p) );
ao12f04 g66016_u1 ( .a(g66016_p), .b(n_675), .c(n_607), .o(n_1393) );
na02f04 g66064_u0 ( .a(n_1508), .b(pci_target_unit_wishbone_master_read_bound), .o(n_2298) );
no02m06 g66065_u0 ( .a(n_208), .b(n_1477), .o(n_1985) );
na02m04 g66066_u0 ( .a(n_1361), .b(wbu_addr_in_251), .o(g66066_p) );
in01f04 g66066_u1 ( .a(g66066_p), .o(n_2225) );
in01m01 g66067_u0 ( .a(n_1965), .o(n_1561) );
na02m04 g66068_u0 ( .a(n_1357), .b(conf_wb_err_addr_in_943), .o(g66068_p) );
in01m02 g66068_u1 ( .a(g66068_p), .o(n_1965) );
na02m02 TIMEBOOST_cell_41698 ( .a(TIMEBOOST_net_13087), .b(wbu_addr_in_265), .o(n_9889) );
na02s01 g66070_u0 ( .a(n_2301), .b(n_3030), .o(n_3217) );
na02s01 g66071_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1213), .o(n_2612) );
no02s02 g66072_u0 ( .a(parchk_pci_ad_reg_in_1208), .b(n_2493), .o(g66072_p) );
in01s04 g66072_u1 ( .a(g66072_p), .o(n_4498) );
na02s01 g66073_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1212), .o(n_2610) );
no02s02 g66074_u0 ( .a(parchk_pci_ad_reg_in_1206), .b(n_2493), .o(g66074_p) );
in01s03 g66074_u1 ( .a(g66074_p), .o(n_4672) );
no02s02 g66075_u0 ( .a(parchk_pci_ad_reg_in_1233), .b(n_2493), .o(g66075_p) );
in01s03 g66075_u1 ( .a(g66075_p), .o(n_4479) );
no02s02 g66076_u0 ( .a(parchk_pci_ad_reg_in), .b(n_2493), .o(g66076_p) );
in01s03 g66076_u1 ( .a(g66076_p), .o(n_4488) );
no02s02 g66077_u0 ( .a(parchk_pci_ad_reg_in_1214), .b(n_2344), .o(g66077_p) );
in01s03 g66077_u1 ( .a(g66077_p), .o(n_3747) );
no02s02 g66078_u0 ( .a(parchk_pci_ad_reg_in_1212), .b(n_2493), .o(g66078_p) );
in01s03 g66078_u1 ( .a(g66078_p), .o(n_4465) );
no02s02 g66079_u0 ( .a(parchk_pci_ad_reg_in_1211), .b(n_2344), .o(g66079_p) );
in01s03 g66079_u1 ( .a(g66079_p), .o(n_3764) );
no02s02 g66080_u0 ( .a(parchk_pci_ad_reg_in_1228), .b(n_2493), .o(g66080_p) );
in01s04 g66080_u1 ( .a(g66080_p), .o(n_4444) );
no02s02 g66081_u0 ( .a(n_2509), .b(n_2344), .o(g66081_p) );
in01s06 g66081_u1 ( .a(FE_OFN335_g66081_p), .o(n_3770) );
no02s02 g66082_u0 ( .a(parchk_pci_ad_reg_in_1213), .b(n_2344), .o(g66082_p) );
in01s03 g66082_u1 ( .a(g66082_p), .o(n_3783) );
na02s02 g66083_u0 ( .a(n_15922), .b(n_2308), .o(g66083_p) );
in01s02 g66083_u1 ( .a(g66083_p), .o(n_2562) );
no02s02 g66084_u0 ( .a(n_1122), .b(wishbone_slave_unit_del_sync_comp_cycle_count_10_), .o(g66084_p) );
in01s01 g66084_u1 ( .a(g66084_p), .o(n_1392) );
no02s01 g66085_u0 ( .a(parchk_pci_ad_reg_in_1229), .b(n_2344), .o(g66085_p) );
in01s06 g66085_u1 ( .a(FE_OFN1938_g66085_p), .o(n_3785) );
no02s02 g66086_u0 ( .a(parchk_pci_ad_reg_in_1235), .b(n_2493), .o(g66086_p) );
in01s04 g66086_u1 ( .a(g66086_p), .o(n_4645) );
no02s02 g66087_u0 ( .a(parchk_pci_ad_reg_in_1216), .b(n_2344), .o(g66087_p) );
in01s06 g66087_u1 ( .a(FE_OFN2061_g66087_p), .o(n_3777) );
na02s01 g66088_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1209), .o(n_2604) );
no02s02 g66089_u0 ( .a(parchk_pci_ad_reg_in_1205), .b(n_2344), .o(g66089_p) );
in01s06 g66089_u1 ( .a(FE_OFN337_g66089_p), .o(n_3774) );
no02s02 g66090_u0 ( .a(parchk_pci_ad_reg_in_1223), .b(n_2493), .o(g66090_p) );
in01s03 g66090_u1 ( .a(g66090_p), .o(n_4447) );
na02s01 g66092_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1207), .o(n_2788) );
no02s02 g66093_u0 ( .a(parchk_pci_ad_reg_in_1225), .b(n_2493), .o(g66093_p) );
in01s03 g66093_u1 ( .a(g66093_p), .o(n_4470) );
no02s02 g66094_u0 ( .a(parchk_pci_ad_reg_in_1217), .b(n_2493), .o(g66094_p) );
in01s04 g66094_u1 ( .a(g66094_p), .o(n_4452) );
no02s01 g66095_u0 ( .a(FE_OFN1781_parchk_pci_ad_reg_in_1221), .b(n_2493), .o(g66095_p) );
in01s06 g66095_u1 ( .a(FE_OFN1940_g66095_p), .o(n_4450) );
na02s02 g66096_u0 ( .a(n_1479), .b(n_1478), .o(g66096_p) );
in01m02 g66096_u1 ( .a(g66096_p), .o(n_2244) );
na02f02 g66097_u0 ( .a(n_2967), .b(n_1390), .o(g66097_p) );
in01m02 g66097_u1 ( .a(g66097_p), .o(n_1391) );
no02s02 g66098_u0 ( .a(parchk_pci_ad_reg_in_1220), .b(n_2344), .o(g66098_p) );
in01s03 g66098_u1 ( .a(g66098_p), .o(n_3744) );
na02s02 g66099_u0 ( .a(n_1378), .b(n_1480), .o(g66099_p) );
in01s02 g66099_u1 ( .a(g66099_p), .o(n_2243) );
no02s02 g66100_u0 ( .a(parchk_pci_ad_reg_in_1232), .b(n_2493), .o(g66100_p) );
in01s03 g66100_u1 ( .a(g66100_p), .o(n_4442) );
in01s01 g66105_u0 ( .a(n_3123), .o(n_2140) );
na02f20 g66106_u0 ( .a(n_1196), .b(pci_target_unit_pci_target_sm_backoff), .o(n_3123) );
no02s02 g66107_u0 ( .a(parchk_pci_ad_reg_in_1210), .b(n_2344), .o(g66107_p) );
in01s03 g66107_u1 ( .a(g66107_p), .o(n_3780) );
no02s02 g66108_u0 ( .a(parchk_pci_ad_reg_in_1218), .b(n_2493), .o(g66108_p) );
in01s03 g66108_u1 ( .a(g66108_p), .o(n_4476) );
na02s01 g66109_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1206), .o(n_2790) );
no02s02 g66110_u0 ( .a(parchk_pci_ad_reg_in_1207), .b(n_2344), .o(g66110_p) );
in01s03 g66110_u1 ( .a(g66110_p), .o(n_3739) );
na02s01 g66111_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1208), .o(n_2732) );
na02s01 g66112_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1210), .o(n_2783) );
na02f02 g66113_u0 ( .a(n_1481), .b(n_1482), .o(g66113_p) );
in01f02 g66113_u1 ( .a(g66113_p), .o(n_2397) );
no02m02 g66114_u0 ( .a(n_1057), .b(n_639), .o(n_2675) );
na02s01 g66117_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1211), .o(n_2606) );
no02s01 g66118_u0 ( .a(n_1124), .b(n_207), .o(g66118_p) );
in01s01 g66118_u1 ( .a(g66118_p), .o(n_1389) );
na02s01 g66119_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1205), .o(n_2779) );
no02m02 g66120_u0 ( .a(n_1435), .b(n_978), .o(n_2415) );
na02m02 g66121_u0 ( .a(n_2435), .b(n_1388), .o(g66121_p) );
in01m02 g66121_u1 ( .a(g66121_p), .o(n_2229) );
no02s01 g66122_u0 ( .a(n_1824), .b(pci_target_unit_pcit_if_req_req_pending_in), .o(g66122_p) );
in01s01 g66122_u1 ( .a(g66122_p), .o(n_1825) );
na02s01 g66123_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in), .o(n_2601) );
no02s02 g66124_u0 ( .a(parchk_pci_ad_reg_in_1231), .b(n_2493), .o(g66124_p) );
in01s04 g66124_u1 ( .a(g66124_p), .o(n_4482) );
no02s01 g66125_u0 ( .a(parchk_pci_ad_reg_in_1215), .b(n_2344), .o(g66125_p) );
in01s03 g66125_u1 ( .a(g66125_p), .o(n_3761) );
no02s02 g66127_u0 ( .a(parchk_pci_ad_reg_in_1227), .b(n_2344), .o(g66127_p) );
in01s03 g66127_u1 ( .a(g66127_p), .o(n_3741) );
no02s02 g66128_u0 ( .a(parchk_pci_ad_reg_in_1226), .b(n_2344), .o(g66128_p) );
in01s03 g66128_u1 ( .a(g66128_p), .o(n_3749) );
no02s02 g66129_u0 ( .a(parchk_pci_ad_reg_in_1224), .b(n_2344), .o(g66129_p) );
in01s03 g66129_u1 ( .a(g66129_p), .o(n_3752) );
no02s02 g66130_u0 ( .a(parchk_pci_ad_reg_in_1219), .b(n_2344), .o(g66130_p) );
in01s03 g66130_u1 ( .a(g66130_p), .o(n_3792) );
na02s02 g66131_u0 ( .a(n_1125), .b(pci_target_unit_del_sync_comp_cycle_count_6_), .o(n_1484) );
no02f04 g66132_u0 ( .a(n_2215), .b(pci_target_unit_wishbone_master_first_wb_data_access), .o(g66132_p) );
in01f02 g66132_u1 ( .a(g66132_p), .o(n_2390) );
no02s02 g66133_u0 ( .a(parchk_pci_ad_reg_in_1209), .b(n_2344), .o(g66133_p) );
in01s03 g66133_u1 ( .a(g66133_p), .o(n_3755) );
no02s02 g66134_u0 ( .a(FE_OFN1777_parchk_pci_ad_reg_in_1222), .b(n_2493), .o(g66134_p) );
in01s04 g66134_u1 ( .a(g66134_p), .o(n_4473) );
na02s02 g66135_u0 ( .a(n_1123), .b(wishbone_slave_unit_del_sync_comp_cycle_count_6_), .o(n_1485) );
no02s02 g66136_u0 ( .a(parchk_pci_ad_reg_in_1230), .b(n_2493), .o(g66136_p) );
in01s06 g66136_u1 ( .a(g66136_p), .o(n_4493) );
no02s01 g66137_u0 ( .a(n_1192), .b(n_5757), .o(n_2303) );
na02m02 g66138_u0 ( .a(n_1227), .b(n_2411), .o(g66138_p) );
in01m02 g66138_u1 ( .a(g66138_p), .o(n_1986) );
no02s02 g66139_u0 ( .a(n_869), .b(n_1019), .o(n_1387) );
no02s01 g66140_u0 ( .a(n_626), .b(n_642), .o(n_1170) );
na02f02 TIMEBOOST_cell_42222 ( .a(TIMEBOOST_net_13349), .b(FE_OFN1400_n_8567), .o(TIMEBOOST_net_12305) );
na02s01 g66142_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__Q), .b(FE_OFN614_n_4501), .o(n_1559) );
no02f02 g66143_u0 ( .a(n_15291), .b(n_2127), .o(g66143_p) );
in01f02 g66143_u1 ( .a(g66143_p), .o(n_3019) );
na02m02 g66145_u0 ( .a(n_1228), .b(n_1229), .o(g66145_p) );
in01m02 g66145_u1 ( .a(g66145_p), .o(n_2753) );
na02s02 g66146_u0 ( .a(FE_OFN996_n_15366), .b(pci_target_unit_pci_target_sm_rd_progress), .o(n_1823) );
no02f03 g66147_u0 ( .a(n_604), .b(n_601), .o(g66147_p) );
in01f03 g66147_u1 ( .a(g66147_p), .o(n_1036) );
na02s01 g66148_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__Q), .b(FE_OFN1795_n_9904), .o(n_1230) );
na02s01 g66150_u0 ( .a(pci_target_unit_pci_target_if_same_read_reg), .b(FE_OFN996_n_15366), .o(n_2371) );
no02s02 g66151_u0 ( .a(n_1091), .b(n_851), .o(n_1486) );
na02s01 g66152_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__Q), .b(FE_OFN1800_n_9690), .o(n_1822) );
no02s01 g66153_u0 ( .a(configuration_rst_inactive), .b(n_2373), .o(g66153_p) );
in01s01 g66153_u1 ( .a(g66153_p), .o(n_1385) );
na02s01 g66154_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__Q), .b(FE_OFN519_n_9697), .o(n_1821) );
na02f02 g66155_u0 ( .a(n_2331), .b(n_16541), .o(g66155_p) );
in01f02 g66155_u1 ( .a(g66155_p), .o(n_3371) );
na02s01 TIMEBOOST_cell_45739 ( .a(n_1906), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__Q), .o(TIMEBOOST_net_15108) );
na02s01 g66158_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__Q), .b(FE_OFN672_n_4505), .o(n_1488) );
na02s01 g66159_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__Q), .b(FE_OFN665_n_4495), .o(n_2138) );
na02f02 g66160_u0 ( .a(n_2560), .b(n_2129), .o(g66160_p) );
in01f02 g66160_u1 ( .a(g66160_p), .o(n_3246) );
na02s01 g66161_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__Q), .b(FE_OFN529_n_9899), .o(n_1820) );
in01s02 g66162_u0 ( .a(FE_OFN780_n_2746), .o(n_2747) );
na02s01 TIMEBOOST_cell_30866 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__Q), .b(pci_target_unit_fifos_pcir_data_in_163), .o(TIMEBOOST_net_9344) );
no02s02 g66164_u0 ( .a(n_620), .b(n_622), .o(n_1169) );
no02f02 g66165_u0 ( .a(n_15276), .b(n_16291), .o(g66165_p) );
in01f02 g66165_u1 ( .a(g66165_p), .o(n_1819) );
no02s02 g66166_u0 ( .a(n_729), .b(n_734), .o(n_1037) );
no02s01 g66167_u0 ( .a(n_1192), .b(FE_OFN999_n_15978), .o(n_2370) );
na02s01 TIMEBOOST_cell_40362 ( .a(TIMEBOOST_net_12419), .b(g65751_db), .o(n_1923) );
na02s01 g66169_u0 ( .a(FE_OFN923_n_4740), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__Q), .o(n_1815) );
na02s01 g66170_u0 ( .a(pci_target_unit_pci_target_sm_rd_from_fifo), .b(FE_OFN996_n_15366), .o(n_2369) );
na02s01 g66171_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__Q), .b(FE_OFN595_n_9694), .o(n_1814) );
no02f10 g66172_u0 ( .a(n_1033), .b(n_863), .o(n_1231) );
no02s01 g66173_u0 ( .a(n_1551), .b(output_backup_trdy_out_reg_Q), .o(n_2137) );
na02s01 g66174_u0 ( .a(pci_target_unit_pci_target_sm_wr_progress), .b(FE_OFN996_n_15366), .o(n_2367) );
no02s01 g66175_u0 ( .a(n_737), .b(n_640), .o(n_1168) );
no02s01 g66176_u0 ( .a(n_3480), .b(n_691), .o(g66176_p) );
in01s01 g66176_u1 ( .a(g66176_p), .o(n_1557) );
no02s02 g66177_u0 ( .a(n_708), .b(n_649), .o(n_1167) );
na02f04 g66178_u0 ( .a(n_1813), .b(n_1812), .o(g66178_p) );
in01f04 g66178_u1 ( .a(g66178_p), .o(n_2447) );
na02s01 g66179_u0 ( .a(n_424), .b(FE_OFN622_n_4409), .o(n_1555) );
na02s01 g66180_u0 ( .a(n_1023), .b(FE_OFN2214_n_15366), .o(n_2366) );
in01s01 g66182_u0 ( .a(n_1554), .o(n_13817) );
no02f04 g66184_u0 ( .a(pci_target_unit_pci_target_sm_backoff), .b(n_1366), .o(g66184_p) );
in01f02 g66184_u1 ( .a(g66184_p), .o(n_1554) );
na02s01 g66185_u0 ( .a(FE_OFN2214_n_15366), .b(n_2078), .o(n_2364) );
na02s01 g66187_u0 ( .a(n_922), .b(n_1383), .o(n_1384) );
na02m02 TIMEBOOST_cell_42223 ( .a(n_9467), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__Q), .o(TIMEBOOST_net_13350) );
na02s01 g66189_u0 ( .a(FE_OFN2214_n_15366), .b(n_15998), .o(n_2363) );
na02m04 g66190_u0 ( .a(n_3194), .b(n_1381), .o(g66190_p) );
in01m02 g66190_u1 ( .a(g66190_p), .o(n_2754) );
na02s01 g66191_u0 ( .a(FE_OFN2214_n_15366), .b(n_16690), .o(n_2362) );
no02f20 g66193_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_), .o(n_313) );
na02s02 g66194_u0 ( .a(wbu_wb_init_complete_in), .b(n_779), .o(g66194_p) );
in01s02 g66194_u1 ( .a(g66194_p), .o(n_2558) );
na02s02 g66195_u0 ( .a(n_1241), .b(n_2433), .o(g66195_p) );
in01s02 g66195_u1 ( .a(g66195_p), .o(n_2236) );
na02s02 g66197_u0 ( .a(n_1479), .b(n_1378), .o(g66197_p) );
in01s02 g66197_u1 ( .a(g66197_p), .o(n_1379) );
no02s01 g66200_u0 ( .a(n_1504), .b(n_695), .o(n_2136) );
na02s01 g66201_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q), .b(FE_OFN1660_n_4490), .o(n_1377) );
na02f02 g66202_u0 ( .a(n_1812), .b(n_2795), .o(g66202_p) );
in01f02 g66202_u1 ( .a(g66202_p), .o(n_3107) );
no02s02 g66203_u0 ( .a(n_1008), .b(n_864), .o(n_1252) );
na02s01 g66204_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__Q), .b(FE_OFN562_n_9895), .o(n_1493) );
na02s01 g66205_u0 ( .a(pci_target_unit_del_sync_bc_in), .b(FE_OFN996_n_15366), .o(n_2361) );
no02s02 g66206_u0 ( .a(n_951), .b(n_1035), .o(n_1253) );
no02s02 g66207_u0 ( .a(n_624), .b(n_613), .o(n_1166) );
na02s01 g66208_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__Q), .b(FE_OFN648_n_4497), .o(n_1553) );
na02s01 g66209_u0 ( .a(pci_target_unit_pci_target_sm_same_read_reg), .b(FE_OFN996_n_15366), .o(n_2359) );
na02s01 g66212_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__Q), .b(FE_OFN577_n_9902), .o(n_1810) );
na02f02 TIMEBOOST_cell_40972 ( .a(TIMEBOOST_net_12724), .b(g57171_sb), .o(n_11585) );
no02s02 g66214_u0 ( .a(n_625), .b(n_610), .o(n_1073) );
no02s01 g66215_u0 ( .a(n_2493), .b(n_3480), .o(g66215_p) );
in01s01 g66215_u1 ( .a(g66215_p), .o(n_3481) );
in01m02 g66216_u0 ( .a(n_1548), .o(n_1549) );
na02m04 g66217_u0 ( .a(n_1269), .b(n_1270), .o(n_1548) );
na02f02 g66219_u0 ( .a(n_1808), .b(n_16159), .o(n_1809) );
na02s02 g66221_u0 ( .a(n_16160), .b(n_16151), .o(n_2966) );
na02s20 g66223_u0 ( .a(wbu_wb_init_complete_in), .b(wbs_cyc_i), .o(g66223_p) );
in01m06 g66223_u1 ( .a(g66223_p), .o(n_2557) );
no02s02 g66224_u0 ( .a(n_616), .b(n_643), .o(n_1080) );
na02s02 g66225_u0 ( .a(n_1374), .b(n_1373), .o(n_1974) );
no02s02 g66226_u0 ( .a(n_615), .b(n_612), .o(n_1207) );
na02s02 g66227_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__Q), .b(FE_OFN1623_n_4438), .o(n_1547) );
no02s01 g66228_u0 ( .a(n_15371), .b(n_2134), .o(n_2135) );
na04s02 TIMEBOOST_cell_34183 ( .a(g63565_da), .b(g63565_db), .c(g61957_sb), .d(g61957_db), .o(n_6958) );
na02f01 g66230_u0 ( .a(n_16160), .b(n_1445), .o(n_3341) );
no02s02 g66231_u0 ( .a(n_2036), .b(n_2297), .o(n_2556) );
no02f04 g66232_u0 ( .a(n_849), .b(n_850), .o(g66232_p) );
in01f02 g66232_u1 ( .a(g66232_p), .o(n_1371) );
na02s01 g66233_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__Q), .b(FE_OFN659_n_4392), .o(n_1546) );
na02m02 g66234_u0 ( .a(n_2431), .b(n_1282), .o(g66234_p) );
in01m02 g66234_u1 ( .a(g66234_p), .o(n_2238) );
no02f06 g66236_u0 ( .a(n_847), .b(n_858), .o(n_1369) );
na02f02 g66237_u0 ( .a(n_15065), .b(wbu_am1_in), .o(g66237_p) );
in01f02 g66237_u1 ( .a(g66237_p), .o(n_2358) );
na02m02 g66239_u0 ( .a(n_2463), .b(n_2596), .o(g66239_p) );
in01m02 g66239_u1 ( .a(g66239_p), .o(n_1969) );
na02s01 g66240_u0 ( .a(n_1120), .b(n_535), .o(n_1545) );
no02s02 g66241_u0 ( .a(n_1012), .b(n_867), .o(n_1365) );
na02s01 g66242_u0 ( .a(n_497), .b(FE_OFN2214_n_15366), .o(n_2356) );
na02s01 TIMEBOOST_cell_44785 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__Q), .b(FE_OFN575_n_9902), .o(TIMEBOOST_net_14631) );
na02s01 g66245_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__Q), .b(FE_OFN601_n_9687), .o(n_1806) );
no02f06 g66246_u0 ( .a(n_1031), .b(n_870), .o(n_1363) );
no02s02 g66247_u0 ( .a(n_617), .b(n_645), .o(n_1208) );
na02s02 g66248_u0 ( .a(n_1361), .b(n_1378), .o(g66248_p) );
in01s02 g66248_u1 ( .a(g66248_p), .o(n_1362) );
in01m02 g66250_u0 ( .a(n_1805), .o(n_2132) );
na02s02 TIMEBOOST_cell_43136 ( .a(TIMEBOOST_net_13806), .b(FE_OFN1246_n_4093), .o(TIMEBOOST_net_12073) );
no02s01 g66252_u0 ( .a(FE_OFN996_n_15366), .b(pci_target_unit_pcit_if_req_req_pending_in), .o(n_2353) );
na02s01 g66253_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__Q), .b(FE_OFN903_n_4736), .o(n_1804) );
na02s01 g66254_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__Q), .b(FE_OFN531_n_9823), .o(n_1542) );
na02s01 g66255_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__Q), .b(FE_OFN1012_n_4734), .o(n_1803) );
na02s01 g66256_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__Q), .b(FE_OFN634_n_4454), .o(n_1642) );
na02s01 TIMEBOOST_cell_42692 ( .a(TIMEBOOST_net_13584), .b(g58182_db), .o(TIMEBOOST_net_10048) );
na02s01 g66258_u0 ( .a(pci_target_unit_pci_target_sm_wr_to_fifo), .b(FE_OFN996_n_15366), .o(n_2352) );
no02s02 g66259_u0 ( .a(n_722), .b(n_658), .o(n_1164) );
na02s01 g66260_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__Q), .b(n_4417), .o(n_2131) );
no02s01 g66261_u0 ( .a(FE_OFN996_n_15366), .b(wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q), .o(n_1802) );
na02s01 g66262_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__Q), .b(FE_OFN554_n_9864), .o(n_1800) );
no02s02 g66264_u0 ( .a(n_641), .b(n_614), .o(n_1209) );
na02s01 g66265_u0 ( .a(n_2314), .b(FE_OFN996_n_15366), .o(n_2351) );
na02s02 TIMEBOOST_cell_17254 ( .a(n_4482), .b(FE_OFN1642_n_4671), .o(TIMEBOOST_net_3884) );
na02m02 g66267_u0 ( .a(n_965), .b(n_2228), .o(g66267_p) );
in01m02 g66267_u1 ( .a(g66267_p), .o(n_1359) );
no02s01 g66268_u0 ( .a(n_2214), .b(n_1808), .o(n_3223) );
na02f01 g66269_u0 ( .a(n_1966), .b(n_1357), .o(g66269_p) );
in01m02 g66269_u1 ( .a(g66269_p), .o(n_1358) );
na02s01 g66270_u0 ( .a(n_1228), .b(n_1355), .o(n_1356) );
na02s01 g66271_u0 ( .a(n_1519), .b(FE_OFN2214_n_15366), .o(n_2349) );
no02s02 g66272_u0 ( .a(n_844), .b(n_838), .o(n_1354) );
na02s01 TIMEBOOST_cell_42693 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q), .b(FE_OFN1657_n_9502), .o(TIMEBOOST_net_13585) );
no02s02 g66274_u0 ( .a(n_1467), .b(n_1034), .o(n_1799) );
no02s02 g66275_u0 ( .a(n_721), .b(n_611), .o(n_1162) );
no02s02 g66276_u0 ( .a(n_609), .b(n_711), .o(n_1161) );
na02f08 g66277_u0 ( .a(n_329), .b(n_1211), .o(n_2430) );
na02f02 g66278_u0 ( .a(n_16541), .b(n_15755), .o(g66278_p) );
in01f02 g66278_u1 ( .a(g66278_p), .o(n_2555) );
in01f02 g66281_u0 ( .a(n_3023), .o(n_3386) );
in01f03 g66282_u0 ( .a(n_2804), .o(n_3023) );
no02f06 g66285_u0 ( .a(n_1306), .b(n_16860), .o(n_2804) );
no02m02 g66286_u0 ( .a(n_1217), .b(n_840), .o(g66286_p) );
in01s02 g66286_u1 ( .a(g66286_p), .o(n_1541) );
na02f02 g66287_u0 ( .a(n_1248), .b(n_15922), .o(g66287_p) );
in01f03 g66287_u1 ( .a(g66287_p), .o(n_2777) );
no02s02 g66288_u0 ( .a(n_742), .b(n_871), .o(n_1352) );
no02s02 g66289_u0 ( .a(n_866), .b(n_960), .o(n_1351) );
na02f06 g66290_dup_u0 ( .a(n_15065), .b(n_2129), .o(g66290_dup_p) );
in01f08 g66290_dup_u1 ( .a(g66290_dup_p), .o(n_15445) );
no02m02 g66291_u0 ( .a(n_1448), .b(pci_target_unit_wbm_sm_pci_tar_read_request), .o(g66291_p) );
in01m02 g66291_u1 ( .a(g66291_p), .o(n_1798) );
in01f04 g66292_u0 ( .a(n_3004), .o(n_3504) );
in01f04 g66293_u0 ( .a(n_3248), .o(n_3004) );
no02f10 g66294_u0 ( .a(n_2553), .b(n_15291), .o(n_3248) );
no02s02 g66295_u0 ( .a(n_2042), .b(n_1754), .o(n_2347) );
no02s02 g66297_u0 ( .a(n_999), .b(n_959), .o(n_1350) );
na02m02 g66298_u0 ( .a(n_16964), .b(n_1347), .o(g66298_p) );
in01s02 g66298_u1 ( .a(g66298_p), .o(n_1349) );
no02f04 g66299_u0 ( .a(n_587), .b(n_952), .o(g66299_p) );
in01f02 g66299_u1 ( .a(g66299_p), .o(n_1346) );
no02s02 g66301_u0 ( .a(n_950), .b(n_855), .o(n_1433) );
no02f02 g66302_u0 ( .a(n_2126), .b(n_2127), .o(g66302_p) );
in01f02 g66302_u1 ( .a(g66302_p), .o(n_4806) );
no02f04 g66303_u0 ( .a(n_2553), .b(n_2552), .o(g66303_p) );
in01f02 g66303_u1 ( .a(g66303_p), .o(n_3018) );
no02f02 g66305_u0 ( .a(n_2126), .b(n_1777), .o(n_3368) );
no02f10 g66309_u0 ( .a(n_2453), .b(n_2552), .o(n_3295) );
no02f04 g66310_u0 ( .a(n_841), .b(n_843), .o(g66310_p) );
in01f02 g66310_u1 ( .a(g66310_p), .o(n_1345) );
na02s01 g66311_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__Q), .b(FE_OFN587_n_9692), .o(n_1540) );
no02s02 g66312_u0 ( .a(n_865), .b(n_744), .o(n_1344) );
no02f10 g66313_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_1_), .o(n_1539) );
no02f08 g66315_u0 ( .a(n_2344), .b(n_2685), .o(g66315_p) );
in01f04 g66315_u1 ( .a(g66315_p), .o(n_2345) );
no02s02 g66316_u0 ( .a(n_839), .b(n_743), .o(n_1343) );
no02s02 g66317_u0 ( .a(n_836), .b(n_747), .o(n_1342) );
na02f02 TIMEBOOST_cell_42224 ( .a(TIMEBOOST_net_13350), .b(FE_OFN1424_n_8567), .o(TIMEBOOST_net_12301) );
no02m02 g66319_u0 ( .a(n_7622), .b(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(n_2343) );
no02s01 g66320_u0 ( .a(n_627), .b(n_623), .o(n_1160) );
no02s02 g66321_u0 ( .a(n_837), .b(n_1007), .o(n_1341) );
no02s01 g66322_u0 ( .a(n_559), .b(wishbone_slave_unit_del_sync_comp_done_reg_main), .o(g66322_p) );
in01s01 g66322_u1 ( .a(g66322_p), .o(n_1696) );
na02s02 g66323_u0 ( .a(n_2125), .b(n_2795), .o(g66323_p) );
in01s02 g66323_u1 ( .a(g66323_p), .o(n_3221) );
no02s02 g66324_u0 ( .a(n_725), .b(n_621), .o(n_1159) );
no02s02 g66325_u0 ( .a(n_1004), .b(n_833), .o(n_1340) );
na02f06 g66327_u0 ( .a(n_2094), .b(n_16424), .o(g66327_p) );
in01f06 g66327_u1 ( .a(g66327_p), .o(n_3231) );
in01f08 g66328_u0 ( .a(n_2768), .o(n_7031) );
in01f08 g66332_u0 ( .a(n_3026), .o(n_2768) );
na02f04 g66336_u0 ( .a(n_2341), .b(n_16036), .o(g66336_p) );
in01f04 g66336_u1 ( .a(g66336_p), .o(n_3026) );
no02s02 g66337_u0 ( .a(n_700), .b(n_648), .o(n_1189) );
na02f01 g66338_u0 ( .a(n_15755), .b(n_16424), .o(g66338_p) );
in01m02 g66338_u1 ( .a(g66338_p), .o(n_2339) );
na02s01 g66339_u0 ( .a(n_2316), .b(FE_OFN2214_n_15366), .o(n_2767) );
na02m02 g66340_u0 ( .a(n_1325), .b(n_15371), .o(n_1538) );
na02s02 TIMEBOOST_cell_41796 ( .a(TIMEBOOST_net_13136), .b(g58387_db), .o(n_9444) );
in01f04 g66346_u0 ( .a(n_1999), .o(n_3250) );
no02f06 g66347_u0 ( .a(n_1808), .b(n_1998), .o(n_1999) );
na02s01 g66348_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__Q), .b(FE_OFN1046_n_16657), .o(n_1795) );
na02s01 g66349_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__Q), .b(FE_OFN682_n_4460), .o(n_1537) );
ao12s02 g66350_u0 ( .a(n_2494), .b(n_716), .c(conf_wb_err_bc_in_846), .o(n_3001) );
ao12s01 g66352_u0 ( .a(configuration_set_pci_err_cs_bit8), .b(configuration_sync_pci_err_cs_8_delayed_del_bit), .c(configuration_sync_pci_err_cs_8_sync_del_bit), .o(n_1191) );
na02f06 g66353_u0 ( .a(pci_target_unit_pci_target_sm_read_completed_reg), .b(n_2337), .o(n_2883) );
ao12s01 g66354_u0 ( .a(n_2031), .b(n_1512), .c(n_15295), .o(n_2547) );
oa12f04 g66356_u0 ( .a(n_1507), .b(n_1220), .c(n_730), .o(n_2000) );
na02f02 g66357_u0 ( .a(n_16541), .b(n_16001), .o(g66357_p) );
in01f02 g66357_u1 ( .a(g66357_p), .o(n_3372) );
na02f04 g66358_u0 ( .a(n_15125), .b(n_1446), .o(g66358_p) );
in01f06 g66358_u1 ( .a(g66358_p), .o(n_3252) );
no02s02 g66359_u0 ( .a(n_930), .b(n_1334), .o(n_1469) );
na02s02 TIMEBOOST_cell_43101 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__Q), .b(n_3654), .o(TIMEBOOST_net_13789) );
ao22s01 g66361_u0 ( .a(n_713), .b(n_345), .c(wishbone_slave_unit_fifos_wbw_outTransactionCount_0_), .d(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q), .o(n_1338) );
ao22s01 g66362_u0 ( .a(n_567), .b(n_362), .c(wishbone_slave_unit_fifos_wbw_inTransactionCount_0_), .d(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q), .o(n_1337) );
ao22s01 g66363_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_956), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_649), .o(n_1794) );
ao22s01 g66365_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_969), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_662), .o(n_1793) );
ao22s01 g66366_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_946), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_639), .o(n_2121) );
na02m02 TIMEBOOST_cell_42225 ( .a(n_9346), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__Q), .o(TIMEBOOST_net_13351) );
ao22s01 g66369_u0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_943), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_636), .o(n_2120) );
ao22s01 g66370_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_951), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_644), .o(n_2119) );
ao22s01 g66371_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_959), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_652), .o(n_2117) );
ao22s02 g66372_u0 ( .a(n_2115), .b(conf_wb_err_addr_in_963), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_656), .o(n_2116) );
ao22s01 g66373_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_971), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_664), .o(n_1790) );
ao22s01 g66374_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_957), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_650), .o(n_2114) );
ao22s01 g66375_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_961), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_654), .o(n_2113) );
ao22m02 g66376_u0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_953), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_646), .o(n_2111) );
ao22s01 g66377_u0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_944), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_637), .o(n_2110) );
na02f02 TIMEBOOST_cell_42226 ( .a(TIMEBOOST_net_13351), .b(FE_OFN1388_n_8567), .o(TIMEBOOST_net_12284) );
ao22s01 g66379_u0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_966), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_659), .o(n_2108) );
ao22s01 g66381_u0 ( .a(n_1787), .b(conf_wb_err_addr_in_967), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_660), .o(n_2106) );
ao22s01 g66382_u0 ( .a(FE_OFN1617_n_1787), .b(wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_665), .o(n_1789) );
ao22s01 g66383_u0 ( .a(n_2046), .b(pci_target_unit_pci_target_if_target_rd_completed), .c(pciu_pciif_bckp_stop_in), .d(output_backup_devsel_out_reg_Q), .o(n_2765) );
ao22s01 g66384_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_968), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_661), .o(n_2105) );
ao22s01 g66385_u0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_962), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_655), .o(n_2104) );
ao22s02 g66386_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_948), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_641), .o(n_1788) );
ao22s01 g66387_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_958), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_651), .o(n_1786) );
ao22s01 g66388_u0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_945), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_638), .o(n_1785) );
ao22s02 g66389_u0 ( .a(n_2115), .b(conf_wb_err_addr_in_947), .c(FE_OFN1612_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_640), .o(n_2103) );
ao22s01 g66390_u0 ( .a(n_2115), .b(conf_wb_err_addr_in_970), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_663), .o(n_2102) );
ao22s02 g66391_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_950), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_643), .o(n_1784) );
ao22s02 g66393_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_964), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_657), .o(n_1782) );
ao22s02 g66394_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_952), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_645), .o(n_2101) );
ao22s01 g66395_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_954), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_647), .o(n_2100) );
ao22s02 g66396_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_955), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_648), .o(n_1781) );
in01s01 g66397_u0 ( .a(FE_OFN2095_n_2520), .o(g66397_sb) );
na02s01 TIMEBOOST_cell_40604 ( .a(TIMEBOOST_net_12540), .b(g62385_sb), .o(n_6830) );
na02f02 TIMEBOOST_cell_43736 ( .a(TIMEBOOST_net_14106), .b(FE_OFN1420_n_8567), .o(TIMEBOOST_net_12812) );
na02s01 TIMEBOOST_cell_32054 ( .a(configuration_pci_err_addr_500), .b(wbm_adr_o_30_), .o(TIMEBOOST_net_9938) );
in01s01 g66398_u0 ( .a(FE_OFN795_n_2520), .o(g66398_sb) );
na02s01 g66398_u2 ( .a(parchk_pci_ad_reg_in_1209), .b(FE_OFN795_n_2520), .o(g66398_db) );
na02s02 TIMEBOOST_cell_40606 ( .a(TIMEBOOST_net_12541), .b(g62972_sb), .o(n_5938) );
in01s01 g66399_u0 ( .a(n_2520), .o(g66399_sb) );
na02s02 TIMEBOOST_cell_43336 ( .a(TIMEBOOST_net_13906), .b(g62365_sb), .o(n_6871) );
na03f02 TIMEBOOST_cell_35253 ( .a(n_9043), .b(g57394_db), .c(g57394_sb), .o(n_10374) );
na02f02 TIMEBOOST_cell_45802 ( .a(TIMEBOOST_net_15139), .b(FE_OFN2185_n_8567), .o(TIMEBOOST_net_14577) );
na02s01 g66400_u2 ( .a(parchk_pci_ad_reg_in_1211), .b(FE_OFN795_n_2520), .o(g66400_db) );
na02s02 TIMEBOOST_cell_40684 ( .a(TIMEBOOST_net_12580), .b(g62891_sb), .o(n_6095) );
na03s02 TIMEBOOST_cell_40685 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__Q), .b(n_3585), .c(FE_OFN1253_n_4143), .o(TIMEBOOST_net_12581) );
na02s01 TIMEBOOST_cell_42709 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__Q), .b(FE_OFN1676_n_4655), .o(TIMEBOOST_net_13593) );
na02s01 TIMEBOOST_cell_40608 ( .a(TIMEBOOST_net_12542), .b(g62669_sb), .o(n_6200) );
in01s01 g66402_u0 ( .a(FE_OFN2096_n_2520), .o(g66402_sb) );
na03s02 TIMEBOOST_cell_40609 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__Q), .b(n_4448), .c(FE_OFN1213_n_4151), .o(TIMEBOOST_net_12543) );
na02m02 TIMEBOOST_cell_43737 ( .a(n_9888), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__Q), .o(TIMEBOOST_net_14107) );
na02s02 TIMEBOOST_cell_40610 ( .a(TIMEBOOST_net_12543), .b(g62464_sb), .o(n_6668) );
in01s01 g66403_u0 ( .a(FE_OFN2096_n_2520), .o(g66403_sb) );
na02s01 TIMEBOOST_cell_16024 ( .a(pci_target_unit_pci_target_if_norm_prf_en), .b(pciu_pref_en_in_320), .o(TIMEBOOST_net_3269) );
na02s02 TIMEBOOST_cell_39165 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_29__Q), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_412), .o(TIMEBOOST_net_11821) );
na02s01 TIMEBOOST_cell_16025 ( .a(TIMEBOOST_net_3269), .b(FE_OFN996_n_15366), .o(TIMEBOOST_net_790) );
na02s01 g66404_u2 ( .a(FE_OFN1780_parchk_pci_ad_reg_in_1221), .b(FE_OFN2096_n_2520), .o(g66404_db) );
na02s02 TIMEBOOST_cell_32053 ( .a(TIMEBOOST_net_9937), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4919) );
na02s02 TIMEBOOST_cell_40784 ( .a(TIMEBOOST_net_12630), .b(g62337_sb), .o(n_6924) );
na02f02 TIMEBOOST_cell_44676 ( .a(TIMEBOOST_net_14576), .b(g57230_sb), .o(n_11524) );
na02s02 TIMEBOOST_cell_45201 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__Q), .b(n_3651), .o(TIMEBOOST_net_14839) );
in01s01 g66406_u0 ( .a(FE_OFN2095_n_2520), .o(g66406_sb) );
na02s02 TIMEBOOST_cell_40786 ( .a(TIMEBOOST_net_12631), .b(g62662_sb), .o(n_6216) );
na02m02 TIMEBOOST_cell_38957 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_21__Q), .o(TIMEBOOST_net_11717) );
na02s02 TIMEBOOST_cell_40612 ( .a(TIMEBOOST_net_12544), .b(g62943_sb), .o(n_5995) );
na02m02 TIMEBOOST_cell_38959 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_3__Q), .o(TIMEBOOST_net_11718) );
na02s02 TIMEBOOST_cell_45004 ( .a(TIMEBOOST_net_14740), .b(g64215_db), .o(n_3954) );
na02s01 TIMEBOOST_cell_40614 ( .a(TIMEBOOST_net_12545), .b(g62951_sb), .o(n_5979) );
na02s01 g66408_u2 ( .a(FE_OFN1778_parchk_pci_ad_reg_in_1222), .b(FE_OFN2096_n_2520), .o(g66408_db) );
na03s02 TIMEBOOST_cell_43027 ( .a(n_3820), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__Q), .c(FE_OFN1119_g64577_p), .o(TIMEBOOST_net_13752) );
na02s01 TIMEBOOST_cell_16035 ( .a(TIMEBOOST_net_3274), .b(FE_OFN2094_n_2520), .o(n_2501) );
na02m02 TIMEBOOST_cell_38961 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_29__Q), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__Q), .o(TIMEBOOST_net_11719) );
na03s02 TIMEBOOST_cell_40615 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__Q), .b(n_3736), .c(FE_OFN1215_n_4151), .o(TIMEBOOST_net_12546) );
na02s01 TIMEBOOST_cell_32052 ( .a(configuration_pci_err_addr_491), .b(wbm_adr_o_21_), .o(TIMEBOOST_net_9937) );
na02s01 g66410_u2 ( .a(parchk_pci_ad_reg_in_1208), .b(FE_OFN795_n_2520), .o(g66410_db) );
na02s01 TIMEBOOST_cell_40616 ( .a(TIMEBOOST_net_12546), .b(g62448_sb), .o(n_6701) );
na03s02 TIMEBOOST_cell_43337 ( .a(n_4254), .b(FE_OFN1272_n_4096), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__Q), .o(TIMEBOOST_net_13907) );
na02s01 g66411_u2 ( .a(n_2648), .b(n_2520), .o(g66411_db) );
na02f02 TIMEBOOST_cell_40422 ( .a(TIMEBOOST_net_12449), .b(g54236_sb), .o(TIMEBOOST_net_10586) );
na02f04 TIMEBOOST_cell_40423 ( .a(n_15598), .b(n_16000), .o(TIMEBOOST_net_12450) );
na02s01 g66412_u2 ( .a(parchk_pci_ad_reg_in_1229), .b(n_2520), .o(g66412_db) );
na02f04 TIMEBOOST_cell_40424 ( .a(TIMEBOOST_net_12450), .b(FE_RN_435_0), .o(TIMEBOOST_net_4375) );
na02s01 TIMEBOOST_cell_16170 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__Q), .b(g65903_sb), .o(TIMEBOOST_net_3342) );
na02s01 g66413_u2 ( .a(n_8511), .b(n_2520), .o(g66413_db) );
na02s01 TIMEBOOST_cell_37852 ( .a(TIMEBOOST_net_11164), .b(g57988_sb), .o(n_9808) );
na02s01 TIMEBOOST_cell_16171 ( .a(TIMEBOOST_net_3342), .b(g65903_db), .o(n_2178) );
na02s01 g66414_u2 ( .a(parchk_pci_ad_reg_in_1214), .b(n_2520), .o(g66414_db) );
na02s01 TIMEBOOST_cell_40425 ( .a(conf_wb_err_addr_in_955), .b(configuration_wb_err_addr_546), .o(TIMEBOOST_net_12451) );
in01s01 g66415_u0 ( .a(FE_OFN795_n_2520), .o(g66415_sb) );
na02m02 TIMEBOOST_cell_38963 ( .a(wbu_sel_in_313), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_34__Q), .o(TIMEBOOST_net_11720) );
na02s02 TIMEBOOST_cell_32051 ( .a(TIMEBOOST_net_9936), .b(FE_OFN1183_n_3476), .o(TIMEBOOST_net_4918) );
na02s02 TIMEBOOST_cell_40618 ( .a(TIMEBOOST_net_12547), .b(g63183_sb), .o(n_5786) );
na02m02 TIMEBOOST_cell_38965 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_18__Q), .o(TIMEBOOST_net_11721) );
na03s02 TIMEBOOST_cell_40619 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__Q), .b(n_4289), .c(FE_OFN1283_n_4097), .o(TIMEBOOST_net_12548) );
na02s01 TIMEBOOST_cell_40426 ( .a(TIMEBOOST_net_12451), .b(FE_OFN1166_n_5615), .o(TIMEBOOST_net_11379) );
na02s01 g66417_u2 ( .a(parchk_pci_ad_reg_in_1206), .b(n_2520), .o(g66417_db) );
na02s01 TIMEBOOST_cell_40427 ( .a(TIMEBOOST_net_4363), .b(g54189_sb), .o(TIMEBOOST_net_12452) );
na02s02 TIMEBOOST_cell_40620 ( .a(TIMEBOOST_net_12548), .b(g62896_sb), .o(n_6085) );
na02s01 TIMEBOOST_cell_39325 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__Q), .b(FE_OFN1803_n_9690), .o(TIMEBOOST_net_11901) );
na02f02 TIMEBOOST_cell_44324 ( .a(TIMEBOOST_net_14400), .b(FE_OFN1387_n_8567), .o(TIMEBOOST_net_13408) );
na02m02 TIMEBOOST_cell_44627 ( .a(n_9671), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__Q), .o(TIMEBOOST_net_14552) );
na02s01 g66419_u2 ( .a(parchk_pci_ad_reg_in_1210), .b(n_2520), .o(g66419_db) );
na02s01 TIMEBOOST_cell_40428 ( .a(TIMEBOOST_net_12452), .b(g54189_db), .o(n_13358) );
na02s01 TIMEBOOST_cell_42710 ( .a(TIMEBOOST_net_13593), .b(n_4479), .o(TIMEBOOST_net_11893) );
na02s01 TIMEBOOST_cell_40503 ( .a(wishbone_slave_unit_pcim_sm_data_in_664), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__Q), .o(TIMEBOOST_net_12490) );
na02m02 TIMEBOOST_cell_42117 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__Q), .b(n_3508), .o(TIMEBOOST_net_13297) );
na02s01 TIMEBOOST_cell_16045 ( .a(TIMEBOOST_net_3279), .b(g63590_sb), .o(n_3315) );
na02s01 g66421_u2 ( .a(parchk_pci_ad_reg_in_1212), .b(FE_OFN795_n_2520), .o(g66421_db) );
na02s02 TIMEBOOST_cell_45123 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__Q), .b(FE_OFN1119_g64577_p), .o(TIMEBOOST_net_14800) );
na02s02 TIMEBOOST_cell_40788 ( .a(TIMEBOOST_net_12632), .b(g63000_sb), .o(n_5882) );
na02s01 TIMEBOOST_cell_40495 ( .a(wishbone_slave_unit_pcim_sm_data_in_637), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__Q), .o(TIMEBOOST_net_12486) );
na02s01 TIMEBOOST_cell_45562 ( .a(TIMEBOOST_net_15019), .b(FE_OFN217_n_9889), .o(n_9696) );
na02s01 g66423_u2 ( .a(parchk_pci_ad_reg_in_1213), .b(n_2520), .o(g66423_db) );
na02s02 TIMEBOOST_cell_30754 ( .a(g54160_sb), .b(wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_9288) );
na02s01 TIMEBOOST_cell_40622 ( .a(TIMEBOOST_net_12549), .b(g62579_sb), .o(n_6395) );
na02s01 TIMEBOOST_cell_40505 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__Q), .b(wishbone_slave_unit_pcim_sm_data_in_635), .o(TIMEBOOST_net_12491) );
na02m04 TIMEBOOST_cell_16050 ( .a(n_1481), .b(n_2914), .o(TIMEBOOST_net_3282) );
na02f02 TIMEBOOST_cell_40429 ( .a(g54312_db), .b(n_12595), .o(TIMEBOOST_net_12453) );
na02s02 TIMEBOOST_cell_40361 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(g65751_sb), .o(TIMEBOOST_net_12419) );
na02f02 TIMEBOOST_cell_40430 ( .a(TIMEBOOST_net_12453), .b(g54312_da), .o(n_13295) );
na02s01 TIMEBOOST_cell_40515 ( .a(wishbone_slave_unit_pcim_sm_data_in_638), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__Q), .o(TIMEBOOST_net_12496) );
na02s01 g66426_u2 ( .a(parchk_pci_ad_reg_in_1207), .b(n_2520), .o(g66426_db) );
na02f02 TIMEBOOST_cell_40974 ( .a(TIMEBOOST_net_12725), .b(g57412_sb), .o(n_11330) );
na03m02 TIMEBOOST_cell_34463 ( .a(n_13218), .b(FE_OFN2070_n_15978), .c(TIMEBOOST_net_9896), .o(n_13512) );
na02s01 g66427_u2 ( .a(n_3030), .b(n_2520), .o(g66427_db) );
na02m02 TIMEBOOST_cell_41655 ( .a(n_1628), .b(n_1384), .o(TIMEBOOST_net_13066) );
na02s01 TIMEBOOST_cell_32050 ( .a(configuration_pci_err_addr_471), .b(wbm_adr_o_1_), .o(TIMEBOOST_net_9936) );
na02m04 TIMEBOOST_cell_16051 ( .a(n_1619), .b(TIMEBOOST_net_3282), .o(TIMEBOOST_net_506) );
na02s02 TIMEBOOST_cell_32049 ( .a(TIMEBOOST_net_9935), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_4917) );
na02m02 TIMEBOOST_cell_38967 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_28__Q), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__Q), .o(TIMEBOOST_net_11722) );
na02s02 TIMEBOOST_cell_45124 ( .a(TIMEBOOST_net_14800), .b(n_3875), .o(TIMEBOOST_net_4637) );
na02s01 TIMEBOOST_cell_32048 ( .a(configuration_pci_err_addr_488), .b(wbm_adr_o_18_), .o(TIMEBOOST_net_9935) );
na02f02 TIMEBOOST_cell_39125 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_10182), .o(TIMEBOOST_net_11801) );
na02s02 TIMEBOOST_cell_40790 ( .a(TIMEBOOST_net_12633), .b(g62975_sb), .o(n_5932) );
in01s01 g66433_u0 ( .a(pci_target_unit_del_sync_req_done_reg), .o(g66433_sb) );
na02s01 g66433_u1 ( .a(pci_target_unit_del_sync_sync_req_comp_pending), .b(g66433_sb), .o(g66433_da) );
na02s01 g66433_u2 ( .a(pci_target_unit_del_sync_req_comp_pending), .b(pci_target_unit_del_sync_req_done_reg), .o(g66433_db) );
na02s01 g66433_u3 ( .a(g66433_da), .b(g66433_db), .o(n_1533) );
oa12s01 g66454_u0 ( .a(n_944), .b(n_1334), .c(n_1263), .o(n_1335) );
in01s01 g66456_u0 ( .a(n_325), .o(g66456_sb) );
no02m02 TIMEBOOST_cell_45563 ( .a(FE_RN_582_0), .b(FE_RN_581_0), .o(TIMEBOOST_net_15020) );
na02s01 g66456_u2 ( .a(wishbone_slave_unit_del_sync_req_comp_pending), .b(n_325), .o(g66456_db) );
na02f02 TIMEBOOST_cell_40976 ( .a(TIMEBOOST_net_12726), .b(g57503_sb), .o(n_11235) );
in01m01 g66457_u0 ( .a(pci_target_unit_pci_target_sm_n_3), .o(g66457_sb) );
na02s01 TIMEBOOST_cell_42713 ( .a(n_3783), .b(g64958_sb), .o(TIMEBOOST_net_13595) );
na02s02 g66457_u2 ( .a(pci_target_unit_pci_target_sm_n_3), .b(pci_target_unit_pci_target_sm_n_2), .o(g66457_db) );
na02m02 TIMEBOOST_cell_42521 ( .a(TIMEBOOST_net_6393), .b(wbu_addr_in_265), .o(TIMEBOOST_net_13499) );
no02s01 g66458_u0 ( .a(wbm_adr_o_2_), .b(wbm_adr_o_3_), .o(g66458_p0) );
ao12s01 g66458_u1 ( .a(g66458_p0), .b(wbm_adr_o_2_), .c(wbm_adr_o_3_), .o(n_740) );
na02s10 g66458_u2 ( .a(wbm_adr_o_3_), .b(wbm_adr_o_2_), .o(g66458_p) );
in01m06 g66458_u3 ( .a(g66458_p), .o(n_1674) );
no02s01 g66459_u0 ( .a(wbu_addr_in_252), .b(wbu_addr_in_251), .o(g66459_p0) );
ao12s01 g66459_u1 ( .a(g66459_p0), .b(wbu_addr_in_252), .c(wbu_addr_in_251), .o(n_739) );
in01s01 g66462_u0 ( .a(n_16030), .o(n_1133) );
no02s04 g66464_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(g66464_p0) );
ao12s02 g66464_u1 ( .a(g66464_p0), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q), .c(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(n_1225) );
na02s06 g66464_u2 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(g66464_p) );
in01s01 g66464_u3 ( .a(g66464_p), .o(n_1224) );
no02s01 g66465_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_), .o(g66465_p0) );
ao12s01 g66465_u1 ( .a(g66465_p0), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_), .o(n_741) );
na02s04 g66465_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_), .o(g66465_p) );
in01s02 g66465_u3 ( .a(g66465_p), .o(n_1418) );
in01m08 g66467_u0 ( .a(n_568), .o(n_1413) );
in01s01 g66470_u0 ( .a(n_1011), .o(n_1175) );
in01s01 g66471_u0 ( .a(n_947), .o(n_566) );
in01s01 g66472_u0 ( .a(n_948), .o(n_733) );
no02s02 g66473_u0 ( .a(n_1332), .b(n_540), .o(g66473_p) );
ao12s02 g66473_u1 ( .a(g66473_p), .b(n_1332), .c(n_540), .o(n_1333) );
no02s02 g66475_u0 ( .a(n_1330), .b(n_558), .o(g66475_p) );
ao12s02 g66475_u1 ( .a(g66475_p), .b(n_1330), .c(n_558), .o(n_1331) );
ao22s01 g66476_u0 ( .a(n_76), .b(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_), .d(n_816), .o(n_1329) );
na02s02 g66477_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__Q), .b(FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source), .o(g66477_da) );
na02s02 g66477_u2 ( .a(n_235), .b(wishbone_slave_unit_pci_initiator_if_data_source), .o(g66477_db) );
na02s02 g66477_u3 ( .a(g66477_da), .b(g66477_db), .o(n_5641) );
in01s01 g66479_u0 ( .a(wishbone_slave_unit_pci_initiator_if_write_req_int), .o(n_1780) );
in01s01 g66483_u0 ( .a(wishbone_slave_unit_del_sync_req_rty_exp_reg), .o(n_1327) );
in01s01 g66497_u0 ( .a(pci_target_unit_del_sync_req_rty_exp_reg), .o(n_249) );
in01s01 g66536_u0 ( .a(pci_target_unit_del_sync_comp_done_reg_main), .o(n_2146) );
in01s01 g66542_u0 ( .a(n_1325), .o(n_1326) );
no02m04 g66543_u0 ( .a(n_943), .b(n_288), .o(n_1325) );
na02m04 g66544_u0 ( .a(n_1107), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(g66544_p) );
in01m02 g66544_u1 ( .a(g66544_p), .o(n_908) );
no02s03 g66547_u0 ( .a(n_914), .b(n_1174), .o(g66547_p) );
in01s02 g66547_u1 ( .a(g66547_p), .o(n_1699) );
no02s02 g66548_u0 ( .a(n_1468), .b(output_backup_trdy_out_reg_Q), .o(n_1126) );
no02f20 g66549_u0 ( .a(n_412), .b(wishbone_slave_unit_wishbone_slave_img_hit_2_), .o(n_931) );
na02s01 g66550_u0 ( .a(n_1173), .b(wishbone_slave_unit_fifos_wbw_whole_waddr), .o(g66550_p) );
in01s01 g66550_u1 ( .a(g66550_p), .o(n_905) );
in01f01 g66551_u0 ( .a(n_1779), .o(n_7622) );
in01f02 g66552_u0 ( .a(n_15055), .o(n_1779) );
na02s02 g66554_u0 ( .a(n_929), .b(n_1263), .o(n_930) );
no02s01 g66555_u0 ( .a(n_2483), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(n_2999) );
no02s06 g66556_u0 ( .a(n_560), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_6_), .o(n_1715) );
no02s02 g66577_u0 ( .a(n_748), .b(wbs_adr_i_4_), .o(g66577_p) );
in01s01 g66577_u1 ( .a(g66577_p), .o(n_1666) );
na02s06 g66579_u0 ( .a(n_1317), .b(n_1293), .o(n_4736) );
no02m02 g66580_u0 ( .a(n_1334), .b(n_221), .o(n_1437) );
in01s01 g66581_u0 ( .a(n_1124), .o(n_1125) );
na02s02 g66582_u0 ( .a(n_937), .b(pci_target_unit_del_sync_comp_cycle_count_7_), .o(n_1124) );
na02s02 g66583_u0 ( .a(n_1294), .b(n_1316), .o(g66583_p) );
in01m02 g66583_u1 ( .a(g66583_p), .o(n_4727) );
na02s06 g66584_u0 ( .a(n_1318), .b(n_1174), .o(g66584_p) );
in01s06 g66584_u1 ( .a(g66584_p), .o(n_2299) );
in01s01 g66585_u0 ( .a(n_1122), .o(n_1123) );
na02s02 g66586_u0 ( .a(n_928), .b(wishbone_slave_unit_del_sync_comp_cycle_count_7_), .o(n_1122) );
in01f04 g66590_u0 ( .a(n_1808), .o(n_4874) );
na02f06 g66591_u0 ( .a(n_993), .b(n_1104), .o(n_1808) );
no02s04 g66592_u0 ( .a(n_915), .b(n_924), .o(n_2872) );
no02s06 g66593_u0 ( .a(n_921), .b(n_900), .o(n_1229) );
no02s06 g66594_u0 ( .a(n_927), .b(n_909), .o(n_1381) );
no02s06 g66595_u0 ( .a(n_926), .b(n_901), .o(n_2756) );
na02s01 g66596_u0 ( .a(configuration_sync_isr_2_delayed_del_bit), .b(configuration_sync_isr_2_sync_del_bit), .o(n_925) );
no02s04 g66597_u0 ( .a(n_877), .b(n_902), .o(n_1480) );
no02f02 g66598_u0 ( .a(n_16291), .b(n_16544), .o(n_2560) );
no02s08 g66599_u0 ( .a(wishbone_slave_unit_del_sync_comp_flush_out), .b(wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg_Q), .o(n_9941) );
in01f02 g66600_u0 ( .a(n_2553), .o(n_2331) );
in01f06 g66602_u0 ( .a(n_2094), .o(n_2553) );
in01f04 g66603_u0 ( .a(n_1777), .o(n_2094) );
na02f08 g66604_u0 ( .a(n_15275), .b(n_15231), .o(n_1777) );
no02s06 g66605_u0 ( .a(n_895), .b(n_904), .o(n_2428) );
na02s01 g66607_u0 ( .a(n_257), .b(n_432), .o(g66607_p) );
in01s02 g66607_u1 ( .a(g66607_p), .o(n_1624) );
na02s01 g66608_u0 ( .a(n_15365), .b(parity_checker_frame_dec2), .o(n_3020) );
no02s06 g66612_u0 ( .a(n_924), .b(n_518), .o(n_2929) );
no02s01 g66613_u0 ( .a(n_2597), .b(n_1774), .o(n_2599) );
no02s01 g66614_u0 ( .a(n_1084), .b(configuration_isr_bit_2975), .o(n_1120) );
no02s08 g66615_u0 ( .a(n_917), .b(n_923), .o(n_2411) );
no02m04 g66616_u0 ( .a(pci_target_unit_pci_target_sm_n_3), .b(n_976), .o(n_922) );
no02s03 g66617_u0 ( .a(n_921), .b(n_911), .o(n_2235) );
no02s02 g66620_u0 ( .a(n_1009), .b(n_1005), .o(g66620_p) );
in01s02 g66620_u1 ( .a(g66620_p), .o(n_4501) );
no02s01 g66621_u0 ( .a(n_16867), .b(n_15680), .o(n_1322) );
no02s02 g66627_u0 ( .a(n_1005), .b(n_538), .o(g66627_p) );
in01s04 g66627_u1 ( .a(g66627_p), .o(n_4490) );
na02s03 g66628_u0 ( .a(n_1118), .b(n_1174), .o(g66628_p) );
in01s02 g66628_u1 ( .a(g66628_p), .o(n_2053) );
in01s01 g66630_u0 ( .a(n_1269), .o(n_1119) );
no02m06 g66631_u0 ( .a(n_886), .b(n_891), .o(n_1269) );
no02s04 g66632_u0 ( .a(n_920), .b(n_919), .o(n_2305) );
no02s06 g66633_u0 ( .a(n_894), .b(n_918), .o(n_1390) );
no02m04 g66634_u0 ( .a(n_956), .b(n_927), .o(n_2237) );
no02s03 g66636_u0 ( .a(n_910), .b(n_941), .o(n_2426) );
no02s04 g66637_u0 ( .a(n_917), .b(n_916), .o(n_1968) );
na02s06 g66638_u0 ( .a(n_1318), .b(n_1117), .o(n_2292) );
in01s01 g66639_u0 ( .a(n_1523), .o(n_1524) );
no02m02 g66640_u0 ( .a(n_790), .b(wishbone_slave_unit_wishbone_slave_c_state), .o(n_1523) );
no02s02 g66641_u0 ( .a(n_888), .b(n_939), .o(n_940) );
na02s03 g66642_u0 ( .a(n_1118), .b(n_1117), .o(n_2047) );
na02f02 TIMEBOOST_cell_42227 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__Q), .b(n_9082), .o(TIMEBOOST_net_13352) );
no02s06 g66644_u0 ( .a(n_916), .b(n_915), .o(n_1227) );
no02s06 g66645_u0 ( .a(n_914), .b(n_1117), .o(n_2248) );
na02f04 g66646_u0 ( .a(n_912), .b(n_913), .o(g66646_p) );
in01f02 g66646_u1 ( .a(g66646_p), .o(n_1481) );
no02s04 g66647_u0 ( .a(n_911), .b(n_910), .o(n_1228) );
no02m02 g66648_u0 ( .a(n_563), .b(n_977), .o(n_1116) );
na02s02 g66649_u0 ( .a(n_1188), .b(n_1115), .o(g66649_p) );
in01s02 g66649_u1 ( .a(g66649_p), .o(n_9528) );
na02s06 g66650_u0 ( .a(n_1317), .b(n_1316), .o(g66650_p) );
in01s06 g66650_u1 ( .a(g66650_p), .o(n_4725) );
no02s03 g66651_u0 ( .a(n_909), .b(n_892), .o(n_2427) );
na02s04 g66652_u0 ( .a(n_1115), .b(n_1290), .o(g66652_p) );
in01s04 g66652_u1 ( .a(g66652_p), .o(n_9502) );
na02s04 g66653_u0 ( .a(n_1288), .b(n_1315), .o(n_9697) );
in01s01 g66655_u0 ( .a(FE_OCPN1875_n_14526), .o(n_1522) );
na02s06 g66658_u0 ( .a(n_1509), .b(n_1210), .o(g66658_p) );
in01s08 g66658_u1 ( .a(g66658_p), .o(n_4669) );
in01f04 g66660_u0 ( .a(n_2127), .o(n_2341) );
na02f06 g66661_u0 ( .a(n_15275), .b(n_15756), .o(n_2127) );
na02s01 g66662_u0 ( .a(n_2763), .b(n_653), .o(g66662_p) );
in01s01 g66662_u1 ( .a(g66662_p), .o(n_2764) );
no02f04 g66663_u0 ( .a(n_16033), .b(n_1291), .o(g66663_p) );
in01f02 g66663_u1 ( .a(g66663_p), .o(n_2126) );
no02s08 g66664_u0 ( .a(n_881), .b(n_885), .o(n_1270) );
in01f04 g66667_u0 ( .a(n_16151), .o(n_2215) );
no02s04 g66669_u0 ( .a(n_1316), .b(n_980), .o(g66669_p) );
in01s04 g66669_u1 ( .a(g66669_p), .o(n_16657) );
no02m01 g66670_u0 ( .a(n_1334), .b(n_906), .o(n_907) );
no02m08 g66671_u0 ( .a(n_884), .b(n_946), .o(n_2306) );
no02m02 g66672_u0 ( .a(n_1316), .b(n_813), .o(g66672_p) );
in01m02 g66672_u1 ( .a(g66672_p), .o(n_4740) );
in01f20 g66701_u0 ( .a(FE_OFN2214_n_15366), .o(n_2301) );
na02s04 g66710_u0 ( .a(n_1289), .b(n_1315), .o(n_9690) );
na02s04 g66711_u0 ( .a(n_1115), .b(n_1315), .o(n_9902) );
no02s06 g66712_u0 ( .a(n_903), .b(n_904), .o(n_1409) );
no02s04 g66713_u0 ( .a(n_902), .b(n_889), .o(n_2681) );
na02f02 g66714_u0 ( .a(n_1198), .b(n_1519), .o(g66714_p) );
in01f02 g66714_u1 ( .a(g66714_p), .o(n_2795) );
no02s04 g66715_u0 ( .a(n_900), .b(n_901), .o(n_2433) );
no02s04 g66716_u0 ( .a(n_899), .b(n_896), .o(n_1373) );
na02s01 g66717_u0 ( .a(n_1334), .b(n_1263), .o(n_944) );
na02f40 g66724_u0 ( .a(n_898), .b(wbm_ack_i), .o(n_1998) );
na02s10 g66726_u0 ( .a(n_791), .b(pci_target_unit_pci_target_sm_master_will_request_read), .o(g66726_p) );
in01s04 g66726_u1 ( .a(g66726_p), .o(n_1824) );
na02f04 g66727_u0 ( .a(n_16867), .b(n_15680), .o(n_1306) );
na02m02 g66728_u0 ( .a(n_1113), .b(n_1107), .o(g66728_p) );
in01m02 g66728_u1 ( .a(g66728_p), .o(n_4655) );
in01m04 g66732_u0 ( .a(n_1435), .o(n_9175) );
na03f40 g66733_u0 ( .a(n_61), .b(pci_target_unit_pci_target_sm_n_2), .c(n_278), .o(n_1435) );
in01s01 g66734_u0 ( .a(n_1304), .o(n_9178) );
na02s02 g66735_u0 ( .a(n_520), .b(n_1628), .o(n_1304) );
no02m06 g66736_u0 ( .a(n_896), .b(n_897), .o(n_2463) );
na02s02 g66737_u0 ( .a(n_2609), .b(n_2742), .o(g66737_p) );
in01s02 g66737_u1 ( .a(g66737_p), .o(n_3222) );
na02m04 g66738_u0 ( .a(n_534), .b(n_912), .o(g66738_p) );
in01m02 g66738_u1 ( .a(g66738_p), .o(n_2982) );
na02s01 g66739_u0 ( .a(FE_OFN1612_n_2122), .b(n_1111), .o(n_1112) );
na02s04 g66742_u0 ( .a(n_1173), .b(n_1288), .o(g66742_p) );
in01s04 g66742_u1 ( .a(g66742_p), .o(n_9428) );
no02f06 g66743_u0 ( .a(n_1519), .b(n_1197), .o(n_1813) );
no02s04 g66744_u0 ( .a(n_945), .b(n_946), .o(n_1282) );
oa12s01 g66745_u0 ( .a(n_1109), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .c(n_8953), .o(n_1110) );
na02s01 g66746_u0 ( .a(FE_OFN1612_n_2122), .b(wishbone_slave_unit_pcim_sm_be_in_558), .o(n_1108) );
no02s08 g66749_u0 ( .a(n_895), .b(n_890), .o(n_3007) );
in01s01 g66751_u0 ( .a(n_6943), .o(n_2134) );
na02f06 g66752_u0 ( .a(n_1432), .b(wishbone_slave_unit_wishbone_slave_c_state_2), .o(g66752_p) );
in01f06 g66752_u1 ( .a(g66752_p), .o(n_6943) );
na02s04 g66753_u0 ( .a(n_1195), .b(n_1107), .o(g66753_p) );
in01m04 g66753_u1 ( .a(g66753_p), .o(n_4671) );
no02s08 g66754_u0 ( .a(n_956), .b(n_957), .o(n_3194) );
no02s04 g66755_u0 ( .a(n_894), .b(n_893), .o(n_1478) );
na02s04 g66756_u0 ( .a(n_1188), .b(n_1440), .o(n_9692) );
no02m02 g66757_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q), .b(n_1014), .o(n_1299) );
na02s04 g66758_u0 ( .a(n_1194), .b(n_1195), .o(n_4392) );
na02s03 g66759_u0 ( .a(n_1017), .b(n_1316), .o(g66759_p) );
in01s04 g66759_u1 ( .a(g66759_p), .o(n_4730) );
no02s06 g66760_u0 ( .a(n_892), .b(n_512), .o(n_3192) );
na02s04 g66761_u0 ( .a(n_1106), .b(n_1107), .o(n_4409) );
in01m01 g66765_u0 ( .a(n_1514), .o(n_1515) );
na02s01 TIMEBOOST_cell_17965 ( .a(TIMEBOOST_net_4239), .b(g65381_da), .o(n_4646) );
no02s06 g66768_u0 ( .a(n_887), .b(n_945), .o(n_2755) );
na02s01 g66769_u0 ( .a(FE_OFN1612_n_2122), .b(wishbone_slave_unit_pcim_sm_be_in_557), .o(n_1105) );
na02s06 g66770_u0 ( .a(n_1290), .b(n_1440), .o(n_9694) );
na02m06 g66771_u0 ( .a(n_16307), .b(n_1774), .o(n_1513) );
no02m06 g66772_u0 ( .a(n_891), .b(n_890), .o(n_2228) );
na02s04 g66773_u0 ( .a(n_1210), .b(n_1201), .o(g66773_p) );
in01m06 g66773_u1 ( .a(g66773_p), .o(n_4677) );
no02s06 g66774_u0 ( .a(n_941), .b(n_549), .o(n_1355) );
no02f06 g66775_u0 ( .a(n_992), .b(n_1104), .o(n_3310) );
na02s06 g66776_u0 ( .a(n_1103), .b(n_1117), .o(n_2055) );
na02s02 g66777_u0 ( .a(n_1173), .b(n_1289), .o(g66777_p) );
in01m02 g66777_u1 ( .a(g66777_p), .o(n_9477) );
no02f04 g66778_u0 ( .a(n_893), .b(n_874), .o(n_964) );
no02s01 g66779_u0 ( .a(n_1739), .b(n_2078), .o(n_2329) );
na02s06 g66780_u0 ( .a(n_1294), .b(n_1293), .o(n_4734) );
no02s04 g66781_u0 ( .a(n_889), .b(n_888), .o(n_2705) );
in01f10 g66783_u0 ( .a(n_1366), .o(n_1196) );
na02f20 g66784_u0 ( .a(n_976), .b(pci_target_unit_pci_target_sm_n_3), .o(n_1366) );
na02s04 g66785_u0 ( .a(n_1315), .b(n_1440), .o(n_9687) );
no02s04 g66786_u0 ( .a(n_530), .b(n_903), .o(n_965) );
no02s04 g66787_u0 ( .a(n_745), .b(n_746), .o(n_2475) );
na02s04 g66788_u0 ( .a(n_1194), .b(n_1210), .o(n_4497) );
na02s03 g66789_u0 ( .a(n_1103), .b(n_1174), .o(g66789_p) );
in01s03 g66789_u1 ( .a(g66789_p), .o(n_2037) );
in01s02 g66794_u0 ( .a(n_1445), .o(n_2214) );
na02s01 g66796_u0 ( .a(FE_OFN1612_n_2122), .b(wishbone_slave_unit_pcim_sm_be_in_559), .o(n_1202) );
in01s01 g66797_u0 ( .a(n_1758), .o(n_1759) );
no02s01 g66798_u0 ( .a(n_1512), .b(n_1505), .o(n_1758) );
no02m06 g66799_u0 ( .a(n_899), .b(n_923), .o(n_2596) );
no02s01 g66800_u0 ( .a(n_2031), .b(output_backup_trdy_out_reg_Q), .o(n_2280) );
no02s01 g66801_u0 ( .a(n_2031), .b(n_15302), .o(n_2729) );
no02m06 g66802_u0 ( .a(n_745), .b(n_533), .o(n_2914) );
no02s06 g66803_u0 ( .a(n_887), .b(n_957), .o(n_2431) );
na02f02 TIMEBOOST_cell_42228 ( .a(TIMEBOOST_net_13352), .b(FE_OFN1394_n_8567), .o(TIMEBOOST_net_12304) );
na02m02 g66805_u0 ( .a(n_812), .b(n_1316), .o(g66805_p) );
in01m02 g66805_u1 ( .a(g66805_p), .o(n_4732) );
in01f01 g66807_u0 ( .a(n_15065), .o(n_2449) );
in01f01 g66811_u0 ( .a(n_1447), .o(n_1448) );
no02f01 g66812_u0 ( .a(n_1200), .b(n_681), .o(n_1447) );
na02s04 g66813_u0 ( .a(n_1210), .b(n_1107), .o(g66813_p) );
in01s04 g66813_u1 ( .a(g66813_p), .o(n_4508) );
na02s08 g66814_u0 ( .a(n_1173), .b(n_1440), .o(n_9904) );
in01m01 g66820_u0 ( .a(n_15370), .o(n_1684) );
na02s08 g66822_u0 ( .a(n_1113), .b(n_1194), .o(n_4460) );
no02f04 g66823_u0 ( .a(n_16291), .b(FE_OCPN1868_n_16289), .o(n_1446) );
na02s02 TIMEBOOST_cell_43102 ( .a(TIMEBOOST_net_13789), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_12056) );
no02m01 g66825_u0 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(n_2685), .o(g66825_p) );
in01s02 g66825_u1 ( .a(g66825_p), .o(n_3480) );
no02s06 g66826_u0 ( .a(n_897), .b(n_977), .o(n_1374) );
na02s01 g66827_u0 ( .a(n_1347), .b(n_16816), .o(g66827_p) );
in01s01 g66827_u1 ( .a(g66827_p), .o(n_1101) );
na02s04 g66829_u0 ( .a(n_1106), .b(n_1201), .o(n_4454) );
na02s01 g66830_u0 ( .a(n_1774), .b(n_5755), .o(n_1100) );
no02m06 g66831_u0 ( .a(n_886), .b(n_885), .o(n_2435) );
no02s04 g66832_u0 ( .a(n_926), .b(n_920), .o(n_1241) );
in01s08 g66852_u0 ( .a(n_2494), .o(n_2493) );
in01m06 g66853_u0 ( .a(n_2344), .o(n_2494) );
na02m20 g66854_u0 ( .a(n_1459), .b(wishbone_slave_unit_pci_initiator_sm_mabort1), .o(g66854_p) );
in01f10 g66854_u1 ( .a(g66854_p), .o(n_2344) );
no02m06 g66855_u0 ( .a(n_1221), .b(n_2742), .o(n_2028) );
na02s04 g66856_u0 ( .a(n_1115), .b(n_1173), .o(g66856_p) );
in01f02 g66856_u1 ( .a(g66856_p), .o(n_9531) );
no02s06 g66857_u0 ( .a(n_528), .b(n_746), .o(n_1442) );
na02m02 g66858_u0 ( .a(FE_OFN1612_n_2122), .b(wishbone_slave_unit_pcim_sm_data_in_635), .o(n_1099) );
na02s04 g66859_u0 ( .a(n_1289), .b(n_1290), .o(n_9864) );
in01f08 g66861_u0 ( .a(n_16001), .o(n_2453) );
na02s06 g66864_u0 ( .a(n_1509), .b(n_1113), .o(n_4417) );
no02m06 g66865_u0 ( .a(n_430), .b(n_884), .o(n_1415) );
no02s01 g66866_u0 ( .a(n_1201), .b(n_1509), .o(g66866_p) );
in01s01 g66866_u1 ( .a(g66866_p), .o(n_1510) );
no02s06 g66868_u0 ( .a(n_374), .b(n_956), .o(n_1378) );
na03s01 TIMEBOOST_cell_33226 ( .a(g65420_da), .b(g65420_db), .c(n_12), .o(TIMEBOOST_net_5437) );
ao12s01 g66870_u0 ( .a(n_1175), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_0_), .c(wishbone_slave_unit_pci_initiator_sm_latency_timer_1_), .o(n_1098) );
na02s04 g66871_u0 ( .a(n_1290), .b(n_1288), .o(n_9899) );
ao12s01 g66872_u0 ( .a(n_987), .b(pci_target_unit_wishbone_master_read_count_1_), .c(pci_target_unit_wishbone_master_read_count_0_), .o(n_988) );
na02s01 TIMEBOOST_cell_43272 ( .a(TIMEBOOST_net_13874), .b(FE_OFN1194_n_6935), .o(TIMEBOOST_net_12530) );
no02s06 g66874_u0 ( .a(n_881), .b(n_232), .o(n_1388) );
no02s01 g66875_u0 ( .a(n_1188), .b(n_1290), .o(g66875_p) );
in01s01 g66875_u1 ( .a(g66875_p), .o(n_1287) );
na02f04 g66876_u0 ( .a(n_411), .b(n_1165), .o(g66876_p) );
in01f04 g66876_u1 ( .a(g66876_p), .o(n_1966) );
na02s02 TIMEBOOST_cell_43103 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__Q), .b(n_4468), .o(TIMEBOOST_net_13790) );
na02m02 TIMEBOOST_cell_42229 ( .a(n_9513), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__Q), .o(TIMEBOOST_net_13353) );
na02s04 g66879_u0 ( .a(n_1113), .b(n_1201), .o(n_4438) );
na02s04 g66880_u0 ( .a(n_1509), .b(n_1195), .o(n_4495) );
ao12s01 g66881_u0 ( .a(n_16860), .b(n_696), .c(n_2092), .o(n_1686) );
na02m04 g66882_u0 ( .a(n_1195), .b(n_1201), .o(n_4505) );
ao12s01 g66883_u0 ( .a(n_703), .b(wishbone_slave_unit_pci_initiator_if_read_count_0_), .c(wishbone_slave_unit_pci_initiator_if_read_count_1_), .o(n_990) );
in01s01 g66884_u0 ( .a(n_2088), .o(n_2328) );
ao12s01 g66885_u0 ( .a(n_2087), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q), .c(n_1041), .o(n_2088) );
no02m04 g66886_u0 ( .a(n_306), .b(n_885), .o(n_1482) );
no02s04 g66887_u0 ( .a(n_918), .b(n_404), .o(n_1479) );
na02m04 g66888_u0 ( .a(n_994), .b(n_375), .o(g66888_p) );
in01m02 g66888_u1 ( .a(g66888_p), .o(n_1357) );
na02m04 g66889_u0 ( .a(n_331), .b(n_994), .o(g66889_p) );
in01m02 g66889_u1 ( .a(g66889_p), .o(n_1414) );
na02s01 g66890_u0 ( .a(n_1283), .b(n_817), .o(n_1284) );
ao12s01 g66891_u0 ( .a(n_546), .b(wishbone_slave_unit_pci_initiator_sm_decode_count_0_), .c(wishbone_slave_unit_pci_initiator_sm_decode_count_1_), .o(n_1204) );
no02s02 g66892_u0 ( .a(n_524), .b(n_939), .o(n_1096) );
na02f02 TIMEBOOST_cell_42230 ( .a(TIMEBOOST_net_13353), .b(FE_OFN1384_n_8567), .o(TIMEBOOST_net_12310) );
ao12s01 g66894_u0 ( .a(n_2046), .b(parchk_pci_trdy_reg_in), .c(pciu_pciif_stop_reg_in), .o(n_2086) );
na02s02 TIMEBOOST_cell_43104 ( .a(TIMEBOOST_net_13790), .b(FE_OFN1285_n_4097), .o(TIMEBOOST_net_12540) );
no02s04 g66896_u0 ( .a(n_304), .b(n_877), .o(n_1971) );
no02s06 g66897_u0 ( .a(n_191), .b(n_957), .o(n_2967) );
ao12s02 g66899_u0 ( .a(pci_target_unit_del_sync_bc_in_203), .b(pci_target_unit_pci_target_if_norm_prf_en), .c(pci_target_unit_del_sync_bc_in_202), .o(n_639) );
no02m04 g66900_u0 ( .a(n_350), .b(n_874), .o(n_1361) );
na02s04 g66901_u0 ( .a(n_1188), .b(n_1288), .o(n_9823) );
no02s01 g66902_u0 ( .a(n_1118), .b(n_1103), .o(g66902_p) );
in01s01 g66902_u1 ( .a(g66902_p), .o(n_7569) );
in01f02 g66903_u0 ( .a(n_1507), .o(n_1508) );
no02f08 g66905_u0 ( .a(n_1221), .b(n_1408), .o(n_2129) );
ao12s02 g66906_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_mabort2), .b(wishbone_slave_unit_pci_initiator_sm_mabort1), .c(wbu_pciif_frame_out_in), .o(n_2803) );
na02s04 g66908_u0 ( .a(n_1188), .b(n_1289), .o(n_9895) );
no02m04 g66909_u0 ( .a(n_405), .b(n_919), .o(n_1412) );
no02s01 g66911_u0 ( .a(pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q), .b(n_996), .o(g66911_p) );
ao12s01 g66911_u1 ( .a(g66911_p), .b(pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q), .c(n_996), .o(n_998) );
no02s01 g66912_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_695), .b(parchk_pci_ad_reg_in_1214), .o(g66912_p) );
ao12s01 g66912_u1 ( .a(g66912_p), .b(pci_target_unit_pcit_if_strd_addr_in_695), .c(parchk_pci_ad_reg_in_1214), .o(n_641) );
no02s02 g66913_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_22__Q), .b(wbu_addr_in_271), .o(g66913_p) );
ao12s02 g66913_u1 ( .a(g66913_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_22__Q), .c(wbu_addr_in_271), .o(n_999) );
no02s01 g66915_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_713), .b(parchk_pci_ad_reg_in_1232), .o(g66915_p) );
ao12s01 g66915_u1 ( .a(g66915_p), .b(pci_target_unit_pcit_if_strd_addr_in_713), .c(parchk_pci_ad_reg_in_1232), .o(n_640) );
ao12f10 g66916_u0 ( .a(n_341), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_2_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_), .o(n_872) );
no02s01 g66917_u0 ( .a(pci_target_unit_pcit_if_strd_bc_in_718), .b(n_2648), .o(g66917_p) );
ao12s01 g66917_u1 ( .a(g66917_p), .b(pci_target_unit_pcit_if_strd_bc_in_718), .c(n_2648), .o(n_2036) );
no02s01 g66918_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_712), .b(parchk_pci_ad_reg_in_1231), .o(g66918_p) );
ao12s01 g66918_u1 ( .a(g66918_p), .b(pci_target_unit_pcit_if_strd_addr_in_712), .c(parchk_pci_ad_reg_in_1231), .o(n_627) );
ao22s01 g66920_u0 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_1_), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_0_), .c(n_345), .d(n_425), .o(n_1095) );
no02s01 g66921_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_714), .b(parchk_pci_ad_reg_in_1233), .o(g66921_p) );
ao12s01 g66921_u1 ( .a(g66921_p), .b(pci_target_unit_pcit_if_strd_addr_in_714), .c(parchk_pci_ad_reg_in_1233), .o(n_695) );
no02s01 g66922_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_710), .b(parchk_pci_ad_reg_in_1229), .o(g66922_p) );
ao12s01 g66922_u1 ( .a(g66922_p), .b(pci_target_unit_pcit_if_strd_addr_in_710), .c(parchk_pci_ad_reg_in_1229), .o(n_626) );
no02s02 g66923_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_16__Q), .b(wbu_addr_in_265), .o(g66923_p) );
ao12s02 g66923_u1 ( .a(g66923_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_16__Q), .c(wbu_addr_in_265), .o(n_871) );
no02s01 g66924_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_706), .b(parchk_pci_ad_reg_in_1225), .o(g66924_p) );
ao12s01 g66924_u1 ( .a(g66924_p), .b(pci_target_unit_pcit_if_strd_addr_in_706), .c(parchk_pci_ad_reg_in_1225), .o(n_700) );
no02s02 g66925_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_6__Q), .b(wbu_addr_in_255), .o(g66925_p) );
ao12s02 g66925_u1 ( .a(g66925_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_6__Q), .c(wbu_addr_in_255), .o(n_1004) );
ao12f08 g66926_u0 ( .a(n_342), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_), .o(n_870) );
no02s01 g66927_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_687), .b(parchk_pci_ad_reg_in_1206), .o(g66927_p) );
ao12s01 g66927_u1 ( .a(g66927_p), .b(pci_target_unit_pcit_if_strd_addr_in_687), .c(parchk_pci_ad_reg_in_1206), .o(n_625) );
ao12s01 g66928_u0 ( .a(n_1266), .b(pci_target_unit_fifos_pcir_whole_waddr_94), .c(n_1174), .o(n_1755) );
no02s02 g66929_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_14__Q), .b(wbu_addr_in_263), .o(g66929_p) );
ao12s02 g66929_u1 ( .a(g66929_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_14__Q), .c(wbu_addr_in_263), .o(n_1007) );
no02s01 g66930_u0 ( .a(n_2651), .b(pci_target_unit_pcit_if_strd_bc_in_717), .o(g66930_p) );
ao12m01 g66930_u1 ( .a(g66930_p), .b(pci_target_unit_pcit_if_strd_bc_in_717), .c(n_2651), .o(n_1754) );
no02s02 g66931_u0 ( .a(wbu_addr_in), .b(wishbone_slave_unit_del_sync_addr_out_reg_0__Q), .o(g66931_p) );
ao12s02 g66931_u1 ( .a(g66931_p), .b(wbu_addr_in), .c(wishbone_slave_unit_del_sync_addr_out_reg_0__Q), .o(n_1008) );
no02s02 g66932_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_23__Q), .b(wbu_addr_in_272), .o(g66932_p) );
ao12s02 g66932_u1 ( .a(g66932_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_23__Q), .c(wbu_addr_in_272), .o(n_950) );
no02s02 g66933_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_27__Q), .b(wbu_addr_in_276), .o(g66933_p) );
ao12s02 g66933_u1 ( .a(g66933_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_27__Q), .c(wbu_addr_in_276), .o(n_869) );
no02s01 g66934_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_690), .b(parchk_pci_ad_reg_in_1209), .o(g66934_p) );
ao12s01 g66934_u1 ( .a(g66934_p), .b(pci_target_unit_pcit_if_strd_addr_in_690), .c(parchk_pci_ad_reg_in_1209), .o(n_708) );
no02s01 g66935_u0 ( .a(n_76), .b(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_), .o(g66935_p) );
ao12s01 g66935_u1 ( .a(g66935_p), .b(n_76), .c(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_), .o(n_868) );
no02s01 g66936_u0 ( .a(pci_target_unit_pcit_if_strd_bc_in_719), .b(n_8511), .o(g66936_p) );
ao12s01 g66936_u1 ( .a(g66936_p), .b(pci_target_unit_pcit_if_strd_bc_in_719), .c(n_8511), .o(n_2042) );
no02s01 g66937_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_699), .b(parchk_pci_ad_reg_in_1218), .o(g66937_p) );
ao12s01 g66937_u1 ( .a(g66937_p), .b(pci_target_unit_pcit_if_strd_addr_in_699), .c(parchk_pci_ad_reg_in_1218), .o(n_624) );
in01s01 g66938_u0 ( .a(FE_OFN197_n_2683), .o(n_2043) );
oa12s02 g66939_u0 ( .a(n_1505), .b(parchk_pci_trdy_en_in), .c(n_34), .o(n_2683) );
no02s02 g66940_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_19__Q), .b(wbu_addr_in_268), .o(g66940_p) );
ao12s01 g66940_u1 ( .a(g66940_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_19__Q), .c(wbu_addr_in_268), .o(n_1012) );
no02s01 g66941_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_715), .b(n_2509), .o(g66941_p) );
ao12s01 g66941_u1 ( .a(g66941_p), .b(pci_target_unit_pcit_if_strd_addr_in_715), .c(n_2509), .o(n_1504) );
no02s02 g66942_u0 ( .a(FE_OCP_RBN2289_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q), .o(g66942_p) );
ao12s02 g66942_u1 ( .a(g66942_p), .b(FE_OCP_RBN2289_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q), .o(n_1217) );
ao12m04 g66943_u0 ( .a(n_433), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_1_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .o(n_952) );
no02s02 g66944_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_11__Q), .b(wbu_addr_in_260), .o(g66944_p) );
ao12s02 g66944_u1 ( .a(g66944_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_11__Q), .c(wbu_addr_in_260), .o(n_951) );
no02s03 g66945_u0 ( .a(wishbone_slave_unit_fifos_wbr_be_in), .b(wbu_sel_in), .o(g66945_p) );
ao12s01 g66945_u1 ( .a(g66945_p), .b(wishbone_slave_unit_fifos_wbr_be_in), .c(wbu_sel_in), .o(n_711) );
no02s02 g66946_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_17__Q), .b(wbu_addr_in_266), .o(g66946_p) );
ao12s01 g66946_u1 ( .a(g66946_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_17__Q), .c(wbu_addr_in_266), .o(n_867) );
no02s01 g66947_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_711), .b(parchk_pci_ad_reg_in_1230), .o(g66947_p) );
ao12s01 g66947_u1 ( .a(g66947_p), .b(pci_target_unit_pcit_if_strd_addr_in_711), .c(parchk_pci_ad_reg_in_1230), .o(n_623) );
no02s01 g66948_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_701), .b(parchk_pci_ad_reg_in_1220), .o(g66948_p) );
ao12s01 g66948_u1 ( .a(g66948_p), .b(pci_target_unit_pcit_if_strd_addr_in_701), .c(parchk_pci_ad_reg_in_1220), .o(n_622) );
no02s02 g66949_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_24__Q), .b(wbu_addr_in_273), .o(g66949_p) );
ao12s02 g66949_u1 ( .a(g66949_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_24__Q), .c(wbu_addr_in_273), .o(n_866) );
oa12s01 g66950_u0 ( .a(n_1093), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_1_), .c(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q), .o(n_1094) );
no02s01 g66951_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in), .b(parchk_pci_ad_reg_in), .o(g66951_p) );
ao12s01 g66951_u1 ( .a(g66951_p), .b(pci_target_unit_pcit_if_strd_addr_in), .c(parchk_pci_ad_reg_in), .o(n_621) );
no02s02 g66952_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_10__Q), .b(wbu_addr_in_259), .o(g66952_p) );
ao12s01 g66952_u1 ( .a(g66952_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_10__Q), .c(wbu_addr_in_259), .o(n_865) );
no02s01 g66953_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_698), .b(parchk_pci_ad_reg_in_1217), .o(g66953_p) );
ao12s01 g66953_u1 ( .a(g66953_p), .b(pci_target_unit_pcit_if_strd_addr_in_698), .c(parchk_pci_ad_reg_in_1217), .o(n_658) );
no02s02 g66954_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_29__Q), .b(n_261), .o(g66954_p) );
ao12s02 g66954_u1 ( .a(g66954_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_29__Q), .c(n_261), .o(n_1467) );
no02s02 g66955_u0 ( .a(wbu_addr_in_250), .b(wishbone_slave_unit_del_sync_addr_out_reg_1__Q), .o(g66955_p) );
ao12s02 g66955_u1 ( .a(g66955_p), .b(wbu_addr_in_250), .c(wishbone_slave_unit_del_sync_addr_out_reg_1__Q), .o(n_864) );
ao12f10 g66956_u0 ( .a(n_377), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_2_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_), .o(n_863) );
no02s03 g66957_u0 ( .a(wishbone_slave_unit_fifos_wbr_be_in_265), .b(wbu_sel_in_313), .o(g66957_p) );
ao12s01 g66957_u1 ( .a(g66957_p), .b(wishbone_slave_unit_fifos_wbr_be_in_265), .c(wbu_sel_in_313), .o(n_721) );
no02s01 g66959_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_697), .b(parchk_pci_ad_reg_in_1216), .o(g66959_p) );
ao12s01 g66959_u1 ( .a(g66959_p), .b(pci_target_unit_pcit_if_strd_addr_in_697), .c(parchk_pci_ad_reg_in_1216), .o(n_722) );
no02s02 g66960_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_31__Q), .b(n_539), .o(g66960_p) );
ao12m01 g66960_u1 ( .a(g66960_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_31__Q), .c(n_539), .o(n_1091) );
ao12f10 g66961_u0 ( .a(n_407), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_0_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_), .o(n_1016) );
oa12s01 g66962_u0 ( .a(n_1088), .b(n_961), .c(FE_OCP_RBN1930_parchk_pci_trdy_reg_in), .o(n_1089) );
no02s01 g66963_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_703), .b(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(g66963_p) );
ao12s01 g66963_u1 ( .a(g66963_p), .b(pci_target_unit_pcit_if_strd_addr_in_703), .c(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(n_620) );
no02s01 g66964_u0 ( .a(n_3030), .b(pci_target_unit_pcit_if_strd_bc_in), .o(g66964_p) );
ao12s01 g66964_u1 ( .a(g66964_p), .b(pci_target_unit_pcit_if_strd_bc_in), .c(n_3030), .o(n_2297) );
no02s02 g66965_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_26__Q), .b(wbu_addr_in_275), .o(g66965_p) );
ao12s02 g66965_u1 ( .a(g66965_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_26__Q), .c(wbu_addr_in_275), .o(n_1019) );
no02s01 g66966_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_709), .b(parchk_pci_ad_reg_in_1228), .o(g66966_p) );
ao12s01 g66966_u1 ( .a(g66966_p), .b(pci_target_unit_pcit_if_strd_addr_in_709), .c(parchk_pci_ad_reg_in_1228), .o(n_642) );
no02s01 g66968_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_691), .b(parchk_pci_ad_reg_in_1210), .o(g66968_p) );
ao12s01 g66968_u1 ( .a(g66968_p), .b(pci_target_unit_pcit_if_strd_addr_in_691), .c(parchk_pci_ad_reg_in_1210), .o(n_643) );
ao12f10 g66970_u0 ( .a(n_335), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_3_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_), .o(n_861) );
no02s01 g66975_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_686), .b(parchk_pci_ad_reg_in_1205), .o(g66975_p) );
ao12s01 g66975_u1 ( .a(g66975_p), .b(pci_target_unit_pcit_if_strd_addr_in_686), .c(parchk_pci_ad_reg_in_1205), .o(n_725) );
ao12f08 g66976_u0 ( .a(n_364), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_), .o(n_858) );
no02s01 g66978_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_707), .b(parchk_pci_ad_reg_in_1226), .o(g66978_p) );
ao12s01 g66978_u1 ( .a(g66978_p), .b(pci_target_unit_pcit_if_strd_addr_in_707), .c(parchk_pci_ad_reg_in_1226), .o(n_617) );
oa12s01 g66982_u0 ( .a(n_1028), .b(n_1280), .c(pci_target_unit_wishbone_master_rty_counter_1_), .o(n_1281) );
no02s01 g66984_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_705), .b(parchk_pci_ad_reg_in_1224), .o(g66984_p) );
ao12s01 g66984_u1 ( .a(g66984_p), .b(pci_target_unit_pcit_if_strd_addr_in_705), .c(parchk_pci_ad_reg_in_1224), .o(n_645) );
no02s01 g66985_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_704), .b(parchk_pci_ad_reg_in_1223), .o(g66985_p) );
ao12s01 g66985_u1 ( .a(g66985_p), .b(pci_target_unit_pcit_if_strd_addr_in_704), .c(parchk_pci_ad_reg_in_1223), .o(n_729) );
no02s01 g66986_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_692), .b(parchk_pci_ad_reg_in_1211), .o(g66986_p) );
ao12s01 g66986_u1 ( .a(g66986_p), .b(pci_target_unit_pcit_if_strd_addr_in_692), .c(parchk_pci_ad_reg_in_1211), .o(n_616) );
no02s01 g66987_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_696), .b(parchk_pci_ad_reg_in_1215), .o(g66987_p) );
ao12s01 g66987_u1 ( .a(g66987_p), .b(pci_target_unit_pcit_if_strd_addr_in_696), .c(parchk_pci_ad_reg_in_1215), .o(n_615) );
no02s02 g66988_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_21__Q), .b(wbu_addr_in_270), .o(g66988_p) );
ao12s01 g66988_u1 ( .a(g66988_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_21__Q), .c(wbu_addr_in_270), .o(n_855) );
no02s01 g66989_u0 ( .a(pci_target_unit_fifos_pciw_inTransactionCount_0_), .b(n_852), .o(g66989_p) );
ao12s01 g66989_u1 ( .a(g66989_p), .b(pci_target_unit_fifos_pciw_inTransactionCount_0_), .c(n_852), .o(n_853) );
no02s02 g66990_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_28__Q), .b(wbu_addr_in_277), .o(g66990_p) );
ao12s02 g66990_u1 ( .a(g66990_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_28__Q), .c(wbu_addr_in_277), .o(n_851) );
ao12f06 g66991_u0 ( .a(n_408), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_1_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .o(n_850) );
ao12f06 g66993_u0 ( .a(n_230), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_0_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .o(n_849) );
ao12f08 g66995_u0 ( .a(n_340), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_), .o(n_847) );
no02s01 g66997_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_694), .b(parchk_pci_ad_reg_in_1213), .o(g66997_p) );
ao12s01 g66997_u1 ( .a(g66997_p), .b(pci_target_unit_pcit_if_strd_addr_in_694), .c(parchk_pci_ad_reg_in_1213), .o(n_614) );
ao12s01 g66999_u0 ( .a(n_1454), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .c(n_1316), .o(n_1752) );
ao12f08 g67000_u0 ( .a(n_409), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_), .o(n_1031) );
no02s01 g67001_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_702), .b(FE_OFN1780_parchk_pci_ad_reg_in_1221), .o(g67001_p) );
ao12s01 g67001_u1 ( .a(g67001_p), .b(pci_target_unit_pcit_if_strd_addr_in_702), .c(FE_OFN1780_parchk_pci_ad_reg_in_1221), .o(n_734) );
ao12f10 g67002_u0 ( .a(n_234), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_1_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_), .o(n_845) );
no02s02 g67003_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_5__Q), .b(wbu_addr_in_254), .o(g67003_p) );
ao12s02 g67003_u1 ( .a(g67003_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_5__Q), .c(wbu_addr_in_254), .o(n_844) );
ao12f10 g67004_u0 ( .a(n_268), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_3_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_), .o(n_1033) );
no02s01 g67005_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_716), .b(parchk_pci_ad_reg_in_1235), .o(g67005_p) );
ao12s01 g67005_u1 ( .a(g67005_p), .b(pci_target_unit_pcit_if_strd_addr_in_716), .c(parchk_pci_ad_reg_in_1235), .o(n_737) );
no02s01 g67006_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_700), .b(parchk_pci_ad_reg_in_1219), .o(g67006_p) );
ao12s01 g67006_u1 ( .a(g67006_p), .b(pci_target_unit_pcit_if_strd_addr_in_700), .c(parchk_pci_ad_reg_in_1219), .o(n_613) );
ao12f06 g67007_u0 ( .a(n_386), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_), .o(n_843) );
no02s01 g67008_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_708), .b(parchk_pci_ad_reg_in_1227), .o(g67008_p) );
ao12s01 g67008_u1 ( .a(g67008_p), .b(pci_target_unit_pcit_if_strd_addr_in_708), .c(parchk_pci_ad_reg_in_1227), .o(n_648) );
no02s01 g67010_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_689), .b(parchk_pci_ad_reg_in_1208), .o(g67010_p) );
ao12s01 g67010_u1 ( .a(g67010_p), .b(pci_target_unit_pcit_if_strd_addr_in_689), .c(parchk_pci_ad_reg_in_1208), .o(n_649) );
no02s01 g67011_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_693), .b(parchk_pci_ad_reg_in_1212), .o(g67011_p) );
ao12s01 g67011_u1 ( .a(g67011_p), .b(pci_target_unit_pcit_if_strd_addr_in_693), .c(parchk_pci_ad_reg_in_1212), .o(n_612) );
ao12f10 g67012_u0 ( .a(n_320), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_1_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_), .o(n_842) );
no02s02 g67014_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_25__Q), .b(wbu_addr_in_274), .o(g67014_p) );
ao12s02 g67014_u1 ( .a(g67014_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_25__Q), .c(wbu_addr_in_274), .o(n_960) );
no02s01 g67015_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_30__Q), .b(wbu_addr_in_279), .o(g67015_p) );
ao12s02 g67015_u1 ( .a(g67015_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_30__Q), .c(wbu_addr_in_279), .o(n_1034) );
ao12f06 g67016_u0 ( .a(n_420), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_), .o(n_841) );
no02s01 g67017_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_), .o(g67017_p) );
ao12m01 g67017_u1 ( .a(g67017_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q), .o(n_840) );
no02s01 g67018_u0 ( .a(n_358), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q), .o(g67018_p) );
ao12s01 g67018_u1 ( .a(g67018_p), .b(n_358), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q), .o(n_1086) );
no02s02 g67019_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_9__Q), .b(wbu_addr_in_258), .o(g67019_p) );
ao12s01 g67019_u1 ( .a(g67019_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_9__Q), .c(wbu_addr_in_258), .o(n_1035) );
no02s02 g67020_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_15__Q), .b(wbu_addr_in_264), .o(g67020_p) );
ao12s01 g67020_u1 ( .a(g67020_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_15__Q), .c(wbu_addr_in_264), .o(n_839) );
no02s01 g67021_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_4__Q), .b(wbu_addr_in_253), .o(g67021_p) );
ao12s01 g67021_u1 ( .a(g67021_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_4__Q), .c(wbu_addr_in_253), .o(n_838) );
no02s02 g67022_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_13__Q), .b(wbu_addr_in_262), .o(g67022_p) );
ao12s02 g67022_u1 ( .a(g67022_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_13__Q), .c(wbu_addr_in_262), .o(n_837) );
no02s02 g67023_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_20__Q), .b(wbu_addr_in_269), .o(g67023_p) );
ao12s02 g67023_u1 ( .a(g67023_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_20__Q), .c(wbu_addr_in_269), .o(n_959) );
no02s03 g67024_u0 ( .a(wishbone_slave_unit_fifos_wbr_be_in_266), .b(wbu_sel_in_314), .o(g67024_p) );
ao12s01 g67024_u1 ( .a(g67024_p), .b(wishbone_slave_unit_fifos_wbr_be_in_266), .c(wbu_sel_in_314), .o(n_611) );
no02s02 g67025_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_2__Q), .b(wbu_addr_in_251), .o(g67025_p) );
ao12s01 g67025_u1 ( .a(g67025_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_2__Q), .c(wbu_addr_in_251), .o(n_836) );
no02s02 g67026_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_18__Q), .b(wbu_addr_in_267), .o(g67026_p) );
ao12s02 g67026_u1 ( .a(g67026_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_18__Q), .c(wbu_addr_in_267), .o(n_742) );
no02s01 g67029_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_688), .b(parchk_pci_ad_reg_in_1207), .o(g67029_p) );
ao12s01 g67029_u1 ( .a(g67029_p), .b(pci_target_unit_pcit_if_strd_addr_in_688), .c(parchk_pci_ad_reg_in_1207), .o(n_610) );
no02s02 g67030_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_8__Q), .b(wbu_addr_in_257), .o(g67030_p) );
ao12s02 g67030_u1 ( .a(g67030_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_8__Q), .c(wbu_addr_in_257), .o(n_744) );
no02s02 g67031_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_12__Q), .b(wbu_addr_in_261), .o(g67031_p) );
ao12s02 g67031_u1 ( .a(g67031_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_12__Q), .c(wbu_addr_in_261), .o(n_743) );
no02s02 g67032_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_7__Q), .b(wbu_addr_in_256), .o(g67032_p) );
ao12s01 g67032_u1 ( .a(g67032_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_7__Q), .c(wbu_addr_in_256), .o(n_833) );
no02s01 g67033_u0 ( .a(wishbone_slave_unit_fifos_wbr_be_in_264), .b(wbu_sel_in_312), .o(g67033_p) );
ao12s02 g67033_u1 ( .a(g67033_p), .b(wishbone_slave_unit_fifos_wbr_be_in_264), .c(wbu_sel_in_312), .o(n_609) );
ao22s01 g67034_u0 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_1_), .b(wishbone_slave_unit_fifos_wbw_inTransactionCount_0_), .c(n_362), .d(n_397), .o(n_1085) );
oa12s01 g67035_u0 ( .a(n_1038), .b(wishbone_slave_unit_fifos_wbw_inTransactionCount_1_), .c(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q), .o(n_1039) );
no02s01 g67036_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_3__Q), .b(wbu_addr_in_252), .o(g67036_p) );
ao12s01 g67036_u1 ( .a(g67036_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_3__Q), .c(wbu_addr_in_252), .o(n_747) );
na02f02 TIMEBOOST_cell_42264 ( .a(TIMEBOOST_net_13370), .b(FE_OFN1404_n_8567), .o(TIMEBOOST_net_12271) );
na02s03 TIMEBOOST_cell_45767 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__Q), .b(n_13161), .o(TIMEBOOST_net_15122) );
in01s01 g67040_u0 ( .a(FE_OFN989_n_574), .o(g67040_sb) );
na02s02 TIMEBOOST_cell_42652 ( .a(TIMEBOOST_net_13564), .b(g64126_da), .o(TIMEBOOST_net_11295) );
na02s01 g67040_u2 ( .a(pci_ad_i_2_), .b(n_574), .o(g67040_db) );
na04m02 TIMEBOOST_cell_34768 ( .a(TIMEBOOST_net_4822), .b(g59800_sb), .c(g52455_sb), .d(g52455_db), .o(n_14834) );
na02s01 TIMEBOOST_cell_15880 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_77), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_3197) );
na02s01 g67041_u2 ( .a(pci_ad_i_20_), .b(n_574), .o(g67041_db) );
na02f02 TIMEBOOST_cell_39094 ( .a(TIMEBOOST_net_11785), .b(FE_OFN1586_n_13736), .o(n_16207) );
in01s01 g67042_u0 ( .a(conf_pci_init_complete_out), .o(g67042_sb) );
na02s01 g67042_u2 ( .a(pci_ad_i_6_), .b(conf_pci_init_complete_out), .o(g67042_db) );
na02s01 TIMEBOOST_cell_42580 ( .a(TIMEBOOST_net_13528), .b(g64139_db), .o(n_4024) );
na02s01 TIMEBOOST_cell_39181 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__Q), .b(g64315_sb), .o(TIMEBOOST_net_11829) );
na02s01 g67043_u2 ( .a(pci_ad_i_8_), .b(conf_pci_init_complete_out), .o(g67043_db) );
na02s01 TIMEBOOST_cell_17659 ( .a(TIMEBOOST_net_4086), .b(g65306_db), .o(n_4274) );
in01s01 g67044_u0 ( .a(parchk_pci_cbe_en_in), .o(g67044_sb) );
na02s01 g67044_u1 ( .a(pci_cbe_i_0_), .b(g67044_sb), .o(g67044_da) );
na02s02 g67044_u2 ( .a(parchk_pci_cbe_out_in), .b(parchk_pci_cbe_en_in), .o(g67044_db) );
na02s03 g67044_u3 ( .a(g67044_da), .b(g67044_db), .o(n_2376) );
na02s02 g67045_u1 ( .a(pci_cbe_i_1_), .b(g57790_sb), .o(g67045_da) );
na02s02 g67045_u2 ( .a(parchk_pci_cbe_out_in_1202), .b(parchk_pci_cbe_en_in), .o(g67045_db) );
na02s03 g67045_u3 ( .a(g67045_da), .b(g67045_db), .o(n_1847) );
in01s01 g67046_u0 ( .a(parchk_pci_cbe_en_in), .o(g67046_sb) );
na02s03 g67046_u1 ( .a(pci_cbe_i_3_), .b(g67046_sb), .o(g67046_da) );
na02s03 g67046_u2 ( .a(parchk_pci_cbe_out_in_1204), .b(parchk_pci_cbe_en_in), .o(g67046_db) );
na02s06 g67046_u3 ( .a(g67046_da), .b(g67046_db), .o(n_2566) );
in01f04 g67047_u0 ( .a(n_1211), .o(n_832) );
in01m10 g67048_u0 ( .a(conf_wb_err_bc_in), .o(g67048_sb) );
na02s01 TIMEBOOST_cell_40351 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__Q), .b(n_8176), .o(TIMEBOOST_net_12414) );
na02f10 g67048_u2 ( .a(conf_wb_err_bc_in), .b(conf_wb_err_bc_in_846), .o(g67048_db) );
na02s01 TIMEBOOST_cell_40364 ( .a(TIMEBOOST_net_12420), .b(g61735_db), .o(n_8349) );
in01s01 g67049_u0 ( .a(conf_pci_init_complete_out), .o(g67049_sb) );
na02f02 TIMEBOOST_cell_42496 ( .a(TIMEBOOST_net_13486), .b(g57175_sb), .o(n_11580) );
na02s01 g67049_u2 ( .a(pci_ad_i_19_), .b(conf_pci_init_complete_out), .o(g67049_db) );
na02s02 TIMEBOOST_cell_17747 ( .a(TIMEBOOST_net_4130), .b(g61754_sb), .o(n_8307) );
na02s02 TIMEBOOST_cell_42134 ( .a(TIMEBOOST_net_13305), .b(g62914_sb), .o(n_6051) );
na02s01 g67050_u2 ( .a(pci_ad_i_31_), .b(conf_pci_init_complete_out), .o(g67050_db) );
na02s01 TIMEBOOST_cell_40366 ( .a(TIMEBOOST_net_12421), .b(g61736_db), .o(n_8346) );
in01s02 g67051_u0 ( .a(FE_OFN989_n_574), .o(g67051_sb) );
na03s02 TIMEBOOST_cell_39355 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__Q), .b(FE_OFN713_n_8140), .c(n_1898), .o(TIMEBOOST_net_11916) );
na02s01 g67051_u2 ( .a(pci_ad_i_24_), .b(n_574), .o(g67051_db) );
no02s02 TIMEBOOST_cell_44770 ( .a(TIMEBOOST_net_14623), .b(n_2430), .o(TIMEBOOST_net_1154) );
no02m02 TIMEBOOST_cell_45564 ( .a(TIMEBOOST_net_15020), .b(FE_RN_578_0), .o(TIMEBOOST_net_2025) );
na02s01 g67052_u2 ( .a(pci_idsel_i), .b(FE_OFN989_n_574), .o(g67052_db) );
na02s01 TIMEBOOST_cell_42605 ( .a(n_3739), .b(g65030_sb), .o(TIMEBOOST_net_13541) );
na03s02 TIMEBOOST_cell_33591 ( .a(TIMEBOOST_net_9552), .b(n_5633), .c(g62106_sb), .o(n_5594) );
na02s01 g67053_u2 ( .a(pci_ad_i_14_), .b(n_574), .o(g67053_db) );
na02s03 TIMEBOOST_cell_45768 ( .a(TIMEBOOST_net_15122), .b(FE_OFN1326_n_13547), .o(TIMEBOOST_net_14957) );
na02s01 TIMEBOOST_cell_45585 ( .a(n_4452), .b(g65036_sb), .o(TIMEBOOST_net_15031) );
na02s01 TIMEBOOST_cell_16643 ( .a(TIMEBOOST_net_3578), .b(g64161_db), .o(n_4004) );
na02s01 g67055_u2 ( .a(pci_ad_i_28_), .b(n_574), .o(g67055_db) );
na03s02 TIMEBOOST_cell_33590 ( .a(TIMEBOOST_net_9553), .b(n_5633), .c(g62133_sb), .o(n_5561) );
na02s01 g67056_u2 ( .a(pci_ad_i_30_), .b(n_2373), .o(g67056_db) );
in01s01 g67057_u0 ( .a(n_2373), .o(g67057_sb) );
na02f02 TIMEBOOST_cell_42348 ( .a(TIMEBOOST_net_13412), .b(g57445_sb), .o(TIMEBOOST_net_12330) );
na03f10 TIMEBOOST_cell_82 ( .a(n_15414), .b(n_16854), .c(n_15417), .o(n_16015) );
na02s02 TIMEBOOST_cell_40432 ( .a(TIMEBOOST_net_12454), .b(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_6228) );
na02s02 TIMEBOOST_cell_38710 ( .a(TIMEBOOST_net_11593), .b(g62446_sb), .o(n_6703) );
na02s01 TIMEBOOST_cell_31286 ( .a(configuration_wb_err_addr_555), .b(conf_wb_err_addr_in_964), .o(TIMEBOOST_net_9554) );
na02s02 TIMEBOOST_cell_40368 ( .a(TIMEBOOST_net_12422), .b(g65709_db), .o(n_1946) );
na02s01 g67059_u2 ( .a(pci_ad_i_9_), .b(n_574), .o(g67059_db) );
na03s02 TIMEBOOST_cell_33589 ( .a(TIMEBOOST_net_9554), .b(n_5633), .c(g62124_sb), .o(n_5572) );
in01m04 g67064_u0 ( .a(n_1551), .o(n_12179) );
na02m02 TIMEBOOST_cell_41667 ( .a(pci_target_unit_fifos_outGreyCount_reg_1__Q), .b(n_996), .o(TIMEBOOST_net_13072) );
na02s01 TIMEBOOST_cell_42581 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__Q), .b(g65935_sb), .o(TIMEBOOST_net_13529) );
na03f02 TIMEBOOST_cell_36192 ( .a(n_12072), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__Q), .c(n_11823), .o(n_12494) );
na02s01 TIMEBOOST_cell_39486 ( .a(TIMEBOOST_net_11981), .b(TIMEBOOST_net_9825), .o(n_7197) );
na04f04 TIMEBOOST_cell_36225 ( .a(n_13046), .b(n_12873), .c(n_12872), .d(n_12781), .o(n_13130) );
na02s02 TIMEBOOST_cell_42136 ( .a(TIMEBOOST_net_13306), .b(g62916_sb), .o(n_6047) );
na02m02 TIMEBOOST_cell_42231 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__Q), .b(n_9578), .o(TIMEBOOST_net_13354) );
in01s01 g67070_u0 ( .a(parchk_pci_cbe_en_in), .o(g67070_sb) );
na02s03 g67070_u1 ( .a(pci_cbe_i_2_), .b(g67070_sb), .o(g67070_da) );
na02s03 g67070_u2 ( .a(parchk_pci_cbe_out_in_1203), .b(parchk_pci_cbe_en_in), .o(g67070_db) );
na02s06 g67070_u3 ( .a(g67070_da), .b(g67070_db), .o(n_2171) );
na02f02 TIMEBOOST_cell_41594 ( .a(FE_OFN1441_n_9372), .b(TIMEBOOST_net_13035), .o(TIMEBOOST_net_11652) );
na02s01 g67071_u2 ( .a(pci_ad_i_16_), .b(FE_OFN989_n_574), .o(g67071_db) );
na02s02 TIMEBOOST_cell_45700 ( .a(TIMEBOOST_net_15088), .b(FE_OFN1248_n_4093), .o(TIMEBOOST_net_13241) );
na03f02 TIMEBOOST_cell_34788 ( .a(n_3290), .b(pciu_bar0_in), .c(n_2905), .o(TIMEBOOST_net_2805) );
na02s01 TIMEBOOST_cell_45565 ( .a(g64207_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__16__Q), .o(TIMEBOOST_net_15021) );
na02s02 TIMEBOOST_cell_43049 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__8__Q), .b(n_4440), .o(TIMEBOOST_net_13763) );
na02s01 TIMEBOOST_cell_41921 ( .a(FE_OFN201_n_9230), .b(g58412_sb), .o(TIMEBOOST_net_13199) );
na02s01 g67073_u2 ( .a(pci_ad_i_3_), .b(n_574), .o(g67073_db) );
na02s02 TIMEBOOST_cell_41932 ( .a(TIMEBOOST_net_13204), .b(g54183_sb), .o(n_13430) );
na02s01 TIMEBOOST_cell_42137 ( .a(TIMEBOOST_net_4276), .b(g64165_db), .o(TIMEBOOST_net_13307) );
na02s01 g67074_u2 ( .a(pci_ad_i_18_), .b(conf_pci_init_complete_out), .o(g67074_db) );
na02s01 TIMEBOOST_cell_42138 ( .a(TIMEBOOST_net_13307), .b(TIMEBOOST_net_10024), .o(n_5513) );
na02s01 TIMEBOOST_cell_41776 ( .a(TIMEBOOST_net_13126), .b(g58194_db), .o(n_9056) );
na02s01 g67075_u2 ( .a(pci_ad_i_11_), .b(conf_pci_init_complete_out), .o(g67075_db) );
na03s03 TIMEBOOST_cell_26 ( .a(output_backup_par_out_reg_Q), .b(g54038_sb), .c(g54038_db), .o(n_13335) );
in01f03 g67080_u0 ( .a(n_1192), .o(n_1436) );
in01m08 g67082_u0 ( .a(parchk_pci_trdy_en_in), .o(g67082_sb) );
na02s02 TIMEBOOST_cell_45566 ( .a(TIMEBOOST_net_15021), .b(g64207_da), .o(TIMEBOOST_net_11274) );
na02s01 TIMEBOOST_cell_16936 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__Q), .b(g65279_sb), .o(TIMEBOOST_net_3725) );
na02s01 TIMEBOOST_cell_16937 ( .a(TIMEBOOST_net_3725), .b(g65279_db), .o(n_3585) );
na02f02 g53412_u0 ( .a(FE_OCP_RBN1962_FE_OFN1591_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__15__Q), .o(n_14060) );
na02s01 g67083_u2 ( .a(pci_ad_i_1_), .b(conf_pci_init_complete_out), .o(g67083_db) );
na03s02 TIMEBOOST_cell_38507 ( .a(TIMEBOOST_net_4090), .b(g65285_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__Q), .o(TIMEBOOST_net_11492) );
na02s02 TIMEBOOST_cell_41931 ( .a(TIMEBOOST_net_9854), .b(FE_OFN1084_n_13221), .o(TIMEBOOST_net_13204) );
na02s01 g67084_u2 ( .a(pci_ad_i_25_), .b(n_574), .o(g67084_db) );
na02s01 TIMEBOOST_cell_45567 ( .a(g60677_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__Q), .o(TIMEBOOST_net_15022) );
na02s01 TIMEBOOST_cell_31284 ( .a(configuration_wb_err_addr_563), .b(wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q), .o(TIMEBOOST_net_9553) );
na02s01 g67085_u2 ( .a(pci_ad_i_21_), .b(conf_pci_init_complete_out), .o(g67085_db) );
na02f02 TIMEBOOST_cell_42232 ( .a(TIMEBOOST_net_13354), .b(FE_OFN1421_n_8567), .o(TIMEBOOST_net_12311) );
na02s01 TIMEBOOST_cell_42606 ( .a(TIMEBOOST_net_13541), .b(g65030_db), .o(n_3627) );
na02s01 TIMEBOOST_cell_39212 ( .a(TIMEBOOST_net_11844), .b(g65010_db), .o(TIMEBOOST_net_4814) );
na02s01 TIMEBOOST_cell_42714 ( .a(TIMEBOOST_net_13595), .b(g64958_db), .o(n_3660) );
na02m02 TIMEBOOST_cell_42233 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__Q), .b(n_9569), .o(TIMEBOOST_net_13355) );
na03s02 TIMEBOOST_cell_35191 ( .a(n_1862), .b(g61907_sb), .c(g61907_db), .o(n_8007) );
na02m02 TIMEBOOST_cell_42139 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__Q), .b(n_9647), .o(TIMEBOOST_net_13308) );
na02s01 TIMEBOOST_cell_30908 ( .a(pci_target_unit_pcit_if_strd_addr_in_712), .b(pci_target_unit_del_sync_addr_in_230), .o(TIMEBOOST_net_9365) );
na02s01 g67088_u2 ( .a(pci_ad_i_23_), .b(n_574), .o(g67088_db) );
na02f02 TIMEBOOST_cell_40978 ( .a(TIMEBOOST_net_12727), .b(g57150_sb), .o(n_11600) );
in01s01 g67089_u0 ( .a(n_1536), .o(n_1450) );
ao22m04 g67090_u0 ( .a(pci_stop_i), .b(n_454), .c(n_205), .d(parchk_pci_trdy_en_in), .o(n_1536) );
na02s02 TIMEBOOST_cell_45568 ( .a(TIMEBOOST_net_15022), .b(g60677_da), .o(TIMEBOOST_net_10633) );
na02s01 g67091_u2 ( .a(pci_ad_i_10_), .b(n_574), .o(g67091_db) );
na02s01 TIMEBOOST_cell_45569 ( .a(FE_OFN229_n_9120), .b(g58184_sb), .o(TIMEBOOST_net_15023) );
na03s02 TIMEBOOST_cell_34465 ( .a(pci_target_unit_wishbone_master_bc_register_reg_0__Q), .b(g52590_sb), .c(TIMEBOOST_net_879), .o(n_14687) );
na02m02 TIMEBOOST_cell_44333 ( .a(n_9038), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__Q), .o(TIMEBOOST_net_14405) );
na02s01 TIMEBOOST_cell_40370 ( .a(TIMEBOOST_net_12423), .b(FE_OFN2079_n_8069), .o(TIMEBOOST_net_11101) );
na02s02 TIMEBOOST_cell_45570 ( .a(TIMEBOOST_net_15023), .b(g58184_db), .o(n_9059) );
na02s01 g67093_u2 ( .a(pci_ad_i_26_), .b(n_574), .o(g67093_db) );
na02s02 TIMEBOOST_cell_45701 ( .a(n_95), .b(n_4487), .o(TIMEBOOST_net_15089) );
na02s01 TIMEBOOST_cell_42938 ( .a(TIMEBOOST_net_13707), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_11197) );
na02s01 g67094_u2 ( .a(pci_ad_i_29_), .b(n_2373), .o(g67094_db) );
na02s01 TIMEBOOST_cell_31282 ( .a(configuration_wb_err_data_575), .b(parchk_pci_ad_out_in_1172), .o(TIMEBOOST_net_9552) );
no02s02 g67095_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(g67095_p) );
ao12s02 g67095_u1 ( .a(g67095_p), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .c(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(n_4939) );
no02m10 g67096_u0 ( .a(parchk_pci_ad_out_in_1180), .b(parchk_pci_ad_out_in_1179), .o(g67096_p) );
ao12f08 g67096_u1 ( .a(g67096_p), .b(parchk_pci_ad_out_in_1180), .c(parchk_pci_ad_out_in_1179), .o(n_652) );
no02m10 g67097_u0 ( .a(parchk_pci_ad_reg_in_1231), .b(parchk_pci_ad_reg_in_1230), .o(g67097_p) );
ao12f06 g67097_u1 ( .a(g67097_p), .b(parchk_pci_ad_reg_in_1231), .c(parchk_pci_ad_reg_in_1230), .o(n_607) );
no02s01 g67098_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_1_), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_), .o(g67098_p) );
ao12s01 g67098_u1 ( .a(g67098_p), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_1_), .c(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_), .o(n_1083) );
no02s01 g67099_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_1_), .b(n_321), .o(g67099_p) );
ao12s01 g67099_u1 ( .a(g67099_p), .b(pci_target_unit_del_sync_comp_cycle_count_1_), .c(n_321), .o(n_963) );
no02m10 g67100_u0 ( .a(parchk_pci_ad_out_in_1190), .b(parchk_pci_ad_out_in_1189), .o(g67100_p) );
ao12f08 g67100_u1 ( .a(g67100_p), .b(parchk_pci_ad_out_in_1190), .c(parchk_pci_ad_out_in_1189), .o(n_606) );
no02m10 g67102_u0 ( .a(parchk_pci_ad_out_in_1198), .b(parchk_pci_ad_out_in_1197), .o(g67102_p) );
ao12f08 g67102_u1 ( .a(g67102_p), .b(parchk_pci_ad_out_in_1198), .c(parchk_pci_ad_out_in_1197), .o(n_605) );
no02s10 g67103_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_1_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_), .o(g67103_p) );
ao12m04 g67103_u1 ( .a(g67103_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_1_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_), .o(n_604) );
no02m10 g67104_u0 ( .a(parchk_pci_ad_out_in_1194), .b(parchk_pci_ad_out_in_1193), .o(g67104_p) );
ao12f08 g67104_u1 ( .a(g67104_p), .b(parchk_pci_ad_out_in_1194), .c(parchk_pci_ad_out_in_1193), .o(n_603) );
no02m08 g67105_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_2_), .o(g67105_p) );
ao12f06 g67105_u1 ( .a(g67105_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_2_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .o(n_602) );
no02s01 g67106_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_), .o(g67106_p) );
ao12s01 g67106_u1 ( .a(g67106_p), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_), .o(n_655) );
no02s04 g67107_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q), .o(g67107_p) );
ao12s02 g67107_u1 ( .a(g67107_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q), .c(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q), .o(n_829) );
no02s01 g67108_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .o(g67108_p) );
ao12s01 g67108_u1 ( .a(g67108_p), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .c(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .o(n_1199) );
no02s06 g67109_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q), .o(g67109_p) );
ao12s01 g67109_u1 ( .a(g67109_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__Q), .c(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q), .o(n_971) );
no02f10 g67110_u0 ( .a(parchk_pci_ad_reg_in_1233), .b(parchk_pci_ad_reg_in_1232), .o(g67110_p) );
ao12f10 g67110_u1 ( .a(g67110_p), .b(parchk_pci_ad_reg_in_1233), .c(parchk_pci_ad_reg_in_1232), .o(n_656) );
no02s01 g67111_u0 ( .a(n_46), .b(n_16071), .o(g67111_p) );
ao12s01 g67111_u1 ( .a(g67111_p), .b(n_46), .c(n_16071), .o(n_969) );
no02s01 g67112_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q), .b(n_160), .o(g67112_p) );
ao12s01 g67112_u1 ( .a(g67112_p), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q), .c(n_160), .o(n_973) );
no02s10 g67113_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_2_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_), .o(g67113_p) );
ao12m04 g67113_u1 ( .a(g67113_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_2_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_), .o(n_601) );
no02s10 g67114_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_0_), .o(g67114_p) );
ao12s10 g67114_u1 ( .a(g67114_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_0_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_), .o(n_659) );
no02f20 g67115_u0 ( .a(parchk_pci_ad_reg_in_1213), .b(parchk_pci_ad_reg_in_1212), .o(g67115_p) );
ao12f10 g67115_u1 ( .a(g67115_p), .b(parchk_pci_ad_reg_in_1213), .c(parchk_pci_ad_reg_in_1212), .o(n_678) );
no02m10 g67116_u0 ( .a(parchk_pci_ad_reg_in_1219), .b(parchk_pci_ad_reg_in_1218), .o(g67116_p) );
ao12f08 g67116_u1 ( .a(g67116_p), .b(parchk_pci_ad_reg_in_1219), .c(parchk_pci_ad_reg_in_1218), .o(n_600) );
no02s01 g67117_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_), .o(g67117_p) );
ao12s01 g67117_u1 ( .a(g67117_p), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_0_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_), .o(n_599) );
no02m10 g67118_u0 ( .a(parchk_pci_ad_reg_in_1227), .b(parchk_pci_ad_reg_in_1226), .o(g67118_p) );
ao12f06 g67118_u1 ( .a(g67118_p), .b(parchk_pci_ad_reg_in_1227), .c(parchk_pci_ad_reg_in_1226), .o(n_674) );
no02s01 g67119_u0 ( .a(conf_wb_err_addr_in_943), .b(conf_wb_err_addr_in_944), .o(g67119_p) );
ao12s01 g67119_u1 ( .a(g67119_p), .b(conf_wb_err_addr_in_943), .c(conf_wb_err_addr_in_944), .o(n_662) );
no02m10 g67120_u0 ( .a(parchk_pci_ad_reg_in_1225), .b(parchk_pci_ad_reg_in_1224), .o(g67120_p) );
ao12f06 g67120_u1 ( .a(g67120_p), .b(parchk_pci_ad_reg_in_1225), .c(parchk_pci_ad_reg_in_1224), .o(n_598) );
no02f20 g67122_u0 ( .a(parchk_pci_ad_reg_in_1211), .b(parchk_pci_ad_reg_in_1210), .o(g67122_p) );
ao12f10 g67122_u1 ( .a(g67122_p), .b(parchk_pci_ad_reg_in_1211), .c(parchk_pci_ad_reg_in_1210), .o(n_597) );
no02f20 g67123_u0 ( .a(parchk_pci_ad_reg_in_1209), .b(parchk_pci_ad_reg_in_1208), .o(g67123_p) );
ao12f10 g67123_u1 ( .a(g67123_p), .b(parchk_pci_ad_reg_in_1209), .c(parchk_pci_ad_reg_in_1208), .o(n_663) );
no02f10 g67125_u0 ( .a(n_15854), .b(n_1061), .o(g67125_p) );
ao12f08 g67125_u1 ( .a(g67125_p), .b(n_15854), .c(n_1061), .o(n_1081) );
no02f20 g67126_u0 ( .a(parchk_pci_ad_reg_in_1215), .b(parchk_pci_ad_reg_in_1214), .o(g67126_p) );
ao12f10 g67126_u1 ( .a(g67126_p), .b(parchk_pci_ad_reg_in_1215), .c(parchk_pci_ad_reg_in_1214), .o(n_664) );
no02m10 g67127_u0 ( .a(parchk_pci_ad_out_in_1192), .b(parchk_pci_ad_out_in_1191), .o(g67127_p) );
ao12f08 g67127_u1 ( .a(g67127_p), .b(parchk_pci_ad_out_in_1192), .c(parchk_pci_ad_out_in_1191), .o(n_666) );
no02s10 g67128_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_), .o(g67128_p) );
ao12m06 g67128_u1 ( .a(g67128_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_), .o(n_596) );
no02s01 g67129_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(g67129_p) );
ao12s01 g67129_u1 ( .a(g67129_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(n_1079) );
no02m10 g67130_u0 ( .a(parchk_pci_ad_out_in_1172), .b(parchk_pci_ad_out_in_1171), .o(g67130_p) );
ao12f08 g67130_u1 ( .a(g67130_p), .b(parchk_pci_ad_out_in_1172), .c(parchk_pci_ad_out_in_1171), .o(n_595) );
no02s01 g67131_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_), .o(g67131_p) );
ao12s01 g67131_u1 ( .a(g67131_p), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_), .o(n_669) );
no02m10 g67132_u0 ( .a(parchk_pci_ad_out_in_1196), .b(parchk_pci_ad_out_in_1195), .o(g67132_p) );
ao12f08 g67132_u1 ( .a(g67132_p), .b(parchk_pci_ad_out_in_1196), .c(parchk_pci_ad_out_in_1195), .o(n_667) );
no02f08 g67133_u0 ( .a(FE_OFN1781_parchk_pci_ad_reg_in_1221), .b(parchk_pci_ad_reg_in_1220), .o(g67133_p) );
ao12f06 g67133_u1 ( .a(g67133_p), .b(FE_OFN1781_parchk_pci_ad_reg_in_1221), .c(parchk_pci_ad_reg_in_1220), .o(n_594) );
no02f10 g67134_u0 ( .a(n_2509), .b(parchk_pci_ad_reg_in_1235), .o(g67134_p) );
ao12f10 g67134_u1 ( .a(g67134_p), .b(n_2509), .c(parchk_pci_ad_reg_in_1235), .o(n_593) );
no02m08 g67135_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_2_), .o(g67135_p) );
ao12m06 g67135_u1 ( .a(g67135_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_2_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .o(n_668) );
no02m10 g67136_u0 ( .a(parchk_pci_ad_out_in_1176), .b(parchk_pci_ad_out_in_1175), .o(g67136_p) );
ao12f08 g67136_u1 ( .a(g67136_p), .b(parchk_pci_ad_out_in_1176), .c(parchk_pci_ad_out_in_1175), .o(n_592) );
no02m10 g67138_u0 ( .a(parchk_pci_ad_reg_in_1205), .b(parchk_pci_ad_reg_in), .o(g67138_p) );
ao12f08 g67138_u1 ( .a(g67138_p), .b(parchk_pci_ad_reg_in_1205), .c(parchk_pci_ad_reg_in), .o(n_588) );
no02m10 g67139_u0 ( .a(parchk_pci_ad_out_in_1182), .b(parchk_pci_ad_out_in_1181), .o(g67139_p) );
ao12f08 g67139_u1 ( .a(g67139_p), .b(parchk_pci_ad_out_in_1182), .c(parchk_pci_ad_out_in_1181), .o(n_670) );
no02m08 g67140_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_0_), .o(g67140_p) );
ao12m04 g67140_u1 ( .a(g67140_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_0_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .o(n_587) );
no02s01 g67141_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q), .b(n_150), .o(g67141_p) );
ao12s01 g67141_u1 ( .a(g67141_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q), .c(n_150), .o(n_826) );
no02s01 g67142_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .o(g67142_p) );
ao12s01 g67142_u1 ( .a(g67142_p), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .c(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .o(n_1465) );
no02m10 g67143_u0 ( .a(parchk_pci_ad_out_in_1170), .b(parchk_pci_ad_out_in_1169), .o(g67143_p) );
ao12f08 g67143_u1 ( .a(g67143_p), .b(parchk_pci_ad_out_in_1170), .c(parchk_pci_ad_out_in_1169), .o(n_586) );
na02s01 TIMEBOOST_cell_40365 ( .a(n_1922), .b(g61736_sb), .o(TIMEBOOST_net_12421) );
no02m10 g67145_u0 ( .a(parchk_pci_ad_out_in_1178), .b(parchk_pci_ad_out_in_1177), .o(g67145_p) );
ao12f08 g67145_u1 ( .a(g67145_p), .b(parchk_pci_ad_out_in_1178), .c(parchk_pci_ad_out_in_1177), .o(n_672) );
no02m10 g67146_u0 ( .a(parchk_pci_ad_reg_in_1217), .b(parchk_pci_ad_reg_in_1216), .o(g67146_p) );
ao12f08 g67146_u1 ( .a(g67146_p), .b(parchk_pci_ad_reg_in_1217), .c(parchk_pci_ad_reg_in_1216), .o(n_673) );
na02s01 TIMEBOOST_cell_42582 ( .a(TIMEBOOST_net_13529), .b(g65935_db), .o(n_2169) );
no02m10 g67148_u0 ( .a(parchk_pci_ad_out_in_1188), .b(parchk_pci_ad_out_in_1187), .o(g67148_p) );
ao12f08 g67148_u1 ( .a(g67148_p), .b(parchk_pci_ad_out_in_1188), .c(parchk_pci_ad_out_in_1187), .o(n_583) );
no02m10 g67149_u0 ( .a(parchk_pci_ad_reg_in_1207), .b(parchk_pci_ad_reg_in_1206), .o(g67149_p) );
ao12f08 g67149_u1 ( .a(g67149_p), .b(parchk_pci_ad_reg_in_1207), .c(parchk_pci_ad_reg_in_1206), .o(n_582) );
no02s01 g67150_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__Q), .b(n_150), .o(g67150_p) );
ao12s01 g67150_u1 ( .a(g67150_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__Q), .c(n_150), .o(n_982) );
no02m10 g67151_u0 ( .a(parchk_pci_ad_out_in_1186), .b(parchk_pci_ad_out_in_1185), .o(g67151_p) );
ao12f08 g67151_u1 ( .a(g67151_p), .b(parchk_pci_ad_out_in_1186), .c(parchk_pci_ad_out_in_1185), .o(n_581) );
no02m10 g67152_u0 ( .a(parchk_pci_ad_out_in_1184), .b(parchk_pci_ad_out_in_1183), .o(g67152_p) );
ao12f08 g67152_u1 ( .a(g67152_p), .b(parchk_pci_ad_out_in_1184), .c(parchk_pci_ad_out_in_1183), .o(n_650) );
no02s01 g67153_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_1_), .b(n_282), .o(g67153_p) );
ao12s01 g67153_u1 ( .a(g67153_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_1_), .c(n_282), .o(n_983) );
no02m10 g67154_u0 ( .a(parchk_pci_ad_reg_in_1229), .b(parchk_pci_ad_reg_in_1228), .o(g67154_p) );
ao12f06 g67154_u1 ( .a(g67154_p), .b(parchk_pci_ad_reg_in_1229), .c(parchk_pci_ad_reg_in_1228), .o(n_675) );
no02s01 g67155_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_1_), .o(g67155_p) );
ao12s01 g67155_u1 ( .a(g67155_p), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_), .c(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_1_), .o(n_580) );
no02s01 g67156_u0 ( .a(parchk_pci_cbe_out_in_1203), .b(parchk_pci_cbe_out_in_1202), .o(g67156_p) );
ao12s01 g67156_u1 ( .a(g67156_p), .b(parchk_pci_cbe_out_in_1203), .c(parchk_pci_cbe_out_in_1202), .o(n_676) );
no02f08 g67157_u0 ( .a(parchk_pci_ad_reg_in_1223), .b(FE_OFN1777_parchk_pci_ad_reg_in_1222), .o(g67157_p) );
ao12f06 g67157_u1 ( .a(g67157_p), .b(parchk_pci_ad_reg_in_1223), .c(FE_OFN1777_parchk_pci_ad_reg_in_1222), .o(n_677) );
in01s03 g67176_u0 ( .a(n_2031), .o(n_2520) );
in01s03 g67185_u0 ( .a(n_2597), .o(n_2031) );
in01m20 g67231_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_mabort2), .o(n_1459) );
in01s01 g67246_u0 ( .a(wishbone_slave_unit_del_sync_sync_comp_req_pending), .o(n_1460) );
in01s01 g67261_u0 ( .a(pci_target_unit_wishbone_master_burst_chopped_delayed), .o(n_824) );
in01s06 g67306_u0 ( .a(n_1009), .o(n_1509) );
na02s10 g67307_u0 ( .a(n_143), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .o(n_1009) );
no02s06 g67308_u0 ( .a(n_689), .b(pci_target_unit_fifos_pcir_whole_waddr_94), .o(n_1118) );
in01s01 g67310_u0 ( .a(n_7426), .o(n_2040) );
na02s01 g67311_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1216), .o(g67311_p) );
in01s01 g67311_u1 ( .a(g67311_p), .o(n_7426) );
in01s01 g67312_u0 ( .a(n_7279), .o(n_2041) );
na02s01 g67313_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1215), .o(g67313_p) );
in01s01 g67313_u1 ( .a(g67313_p), .o(n_7279) );
no02m03 g67314_u0 ( .a(n_242), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(n_1195) );
in01s01 g67317_u0 ( .a(n_2464), .o(n_7802) );
na02m01 g67318_u0 ( .a(FE_OCPN1854_n_2071), .b(parchk_pci_ad_reg_in_1205), .o(n_2464) );
no02m08 g67319_u0 ( .a(pciu_pciif_stop_reg_in), .b(n_707), .o(n_2685) );
in01s01 g67320_u0 ( .a(n_1014), .o(n_1826) );
na02f10 g67322_u0 ( .a(wishbone_slave_unit_del_sync_req_comp_pending), .b(n_709), .o(n_1014) );
in01s01 g67323_u0 ( .a(n_7269), .o(n_2084) );
na02s01 g67324_u0 ( .a(n_2044), .b(FE_OFN1780_parchk_pci_ad_reg_in_1221), .o(g67324_p) );
in01s02 g67324_u1 ( .a(g67324_p), .o(n_7269) );
na02s01 g67325_u0 ( .a(FE_OCPN1855_n_2071), .b(parchk_pci_ad_reg_in_1211), .o(n_3265) );
in01s01 g67326_u0 ( .a(n_7244), .o(n_2083) );
na02s01 g67327_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1229), .o(g67327_p) );
in01s01 g67327_u1 ( .a(g67327_p), .o(n_7244) );
in01s01 g67328_u0 ( .a(n_7285), .o(n_2286) );
na02s01 g67329_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1230), .o(g67329_p) );
in01s01 g67329_u1 ( .a(g67329_p), .o(n_7285) );
in01s01 g67331_u0 ( .a(n_2046), .o(n_2287) );
na02s02 g67332_u0 ( .a(n_565), .b(n_15302), .o(n_2046) );
in01s01 g67333_u0 ( .a(n_1290), .o(n_1218) );
no02m06 g67335_u0 ( .a(n_349), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .o(n_1290) );
no02s10 g67336_u0 ( .a(n_143), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .o(n_1201) );
na02s01 g67337_u0 ( .a(pciu_pciif_bckp_stop_in), .b(output_backup_trdy_out_reg_Q), .o(n_1512) );
in01s01 g67339_u0 ( .a(n_7287), .o(n_2082) );
na02s01 g67340_u0 ( .a(n_2044), .b(parchk_pci_ad_reg_in_1226), .o(g67340_p) );
in01s02 g67340_u1 ( .a(g67340_p), .o(n_7287) );
na02f10 g67341_u0 ( .a(n_1104), .b(n_16906), .o(n_819) );
na02f10 g67342_u0 ( .a(n_15924), .b(n_15998), .o(n_1408) );
in01s01 g67350_u0 ( .a(n_8540), .o(n_6996) );
na02s02 g67351_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1235), .o(n_8540) );
in01s01 g67352_u0 ( .a(n_7424), .o(n_1746) );
na02s01 g67353_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1217), .o(g67353_p) );
in01s01 g67353_u1 ( .a(g67353_p), .o(n_7424) );
in01s01 g67354_u0 ( .a(n_7806), .o(n_8517) );
na02s01 g67355_u0 ( .a(FE_OCPN1854_n_2071), .b(parchk_pci_ad_reg_in), .o(g67355_p) );
in01s01 g67355_u1 ( .a(g67355_p), .o(n_7806) );
no02s01 g67356_u0 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_0_), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q), .o(n_713) );
in01s01 g67358_u0 ( .a(n_2080), .o(n_7239) );
na02s01 g67359_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1231), .o(n_2080) );
na02s02 g67360_u0 ( .a(n_715), .b(conf_wb_err_bc_in_848), .o(g67360_p) );
in01s02 g67360_u1 ( .a(g67360_p), .o(n_716) );
in01s01 g67362_u0 ( .a(n_2079), .o(n_7234) );
na02s01 g67363_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1232), .o(n_2079) );
na02m01 g67364_u0 ( .a(n_763), .b(n_2078), .o(g67364_p) );
in01m02 g67364_u1 ( .a(g67364_p), .o(n_2609) );
in01s01 g67365_u0 ( .a(n_816), .o(n_817) );
no02s01 g67366_u0 ( .a(n_148), .b(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_), .o(n_816) );
na02s01 g67367_u0 ( .a(FE_OCPN1855_n_2071), .b(parchk_pci_ad_reg_in_1207), .o(n_3277) );
na02m04 g67369_u0 ( .a(n_653), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(g67369_p) );
in01m02 g67369_u1 ( .a(g67369_p), .o(n_1615) );
in01s01 g67370_u0 ( .a(n_1265), .o(n_1266) );
no02s01 g67371_u0 ( .a(pci_target_unit_fifos_pcir_whole_waddr_94), .b(n_1174), .o(g67371_p) );
in01s01 g67371_u1 ( .a(g67371_p), .o(n_1265) );
na02s01 g67372_u0 ( .a(n_148), .b(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_), .o(n_1283) );
in01s01 g67375_u0 ( .a(n_3280), .o(n_7289) );
na02s01 g67376_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1212), .o(n_3280) );
in01f02 g67377_u0 ( .a(n_1219), .o(n_1220) );
no02f10 g67378_u0 ( .a(n_815), .b(pci_target_unit_pcit_if_strd_bc_in), .o(n_1219) );
na02s01 g67379_u0 ( .a(n_1263), .b(n_705), .o(n_1264) );
in01m03 g67380_u0 ( .a(n_1017), .o(n_980) );
no02s08 g67382_u0 ( .a(n_573), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .o(n_1017) );
na02s01 g67383_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_7_), .b(n_705), .o(n_1261) );
in01s01 g67385_u0 ( .a(n_7265), .o(n_2077) );
na02s01 g67386_u0 ( .a(n_2044), .b(parchk_pci_ad_reg_in_1224), .o(g67386_p) );
in01s02 g67386_u1 ( .a(g67386_p), .o(n_7265) );
na02s01 g67387_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_6_), .b(n_705), .o(n_1260) );
in01s01 g67388_u0 ( .a(n_7254), .o(n_2076) );
na02s01 g67389_u0 ( .a(n_2044), .b(parchk_pci_ad_reg_in_1227), .o(g67389_p) );
in01s02 g67389_u1 ( .a(g67389_p), .o(n_7254) );
na02s08 g67390_u0 ( .a(n_242), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(g67390_p) );
in01s08 g67390_u1 ( .a(g67390_p), .o(n_1113) );
in01s01 g67391_u0 ( .a(n_7267), .o(n_2075) );
na02s01 g67392_u0 ( .a(n_2044), .b(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(g67392_p) );
in01s02 g67392_u1 ( .a(g67392_p), .o(n_7267) );
in01s01 g67393_u0 ( .a(n_7272), .o(n_2074) );
na02s01 g67394_u0 ( .a(n_2044), .b(parchk_pci_ad_reg_in_1220), .o(g67394_p) );
in01s02 g67394_u1 ( .a(g67394_p), .o(n_7272) );
na02s08 g67396_u0 ( .a(n_349), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .o(g67396_p) );
in01s06 g67396_u1 ( .a(g67396_p), .o(n_1188) );
na02s01 g67397_u0 ( .a(FE_OCPN1854_n_2071), .b(parchk_pci_ad_reg_in_1210), .o(g67397_p) );
in01s01 g67397_u1 ( .a(g67397_p), .o(n_7792) );
no02s10 g67398_u0 ( .a(n_2), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .o(n_1288) );
in01s01 g67400_u0 ( .a(n_2072), .o(n_7295) );
na02s01 g67401_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1233), .o(n_2072) );
in01s01 g67402_u0 ( .a(n_7282), .o(n_1743) );
na02s01 g67403_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1214), .o(g67403_p) );
in01s01 g67403_u1 ( .a(g67403_p), .o(n_7282) );
in01f02 g67404_u0 ( .a(n_1197), .o(n_1198) );
no02f06 g67405_u0 ( .a(n_1023), .b(n_551), .o(g67405_p) );
in01f04 g67405_u1 ( .a(g67405_p), .o(n_1197) );
no02s01 g67406_u0 ( .a(n_85), .b(pci_target_unit_pcit_if_strd_bc_in_718), .o(n_661) );
na02s01 g67407_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_5_), .b(n_705), .o(n_1077) );
in01s01 g67409_u0 ( .a(n_2319), .o(n_7800) );
na02m01 g67410_u0 ( .a(FE_OCPN1854_n_2071), .b(parchk_pci_ad_reg_in_1206), .o(n_2319) );
na02f01 g67411_u0 ( .a(n_16685), .b(n_15998), .o(g67411_p) );
in01s02 g67411_u1 ( .a(g67411_p), .o(n_1742) );
na02s01 g67412_u0 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_1_), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q), .o(n_1093) );
na02s01 g67413_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_3_), .b(n_705), .o(n_1259) );
in01s01 g67415_u0 ( .a(n_2070), .o(n_7291) );
na02s01 g67416_u0 ( .a(n_1061), .b(n_2509), .o(n_2070) );
in01m06 g67419_u0 ( .a(n_2337), .o(n_8498) );
na02f10 g67421_u0 ( .a(pci_target_unit_del_sync_req_comp_pending), .b(n_373), .o(g67421_p) );
in01m03 g67421_u1 ( .a(g67421_p), .o(n_2337) );
no02s01 g67422_u0 ( .a(n_181), .b(pci_target_unit_pcit_if_strd_bc_in_718), .o(n_671) );
in01s02 g67423_u0 ( .a(n_812), .o(n_813) );
na02s06 g67425_u0 ( .a(n_573), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .o(g67425_p) );
in01s04 g67425_u1 ( .a(g67425_p), .o(n_812) );
in01m02 g67426_u0 ( .a(n_16326), .o(n_1074) );
in01s01 g67429_u0 ( .a(n_7440), .o(n_1740) );
na02s01 g67430_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1219), .o(g67430_p) );
in01s01 g67430_u1 ( .a(g67430_p), .o(n_7440) );
in01s01 g67431_u0 ( .a(n_7259), .o(n_2069) );
na02s01 g67432_u0 ( .a(n_2044), .b(parchk_pci_ad_reg_in_1225), .o(g67432_p) );
in01s02 g67432_u1 ( .a(g67432_p), .o(n_7259) );
in01s01 g67433_u0 ( .a(n_1027), .o(n_1028) );
na02f20 g67434_u0 ( .a(n_1280), .b(pci_target_unit_wishbone_master_rty_counter_1_), .o(g67434_p) );
in01f08 g67434_u1 ( .a(g67434_p), .o(n_1027) );
in01f02 g67435_u0 ( .a(n_16033), .o(n_1072) );
na02s08 g67437_u0 ( .a(n_2), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .o(g67437_p) );
in01s06 g67437_u1 ( .a(g67437_p), .o(n_1289) );
na02s01 g67438_u0 ( .a(FE_OCPN1855_n_2071), .b(parchk_pci_ad_reg_in_1209), .o(n_3275) );
in01s01 g67442_u0 ( .a(n_2068), .o(n_7249) );
na02s01 g67443_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1228), .o(n_2068) );
na02s01 g67444_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_4_), .b(n_705), .o(n_1475) );
in01s01 g67445_u0 ( .a(n_7241), .o(n_2067) );
na02s01 g67446_u0 ( .a(n_2044), .b(parchk_pci_ad_reg_in_1223), .o(g67446_p) );
in01s02 g67446_u1 ( .a(g67446_p), .o(n_7241) );
no02m02 g67447_u0 ( .a(n_2742), .b(n_2316), .o(n_2778) );
in01f04 g67448_u0 ( .a(n_15757), .o(n_1221) );
no02s01 g67452_u0 ( .a(n_5755), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(n_1069) );
na02s06 g67453_u0 ( .a(n_689), .b(pci_target_unit_fifos_pcir_whole_waddr_94), .o(g67453_p) );
in01s04 g67453_u1 ( .a(g67453_p), .o(n_1103) );
no02s01 g67454_u0 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_0_), .b(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q), .o(n_567) );
no02s01 g67456_u0 ( .a(configuration_set_isr_bit2), .b(configuration_sync_isr_2_del_bit_reg_Q), .o(n_1084) );
no02s01 g67457_u0 ( .a(n_16685), .b(n_15998), .o(g67457_p) );
in01s01 g67457_u1 ( .a(g67457_p), .o(n_1739) );
in01s01 g67458_u0 ( .a(n_1453), .o(n_1454) );
no02s01 g67459_u0 ( .a(pci_target_unit_fifos_pciw_whole_waddr_47), .b(n_1316), .o(g67459_p) );
in01s01 g67459_u1 ( .a(g67459_p), .o(n_1453) );
in01f02 g67460_u0 ( .a(n_992), .o(n_993) );
na02f08 g67461_u0 ( .a(n_681), .b(n_16904), .o(n_992) );
in01s01 g67462_u0 ( .a(n_7231), .o(n_1737) );
na02s01 g67463_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1213), .o(g67463_p) );
in01s01 g67463_u1 ( .a(g67463_p), .o(n_7231) );
no02s01 g67464_u0 ( .a(configuration_set_pci_err_cs_bit8), .b(configuration_sync_pci_err_cs_8_del_bit_reg_Q), .o(n_736) );
no02s01 g67466_u0 ( .a(n_2314), .b(n_1724), .o(n_2315) );
in01s01 g67467_u0 ( .a(n_7422), .o(n_2052) );
na02s01 g67468_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1218), .o(g67468_p) );
in01s01 g67468_u1 ( .a(g67468_p), .o(n_7422) );
na02s03 g67469_u0 ( .a(wishbone_slave_unit_pcim_sm_be_in_558), .b(n_57), .o(n_564) );
in01s06 g67479_u0 ( .a(n_1258), .o(n_2115) );
in01m04 g67480_u0 ( .a(FE_OFN1619_n_1787), .o(n_1258) );
no02m10 g67481_u0 ( .a(n_504), .b(n_541), .o(n_1787) );
na02s01 g67483_u0 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_1_), .b(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q), .o(n_1038) );
no02s01 g67484_u0 ( .a(n_763), .b(n_2078), .o(n_3108) );
na02s01 g67485_u0 ( .a(FE_OCPN1855_n_2071), .b(parchk_pci_ad_reg_in_1208), .o(n_3273) );
na02s01 g67486_u0 ( .a(n_123), .b(pci_rst_i), .o(wb_rst_o) );
na02s06 g67487_u0 ( .a(wbu_addr_in_265), .b(wbu_addr_in_262), .o(n_191) );
in01s01 g67488_u0 ( .a(n_560), .o(n_561) );
no02s06 g67489_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_4_), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_5_), .o(g67489_p) );
in01s04 g67489_u1 ( .a(g67489_p), .o(n_560) );
no02f20 g67490_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_3_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_), .o(n_335) );
na02m03 g67491_u0 ( .a(wbu_addr_in_274), .b(wbu_addr_in_275), .o(n_888) );
in01s04 g67492_u0 ( .a(n_1005), .o(n_1106) );
no02m03 g67493_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(g67493_p) );
in01s06 g67493_u1 ( .a(g67493_p), .o(n_1005) );
na02m10 g67494_u0 ( .a(pciu_am1_in_535), .b(parchk_pci_ad_reg_in_1230), .o(n_336) );
na02m20 g67495_u0 ( .a(pciu_bar1_in_387), .b(pciu_am1_in_525), .o(g67495_p) );
in01f08 g67495_u1 ( .a(g67495_p), .o(n_3404) );
na02s03 g67496_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(n_808) );
na02m06 g67497_u0 ( .a(wbm_adr_o_16_), .b(wbm_adr_o_15_), .o(n_923) );
no02s03 g67498_u0 ( .a(wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q), .b(wishbone_slave_unit_del_sync_comp_rty_exp_reg), .o(g67498_p) );
in01s01 g67498_u1 ( .a(g67498_p), .o(n_559) );
na02s10 g67499_u0 ( .a(conf_wb_err_addr_in_961), .b(conf_wb_err_addr_in_962), .o(n_895) );
na02m03 g67500_u0 ( .a(pci_target_unit_fifos_pcir_whole_waddr_94), .b(pci_target_unit_fifos_pcir_whole_waddr), .o(n_914) );
na02s10 g67501_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_0_), .b(pci_target_unit_wishbone_master_rty_counter_1_), .o(n_1334) );
na02s20 g67502_u0 ( .a(conf_wb_err_addr_in_947), .b(conf_wb_err_addr_in_946), .o(g67502_p) );
in01m08 g67502_u1 ( .a(g67502_p), .o(n_994) );
na02m02 g67503_u0 ( .a(n_539), .b(wbu_am1_in), .o(n_558) );
na02m10 g67504_u0 ( .a(pciu_am1_in_530), .b(parchk_pci_ad_reg_in_1225), .o(n_204) );
na02m20 g67505_u0 ( .a(pciu_bar1_in_394), .b(pciu_am1_in_532), .o(g67505_p) );
in01f08 g67505_u1 ( .a(g67505_p), .o(n_3078) );
na02s01 g67506_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_11_), .b(pci_target_unit_del_sync_comp_cycle_count_12_), .o(g67506_p) );
in01s01 g67506_u1 ( .a(g67506_p), .o(n_1989) );
na02s01 g67507_u0 ( .a(pci_target_unit_pci_target_sm_rd_progress), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(g67507_p) );
in01s01 g67507_u1 ( .a(g67507_p), .o(n_7530) );
na02m10 g67510_u0 ( .a(pciu_am1_in_525), .b(parchk_pci_ad_reg_in_1220), .o(n_290) );
no02m10 g67511_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_), .o(n_340) );
na02m03 g67512_u0 ( .a(wbm_adr_o_22_), .b(wbm_adr_o_21_), .o(n_915) );
no02s06 g67514_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_0_), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_1_), .o(g67514_p) );
in01s04 g67514_u1 ( .a(g67514_p), .o(n_1011) );
no02f20 g67515_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_2_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_), .o(n_341) );
in01s02 g67518_u0 ( .a(n_562), .o(n_563) );
na02s10 g67519_u0 ( .a(wbm_adr_o_6_), .b(wbm_adr_o_5_), .o(g67519_p) );
in01m04 g67519_u1 ( .a(g67519_p), .o(n_562) );
no02f02 g67520_u0 ( .a(n_16690), .b(n_15998), .o(n_1812) );
na02m03 g67521_u0 ( .a(wbu_addr_in_260), .b(wbu_addr_in_259), .o(n_945) );
na02s08 g67522_u0 ( .a(wbu_addr_in_253), .b(wbu_addr_in_254), .o(n_430) );
na02m03 g67523_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .o(g67523_p) );
in01s06 g67523_u1 ( .a(g67523_p), .o(n_1115) );
na02f04 g67526_u0 ( .a(pciu_am1_in_526), .b(FE_OFN1780_parchk_pci_ad_reg_in_1221), .o(n_287) );
na02s01 g67527_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_), .o(n_554) );
no02s10 g67528_u0 ( .a(parchk_pci_ad_reg_in), .b(parchk_pci_ad_reg_in_1205), .o(n_343) );
na02s08 g67530_u0 ( .a(wbu_addr_in_252), .b(wbu_addr_in_253), .o(n_350) );
na02s03 g67531_u0 ( .a(wbm_adr_o_27_), .b(wbm_adr_o_28_), .o(g67531_p) );
in01s01 g67531_u1 ( .a(g67531_p), .o(n_879) );
na02m04 g67532_u0 ( .a(n_1628), .b(pci_target_unit_pci_target_sm_n_2), .o(n_1383) );
na02m03 g67533_u0 ( .a(wbu_addr_in_255), .b(wbu_addr_in_254), .o(n_874) );
na02m20 g67534_u0 ( .a(pciu_bar1_in_384), .b(pciu_am1_in_522), .o(g67534_p) );
in01f08 g67534_u1 ( .a(g67534_p), .o(n_2812) );
na02s03 g67535_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_5_), .b(pci_target_unit_del_sync_comp_cycle_count_6_), .o(g67535_p) );
in01s03 g67535_u1 ( .a(g67535_p), .o(n_1690) );
na02m20 g67536_u0 ( .a(pciu_bar1_in_382), .b(pciu_am1_in_520), .o(g67536_p) );
in01f08 g67536_u1 ( .a(g67536_p), .o(n_2818) );
na02s10 g67537_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .o(g67537_p) );
in01s08 g67537_u1 ( .a(g67537_p), .o(n_1173) );
no02s01 g67538_u0 ( .a(configuration_cache_line_size_reg), .b(configuration_cache_line_size_reg_2996), .o(g67538_p) );
in01s01 g67538_u1 ( .a(g67538_p), .o(n_434) );
na02f10 g67539_u0 ( .a(n_16695), .b(n_551), .o(n_1291) );
na02s10 g67540_u0 ( .a(conf_wb_err_addr_in_963), .b(conf_wb_err_addr_in_962), .o(n_745) );
na02m10 g67542_u0 ( .a(pciu_am1_in_529), .b(parchk_pci_ad_reg_in_1224), .o(n_419) );
no02f02 g67543_u0 ( .a(n_1519), .b(n_15998), .o(n_2016) );
na02m20 g67544_u0 ( .a(pciu_bar1_in_388), .b(pciu_am1_in_526), .o(g67544_p) );
in01f08 g67544_u1 ( .a(g67544_p), .o(n_2869) );
na02m03 g67545_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(g67545_p) );
in01s06 g67545_u1 ( .a(g67545_p), .o(n_1210) );
in01s01 g67546_u0 ( .a(n_549), .o(n_550) );
na02m03 g67547_u0 ( .a(wbm_adr_o_24_), .b(wbm_adr_o_25_), .o(n_549) );
no02s02 g67548_u0 ( .a(wishbone_slave_unit_pcim_if_del_burst_in), .b(wishbone_slave_unit_fifos_wbr_be_in_264), .o(n_235) );
na02s06 g67549_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_1_), .b(pci_target_unit_del_sync_comp_cycle_count_0_), .o(g67549_p) );
in01s03 g67549_u1 ( .a(g67549_p), .o(n_948) );
na02m03 g67550_u0 ( .a(wbm_adr_o_23_), .b(wbm_adr_o_24_), .o(n_924) );
na02m10 g67551_u0 ( .a(parchk_pci_ad_reg_in_1227), .b(pciu_am1_in_532), .o(n_357) );
na02m10 g67553_u0 ( .a(pciu_am1_in_528), .b(parchk_pci_ad_reg_in_1223), .o(n_360) );
na02s10 g67554_u0 ( .a(wbu_addr_in_265), .b(wbu_addr_in_266), .o(n_956) );
na02m03 g67556_u0 ( .a(wbu_addr_in_271), .b(wbu_addr_in_272), .o(n_892) );
no02s01 g67557_u0 ( .a(n_2629), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(n_2313) );
na02m03 g67558_u0 ( .a(wbm_adr_o_15_), .b(wbm_adr_o_14_), .o(n_900) );
na02m20 g67559_u0 ( .a(pciu_bar1_in_402), .b(pciu_am1_in_540), .o(g67559_p) );
in01f08 g67559_u1 ( .a(g67559_p), .o(n_3592) );
no02s01 g67560_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_11_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_12_), .o(n_1993) );
no02m03 g67562_u0 ( .a(pci_target_unit_fifos_pcir_whole_waddr_94), .b(pci_target_unit_fifos_pcir_whole_waddr), .o(n_1318) );
na02s01 g67563_u0 ( .a(wishbone_slave_unit_pci_initiator_if_read_bound), .b(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(n_4869) );
na02m03 g67564_u0 ( .a(wbu_addr_in_267), .b(wbu_addr_in_268), .o(n_927) );
na02m03 g67565_u0 ( .a(wbm_adr_o_10_), .b(wbm_adr_o_11_), .o(n_926) );
in01s01 g67568_u0 ( .a(n_546), .o(n_547) );
no02s01 g67569_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_decode_count_0_), .b(wishbone_slave_unit_pci_initiator_sm_decode_count_1_), .o(n_546) );
in01m04 g67570_u0 ( .a(n_544), .o(n_545) );
na02m20 g67571_u0 ( .a(conf_wb_err_bc_in_847), .b(conf_wb_err_bc_in_848), .o(n_544) );
in01s01 g67573_u0 ( .a(n_703), .o(n_660) );
no02s01 g67574_u0 ( .a(wishbone_slave_unit_pci_initiator_if_read_count_0_), .b(wishbone_slave_unit_pci_initiator_if_read_count_1_), .o(n_703) );
in01m01 g67576_u0 ( .a(n_15859), .o(n_2354) );
na02s01 g67579_u0 ( .a(configuration_wb_err_cs_bit0), .b(configuration_icr_bit_2961), .o(n_369) );
no02s01 g67580_u0 ( .a(wbu_cache_line_size_in_206), .b(wbu_cache_line_size_in_207), .o(n_802) );
na02s03 g67581_u0 ( .a(wbm_adr_o_26_), .b(wbm_adr_o_27_), .o(g67581_p) );
in01s01 g67581_u1 ( .a(g67581_p), .o(n_875) );
na02s08 g67582_u0 ( .a(conf_wb_err_addr_in_948), .b(conf_wb_err_addr_in_945), .o(g67582_p) );
in01m02 g67582_u1 ( .a(g67582_p), .o(n_331) );
na02f08 g67583_u0 ( .a(n_324), .b(n_541), .o(g67583_p) );
in01f06 g67583_u1 ( .a(g67583_p), .o(n_2122) );
no02s01 g67584_u0 ( .a(pci_target_unit_wishbone_master_read_count_0_), .b(pci_target_unit_wishbone_master_read_count_reg_2__Q), .o(n_3164) );
no02f40 g67585_u0 ( .a(wishbone_slave_unit_wishbone_slave_img_hit_4_), .b(wishbone_slave_unit_wishbone_slave_img_hit_3_), .o(n_370) );
no02f80 g67586_u0 ( .a(wbm_rty_i), .b(wbm_err_i), .o(n_898) );
no02m02 g67588_u0 ( .a(n_629), .b(n_2078), .o(n_3503) );
in01f04 g67589_u0 ( .a(n_730), .o(n_731) );
na02f10 g67590_u0 ( .a(pci_target_unit_pcit_if_strd_bc_in_718), .b(pci_target_unit_pcit_if_strd_bc_in_719), .o(n_730) );
na02m03 g67591_u0 ( .a(wbm_adr_o_9_), .b(wbm_adr_o_8_), .o(n_920) );
na02m08 g67592_u0 ( .a(conf_wb_err_addr_in_944), .b(conf_wb_err_addr_in_945), .o(g67592_p) );
in01m04 g67592_u1 ( .a(g67592_p), .o(n_375) );
na02s10 g67593_u0 ( .a(conf_wb_err_addr_in_955), .b(conf_wb_err_addr_in_956), .o(n_886) );
na02m02 g67594_u0 ( .a(wbu_am2_in), .b(n_539), .o(n_540) );
in01s06 g67595_u0 ( .a(n_538), .o(n_1194) );
no02m03 g67596_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .o(g67596_p) );
in01s06 g67596_u1 ( .a(g67596_p), .o(n_538) );
na02s03 g67598_u0 ( .a(wbu_addr_in_266), .b(wbu_addr_in_267), .o(n_304) );
no02f20 g67599_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_1_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_), .o(n_234) );
na02m10 g67600_u0 ( .a(pciu_am1_in_540), .b(parchk_pci_ad_reg_in_1235), .o(g67600_p) );
in01f04 g67600_u1 ( .a(g67600_p), .o(n_372) );
na02s06 g67601_u0 ( .a(wbu_addr_in_267), .b(wbu_addr_in_264), .o(n_374) );
na02m03 g67602_u0 ( .a(wbu_addr_in_269), .b(wbu_addr_in_270), .o(n_909) );
na02s08 g67603_u0 ( .a(conf_wb_err_addr_in_968), .b(conf_wb_err_addr_in_969), .o(g67603_p) );
in01s04 g67603_u1 ( .a(g67603_p), .o(n_1441) );
na02s01 g67604_u0 ( .a(wbs_bte_i_0_), .b(wbs_bte_i_1_), .o(n_382) );
na02m20 g67605_u0 ( .a(pciu_bar1_in_396), .b(pciu_am1_in_534), .o(g67605_p) );
in01f08 g67605_u1 ( .a(g67605_p), .o(n_2833) );
no02f20 g67606_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_3_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_), .o(n_268) );
no02s01 g67607_u0 ( .a(wbm_ack_i), .b(wbm_err_i), .o(TIMEBOOST_net_10356) );
na02s10 g67608_u0 ( .a(conf_wb_err_addr_in_957), .b(conf_wb_err_addr_in_958), .o(n_891) );
na02m20 g67610_u0 ( .a(pciu_bar1_in_399), .b(pciu_am1_in_537), .o(g67610_p) );
in01f08 g67610_u1 ( .a(g67610_p), .o(n_2825) );
na02m10 g67611_u0 ( .a(pciu_am1_in), .b(parchk_pci_ad_reg_in_1212), .o(n_376) );
na02m20 g67613_u0 ( .a(pciu_bar1_in_381), .b(pciu_am1_in_519), .o(g67613_p) );
in01f08 g67613_u1 ( .a(g67613_p), .o(n_2822) );
na02s20 g67614_u0 ( .a(wbu_addr_in_264), .b(wbu_addr_in_263), .o(n_957) );
in01s01 g67616_u0 ( .a(n_535), .o(n_536) );
na02s01 g67617_u0 ( .a(wb_int_i), .b(configuration_icr_bit2_0), .o(n_535) );
na02s10 g67618_u0 ( .a(conf_wb_err_addr_in_964), .b(conf_wb_err_addr_in_965), .o(n_746) );
na02f40 g67619_u0 ( .a(wishbone_slave_unit_wishbone_slave_c_state_1), .b(wishbone_slave_unit_wishbone_slave_c_state), .o(n_943) );
na02m03 g67620_u0 ( .a(wbm_adr_o_13_), .b(wbm_adr_o_12_), .o(n_901) );
no02f20 g67621_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_2_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_), .o(n_377) );
na02s08 g67624_u0 ( .a(pci_target_unit_fifos_pciw_whole_waddr), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .o(g67624_p) );
in01m04 g67624_u1 ( .a(g67624_p), .o(n_1317) );
na02m10 g67625_u0 ( .a(pciu_am1_in_539), .b(n_2509), .o(g67625_p) );
in01f06 g67625_u1 ( .a(g67625_p), .o(n_233) );
na02m20 g67626_u0 ( .a(pciu_bar1_in_398), .b(pciu_am1_in_536), .o(g67626_p) );
in01f08 g67626_u1 ( .a(g67626_p), .o(n_2841) );
na02m10 g67627_u0 ( .a(pciu_am1_in_519), .b(parchk_pci_ad_reg_in_1214), .o(n_439) );
no02s01 g67628_u0 ( .a(n_2308), .b(n_2316), .o(n_2995) );
na02m03 g67629_u0 ( .a(wbm_adr_o_6_), .b(wbm_adr_o_7_), .o(n_919) );
na02m03 g67630_u0 ( .a(conf_wb_err_addr_in_950), .b(conf_wb_err_addr_in_949), .o(n_232) );
na02s10 g67631_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .o(g67631_p) );
in01m06 g67631_u1 ( .a(g67631_p), .o(n_1107) );
no02s02 g67632_u0 ( .a(wishbone_slave_unit_pcim_if_del_burst_in), .b(wishbone_slave_unit_fifos_wbr_be_in_266), .o(n_398) );
no02s01 g67633_u0 ( .a(wbs_cti_i_0_), .b(wbs_cti_i_2_), .o(n_272) );
na02m03 g67634_u0 ( .a(wbm_adr_o_18_), .b(wbm_adr_o_19_), .o(n_911) );
na02s10 g67635_u0 ( .a(wbu_addr_in_256), .b(wbu_addr_in_257), .o(n_893) );
in01m02 g67638_u0 ( .a(n_533), .o(n_534) );
na02s10 g67639_u0 ( .a(conf_wb_err_addr_in_961), .b(conf_wb_err_addr_in_960), .o(n_533) );
in01m06 g67640_u0 ( .a(n_16052), .o(n_1774) );
na02m10 g67642_u0 ( .a(pciu_am1_in_536), .b(parchk_pci_ad_reg_in_1231), .o(n_385) );
na02f20 g67644_u0 ( .a(n_16906), .b(n_391), .o(n_1200) );
no02s01 g67645_u0 ( .a(wbu_cache_line_size_in_211), .b(wbu_cache_line_size_in_210), .o(n_257) );
no02f08 g67646_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_), .o(n_386) );
na02s06 g67647_u0 ( .a(wbu_addr_in_277), .b(wbu_addr_in_276), .o(n_939) );
in01m03 g67651_u0 ( .a(n_1468), .o(n_13354) );
in01m10 g67654_u0 ( .a(n_1468), .o(n_7552) );
in01m06 g67657_u0 ( .a(n_1468), .o(n_7822) );
in01m10 g67662_u0 ( .a(n_1468), .o(n_12595) );
in01m20 g67663_u0 ( .a(n_532), .o(n_1468) );
no02f40 g67666_u0 ( .a(pci_target_unit_pci_target_sm_cnf_progress), .b(n_2314), .o(n_532) );
na02m03 g67667_u0 ( .a(wbm_adr_o_17_), .b(wbm_adr_o_16_), .o(n_921) );
na02m08 g67668_u0 ( .a(pciu_am1_in_520), .b(parchk_pci_ad_reg_in_1215), .o(n_231) );
no02s01 g67669_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_decode_count_1_), .b(wishbone_slave_unit_pci_initiator_sm_decode_count_2_), .o(n_1471) );
na02m10 g67670_u0 ( .a(pciu_am1_in_522), .b(parchk_pci_ad_reg_in_1217), .o(n_389) );
na02m10 g67671_u0 ( .a(pciu_am1_in_538), .b(parchk_pci_ad_reg_in_1233), .o(g67671_p) );
in01f06 g67671_u1 ( .a(g67671_p), .o(n_277) );
na02m10 g67672_u0 ( .a(conf_wb_err_addr_in_957), .b(conf_wb_err_addr_in_956), .o(g67672_p) );
in01m06 g67672_u1 ( .a(g67672_p), .o(n_913) );
no02f06 g67673_u0 ( .a(wishbone_slave_unit_wishbone_slave_c_state_1), .b(wishbone_slave_unit_wishbone_slave_c_state), .o(n_1432) );
na02m20 g67675_u0 ( .a(pciu_bar1_in_389), .b(pciu_am1_in_527), .o(g67675_p) );
in01f08 g67675_u1 ( .a(g67675_p), .o(n_2866) );
no02m03 g67676_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_2_), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_3_), .o(n_1416) );
na02s06 g67677_u0 ( .a(wbu_addr_in_273), .b(wbu_addr_in_272), .o(n_889) );
no02s01 g67678_u0 ( .a(n_1724), .b(n_2311), .o(n_2763) );
na02s10 g67680_u0 ( .a(wbu_bar2_in), .b(wbu_am2_in), .o(g67680_p) );
in01m04 g67680_u1 ( .a(g67680_p), .o(n_1332) );
na02m03 g67682_u0 ( .a(wbu_addr_in_262), .b(wbu_addr_in_261), .o(n_887) );
no02m08 g67684_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .o(n_230) );
in01s04 g67685_u0 ( .a(n_530), .o(n_531) );
na02m03 g67686_u0 ( .a(conf_wb_err_addr_in_967), .b(conf_wb_err_addr_in_968), .o(n_530) );
na02s08 g67688_u0 ( .a(wbu_bar1_in), .b(wbu_am1_in), .o(g67688_p) );
in01s04 g67688_u1 ( .a(g67688_p), .o(n_1330) );
na02m20 g67689_u0 ( .a(pciu_bar1_in_392), .b(pciu_am1_in_530), .o(g67689_p) );
in01f08 g67689_u1 ( .a(g67689_p), .o(n_2828) );
no02f08 g67690_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_), .o(n_420) );
na02s10 g67691_u0 ( .a(wbu_addr_in_258), .b(wbu_addr_in_259), .o(n_894) );
no02f02 g67692_u0 ( .a(n_497), .b(n_1023), .o(n_798) );
no02m01 g67694_u0 ( .a(n_15302), .b(n_978), .o(n_1251) );
no02m06 g67695_u0 ( .a(wbs_err_o), .b(wbs_rty_o), .o(n_3083) );
no02m06 g67698_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .o(n_1440) );
na02m20 g67699_u0 ( .a(conf_wb_err_addr_in_948), .b(conf_wb_err_addr_in_949), .o(g67699_p) );
in01f08 g67699_u1 ( .a(g67699_p), .o(n_1165) );
in01s02 g67700_u0 ( .a(n_528), .o(n_529) );
na02s10 g67701_u0 ( .a(conf_wb_err_addr_in_967), .b(conf_wb_err_addr_in_966), .o(n_528) );
na02f20 g67702_u0 ( .a(n_1263), .b(pci_target_unit_wishbone_master_rty_counter_3_), .o(n_906) );
no02s02 g67703_u0 ( .a(wishbone_slave_unit_pcim_if_del_burst_in), .b(wishbone_slave_unit_fifos_wbr_be_in), .o(n_294) );
na02m03 g67704_u0 ( .a(wbm_adr_o_20_), .b(wbm_adr_o_21_), .o(n_910) );
na02m06 g67705_u0 ( .a(wbm_adr_o_10_), .b(wbm_adr_o_9_), .o(n_897) );
no02m10 g67706_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_), .o(n_409) );
na02m20 g67707_u0 ( .a(pciu_bar1_in_397), .b(pciu_am1_in_535), .o(g67707_p) );
in01f08 g67707_u1 ( .a(g67707_p), .o(n_2856) );
no02s01 g67709_u0 ( .a(n_526), .b(wishbone_slave_unit_del_sync_bc_out_reg_1__Q), .o(g67709_p) );
in01s01 g67709_u1 ( .a(g67709_p), .o(n_527) );
na02f03 g67710_u0 ( .a(conf_wb_err_addr_in_953), .b(conf_wb_err_addr_in_954), .o(n_885) );
na02m20 g67712_u0 ( .a(pciu_bar1_in_391), .b(pciu_am1_in_529), .o(g67712_p) );
in01f08 g67712_u1 ( .a(g67712_p), .o(n_2835) );
na02m10 g67713_u0 ( .a(pciu_am1_in_518), .b(parchk_pci_ad_reg_in_1213), .o(n_298) );
na02m03 g67714_u0 ( .a(wbm_adr_o_7_), .b(wbm_adr_o_8_), .o(n_977) );
na02s06 g67715_u0 ( .a(wbu_addr_in_262), .b(wbu_addr_in_263), .o(n_404) );
na02s04 g67716_u0 ( .a(wbm_adr_o_4_), .b(wbm_adr_o_5_), .o(n_405) );
na02m03 g67717_u0 ( .a(wbm_adr_o_18_), .b(wbm_adr_o_17_), .o(n_917) );
no02f20 g67720_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_), .o(n_407) );
no02s02 g67721_u0 ( .a(wbs_adr_i_2_), .b(wbs_adr_i_3_), .o(g67721_p) );
in01s01 g67721_u1 ( .a(g67721_p), .o(n_748) );
na02m10 g67722_u0 ( .a(pciu_am1_in_533), .b(parchk_pci_ad_reg_in_1228), .o(g67722_p) );
in01f06 g67722_u1 ( .a(g67722_p), .o(n_227) );
in01s01 g67723_u0 ( .a(n_8486), .o(n_2483) );
no02s01 g67724_u0 ( .a(n_2314), .b(n_2629), .o(n_8486) );
na02m06 g67725_u0 ( .a(wbs_stb_i), .b(wbs_cyc_i), .o(g67725_p) );
in01s04 g67725_u1 ( .a(g67725_p), .o(n_1347) );
na02s03 g67726_u0 ( .a(wbu_addr_in_279), .b(n_261), .o(n_524) );
no02m08 g67727_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .o(n_408) );
no02m10 g67730_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_), .o(n_364) );
na02s03 g67731_u0 ( .a(wbu_addr_in_276), .b(wbu_addr_in_275), .o(g67731_p) );
in01s01 g67731_u1 ( .a(g67731_p), .o(n_1285) );
no02m10 g67734_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_), .o(n_342) );
na02s06 g67735_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_5_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_6_), .o(g67735_p) );
in01s03 g67735_u1 ( .a(g67735_p), .o(n_1689) );
in01s01 g67736_u0 ( .a(n_522), .o(n_523) );
na02s01 g67737_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_12_), .b(pci_target_unit_del_sync_comp_cycle_count_13_), .o(n_522) );
na02m20 g67739_u0 ( .a(pciu_bar1_in_395), .b(pciu_am1_in_533), .o(g67739_p) );
in01f08 g67739_u1 ( .a(g67739_p), .o(n_2815) );
in01s04 g67741_u0 ( .a(n_881), .o(n_521) );
na02s40 g67742_u0 ( .a(conf_wb_err_addr_in_952), .b(conf_wb_err_addr_in_951), .o(n_881) );
no02s08 g67744_u0 ( .a(conf_wb_err_bc_in_847), .b(conf_wb_err_bc_in_848), .o(n_329) );
na02f10 g67745_u0 ( .a(n_653), .b(n_1724), .o(g67745_p) );
in01f08 g67745_u1 ( .a(g67745_p), .o(n_7044) );
na02m20 g67746_u0 ( .a(pciu_bar1_in_386), .b(pciu_am1_in_524), .o(g67746_p) );
in01f08 g67746_u1 ( .a(g67746_p), .o(n_2831) );
na02m20 g67747_u0 ( .a(pciu_bar1_in_401), .b(pciu_am1_in_539), .o(g67747_p) );
in01f08 g67747_u1 ( .a(g67747_p), .o(n_2851) );
na02m06 g67748_u0 ( .a(wbu_addr_in_258), .b(wbu_addr_in_257), .o(n_946) );
no02s02 g67749_u0 ( .a(pci_target_unit_wishbone_master_read_count_1_), .b(pci_target_unit_wishbone_master_read_count_0_), .o(n_987) );
no02f20 g67750_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_1_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_), .o(n_320) );
no02m06 g67751_u0 ( .a(pci_target_unit_pci_target_sm_n_3), .b(pci_target_unit_pci_target_sm_n_2), .o(n_520) );
na02s20 g67752_u0 ( .a(wbu_addr_in_256), .b(wbu_addr_in_255), .o(n_884) );
na02s06 g67753_u0 ( .a(wbu_addr_in_271), .b(wbu_addr_in_270), .o(n_902) );
na02m08 g67754_u0 ( .a(conf_wb_err_addr_in_950), .b(conf_wb_err_addr_in_951), .o(g67754_p) );
in01m04 g67754_u1 ( .a(g67754_p), .o(n_411) );
na02f04 g67755_u0 ( .a(pciu_am1_in_527), .b(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(n_300) );
na02m03 g67756_u0 ( .a(wbm_adr_o_20_), .b(wbm_adr_o_19_), .o(n_916) );
na02m10 g67757_u0 ( .a(conf_wb_err_addr_in_958), .b(conf_wb_err_addr_in_959), .o(g67757_p) );
in01m06 g67757_u1 ( .a(g67757_p), .o(n_912) );
na02s01 g67758_u0 ( .a(conf_pci_init_complete_out), .b(configuration_sync_command_bit6), .o(g67758_p) );
in01s01 g67758_u1 ( .a(g67758_p), .o(n_13766) );
na02m10 g67759_u0 ( .a(pciu_am1_in_523), .b(parchk_pci_ad_reg_in_1218), .o(n_413) );
in01s01 g67760_u0 ( .a(n_518), .o(n_519) );
na02m03 g67761_u0 ( .a(wbm_adr_o_25_), .b(wbm_adr_o_26_), .o(n_518) );
no02f20 g67762_u0 ( .a(n_1628), .b(pci_target_unit_pci_target_sm_n_2), .o(n_976) );
no02f20 g67763_u0 ( .a(wishbone_slave_unit_wishbone_slave_img_hit_1_), .b(wishbone_slave_unit_wishbone_slave_img_hit_0_), .o(g67763_p) );
in01f10 g67763_u1 ( .a(g67763_p), .o(n_412) );
no02s08 g67764_u0 ( .a(n_657), .b(pci_target_unit_pcit_if_req_req_pending_in), .o(n_791) );
na02m20 g67765_u0 ( .a(pciu_bar1_in_393), .b(pciu_am1_in_531), .o(g67765_p) );
in01f08 g67765_u1 ( .a(g67765_p), .o(n_2864) );
no02f01 g67766_u0 ( .a(n_16690), .b(n_2078), .o(n_1248) );
na02s02 g67768_u0 ( .a(n_440), .b(n_16070), .o(n_1215) );
na02s01 g67770_u0 ( .a(parchk_pci_trdy_en_in), .b(output_backup_devsel_out_reg_Q), .o(n_1505) );
no02m03 g67771_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .o(n_1315) );
no02s01 g67772_u0 ( .a(n_961), .b(n_333), .o(n_727) );
na02m02 g67773_u0 ( .a(wishbone_slave_unit_wishbone_slave_c_state_1), .b(wishbone_slave_unit_wishbone_slave_c_state_2), .o(n_790) );
no02s01 g67774_u0 ( .a(wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q), .b(wishbone_slave_unit_wishbone_slave_pref_en_reg_Q), .o(n_665) );
na02m10 g67775_u0 ( .a(pciu_am1_in_521), .b(parchk_pci_ad_reg_in_1216), .o(n_297) );
na02m20 g67778_u0 ( .a(pciu_bar1_in_380), .b(pciu_am1_in_518), .o(g67778_p) );
in01f08 g67778_u1 ( .a(g67778_p), .o(n_2838) );
na02s06 g67779_u0 ( .a(wbu_addr_in_269), .b(wbu_addr_in_268), .o(n_877) );
na02s10 g67780_u0 ( .a(wbu_addr_in_260), .b(wbu_addr_in_261), .o(n_918) );
na02m10 g67783_u0 ( .a(pciu_am1_in_537), .b(parchk_pci_ad_reg_in_1232), .o(g67783_p) );
in01f06 g67783_u1 ( .a(g67783_p), .o(n_302) );
na02m03 g67785_u0 ( .a(wbm_adr_o_12_), .b(wbm_adr_o_11_), .o(n_896) );
no02s01 g67786_u0 ( .a(wbu_cache_line_size_in_209), .b(wbu_cache_line_size_in_208), .o(n_432) );
no02s04 g67787_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_8_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_9_), .o(n_928) );
na02m10 g67788_u0 ( .a(pciu_am1_in_524), .b(parchk_pci_ad_reg_in_1219), .o(n_303) );
na02s02 g67791_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_3_), .b(pci_target_unit_wishbone_master_rty_counter_4_), .o(g67791_p) );
in01s02 g67791_u1 ( .a(g67791_p), .o(n_929) );
na02m03 g67792_u0 ( .a(wbm_adr_o_22_), .b(wbm_adr_o_23_), .o(n_941) );
in01s01 g67793_u0 ( .a(n_512), .o(n_513) );
na02m03 g67794_u0 ( .a(wbu_addr_in_274), .b(wbu_addr_in_273), .o(n_512) );
in01m01 g67797_u0 ( .a(n_16307), .o(n_1057) );
na02m20 g67799_u0 ( .a(pciu_bar1_in_400), .b(pciu_am1_in_538), .o(g67799_p) );
in01f08 g67799_u1 ( .a(g67799_p), .o(n_2854) );
no02s02 g67800_u0 ( .a(wishbone_slave_unit_pcim_if_del_burst_in), .b(wishbone_slave_unit_fifos_wbr_be_in_265), .o(n_236) );
no02s01 g67801_u0 ( .a(n_16685), .b(n_15746), .o(n_2125) );
na02s03 g67802_u0 ( .a(n_1111), .b(wishbone_slave_unit_pcim_sm_be_in_557), .o(g67802_p) );
in01s01 g67802_u1 ( .a(g67802_p), .o(n_1013) );
na02s20 g67803_u0 ( .a(conf_wb_err_addr_in_943), .b(conf_wb_err_addr_in_944), .o(n_568) );
na02s02 g67804_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_3_), .b(pci_target_unit_del_sync_comp_cycle_count_4_), .o(g67804_p) );
in01s02 g67804_u1 ( .a(g67804_p), .o(n_1187) );
na02s08 g67805_u0 ( .a(conf_wb_err_addr_in_955), .b(conf_wb_err_addr_in_952), .o(n_306) );
na02s03 g67806_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_3_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_4_), .o(g67806_p) );
in01s02 g67806_u1 ( .a(g67806_p), .o(n_1186) );
na02s10 g67807_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_1_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_0_), .o(g67807_p) );
in01s06 g67807_u1 ( .a(g67807_p), .o(n_947) );
in01s01 g67808_u0 ( .a(n_784), .o(n_785) );
na02s02 g67809_u0 ( .a(n_206), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q), .o(n_784) );
no02m08 g67810_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_1_), .o(n_433) );
na02m06 g67811_u0 ( .a(conf_wb_err_addr_in_964), .b(conf_wb_err_addr_in_963), .o(n_904) );
na02m03 g67812_u0 ( .a(conf_wb_err_addr_in_965), .b(conf_wb_err_addr_in_966), .o(n_903) );
no02s06 g67813_u0 ( .a(n_3415), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .o(n_1294) );
na02s04 g67814_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_8_), .b(pci_target_unit_del_sync_comp_cycle_count_9_), .o(g67814_p) );
in01s02 g67814_u1 ( .a(g67814_p), .o(n_937) );
na02s01 g67817_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .b(wishbone_slave_unit_fifos_wbw_whole_waddr), .o(n_1109) );
no02m02 g67818_u0 ( .a(n_763), .b(n_15932), .o(n_2392) );
na02s20 g67820_u0 ( .a(conf_wb_err_addr_in_959), .b(conf_wb_err_addr_in_960), .o(n_890) );
na02m03 g67822_u0 ( .a(wbm_adr_o_13_), .b(wbm_adr_o_14_), .o(n_899) );
na02m10 g67823_u0 ( .a(pciu_am1_in_531), .b(parchk_pci_ad_reg_in_1226), .o(n_436) );
na02m10 g67824_u0 ( .a(parchk_pci_ad_reg_in_1229), .b(pciu_am1_in_534), .o(n_307) );
no02m04 g67826_u0 ( .a(wbs_ack_o), .b(n_16635), .o(n_783) );
na02f20 g67827_u0 ( .a(wishbone_slave_unit_wishbone_slave_del_addr_hit), .b(wishbone_slave_unit_wishbone_slave_del_completion_allow), .o(n_319) );
na02m10 g67828_u0 ( .a(pciu_bar1_in), .b(pciu_am1_in), .o(g67828_p) );
in01f06 g67828_u1 ( .a(g67828_p), .o(n_2844) );
in01s01 g67832_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__260), .o(n_4403) );
in01f80 g67857_u0 ( .a(wbm_rty_i), .o(n_705) );
in01m03 g67868_u0 ( .a(n_1111), .o(n_2263) );
in01s01 g67877_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__243), .o(n_3636) );
in01s01 g67885_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13_), .o(n_4280) );
in01s01 g67936_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__487), .o(n_28) );
in01s06 g67939_u0 ( .a(wishbone_slave_unit_pcim_sm_last_in), .o(n_5757) );
in01s01 g67945_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__258), .o(n_156) );
in01s01 g67948_u0 ( .a(wishbone_slave_unit_pci_initiator_if_read_count_2_), .o(n_9) );
in01s01 g67969_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__70), .o(n_4312) );
in01s03 g67991_u0 ( .a(n_689), .o(n_8876) );
in01s10 g67993_u0 ( .a(pci_target_unit_fifos_pcir_whole_waddr), .o(n_689) );
in01s01 g68021_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__46), .o(n_3763) );
in01s01 g68029_u0 ( .a(n_1263), .o(n_221) );
in01s01 g68042_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__236), .o(n_4399) );
in01f40 g68103_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_0_), .o(n_1280) );
in01s01 g68110_u0 ( .a(wbu_pci_drcomp_pending_in), .o(n_1816) );
in01s20 g68132_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_rdata_selector), .o(n_541) );
in01s01 g68160_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_0_), .o(n_321) );
in01s01 g68163_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_14__582), .o(n_317) );
in01m01 g68172_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_mabort1), .o(n_188) );
in01s01 g68212_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_7__310), .o(n_7373) );
in01s01 g68217_u0 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_1_), .o(n_362) );
in01m20 g68225_u0 ( .a(n_324), .o(n_13447) );
in01m10 g68229_u0 ( .a(n_324), .o(n_504) );
in01m40 g68230_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_rdata_selector_14), .o(n_324) );
in01s01 g68239_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_15__622), .o(n_323) );
in01s01 g68251_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__43), .o(n_95) );
in01s01 g68277_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_0_), .o(n_276) );
in01s02 g68284_u0 ( .a(wbu_pciif_frame_out_in), .o(n_3022) );
in01s01 g68315_u0 ( .a(pci_target_unit_del_sync_addr_in_204), .o(n_2598) );
in01s01 g68318_u0 ( .a(wishbone_slave_unit_del_sync_req_done_reg), .o(n_325) );
in01s01 g68325_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_2__6), .o(n_75) );
in01s01 g68332_u0 ( .a(pci_target_unit_fifos_inGreyCount_0_), .o(n_42) );
in01s01 g68346_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__380), .o(n_74) );
in01s01 g68356_u0 ( .a(pci_frame_o), .o(n_67) );
in01m01 g68368_u0 ( .a(wbs_ack_o), .o(n_779) );
in01m02 g68369_u0 ( .a(n_326), .o(wbs_ack_o) );
in01m20 g68370_u0 ( .a(wbs_ack_o_1307), .o(n_326) );
in01s20 g68381_u0 ( .a(wishbone_slave_unit_wbs_sm_del_req_pending_in), .o(n_709) );
in01s01 g68389_u0 ( .a(pci_target_unit_del_sync_addr_in_209), .o(n_2512) );
in01s01 g68393_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__183), .o(n_6) );
in01s01 g68398_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__238), .o(n_4396) );
in01s01 g68401_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__377), .o(n_139) );
in01s01 g68410_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__376), .o(n_3665) );
in01m10 g68420_u0 ( .a(n_525), .o(n_1023) );
in01f80 g68421_u0 ( .a(conf_w_addr_in_939), .o(n_525) );
in01m06 g68423_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr), .o(n_2) );
in01s01 g68426_u0 ( .a(n_2), .o(n_8953) );
in01s01 g68439_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_0_), .o(n_282) );
in01s03 g68448_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_11_), .o(n_193) );
in01s01 g68452_u0 ( .a(configuration_set_isr_bit2), .o(n_72) );
in01s01 g68454_u0 ( .a(pci_target_unit_del_sync_addr_in_210), .o(n_2541) );
in01s01 g68465_u0 ( .a(pci_target_unit_del_sync_addr_in_212), .o(n_2503) );
in01m08 g68472_u0 ( .a(n_2314), .o(n_5755) );
in01m20 g68485_u0 ( .a(n_1061), .o(n_8511) );
in01s01 g68501_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__247), .o(n_4410) );
in01f06 g68509_u0 ( .a(wbu_pciif_devsel_reg_in), .o(n_707) );
in01s02 g68515_u0 ( .a(n_551), .o(n_497) );
in01f10 g68516_u0 ( .a(conf_w_addr_in_938), .o(n_551) );
in01s01 g68522_u0 ( .a(n_333), .o(n_447) );
in01s01 g68523_u0 ( .a(parchk_pci_frame_en_in), .o(n_333) );
in01s01 g68548_u0 ( .a(configuration_pci_err_cs_bit0), .o(n_200) );
in01m06 g68550_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_), .o(n_160) );
in01m06 g68572_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .o(n_349) );
in01s02 g68604_u0 ( .a(pci_target_unit_fifos_outGreyCount_0_), .o(n_202) );
in01s01 g68613_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__237), .o(n_3738) );
in01s01 g68616_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_11__466), .o(n_351) );
in01s01 g68622_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__248), .o(n_0) );
in01m10 g68642_u0 ( .a(wbu_addr_in_280), .o(n_539) );
in01s08 g68652_u0 ( .a(pciu_pciif_bckp_stop_in), .o(n_205) );
in01f20 g68658_u0 ( .a(wishbone_slave_unit_wishbone_slave_c_state_1), .o(n_279) );
in01s06 g68674_u0 ( .a(parchk_pci_irdy_en_in), .o(n_961) );
in01s01 g68681_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__51), .o(n_17) );
in01s01 g68683_u0 ( .a(wbs_bte_i_0_), .o(n_23) );
in01s01 g68703_u0 ( .a(pci_target_unit_del_sync_addr_in), .o(n_2671) );
in01s01 g68707_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__309), .o(n_337) );
in01s01 g68759_u0 ( .a(pci_target_unit_del_sync_addr_in_211), .o(n_2507) );
in01s06 g68771_u0 ( .a(wbm_adr_o_2_), .o(n_208) );
in01s01 g68773_u0 ( .a(pci_target_unit_fifos_pciw_outTransactionCount_1_), .o(n_996) );
in01s02 g68776_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_12_), .o(n_206) );
in01s06 g68778_u0 ( .a(n_691), .o(n_692) );
in01m02 g68787_u0 ( .a(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(n_691) );
in01s01 g68814_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__358), .o(n_40) );
in01f10 g68832_u0 ( .a(n_2071), .o(n_3030) );
in01s01 g68839_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__544), .o(n_263) );
in01s02 g68852_u0 ( .a(n_2648), .o(n_2044) );
in01f10 g68853_u0 ( .a(n_15854), .o(n_2648) );
in01s06 g68866_u0 ( .a(n_573), .o(n_3415) );
in01s20 g68867_u0 ( .a(pci_target_unit_fifos_pciw_whole_waddr), .o(n_573) );
in01s01 g68882_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_), .o(n_148) );
in01s01 g68888_u0 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_1_), .o(n_345) );
in01s01 g68917_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_13__543), .o(n_354) );
in01s03 g68929_u0 ( .a(n_285), .o(n_574) );
in01s02 g68941_u0 ( .a(n_285), .o(n_2373) );
in01s01 g68942_u0 ( .a(conf_pci_init_complete_out), .o(n_285) );
in01s01 g68949_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in), .o(n_181) );
in01s01 g68961_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__359), .o(n_4323) );
in01s01 g68971_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_2__231), .o(n_366) );
in01s01 g68991_u0 ( .a(n_15856), .o(n_2087) );
na02f04 g68_u0 ( .a(n_16566), .b(n_16105), .o(g68_p) );
in01f06 g68_u1 ( .a(g68_p), .o(n_16992) );
in01s01 g69007_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__360), .o(n_119) );
in01m10 g69013_u0 ( .a(pci_target_unit_pci_target_if_keep_desconnect_wo_data_set), .o(n_8728) );
in01f20 g69023_u0 ( .a(pci_target_unit_wishbone_master_addr_into_cnt_reg), .o(n_168) );
in01f20 g69033_u0 ( .a(n_1628), .o(n_278) );
in01s01 g69050_u0 ( .a(pci_target_unit_del_sync_addr_in_205), .o(n_2515) );
in01m04 g69063_u0 ( .a(wishbone_slave_unit_wishbone_slave_c_state_2), .o(n_288) );
in01m02 g69074_u0 ( .a(n_15249), .o(n_7114) );
in01s01 g69089_u0 ( .a(pci_target_unit_del_sync_addr_in_207), .o(n_2526) );
in01s01 g69092_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__484), .o(n_83) );
in01s02 g69098_u0 ( .a(pci_target_unit_pci_target_sm_wr_progress), .o(n_2311) );
in01f20 g69104_u0 ( .a(pci_target_unit_pcit_if_req_req_pending_in), .o(n_373) );
in01s08 g69114_u0 ( .a(wbu_addr_in_278), .o(n_261) );
in01s03 g69135_u0 ( .a(pciu_pciif_stop_reg_in), .o(n_378) );
in01m08 g69146_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_), .o(n_440) );
in01f20 g69180_u0 ( .a(pci_target_unit_pci_target_sm_n_3), .o(n_61) );
in01f20 g69207_u0 ( .a(wishbone_slave_unit_wishbone_slave_map), .o(n_1323) );
in01f06 g69209_u0 ( .a(n_15331), .o(n_2092) );
in01s01 g69218_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__67), .o(n_38) );
in01s01 g69220_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__177), .o(n_18) );
in01s01 g69230_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__265), .o(n_50) );
in01s01 g69252_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_3__270), .o(n_271) );
in01s01 g69259_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_), .o(n_76) );
in01f08 g69271_u0 ( .a(n_16284), .o(n_1519) );
in01s01 g69285_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_686), .o(n_85) );
in01s01 g69321_u0 ( .a(pci_target_unit_pci_target_sm_rd_progress), .o(n_243) );
in01m01 g69337_u0 ( .a(wishbone_slave_unit_pcim_sm_be_in_559), .o(n_57) );
in01f10 g69362_u0 ( .a(pci_target_unit_wbm_sm_pci_tar_burst_ok), .o(n_815) );
in01s01 g69364_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__365), .o(n_4429) );
in01s01 g69369_u0 ( .a(wishbone_slave_unit_pcim_if_del_req_in), .o(n_169) );
in01s01 g69378_u0 ( .a(pci_target_unit_del_sync_comp_rty_exp_reg), .o(n_1817) );
in01s01 g69418_u0 ( .a(wishbone_slave_unit_pcim_if_del_bc_in_382), .o(n_213) );
in01m06 g69428_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .o(n_242) );
in01s01 g69431_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_8_), .o(n_882) );
in01s01 g69436_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__522), .o(n_12) );
in01s01 g69457_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__249), .o(n_3691) );
in01s01 g69489_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_9_), .o(n_1992) );
in01s01 g69505_u0 ( .a(pci_target_unit_del_sync_addr_in_206), .o(n_2499) );
in01f40 g69532_u0 ( .a(n_657), .o(n_565) );
in01s01 g69534_u0 ( .a(pci_resi_conf_soft_res_in), .o(n_123) );
in01s01 g69550_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_0__153), .o(n_384) );
in01f01 g69558_u0 ( .a(n_763), .o(n_2316) );
in01f08 g69561_u0 ( .a(n_629), .o(n_763) );
in01f20 g69562_u0 ( .a(n_16285), .o(n_629) );
in01s01 g69576_u0 ( .a(wishbone_slave_unit_pcim_if_del_bc_in_383), .o(n_211) );
in01s01 g69593_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_), .o(n_11) );
in01s01 g69609_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__374), .o(n_65) );
in01s01 g69632_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__509), .o(n_14) );
in01s01 g69640_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__178), .o(n_27) );
in01s01 g69643_u0 ( .a(wbu_cache_line_size_in_207), .o(n_292) );
in01f08 g69650_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_3_), .o(n_135) );
in01s01 g69652_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__342), .o(n_84) );
in01s01 g69673_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__330), .o(n_26) );
in01s01 g69686_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_1_), .o(n_150) );
in01f10 g69707_u0 ( .a(n_391), .o(n_1104) );
in01f40 g69708_u0 ( .a(pci_target_unit_wishbone_master_c_state_0_), .o(n_391) );
in01m01 g69724_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_1_), .o(n_247) );
in01s01 g69746_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_15__621), .o(n_393) );
in01s01 g69749_u0 ( .a(wbs_err_o), .o(n_471) );
in01s03 g69750_u0 ( .a(n_15204), .o(wbs_err_o) );
in01m06 g69754_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .o(n_143) );
in01s10 g69761_u0 ( .a(n_1293), .o(n_1316) );
in01f10 g69775_u0 ( .a(n_2509), .o(n_396) );
in01s01 g69786_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_14__583), .o(n_395) );
in01s01 g69794_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_decode_count_0_), .o(n_401) );
in01s01 g69797_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__532), .o(n_15) );
in01s06 g69799_u0 ( .a(wishbone_slave_unit_pcim_if_del_we_in), .o(n_4078) );
in01s01 g69804_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_11__465), .o(n_251) );
in01m08 g69834_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_0_), .o(n_46) );
in01s01 g69845_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__56), .o(n_4394) );
in01s01 g69855_u0 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_0_), .o(n_397) );
in01s01 g69856_u0 ( .a(configuration_wb_err_cs_bit0), .o(n_24) );
in01s03 g69886_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_10_), .o(n_245) );
in01s01 g69888_u0 ( .a(wishbone_slave_unit_fifos_inGreyCount_0_), .o(n_22) );
in01s01 g69901_u0 ( .a(pci_target_unit_pci_target_if_same_read_reg), .o(n_152) );
in01m03 g69904_u0 ( .a(pci_gnt_i), .o(n_47) );
in01s01 g69937_u0 ( .a(pci_devsel_i), .o(n_34) );
in01s01 g69939_u0 ( .a(wbm_cti_o_1_), .o(n_112) );
in01m04 g69962_u0 ( .a(n_2308), .o(n_2742) );
in01s40 g69963_u0 ( .a(n_15924), .o(n_2308) );
in01s01 g70007_u0 ( .a(pci_target_unit_del_sync_addr_in_208), .o(n_2544) );
in01s10 g70023_u0 ( .a(n_1117), .o(n_1174) );
in01s01 g70029_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_10_), .o(n_207) );
in01s06 g70054_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_7_), .o(n_104) );
in01s01 g70062_u0 ( .a(n_16175), .o(n_13608) );
in01f20 g70068_u0 ( .a(pci_target_unit_pci_target_sm_cnf_progress), .o(n_653) );
in01m10 g70083_u0 ( .a(n_1724), .o(n_2629) );
in01f40 g70086_u0 ( .a(n_978), .o(n_1724) );
in01s01 g70097_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_1__192), .o(n_255) );
in01s01 g70100_u0 ( .a(wishbone_slave_unit_pci_initiator_if_read_count_3_), .o(n_416) );
in01s01 g70132_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__536), .o(n_4273) );
in01s01 g70154_u0 ( .a(wbm_ack_i), .o(n_1183) );
in01f40 g70183_u0 ( .a(pci_target_unit_wishbone_master_c_state_2_), .o(n_681) );
in01s01 g70191_u0 ( .a(FE_OCP_RBN2277_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_), .o(n_358) );
in01s01 g70203_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__379), .o(n_4343) );
in01s01 g70209_u0 ( .a(pci_target_unit_fifos_pciw_inTransactionCount_1_), .o(n_852) );
in01f08 g70215_u0 ( .a(n_15330), .o(n_696) );
in01s01 g70227_u0 ( .a(wishbone_slave_unit_pcim_if_del_burst_in), .o(n_21) );
in01s01 g70251_u0 ( .a(wishbone_slave_unit_pcim_if_del_bc_in), .o(n_526) );
in01m10 g70258_u0 ( .a(conf_wb_err_bc_in_847), .o(n_715) );
in01s01 g70269_u0 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_0_), .o(n_425) );
in01s01 g70281_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__271), .o(n_424) );
in01m01 g70305_u0 ( .a(n_1698), .o(n_2651) );
in01f10 g70310_u0 ( .a(parchk_pci_cbe_reg_in_1236), .o(n_1698) );
in01s01 g70414_u0 ( .a(pci_target_unit_pci_target_sm_rd_request), .o(n_177) );
in01s01 g70418_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__62), .o(n_3608) );
in01s01 g70425_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__363), .o(n_3672) );
in01s01 g70441_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__47), .o(n_36) );
in01s01 g70451_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__59), .o(n_3616) );
in01m02 g70465_u0 ( .a(parchk_pci_trdy_en_in), .o(n_454) );
na02f02 g70_u0 ( .a(n_16566), .b(n_8860), .o(g70_p) );
in01f03 g70_u1 ( .a(g70_p), .o(n_15534) );
no02f02 g71_u0 ( .a(n_12151), .b(n_10669), .o(n_15527) );
in01m01 g73860_u0 ( .a(n_14967), .o(n_14965) );
in01f06 g73876_u0 ( .a(FE_OCPN1827_n_14995), .o(n_15001) );
na02s02 TIMEBOOST_cell_40624 ( .a(TIMEBOOST_net_12550), .b(g62691_sb), .o(n_6164) );
na02s01 TIMEBOOST_cell_45571 ( .a(g64785_db), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__Q), .o(TIMEBOOST_net_15024) );
no02f08 g73934_u0 ( .a(n_16287), .b(n_1408), .o(n_15125) );
no02f06 g73935_u0 ( .a(n_16291), .b(n_16033), .o(n_15128) );
na02f02 g73947_u0 ( .a(n_16156), .b(n_15388), .o(n_15142) );
oa12m02 g73970_u0 ( .a(n_15196), .b(n_15187), .c(FE_OFN2164_n_16301), .o(n_15197) );
ao12f02 g73971_u0 ( .a(n_14730), .b(n_14800), .c(wbm_dat_o_10_), .o(n_15187) );
na02s02 TIMEBOOST_cell_43597 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__Q), .b(n_3734), .o(TIMEBOOST_net_14037) );
na02f02 g73977_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_10_), .o(n_15196) );
in01f40 g73986_u0 ( .a(wbs_err_o_1309), .o(n_15204) );
no02f08 g73989_u0 ( .a(n_16284), .b(n_16285), .o(g73989_p) );
in01f06 g73989_u1 ( .a(g73989_p), .o(n_15210) );
in01f02 g73996_u0 ( .a(n_15389), .o(n_15217) );
in01f20 g74023_u0 ( .a(n_16501), .o(n_15249) );
na02s04 g74027_u0 ( .a(n_15260), .b(wishbone_slave_unit_pci_initiator_if_posted_write_req), .o(n_15261) );
na02f08 g74028_u0 ( .a(n_4718), .b(n_15805), .o(g74028_p) );
in01f06 g74028_u1 ( .a(g74028_p), .o(n_15260) );
in01f02 g74031_u0 ( .a(n_15260), .o(n_15262) );
na02f02 g74037_u0 ( .a(n_15994), .b(n_15275), .o(n_15276) );
in01f08 g74038_u0 ( .a(n_16287), .o(n_15275) );
in01f04 g74050_u0 ( .a(n_16002), .o(n_15291) );
na02f02 g74053_u0 ( .a(n_3452), .b(n_1251), .o(n_15292) );
na02f02 g74059_u0 ( .a(n_15614), .b(n_15292), .o(n_15301) );
in01f03 g74061_u0 ( .a(n_15295), .o(n_15302) );
na03s02 TIMEBOOST_cell_5791 ( .a(n_3785), .b(g65041_sb), .c(g65041_db), .o(n_3624) );
no02f20 g74074_u0 ( .a(n_16964), .b(n_15313), .o(n_15314) );
in01f40 g74075_u0 ( .a(wbs_stb_i), .o(n_15313) );
na02s02 TIMEBOOST_cell_43014 ( .a(TIMEBOOST_net_13745), .b(g63101_sb), .o(n_5052) );
na02f06 g74082_u0 ( .a(n_2447), .b(n_2392), .o(n_15324) );
in01f10 g74087_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_cur_state_1_), .o(n_15330) );
in01f08 g74088_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_cur_state_0_), .o(n_15331) );
no02f20 g74121_u0 ( .a(parchk_pci_frame_reg_in), .b(parchk_pci_frame_en_in), .o(n_15365) );
in01f10 g74122_u0 ( .a(parchk_pci_frame_reg_in), .o(n_15295) );
na02f02 g74124_u0 ( .a(n_16560), .b(n_15372), .o(n_15373) );
no02f06 g74126_u0 ( .a(n_15370), .b(n_15371), .o(n_15372) );
in01f02 g74129_u0 ( .a(n_15371), .o(n_15376) );
na02f20 g74140_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_5_), .b(pci_target_unit_wishbone_master_rty_counter_7_), .o(g74140_p) );
in01f08 g74140_u1 ( .a(g74140_p), .o(n_15385) );
na02f06 g74141_u0 ( .a(n_16980), .b(n_1445), .o(n_15388) );
na02f03 g74142_u0 ( .a(n_16154), .b(n_16150), .o(n_15390) );
in01f06 g74147_u0 ( .a(n_16495), .o(n_15397) );
na02m01 g74153_u0 ( .a(pci_target_unit_pci_target_sm_same_read_reg), .b(n_1724), .o(g74153_p) );
in01s02 g74153_u1 ( .a(g74153_p), .o(n_15405) );
na02f04 g74154_u0 ( .a(pci_target_unit_pci_target_sm_rd_from_fifo), .b(FE_OCPN1836_n_16798), .o(g74154_p) );
in01f02 g74154_u1 ( .a(g74154_p), .o(n_15406) );
no02f02 g74155_u0 ( .a(n_1435), .b(pci_target_unit_pci_target_sm_cnf_progress), .o(n_15407) );
na02f08 g74162_dup_u0 ( .a(n_16949), .b(n_16635), .o(g74162_dup_p) );
in01f06 g74162_dup_u1 ( .a(g74162_dup_p), .o(n_16855) );
na02s01 TIMEBOOST_cell_38540 ( .a(TIMEBOOST_net_11508), .b(g62044_sb), .o(n_7768) );
no02f04 g74173_u0 ( .a(n_15446), .b(n_15467), .o(n_15442) );
na02f06 g74174_u0 ( .a(n_15065), .b(n_2129), .o(g74174_p) );
in01f08 g74174_u1 ( .a(g74174_p), .o(n_15444) );
na02f02 TIMEBOOST_cell_22161 ( .a(TIMEBOOST_net_6337), .b(FE_OFN1600_n_13995), .o(n_14467) );
na02m04 TIMEBOOST_cell_36831 ( .a(n_4160), .b(FE_OFN1700_n_5751), .o(TIMEBOOST_net_10654) );
in01f04 g74183_u0 ( .a(n_16160), .o(n_15456) );
na02f04 g74191_u0 ( .a(n_15918), .b(n_15908), .o(n_15467) );
no02f08 g74197_u0 ( .a(n_15924), .b(n_15998), .o(n_15474) );
no02f02 g74218_u0 ( .a(n_15514), .b(n_15515), .o(n_15516) );
no02f02 g74220_u0 ( .a(n_15512), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_1_), .o(n_15513) );
na02f08 g74221_u0 ( .a(n_8653), .b(n_8657), .o(n_15515) );
in01f04 g74222_u0 ( .a(n_15514), .o(n_15517) );
in01f10 g74224_u0 ( .a(n_15518), .o(n_8747) );
no02f08 g74225_u0 ( .a(n_15397), .b(n_15403), .o(n_15518) );
ao12f02 g74239_u0 ( .a(n_15553), .b(n_14918), .c(n_16810), .o(n_16853) );
na02f02 g74240_u0 ( .a(n_15549), .b(n_15552), .o(n_15553) );
ao22f02 g74241_u0 ( .a(n_2831), .b(FE_OCPN1845_n_16427), .c(FE_OFN1063_n_15808), .d(configuration_pci_err_data_516), .o(n_15549) );
ao12f02 g74242_u0 ( .a(n_15551), .b(FE_OFN1069_n_15729), .c(configuration_wb_err_data_585), .o(n_15552) );
na02f04 g74243_u0 ( .a(n_16791), .b(pciu_bar0_in_363), .o(g74243_p) );
in01f02 g74243_u1 ( .a(g74243_p), .o(n_15551) );
no02f02 g74245_u0 ( .a(n_15594), .b(n_11739), .o(g74245_p) );
in01f02 g74245_u1 ( .a(g74245_p), .o(n_15565) );
oa22f01 g74248_u0 ( .a(n_15560), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_6__252), .c(n_16572), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__291), .o(n_15562) );
in01f06 g74249_u0 ( .a(FE_OFN1502_n_15558), .o(n_15560) );
in01f06 g74251_u0 ( .a(n_16572), .o(n_15566) );
in01f06 g74252_u0 ( .a(n_15560), .o(n_15568) );
na02f02 g74266_u0 ( .a(n_9305), .b(n_15584), .o(n_15585) );
na02f02 g74267_u0 ( .a(FE_OFN1529_n_10853), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__Q), .o(n_15584) );
in01f04 g74268_u0 ( .a(FE_OFN1508_n_15587), .o(n_15589) );
na02f02 g74270_u0 ( .a(n_8867), .b(n_8866), .o(g74270_p) );
in01f02 g74270_u1 ( .a(g74270_p), .o(n_15587) );
na02f02 g74272_u0 ( .a(n_10728), .b(n_10144), .o(n_15592) );
na02m08 g74283_u0 ( .a(n_978), .b(n_15295), .o(g74283_p) );
in01m04 g74283_u1 ( .a(g74283_p), .o(n_15607) );
oa12f01 g74287_u0 ( .a(n_15607), .b(n_8819), .c(n_1513), .o(n_15614) );
in01f02 g74313_u0 ( .a(n_15373), .o(n_15638) );
in01m06 g74317_u0 ( .a(n_16560), .o(n_15645) );
na02f20 g74343_u0 ( .a(n_16864), .b(n_16871), .o(n_16940) );
no02f40 g74346_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_cur_state_1_), .b(wishbone_slave_unit_pci_initiator_sm_cur_state_0_), .o(n_15680) );
no02f01 g74357_u0 ( .a(n_15919), .b(n_16911), .o(n_15689) );
ao12f02 g74359_u0 ( .a(n_15698), .b(n_14917), .c(n_16810), .o(n_15699) );
na02s01 TIMEBOOST_cell_44786 ( .a(TIMEBOOST_net_14631), .b(g58071_sb), .o(TIMEBOOST_net_13163) );
ao12f02 g74361_u0 ( .a(n_15694), .b(FE_OFN1069_n_15729), .c(configuration_wb_err_data_584), .o(n_15695) );
na02f02 g74363_u0 ( .a(n_16791), .b(pciu_bar0_in_362), .o(g74363_p) );
in01f02 g74363_u1 ( .a(g74363_p), .o(n_15694) );
na02s01 TIMEBOOST_cell_36399 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__Q), .b(g65850_sb), .o(TIMEBOOST_net_10438) );
na02s01 TIMEBOOST_cell_9198 ( .a(pci_target_unit_fifos_pcir_data_in_165), .b(g65774_sb), .o(TIMEBOOST_net_1166) );
in01f02 g74388_u0 ( .a(n_15732), .o(n_15733) );
na02s01 TIMEBOOST_cell_45005 ( .a(pci_target_unit_fifos_pciw_addr_data_in_132), .b(g64204_sb), .o(TIMEBOOST_net_14741) );
na02s01 TIMEBOOST_cell_37271 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__14__Q), .b(FE_OFN671_n_4505), .o(TIMEBOOST_net_10874) );
na02f02 TIMEBOOST_cell_40980 ( .a(TIMEBOOST_net_12728), .b(g57132_sb), .o(n_11616) );
no02f06 g74406_u0 ( .a(n_1828), .b(n_1829), .o(n_15736) );
no02f06 g74407_u0 ( .a(n_15859), .b(n_15738), .o(n_15739) );
no02f20 g74408_u0 ( .a(wishbone_slave_unit_pci_initiator_if_del_read_req), .b(wishbone_slave_unit_pci_initiator_if_err_recovery), .o(g74408_p) );
in01f08 g74408_u1 ( .a(g74408_p), .o(n_15738) );
in01s01 g74409_u0 ( .a(wishbone_slave_unit_pci_initiator_if_err_recovery), .o(n_15741) );
na02f40 g74416_u0 ( .a(n_525), .b(n_2078), .o(n_15744) );
in01f04 g74423_u0 ( .a(n_15754), .o(n_15756) );
in01f08 g74424_u0 ( .a(n_15744), .o(n_15757) );
in01f04 g74428_u0 ( .a(n_8820), .o(n_15758) );
na02f02 g74429_u0 ( .a(n_4635), .b(n_3810), .o(g74429_p) );
in01f02 g74429_u1 ( .a(g74429_p), .o(n_15759) );
in01m02 g74430_u0 ( .a(n_2416), .o(n_15760) );
no02m06 g74433_u0 ( .a(n_1536), .b(n_1436), .o(n_15762) );
in01s04 g74434_u0 ( .a(parchk_pci_frame_en_in), .o(g74434_sb) );
na02s08 g74434_u1 ( .a(pci_frame_i), .b(g74434_sb), .o(g74434_da) );
na02s08 g74434_u2 ( .a(parchk_pci_frame_en_in), .b(wbu_pciif_frame_out_in), .o(g74434_db) );
na02s10 g74434_u3 ( .a(g74434_da), .b(g74434_db), .o(n_1551) );
na02m02 TIMEBOOST_cell_32594 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__30__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__Q), .o(TIMEBOOST_net_10208) );
in01f01 g74437_u0 ( .a(n_15758), .o(n_15769) );
no02s01 g74455_u0 ( .a(n_3320), .b(n_16512), .o(n_15788) );
no02f20 g74470_u0 ( .a(n_16763), .b(wishbone_slave_unit_pcim_sm_rdy_in), .o(g74470_p) );
in01f08 g74470_u1 ( .a(g74470_p), .o(n_15802) );
no02f08 g74471_u0 ( .a(wbu_pciif_devsel_reg_in), .b(parchk_pci_trdy_reg_in), .o(n_15805) );
no02f10 g74472_u0 ( .a(n_15988), .b(n_16936), .o(n_4718) );
na02f06 g74475_u0 ( .a(n_15128), .b(n_15125), .o(g74475_p) );
in01f06 g74475_u1 ( .a(g74475_p), .o(n_15808) );
na03s02 TIMEBOOST_cell_41979 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__Q), .b(n_4251), .c(FE_OFN1283_n_4097), .o(TIMEBOOST_net_13228) );
in01f20 g74518_u0 ( .a(parchk_pci_cbe_reg_in_1237), .o(n_15854) );
na02s10 g74520_u0 ( .a(n_1238), .b(n_15856), .o(n_15859) );
in01f20 g74522_u0 ( .a(wishbone_slave_unit_pci_initiator_if_del_write_req), .o(n_15856) );
na02f08 g74553_u0 ( .a(n_16462), .b(n_15824), .o(g74553_p) );
in01f08 g74553_u1 ( .a(g74553_p), .o(n_16599) );
na02f02 TIMEBOOST_cell_41164 ( .a(TIMEBOOST_net_12820), .b(g57392_sb), .o(n_11350) );
in01f02 g74563_u1 ( .a(g74563_p), .o(n_15910) );
na02f06 g74573_u0 ( .a(n_319), .b(FE_OCP_RBN2222_n_15347), .o(n_15918) );
na02f04 g74575_u0 ( .a(n_16015), .b(n_16016), .o(n_15920) );
na02f06 g74576_u0 ( .a(n_15928), .b(n_4743), .o(g74576_p) );
in01f10 g74576_u1 ( .a(g74576_p), .o(n_15931) );
na02s02 TIMEBOOST_cell_32047 ( .a(TIMEBOOST_net_9934), .b(FE_OFN1179_n_3476), .o(TIMEBOOST_net_4916) );
na02s02 TIMEBOOST_cell_41904 ( .a(TIMEBOOST_net_13190), .b(n_4061), .o(n_5503) );
in01s01 TIMEBOOST_cell_45872 ( .a(TIMEBOOST_net_15178), .o(TIMEBOOST_net_15179) );
na02f02 g74580_u0 ( .a(n_2016), .b(n_798), .o(g74580_p) );
in01f02 g74580_u1 ( .a(g74580_p), .o(n_15922) );
no02m06 g74581_u0 ( .a(n_16690), .b(n_629), .o(n_15923) );
in01f80 g74583_u0 ( .a(conf_w_addr_in_932), .o(n_15924) );
na02f02 TIMEBOOST_cell_42234 ( .a(TIMEBOOST_net_13355), .b(FE_OFN1384_n_8567), .o(TIMEBOOST_net_12308) );
in01s01 g74586_u0 ( .a(n_2078), .o(n_15932) );
na02f02 g74592_u0 ( .a(FE_OFN1559_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__Q), .o(n_15936) );
no02f04 g74593_u0 ( .a(n_15939), .b(n_12716), .o(n_15940) );
in01f02 g74594_u0 ( .a(n_12924), .o(n_15939) );
no02f02 g74595_u0 ( .a(n_12717), .b(n_12461), .o(n_15941) );
na02f04 g74612_u0 ( .a(n_16334), .b(FE_OCP_RBN2227_g75174_p), .o(n_15969) );
ao12f06 g74627_u0 ( .a(n_1238), .b(n_15982), .c(n_15980), .o(n_15985) );
na02f08 g74628_u0 ( .a(n_15802), .b(wishbone_slave_unit_pci_initiator_if_write_req_int), .o(g74628_p) );
in01f04 g74628_u1 ( .a(g74628_p), .o(n_15980) );
in01f40 g74632_u0 ( .a(wishbone_slave_unit_pci_initiator_if_posted_write_req), .o(n_1238) );
in01s03 g74633_u0 ( .a(FE_OCPN1839_n_1238), .o(n_1041) );
in01f06 g74634_u0 ( .a(n_15981), .o(n_15988) );
in01f01 g74640_u0 ( .a(n_16290), .o(n_15994) );
na02f10 g74642_u0 ( .a(n_15996), .b(parchk_pci_cbe_reg_in_1236), .o(n_16326) );
in01f10 g74643_u0 ( .a(parchk_pci_cbe_reg_in_1237), .o(n_15996) );
no02f10 g74644_u0 ( .a(n_15744), .b(n_15924), .o(g74644_p) );
in01f10 g74644_u1 ( .a(g74644_p), .o(n_15999) );
no02f08 g74645_u0 ( .a(n_1291), .b(n_16289), .o(n_16002) );
in01f10 g74646_u0 ( .a(n_15998), .o(n_16003) );
na02s02 TIMEBOOST_cell_42961 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_69), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_13719) );
na02f10 g74660_u0 ( .a(n_16942), .b(n_16635), .o(g74660_p) );
in01f08 g74660_u1 ( .a(g74660_p), .o(n_16016) );
na02f06 g74661_u0 ( .a(n_16914), .b(n_16021), .o(g74661_p) );
in01f02 g74661_u1 ( .a(g74661_p), .o(n_16022) );
in01f20 g74667_u0 ( .a(conf_w_addr_in_931), .o(n_16027) );
in01f04 g74668_u0 ( .a(n_16351), .o(n_16030) );
na02f20 g74673_u0 ( .a(n_629), .b(n_16284), .o(n_16033) );
in01f02 g74674_u0 ( .a(n_16034), .o(n_16036) );
no02f08 g74686_u0 ( .a(n_16048), .b(pci_target_unit_del_sync_bc_in_202), .o(n_16049) );
na02f10 g74687_u0 ( .a(n_16047), .b(pci_target_unit_del_sync_bc_in_201), .o(n_16048) );
in01f10 g74688_u0 ( .a(pci_target_unit_del_sync_bc_in_203), .o(n_16047) );
na02s01 g74689_u0 ( .a(FE_OFN2214_n_15366), .b(pci_target_unit_del_sync_bc_in_201), .o(g74689_p) );
no02m20 g74690_u0 ( .a(pci_target_unit_del_sync_bc_in_203), .b(pci_target_unit_del_sync_bc_in_202), .o(n_16052) );
na02s02 TIMEBOOST_cell_44854 ( .a(TIMEBOOST_net_14665), .b(g64969_db), .o(n_4372) );
na02f10 g74704_u0 ( .a(n_16066), .b(FE_OCPN1841_n_16089), .o(n_13221) );
in01m06 g74705_u0 ( .a(n_16486), .o(n_16066) );
in01m10 g74709_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_1_), .o(n_16070) );
no02f02 g74733_u0 ( .a(n_16573), .b(n_16577), .o(n_16105) );
no02f02 g74739_u0 ( .a(n_14981), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_), .o(g74739_p) );
in01f02 g74739_u1 ( .a(g74739_p), .o(n_16101) );
na02f04 g74740_u0 ( .a(n_14981), .b(n_16102), .o(n_16103) );
in01s10 g74741_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_), .o(n_16102) );
na02f10 g74749_u0 ( .a(n_16980), .b(n_16157), .o(g74749_p) );
na02s02 TIMEBOOST_cell_45694 ( .a(TIMEBOOST_net_15085), .b(FE_OFN1268_n_4095), .o(TIMEBOOST_net_12520) );
no02f04 g74785_u0 ( .a(n_16152), .b(pci_target_unit_wbm_sm_pciw_fifo_control_in_86), .o(n_16153) );
na02f06 g74786_u0 ( .a(n_16150), .b(n_16151), .o(n_16152) );
na02f08 g74787_u0 ( .a(n_15385), .b(pci_target_unit_wishbone_master_rty_counter_6_), .o(g74787_p) );
in01f04 g74787_u1 ( .a(g74787_p), .o(n_16150) );
no03f40 g74788_u0 ( .a(n_705), .b(wbm_err_i), .c(wbm_ack_i), .o(n_16151) );
na02s02 TIMEBOOST_cell_43338 ( .a(TIMEBOOST_net_13907), .b(g62993_sb), .o(n_5896) );
in01f10 g74793_u0 ( .a(n_1998), .o(n_16159) );
no02f10 g74794_u0 ( .a(pci_target_unit_wishbone_master_c_state_2_), .b(n_819), .o(n_16160) );
oa12f02 g74795_u0 ( .a(n_16160), .b(n_4642), .c(n_2387), .o(n_16162) );
ao12f04 g74796_u0 ( .a(n_16164), .b(n_2702), .c(n_4874), .o(n_16165) );
in01f02 g74797_u0 ( .a(n_16163), .o(n_16164) );
na02f06 g74798_u0 ( .a(n_16738), .b(n_16474), .o(n_16163) );
na03s02 TIMEBOOST_cell_33588 ( .a(TIMEBOOST_net_9555), .b(n_5633), .c(g62095_sb), .o(n_5609) );
in01m01 g74800_u0 ( .a(n_16160), .o(n_16168) );
no02f02 g74802_u0 ( .a(n_16169), .b(n_14419), .o(n_16170) );
na02f02 g74803_u0 ( .a(n_13871), .b(n_14025), .o(n_16169) );
in01f20 g74810_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_1_), .o(n_16175) );
no02f06 g74818_u0 ( .a(n_16326), .b(n_16350), .o(n_16183) );
na03f02 g74828_u0 ( .a(n_16205), .b(n_16970), .c(n_16967), .o(n_16206) );
na02f02 g74838_u0 ( .a(n_16212), .b(n_16209), .o(n_16213) );
no02f02 g74839_u0 ( .a(n_16207), .b(n_16208), .o(n_16209) );
na02s01 TIMEBOOST_cell_32046 ( .a(configuration_pci_err_addr_486), .b(wbm_adr_o_16_), .o(TIMEBOOST_net_9934) );
na02f02 g74841_u0 ( .a(n_14186), .b(n_14185), .o(n_16208) );
no02f02 g74842_u0 ( .a(n_16211), .b(n_16210), .o(n_16212) );
na02f02 TIMEBOOST_cell_36272 ( .a(TIMEBOOST_net_10374), .b(n_2214), .o(TIMEBOOST_net_100) );
na02f02 g74850_u0 ( .a(n_16223), .b(n_16221), .o(n_16224) );
in01f02 g74851_u0 ( .a(n_16220), .o(n_16221) );
in01f02 g74853_u0 ( .a(n_16222), .o(n_16223) );
no02f02 g74856_u0 ( .a(n_16225), .b(n_16226), .o(n_16227) );
na02s02 TIMEBOOST_cell_38102 ( .a(TIMEBOOST_net_11289), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_4625) );
na02f02 g74858_u0 ( .a(n_14211), .b(n_14212), .o(n_16226) );
na02s01 TIMEBOOST_cell_37854 ( .a(TIMEBOOST_net_11165), .b(FE_OFN1689_n_9528), .o(TIMEBOOST_net_4321) );
in01f02 g74859_u1 ( .a(g74859_p), .o(n_16228) );
in01f02 g74860_u0 ( .a(n_16229), .o(n_16230) );
na02m02 TIMEBOOST_cell_32382 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__Q), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_19__Q), .o(TIMEBOOST_net_10102) );
na02f02 TIMEBOOST_cell_40982 ( .a(TIMEBOOST_net_12729), .b(g57233_sb), .o(n_11521) );
no02f02 g74866_u0 ( .a(n_16235), .b(n_16236), .o(n_16237) );
in01f02 g74867_u0 ( .a(n_13868), .o(n_16235) );
in01f02 g74868_u0 ( .a(n_14022), .o(n_16236) );
in01f02 g74869_u0 ( .a(n_16238), .o(n_16239) );
na02m02 TIMEBOOST_cell_32380 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_17__Q), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__Q), .o(TIMEBOOST_net_10101) );
na02f02 TIMEBOOST_cell_40906 ( .a(TIMEBOOST_net_12691), .b(g57396_sb), .o(n_11345) );
in01f02 g74872_u1 ( .a(g74872_p), .o(n_16241) );
no02f03 g74873_u0 ( .a(n_16243), .b(n_16242), .o(n_16244) );
na02s01 TIMEBOOST_cell_30872 ( .a(pci_target_unit_pcit_if_strd_addr_in_704), .b(pci_target_unit_del_sync_addr_in_222), .o(TIMEBOOST_net_9347) );
na02m02 TIMEBOOST_cell_32378 ( .a(wbs_wbb3_2_wbb2_dat_o_i_121), .b(wbs_dat_o_22_), .o(TIMEBOOST_net_10100) );
in01f02 g74879_u1 ( .a(g74879_p), .o(n_16248) );
no02f02 g74880_u0 ( .a(n_16250), .b(n_16249), .o(n_16251) );
na02s01 TIMEBOOST_cell_36360 ( .a(TIMEBOOST_net_10418), .b(FE_OFN2094_n_2520), .o(n_3000) );
na02m02 TIMEBOOST_cell_32450 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__12__Q), .o(TIMEBOOST_net_10136) );
in01f02 g74883_u0 ( .a(n_16252), .o(n_16253) );
na02f02 TIMEBOOST_cell_40908 ( .a(TIMEBOOST_net_12692), .b(g57549_sb), .o(n_11196) );
na04m02 TIMEBOOST_cell_34393 ( .a(n_14671), .b(n_14839), .c(n_3426), .d(g52452_sb), .o(n_14807) );
in01f02 g74886_u1 ( .a(g74886_p), .o(n_16255) );
no02f02 g74887_u0 ( .a(n_16257), .b(n_16256), .o(n_16258) );
na02s01 TIMEBOOST_cell_32044 ( .a(configuration_pci_err_cs_bit_466), .b(pci_target_unit_wishbone_master_bc_register_reg_3__Q), .o(TIMEBOOST_net_9933) );
na02f02 g74889_u0 ( .a(n_14018), .b(n_13865), .o(n_16257) );
in01f02 g74890_u0 ( .a(n_16259), .o(n_16260) );
na02m02 TIMEBOOST_cell_32376 ( .a(wbs_wbb3_2_wbb2_dat_o_i_130), .b(wbs_dat_o_31_), .o(TIMEBOOST_net_10099) );
no02f08 g74892_u0 ( .a(n_16264), .b(n_16262), .o(n_16265) );
na02f20 g74893_u0 ( .a(n_15249), .b(pci_target_unit_wbm_sm_pci_tar_read_request), .o(n_16262) );
no02f40 g74894_u0 ( .a(FE_OCP_RBN2269_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_), .o(n_16264) );
in01m01 g74902_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_), .o(n_16271) );
na02s01 TIMEBOOST_cell_36362 ( .a(TIMEBOOST_net_10419), .b(g66399_sb), .o(n_2524) );
no02f40 g74907_u0 ( .a(pci_target_unit_pcit_if_strd_bc_in), .b(pci_target_unit_pcit_if_strd_bc_in_717), .o(n_16275) );
na02s02 TIMEBOOST_cell_43042 ( .a(TIMEBOOST_net_13759), .b(g58365_sb), .o(n_9210) );
in01f40 g74916_u0 ( .a(conf_w_addr_in_937), .o(n_16284) );
in01f40 g74917_u0 ( .a(conf_w_addr_in_933), .o(n_16285) );
no02f08 g74920_u0 ( .a(n_16003), .b(n_15924), .o(g74920_p) );
in01f06 g74920_u1 ( .a(g74920_p), .o(n_16290) );
na02f10 g74921_u0 ( .a(n_16690), .b(conf_w_addr_in_938), .o(n_16291) );
na02f08 g74929_u0 ( .a(n_16293), .b(n_168), .o(n_13363) );
no02f02 g74930_u0 ( .a(n_14837), .b(n_12858), .o(g74930_p) );
in01f02 g74930_u1 ( .a(g74930_p), .o(n_16293) );
in01f08 g74932_u0 ( .a(n_16300), .o(n_16301) );
in01f06 g74933_u0 ( .a(n_16299), .o(n_16300) );
in01f01 g74935_u0 ( .a(n_16300), .o(n_16305) );
in01f08 g74936_u0 ( .a(n_13363), .o(n_16306) );
oa12f06 g74939_u0 ( .a(n_16354), .b(n_15958), .c(n_15960), .o(n_16309) );
na02s01 TIMEBOOST_cell_45572 ( .a(TIMEBOOST_net_15024), .b(TIMEBOOST_net_3385), .o(TIMEBOOST_net_4797) );
no02m01 g74961_u0 ( .a(n_2440), .b(FE_OFN996_n_15366), .o(g74961_p) );
in01m02 g74961_u1 ( .a(g74961_p), .o(n_16330) );
in01f01 g74962_u0 ( .a(n_16325), .o(n_16332) );
na02f02 g74963_u0 ( .a(FE_OFN1751_n_12086), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__Q), .o(n_16338) );
na02f02 g74965_u0 ( .a(n_16334), .b(n_16364), .o(n_11767) );
na02f02 g74967_u0 ( .a(n_16550), .b(n_16368), .o(g74967_p) );
in01f02 g74967_u1 ( .a(g74967_p), .o(n_16334) );
na02f06 g74981_u0 ( .a(n_16351), .b(conf_w_addr_in), .o(g74981_p) );
in01f02 g74981_u1 ( .a(g74981_p), .o(n_16352) );
in01f40 g74983_u0 ( .a(parchk_pci_cbe_reg_in), .o(n_16350) );
in01f40 g74984_u0 ( .a(n_16354), .o(n_2071) );
in01f40 g74985_u0 ( .a(n_16350), .o(n_16354) );
na02f06 g74989_u0 ( .a(n_16474), .b(pci_target_unit_wbm_sm_pci_tar_burst_ok), .o(n_16358) );
no02f06 g74995_u0 ( .a(n_16076), .b(n_16444), .o(n_16364) );
na02f04 g74996_u0 ( .a(n_16368), .b(n_16554), .o(g74996_p) );
in01f04 g75021_u0 ( .a(n_16183), .o(n_16389) );
in01f20 g75022_u0 ( .a(conf_w_addr_in), .o(n_16390) );
na02s01 TIMEBOOST_cell_17276 ( .a(n_3792), .b(FE_OFN651_n_4508), .o(TIMEBOOST_net_3895) );
in01f08 g75024_u0 ( .a(conf_w_addr_in), .o(g75024_sb) );
na02s02 TIMEBOOST_cell_43491 ( .a(n_4428), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__Q), .o(TIMEBOOST_net_13984) );
na03s02 TIMEBOOST_cell_42985 ( .a(g64221_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__Q), .c(FE_OFN882_g64577_p), .o(TIMEBOOST_net_13731) );
na02f02 TIMEBOOST_cell_45780 ( .a(TIMEBOOST_net_15128), .b(TIMEBOOST_net_5445), .o(n_14828) );
no02f02 g75025_u0 ( .a(n_16400), .b(n_16398), .o(n_16401) );
in01f02 g75027_u0 ( .a(n_12600), .o(n_16395) );
no02f02 g75028_u0 ( .a(n_16396), .b(n_12597), .o(n_16397) );
in01f02 g75029_u0 ( .a(n_11887), .o(n_16396) );
in01f02 g75030_u0 ( .a(n_16399), .o(n_16400) );
no02f02 g75031_u0 ( .a(n_12599), .b(n_12598), .o(n_16399) );
na02f02 TIMEBOOST_cell_42140 ( .a(TIMEBOOST_net_13308), .b(g57285_sb), .o(TIMEBOOST_net_11634) );
in01f02 g75034_u0 ( .a(n_12754), .o(n_16402) );
in01f02 g75036_u0 ( .a(n_12752), .o(n_16404) );
no02f02 g75038_u0 ( .a(n_16408), .b(n_16412), .o(n_16413) );
na02f02 g75039_u0 ( .a(n_12465), .b(n_12383), .o(n_16408) );
na03f02 g75040_u0 ( .a(n_16411), .b(n_16410), .c(n_16409), .o(n_16412) );
no02f02 g75041_u0 ( .a(n_12507), .b(n_12685), .o(n_16409) );
in01f02 g75042_u0 ( .a(n_12686), .o(n_16410) );
na02f01 g75054_u0 ( .a(n_16427), .b(n_16428), .o(n_16429) );
in01f02 g75056_u0 ( .a(n_16425), .o(n_16427) );
no02f10 g75058_u0 ( .a(n_16538), .b(n_16289), .o(n_16424) );
na02m20 g75059_u0 ( .a(pciu_bar1_in_383), .b(pciu_am1_in_521), .o(g75059_p) );
in01f08 g75059_u1 ( .a(g75059_p), .o(n_16428) );
na02f40 g75061_u0 ( .a(FE_OCP_RBN2269_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_), .o(g75061_p) );
na02f01 g75066_u0 ( .a(n_16437), .b(n_16438), .o(n_16439) );
no02f02 g75067_u0 ( .a(n_16435), .b(n_16436), .o(g75067_p) );
in01f02 g75067_u1 ( .a(g75067_p), .o(n_16437) );
na02f08 g75069_u0 ( .a(n_7398), .b(n_6943), .o(n_16436) );
no02f04 g75071_u0 ( .a(n_16444), .b(n_16441), .o(n_16445) );
in01f02 g75072_u0 ( .a(n_16523), .o(g75072_sb) );
na02s01 TIMEBOOST_cell_37201 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__Q), .b(FE_OFN600_n_9687), .o(TIMEBOOST_net_10839) );
na02f02 g75072_u2 ( .a(n_16523), .b(n_16071), .o(g75072_db) );
na02s01 TIMEBOOST_cell_37210 ( .a(TIMEBOOST_net_10843), .b(n_14070), .o(TIMEBOOST_net_614) );
na02f06 g75073_u0 ( .a(n_16564), .b(n_16442), .o(n_16444) );
na02f02 TIMEBOOST_cell_32593 ( .a(FE_OFN1553_n_12104), .b(TIMEBOOST_net_10207), .o(TIMEBOOST_net_6499) );
na02s01 TIMEBOOST_cell_37786 ( .a(TIMEBOOST_net_11131), .b(g61912_sb), .o(TIMEBOOST_net_9784) );
in01f02 g75081_u1 ( .a(g75081_p), .o(n_16459) );
no04f06 TIMEBOOST_cell_34394 ( .a(n_7216), .b(wishbone_slave_unit_wbs_sm_wbr_control_in_190), .c(n_16455), .d(n_16456), .o(g75081_p) );
no02f04 g75083_u0 ( .a(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .b(n_1779), .o(n_16451) );
na02f02 g75084_u0 ( .a(n_15014), .b(n_16021), .o(g75084_p) );
in01f04 g75084_u1 ( .a(g75084_p), .o(n_16452) );
no02f20 g75086_u0 ( .a(n_943), .b(wishbone_slave_unit_wishbone_slave_c_state_2), .o(n_14526) );
na02s02 TIMEBOOST_cell_36826 ( .a(TIMEBOOST_net_10651), .b(g54172_sb), .o(TIMEBOOST_net_9875) );
na02f02 g75088_u0 ( .a(n_7398), .b(n_6989), .o(g75088_p) );
in01f02 g75088_u1 ( .a(g75088_p), .o(n_16456) );
na02m02 TIMEBOOST_cell_36828 ( .a(TIMEBOOST_net_10652), .b(g54169_sb), .o(TIMEBOOST_net_9874) );
in01f10 g75090_u0 ( .a(n_14526), .o(n_16460) );
na02f08 g75114_u0 ( .a(n_16485), .b(n_16486), .o(n_16487) );
no02f06 g75115_u0 ( .a(n_15985), .b(n_15979), .o(n_16485) );
na02m02 TIMEBOOST_cell_32592 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q), .o(TIMEBOOST_net_10207) );
na02f10 g75117_u0 ( .a(n_1434), .b(n_1231), .o(n_16089) );
na02f10 g75119_u0 ( .a(n_16495), .b(n_16496), .o(n_16497) );
ao12f08 g75121_u0 ( .a(n_1539), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_2_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_), .o(n_16490) );
ao12m06 g75122_u0 ( .a(n_16491), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_0_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_), .o(n_16492) );
no02f10 g75123_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_2_), .o(n_16491) );
ao12f08 g75124_u0 ( .a(n_16493), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_1_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_), .o(n_16494) );
no02f10 g75125_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_0_), .o(n_16493) );
na02f10 g75126_u0 ( .a(n_2597), .b(n_565), .o(g75126_p) );
in01f08 g75126_u1 ( .a(g75126_p), .o(n_16496) );
in01f02 g75131_u0 ( .a(n_16503), .o(n_16504) );
no02s01 TIMEBOOST_cell_41699 ( .a(n_382), .b(wbs_adr_i_5_), .o(TIMEBOOST_net_13088) );
na02f06 g75138_u0 ( .a(n_16280), .b(pciu_cache_lsize_not_zero_in), .o(n_16507) );
in01s01 g75140_u0 ( .a(n_16507), .o(n_16512) );
in01f20 g75146_u0 ( .a(pci_target_unit_wishbone_master_retried), .o(n_16516) );
na02f08 g75147_u0 ( .a(n_16521), .b(FE_OCPN1823_n_16560), .o(n_16523) );
na02f06 g75148_u0 ( .a(n_16520), .b(n_16524), .o(n_16521) );
na02f08 g75151_u0 ( .a(FE_OCP_RBN2223_n_15347), .b(n_15638), .o(n_16524) );
no02f04 g75159_u0 ( .a(n_16533), .b(n_16534), .o(n_16535) );
in01f02 g75160_u0 ( .a(n_14981), .o(g75160_sb) );
na04m02 TIMEBOOST_cell_34803 ( .a(g52404_db), .b(g52404_sb), .c(n_3472), .d(TIMEBOOST_net_596), .o(n_14815) );
na02f04 g75160_u2 ( .a(n_14981), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_), .o(g75160_db) );
na03s02 TIMEBOOST_cell_34798 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .b(g63197_sb), .c(g63197_db), .o(n_5770) );
in01f02 g75162_u0 ( .a(n_14981), .o(g75162_sb) );
na02s01 TIMEBOOST_cell_45125 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__Q), .b(n_3986), .o(TIMEBOOST_net_14801) );
na02f04 g75162_u2 ( .a(n_14981), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_0_), .o(g75162_db) );
na02s01 TIMEBOOST_cell_40372 ( .a(TIMEBOOST_net_12424), .b(FE_OFN2079_n_8069), .o(TIMEBOOST_net_11063) );
in01f02 g75163_u0 ( .a(n_16534), .o(n_16536) );
in01f06 g75164_u0 ( .a(n_16533), .o(n_16537) );
na02f08 g75165_u0 ( .a(n_16541), .b(n_16542), .o(g75165_p) );
in01f08 g75165_u1 ( .a(g75165_p), .o(n_16543) );
in01f06 g75166_u0 ( .a(n_16540), .o(n_16541) );
in01f06 g75168_u0 ( .a(FE_OCPN1852_n_16538), .o(n_16539) );
na02f40 g75169_u0 ( .a(n_16695), .b(conf_w_addr_in_938), .o(n_16538) );
no02f04 g75170_u0 ( .a(n_16290), .b(n_15744), .o(n_16542) );
na02f01 g75171_u0 ( .a(n_763), .b(n_1519), .o(n_16544) );
na02f02 g75173_u0 ( .a(FE_OCP_RBN2226_g75174_p), .b(n_16552), .o(n_16553) );
na02f04 g75174_u0 ( .a(n_16444), .b(n_16441), .o(g75174_p) );
na02m02 TIMEBOOST_cell_21980 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__Q), .o(TIMEBOOST_net_6247) );
na02s02 TIMEBOOST_cell_37972 ( .a(TIMEBOOST_net_11224), .b(FE_OFN712_n_8140), .o(TIMEBOOST_net_4290) );
na02s02 TIMEBOOST_cell_19295 ( .a(TIMEBOOST_net_4904), .b(g60605_sb), .o(n_4849) );
na02f02 TIMEBOOST_cell_32563 ( .a(n_12313), .b(TIMEBOOST_net_10192), .o(TIMEBOOST_net_6566) );
na02f03 g75178_u2 ( .a(n_16273), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_), .o(g75178_db) );
no03f02 TIMEBOOST_cell_14209 ( .a(TIMEBOOST_net_2025), .b(FE_RN_584_0), .c(FE_OFN1710_n_4868), .o(TIMEBOOST_net_2890) );
na02f02 g75181_u1 ( .a(FE_OCP_RBN2233_n_16273), .b(n_16271), .o(g75181_da) );
na02f02 g75181_u2 ( .a(n_16273), .b(n_160), .o(g75181_db) );
na02f04 g75181_u3 ( .a(g75181_db), .b(g75181_da), .o(n_16554) );
na02s02 TIMEBOOST_cell_45209 ( .a(n_4332), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__Q), .o(TIMEBOOST_net_14843) );
na02f04 g75194_u0 ( .a(n_16579), .b(n_16566), .o(n_16572) );
no02f08 g75195_u0 ( .a(n_16536), .b(n_16537), .o(n_16566) );
na02f02 g75200_u0 ( .a(n_16573), .b(n_16578), .o(g75200_p) );
in01f02 g75200_u1 ( .a(g75200_p), .o(n_16579) );
na02f08 g75201_u0 ( .a(n_16103), .b(n_16101), .o(n_16573) );
na02f08 g75205_u0 ( .a(n_16487), .b(n_16089), .o(n_14981) );
in01f08 g75221_u0 ( .a(n_9256), .o(n_16637) );
in01f01 g75235_u0 ( .a(n_16690), .o(n_16685) );
in01f10 g75244_u0 ( .a(n_16695), .o(n_16690) );
in01f06 g75246_u0 ( .a(n_16695), .o(n_16696) );
in01f80 g75247_u0 ( .a(conf_w_addr_in_935), .o(n_16695) );
in01f02 g75259_u0 ( .a(n_8940), .o(n_16698) );
in01f04 g75272_u0 ( .a(FE_OCP_RBN2003_FE_OFN1026_n_16760), .o(n_16738) );
in01f03 g75277_u0 ( .a(n_16738), .o(n_16748) );
in01f02 g75295_u0 ( .a(n_9170), .o(n_16779) );
in01s01 g75316_u0 ( .a(n_16818), .o(n_16816) );
na02f10 g75332_u0 ( .a(n_16952), .b(n_16635), .o(g75332_p) );
in01f08 g75332_u1 ( .a(g75332_p), .o(n_16854) );
in01f02 g75337_u0 ( .a(n_16864), .o(n_16860) );
in01f20 g75341_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_cur_state_3_), .o(n_16864) );
in01f03 g75343_u0 ( .a(n_16871), .o(n_16867) );
in01f20 g75350_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_cur_state_2_), .o(n_16871) );
in01s01 g75351_u0 ( .a(n_16980), .o(n_16876) );
in01f03 g75362_u0 ( .a(n_16888), .o(n_16891) );
in01f08 g75365_u0 ( .a(n_16906), .o(n_16904) );
in01f40 g75367_u0 ( .a(pci_target_unit_wishbone_master_c_state_1_), .o(n_16906) );
in01s03 g75368_u0 ( .a(n_16910), .o(wbs_rty_o) );
in01f40 g75371_u0 ( .a(wbs_rty_o_1308), .o(n_16910) );
in01s01 g75372_u0 ( .a(n_16914), .o(n_16911) );
in01f08 g75386_u0 ( .a(n_16940), .o(n_16936) );
in01s02 g75393_u0 ( .a(FE_OCPN1832_n_16949), .o(n_16945) );
in01f06 g75399_u0 ( .a(n_16942), .o(n_16949) );
in01f20 g75400_u0 ( .a(n_16952), .o(n_16942) );
in01f40 g75401_u0 ( .a(wbu_we_in), .o(n_16952) );
na02f04 g75413_u2 ( .a(n_16981), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q), .o(g75413_db) );
na02f06 g75416_u1 ( .a(FE_OCP_RBN1956_n_16981), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(g75416_da) );
na02f04 g75416_u2 ( .a(n_16981), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__Q), .o(g75416_db) );
na02f08 g75416_u3 ( .a(g75416_db), .b(g75416_da), .o(n_16970) );
na02f06 g75418_u1 ( .a(FE_OCP_RBN1956_n_16981), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q), .o(g75418_da) );
na02f04 g75418_u2 ( .a(n_16981), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q), .o(g75418_db) );
na02f08 g75420_u0 ( .a(n_16131), .b(n_16980), .o(n_16981) );
na02f02 TIMEBOOST_cell_41090 ( .a(TIMEBOOST_net_12783), .b(g57068_sb), .o(n_11674) );
no02f04 g75423_u0 ( .a(n_3421), .b(n_15117), .o(n_16977) );
na02f02 g75_u0 ( .a(n_8867), .b(n_16579), .o(g75_p) );
in01f02 g75_u1 ( .a(g75_p), .o(n_15558) );
in01s01 g78_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__291), .o(n_15567) );
in01s01 g79_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_6__252), .o(n_15569) );
na02f20 g7_u0 ( .a(n_16635), .b(n_16818), .o(n_15371) );
no02f40 g9_u0 ( .a(n_16963), .b(FE_OCP_RBN1918_wbs_cti_i_1_), .o(n_16964) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg_u0 ( .ck(ispd_clk), .d(n_10441), .o(wbs_ack_o_1307) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_0__u0 ( .ck(ispd_clk), .d(n_4106), .o(wbu_addr_in) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_10__u0 ( .ck(ispd_clk), .d(n_11876), .o(wbu_addr_in_259) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_11__u0 ( .ck(ispd_clk), .d(n_11878), .o(wbu_addr_in_260) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_12__u0 ( .ck(ispd_clk), .d(n_11875), .o(wbu_addr_in_261) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_13__u0 ( .ck(ispd_clk), .d(n_11874), .o(wbu_addr_in_262) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_14__u0 ( .ck(ispd_clk), .d(n_11872), .o(wbu_addr_in_263) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_15__u0 ( .ck(ispd_clk), .d(n_11873), .o(wbu_addr_in_264) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_16__u0 ( .ck(ispd_clk), .d(n_11871), .o(wbu_addr_in_265) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_17__u0 ( .ck(ispd_clk), .d(n_11870), .o(wbu_addr_in_266) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_18__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15177), .o(wbu_addr_in_267) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_19__u0 ( .ck(ispd_clk), .d(n_11868), .o(wbu_addr_in_268) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_1__u0 ( .ck(ispd_clk), .d(n_4105), .o(wbu_addr_in_250) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_20__u0 ( .ck(ispd_clk), .d(n_11867), .o(wbu_addr_in_269) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_21__u0 ( .ck(ispd_clk), .d(n_11866), .o(wbu_addr_in_270) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_22__u0 ( .ck(ispd_clk), .d(n_11865), .o(wbu_addr_in_271) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_23__u0 ( .ck(ispd_clk), .d(n_11864), .o(wbu_addr_in_272) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_24__u0 ( .ck(ispd_clk), .d(n_11863), .o(wbu_addr_in_273) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_25__u0 ( .ck(ispd_clk), .d(n_11862), .o(wbu_addr_in_274) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_26__u0 ( .ck(ispd_clk), .d(n_11861), .o(wbu_addr_in_275) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_27__u0 ( .ck(ispd_clk), .d(n_11860), .o(wbu_addr_in_276) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_28__u0 ( .ck(ispd_clk), .d(n_11859), .o(wbu_addr_in_277) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_29__u0 ( .ck(ispd_clk), .d(n_11856), .o(i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_29__Q) );
in01s10 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_29__u1 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_29__Q), .o(wbu_addr_in_278) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_2__u0 ( .ck(ispd_clk), .d(n_11858), .o(wbu_addr_in_251) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_30__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15179), .o(wbu_addr_in_279) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_31__u0 ( .ck(ispd_clk), .d(n_11855), .o(i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_31__Q) );
in01m20 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_31__u1 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_31__Q), .o(wbu_addr_in_280) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_3__u0 ( .ck(ispd_clk), .d(n_11854), .o(wbu_addr_in_252) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_4__u0 ( .ck(ispd_clk), .d(n_11853), .o(wbu_addr_in_253) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_5__u0 ( .ck(ispd_clk), .d(n_11852), .o(wbu_addr_in_254) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_6__u0 ( .ck(ispd_clk), .d(n_11851), .o(wbu_addr_in_255) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_7__u0 ( .ck(ispd_clk), .d(n_11850), .o(wbu_addr_in_256) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_8__u0 ( .ck(ispd_clk), .d(n_11848), .o(wbu_addr_in_257) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_9__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15181), .o(wbu_addr_in_258) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg_u0 ( .ck(ispd_clk), .d(n_5723), .o(n_16818) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg_u0 ( .ck(ispd_clk), .d(n_12169), .o(n_16635) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__u0 ( .ck(ispd_clk), .d(n_7147), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__u0 ( .ck(ispd_clk), .d(n_7145), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__u0 ( .ck(ispd_clk), .d(n_7193), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__u0 ( .ck(ispd_clk), .d(n_7191), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__u0 ( .ck(ispd_clk), .d(n_7189), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__u0 ( .ck(ispd_clk), .d(n_7143), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__u0 ( .ck(ispd_clk), .d(n_7151), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__u0 ( .ck(ispd_clk), .d(n_7177), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__u0 ( .ck(ispd_clk), .d(n_7187), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__u0 ( .ck(ispd_clk), .d(n_7149), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__u0 ( .ck(ispd_clk), .d(n_7157), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__u0 ( .ck(ispd_clk), .d(n_7197), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__u0 ( .ck(ispd_clk), .d(n_7141), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__u0 ( .ck(ispd_clk), .d(n_7185), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__u0 ( .ck(ispd_clk), .d(n_7139), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__u0 ( .ck(ispd_clk), .d(n_7195), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__u0 ( .ck(ispd_clk), .d(n_7182), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__u0 ( .ck(ispd_clk), .d(n_7203), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__u0 ( .ck(ispd_clk), .d(n_7205), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__u0 ( .ck(ispd_clk), .d(n_7180), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__u0 ( .ck(ispd_clk), .d(n_7207), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15183), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__u0 ( .ck(ispd_clk), .d(n_7171), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__u0 ( .ck(ispd_clk), .d(n_7168), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__u0 ( .ck(ispd_clk), .d(n_7165), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__u0 ( .ck(ispd_clk), .d(n_7163), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__u0 ( .ck(ispd_clk), .d(n_7161), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__u0 ( .ck(ispd_clk), .d(n_7159), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__u0 ( .ck(ispd_clk), .d(n_7209), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__u0 ( .ck(ispd_clk), .d(n_7155), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__u0 ( .ck(ispd_clk), .d(n_7200), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__u0 ( .ck(ispd_clk), .d(n_7153), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg_u0 ( .ck(ispd_clk), .d(n_11844), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_0__u0 ( .ck(ispd_clk), .d(n_13727), .o(wbs_dat_o_0_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_10__u0 ( .ck(ispd_clk), .d(n_13823), .o(wbs_dat_o_10_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_11__u0 ( .ck(ispd_clk), .d(n_13822), .o(wbs_dat_o_11_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_12__u0 ( .ck(ispd_clk), .d(n_13724), .o(wbs_dat_o_12_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_13__u0 ( .ck(ispd_clk), .d(n_13719), .o(wbs_dat_o_13_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_14__u0 ( .ck(ispd_clk), .d(n_13717), .o(wbs_dat_o_14_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_15__u0 ( .ck(ispd_clk), .d(n_13744), .o(wbs_dat_o_15_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_16__u0 ( .ck(ispd_clk), .d(n_13816), .o(wbs_dat_o_16_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_17__u0 ( .ck(ispd_clk), .d(n_13712), .o(wbs_dat_o_17_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_18__u0 ( .ck(ispd_clk), .d(n_13815), .o(wbs_dat_o_18_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_19__u0 ( .ck(ispd_clk), .d(n_13812), .o(wbs_dat_o_19_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_1__u0 ( .ck(ispd_clk), .d(n_13809), .o(wbs_dat_o_1_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_20__u0 ( .ck(ispd_clk), .d(n_13709), .o(wbs_dat_o_20_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_21__u0 ( .ck(ispd_clk), .d(n_13806), .o(wbs_dat_o_21_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_22__u0 ( .ck(ispd_clk), .d(n_13798), .o(wbs_dat_o_22_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_23__u0 ( .ck(ispd_clk), .d(n_13705), .o(wbs_dat_o_23_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_24__u0 ( .ck(ispd_clk), .d(n_13740), .o(wbs_dat_o_24_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_25__u0 ( .ck(ispd_clk), .d(n_13738), .o(wbs_dat_o_25_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_26__u0 ( .ck(ispd_clk), .d(n_13698), .o(wbs_dat_o_26_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_27__u0 ( .ck(ispd_clk), .d(n_13735), .o(wbs_dat_o_27_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_28__u0 ( .ck(ispd_clk), .d(n_13697), .o(wbs_dat_o_28_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_29__u0 ( .ck(ispd_clk), .d(n_13696), .o(wbs_dat_o_29_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_2__u0 ( .ck(ispd_clk), .d(n_13734), .o(wbs_dat_o_2_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_30__u0 ( .ck(ispd_clk), .d(n_13794), .o(wbs_dat_o_30_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_31__u0 ( .ck(ispd_clk), .d(n_13694), .o(wbs_dat_o_31_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_3__u0 ( .ck(ispd_clk), .d(n_13693), .o(wbs_dat_o_3_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_4__u0 ( .ck(ispd_clk), .d(n_13688), .o(wbs_dat_o_4_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_5__u0 ( .ck(ispd_clk), .d(n_13793), .o(wbs_dat_o_5_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_6__u0 ( .ck(ispd_clk), .d(n_13792), .o(wbs_dat_o_6_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_7__u0 ( .ck(ispd_clk), .d(n_13687), .o(wbs_dat_o_7_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_8__u0 ( .ck(ispd_clk), .d(n_13686), .o(wbs_dat_o_8_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_9__u0 ( .ck(ispd_clk), .d(n_13685), .o(wbs_dat_o_9_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg_u0 ( .ck(ispd_clk), .d(n_8874), .o(wbs_err_o_1309) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg_u0 ( .ck(ispd_clk), .d(n_8583), .o(wbs_rty_o_1308) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg_0__u0 ( .ck(ispd_clk), .d(n_4104), .o(wbu_sel_in) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg_1__u0 ( .ck(ispd_clk), .d(n_4103), .o(wbu_sel_in_312) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg_2__u0 ( .ck(ispd_clk), .d(n_4102), .o(wbu_sel_in_313) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg_3__u0 ( .ck(ispd_clk), .d(n_4101), .o(wbu_sel_in_314) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg_u0 ( .ck(ispd_clk), .d(n_4100), .o(wbu_we_in) );
ms00f80 input_register_pci_ad_reg_out_reg_0__u0 ( .ck(ispd_clk), .d(n_1654), .o(parchk_pci_ad_reg_in) );
ms00f80 input_register_pci_ad_reg_out_reg_10__u0 ( .ck(ispd_clk), .d(n_1497), .o(parchk_pci_ad_reg_in_1214) );
ms00f80 input_register_pci_ad_reg_out_reg_11__u0 ( .ck(ispd_clk), .d(n_1429), .o(parchk_pci_ad_reg_in_1215) );
ms00f80 input_register_pci_ad_reg_out_reg_12__u0 ( .ck(ispd_clk), .d(n_1647), .o(parchk_pci_ad_reg_in_1216) );
ms00f80 input_register_pci_ad_reg_out_reg_13__u0 ( .ck(ispd_clk), .d(n_1685), .o(parchk_pci_ad_reg_in_1217) );
ms00f80 input_register_pci_ad_reg_out_reg_14__u0 ( .ck(ispd_clk), .d(n_1502), .o(parchk_pci_ad_reg_in_1218) );
ms00f80 input_register_pci_ad_reg_out_reg_15__u0 ( .ck(ispd_clk), .d(n_1634), .o(parchk_pci_ad_reg_in_1219) );
ms00f80 input_register_pci_ad_reg_out_reg_16__u0 ( .ck(ispd_clk), .d(n_1499), .o(parchk_pci_ad_reg_in_1220) );
ms00f80 input_register_pci_ad_reg_out_reg_17__u0 ( .ck(ispd_clk), .d(n_1652), .o(parchk_pci_ad_reg_in_1221) );
ms00f80 input_register_pci_ad_reg_out_reg_18__u0 ( .ck(ispd_clk), .d(n_1428), .o(parchk_pci_ad_reg_in_1222) );
ms00f80 input_register_pci_ad_reg_out_reg_19__u0 ( .ck(ispd_clk), .d(n_1274), .o(parchk_pci_ad_reg_in_1223) );
ms00f80 input_register_pci_ad_reg_out_reg_1__u0 ( .ck(ispd_clk), .d(n_1272), .o(parchk_pci_ad_reg_in_1205) );
ms00f80 input_register_pci_ad_reg_out_reg_20__u0 ( .ck(ispd_clk), .d(n_1495), .o(parchk_pci_ad_reg_in_1224) );
ms00f80 input_register_pci_ad_reg_out_reg_21__u0 ( .ck(ispd_clk), .d(n_1431), .o(parchk_pci_ad_reg_in_1225) );
ms00f80 input_register_pci_ad_reg_out_reg_22__u0 ( .ck(ispd_clk), .d(n_1474), .o(parchk_pci_ad_reg_in_1226) );
ms00f80 input_register_pci_ad_reg_out_reg_23__u0 ( .ck(ispd_clk), .d(n_1681), .o(parchk_pci_ad_reg_in_1227) );
ms00f80 input_register_pci_ad_reg_out_reg_24__u0 ( .ck(ispd_clk), .d(n_1503), .o(parchk_pci_ad_reg_in_1228) );
ms00f80 input_register_pci_ad_reg_out_reg_25__u0 ( .ck(ispd_clk), .d(n_1704), .o(parchk_pci_ad_reg_in_1229) );
ms00f80 input_register_pci_ad_reg_out_reg_26__u0 ( .ck(ispd_clk), .d(n_1444), .o(parchk_pci_ad_reg_in_1230) );
ms00f80 input_register_pci_ad_reg_out_reg_27__u0 ( .ck(ispd_clk), .d(n_1483), .o(parchk_pci_ad_reg_in_1231) );
ms00f80 input_register_pci_ad_reg_out_reg_28__u0 ( .ck(ispd_clk), .d(n_1501), .o(parchk_pci_ad_reg_in_1232) );
ms00f80 input_register_pci_ad_reg_out_reg_29__u0 ( .ck(ispd_clk), .d(n_1677), .o(parchk_pci_ad_reg_in_1233) );
ms00f80 input_register_pci_ad_reg_out_reg_2__u0 ( .ck(ispd_clk), .d(n_1277), .o(parchk_pci_ad_reg_in_1206) );
ms00f80 input_register_pci_ad_reg_out_reg_30__u0 ( .ck(ispd_clk), .d(n_1640), .o(n_2509) );
ms00f80 input_register_pci_ad_reg_out_reg_31__u0 ( .ck(ispd_clk), .d(n_1470), .o(parchk_pci_ad_reg_in_1235) );
ms00f80 input_register_pci_ad_reg_out_reg_3__u0 ( .ck(ispd_clk), .d(n_1649), .o(parchk_pci_ad_reg_in_1207) );
ms00f80 input_register_pci_ad_reg_out_reg_4__u0 ( .ck(ispd_clk), .d(n_1683), .o(parchk_pci_ad_reg_in_1208) );
ms00f80 input_register_pci_ad_reg_out_reg_5__u0 ( .ck(ispd_clk), .d(n_1411), .o(parchk_pci_ad_reg_in_1209) );
ms00f80 input_register_pci_ad_reg_out_reg_6__u0 ( .ck(ispd_clk), .d(n_1276), .o(parchk_pci_ad_reg_in_1210) );
ms00f80 input_register_pci_ad_reg_out_reg_7__u0 ( .ck(ispd_clk), .d(n_1614), .o(parchk_pci_ad_reg_in_1211) );
ms00f80 input_register_pci_ad_reg_out_reg_8__u0 ( .ck(ispd_clk), .d(n_1275), .o(parchk_pci_ad_reg_in_1212) );
ms00f80 input_register_pci_ad_reg_out_reg_9__u0 ( .ck(ispd_clk), .d(n_1641), .o(parchk_pci_ad_reg_in_1213) );
ms00f80 input_register_pci_cbe_reg_out_reg_0__u0 ( .ck(ispd_clk), .d(n_3118), .o(parchk_pci_cbe_reg_in) );
ms00f80 input_register_pci_cbe_reg_out_reg_1__u0 ( .ck(ispd_clk), .d(n_2564), .o(parchk_pci_cbe_reg_in_1236) );
ms00f80 input_register_pci_cbe_reg_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2568), .o(parchk_pci_cbe_reg_in_1237) );
ms00f80 input_register_pci_cbe_reg_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2567), .o(parchk_pci_cbe_reg_in_1238) );
ms00f80 input_register_pci_devsel_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_2374), .o(wbu_pciif_devsel_reg_in) );
ms00f80 input_register_pci_frame_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_2372), .o(parchk_pci_frame_reg_in) );
ms00f80 input_register_pci_idsel_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_1452), .o(pciu_pciif_idsel_reg_in) );
ms00f80 input_register_pci_irdy_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_2471), .o(n_657) );
ms00f80 input_register_pci_stop_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_2147), .o(pciu_pciif_stop_reg_in) );
ms00f80 input_register_pci_trdy_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_2718), .o(parchk_pci_trdy_reg_in) );
ms00f80 output_backup_ad_out_reg_0__u0 ( .ck(ispd_clk), .d(n_13908), .o(parchk_pci_ad_out_in) );
ms00f80 output_backup_ad_out_reg_10__u0 ( .ck(ispd_clk), .d(n_14320), .o(parchk_pci_ad_out_in_1177) );
ms00f80 output_backup_ad_out_reg_11__u0 ( .ck(ispd_clk), .d(n_14316), .o(parchk_pci_ad_out_in_1178) );
ms00f80 output_backup_ad_out_reg_12__u0 ( .ck(ispd_clk), .d(n_14318), .o(parchk_pci_ad_out_in_1179) );
ms00f80 output_backup_ad_out_reg_13__u0 ( .ck(ispd_clk), .d(n_14314), .o(parchk_pci_ad_out_in_1180) );
ms00f80 output_backup_ad_out_reg_14__u0 ( .ck(ispd_clk), .d(n_14312), .o(parchk_pci_ad_out_in_1181) );
ms00f80 output_backup_ad_out_reg_15__u0 ( .ck(ispd_clk), .d(n_14310), .o(parchk_pci_ad_out_in_1182) );
ms00f80 output_backup_ad_out_reg_16__u0 ( .ck(ispd_clk), .d(n_14383), .o(parchk_pci_ad_out_in_1183) );
ms00f80 output_backup_ad_out_reg_17__u0 ( .ck(ispd_clk), .d(n_14382), .o(parchk_pci_ad_out_in_1184) );
ms00f80 output_backup_ad_out_reg_18__u0 ( .ck(ispd_clk), .d(n_14381), .o(parchk_pci_ad_out_in_1185) );
ms00f80 output_backup_ad_out_reg_19__u0 ( .ck(ispd_clk), .d(n_14380), .o(parchk_pci_ad_out_in_1186) );
ms00f80 output_backup_ad_out_reg_1__u0 ( .ck(ispd_clk), .d(n_14094), .o(parchk_pci_ad_out_in_1168) );
ms00f80 output_backup_ad_out_reg_20__u0 ( .ck(ispd_clk), .d(n_14379), .o(parchk_pci_ad_out_in_1187) );
ms00f80 output_backup_ad_out_reg_21__u0 ( .ck(ispd_clk), .d(n_14093), .o(parchk_pci_ad_out_in_1188) );
ms00f80 output_backup_ad_out_reg_22__u0 ( .ck(ispd_clk), .d(n_14378), .o(parchk_pci_ad_out_in_1189) );
ms00f80 output_backup_ad_out_reg_23__u0 ( .ck(ispd_clk), .d(n_14377), .o(parchk_pci_ad_out_in_1190) );
ms00f80 output_backup_ad_out_reg_24__u0 ( .ck(ispd_clk), .d(n_14376), .o(parchk_pci_ad_out_in_1191) );
ms00f80 output_backup_ad_out_reg_25__u0 ( .ck(ispd_clk), .d(n_13831), .o(parchk_pci_ad_out_in_1192) );
ms00f80 output_backup_ad_out_reg_26__u0 ( .ck(ispd_clk), .d(n_14078), .o(parchk_pci_ad_out_in_1193) );
ms00f80 output_backup_ad_out_reg_27__u0 ( .ck(ispd_clk), .d(n_14375), .o(parchk_pci_ad_out_in_1194) );
ms00f80 output_backup_ad_out_reg_28__u0 ( .ck(ispd_clk), .d(n_14374), .o(parchk_pci_ad_out_in_1195) );
ms00f80 output_backup_ad_out_reg_29__u0 ( .ck(ispd_clk), .d(n_14373), .o(parchk_pci_ad_out_in_1196) );
ms00f80 output_backup_ad_out_reg_2__u0 ( .ck(ispd_clk), .d(n_14372), .o(parchk_pci_ad_out_in_1169) );
ms00f80 output_backup_ad_out_reg_30__u0 ( .ck(ispd_clk), .d(n_14088), .o(parchk_pci_ad_out_in_1197) );
ms00f80 output_backup_ad_out_reg_31__u0 ( .ck(ispd_clk), .d(n_14531), .o(parchk_pci_ad_out_in_1198) );
ms00f80 output_backup_ad_out_reg_3__u0 ( .ck(ispd_clk), .d(n_14371), .o(parchk_pci_ad_out_in_1170) );
ms00f80 output_backup_ad_out_reg_4__u0 ( .ck(ispd_clk), .d(n_14370), .o(parchk_pci_ad_out_in_1171) );
ms00f80 output_backup_ad_out_reg_5__u0 ( .ck(ispd_clk), .d(n_14369), .o(parchk_pci_ad_out_in_1172) );
ms00f80 output_backup_ad_out_reg_6__u0 ( .ck(ispd_clk), .d(n_14368), .o(parchk_pci_ad_out_in_1173) );
ms00f80 output_backup_ad_out_reg_7__u0 ( .ck(ispd_clk), .d(n_14367), .o(parchk_pci_ad_out_in_1174) );
ms00f80 output_backup_ad_out_reg_8__u0 ( .ck(ispd_clk), .d(n_14366), .o(parchk_pci_ad_out_in_1175) );
ms00f80 output_backup_ad_out_reg_9__u0 ( .ck(ispd_clk), .d(n_14365), .o(parchk_pci_ad_out_in_1176) );
ms00f80 output_backup_cbe_en_out_reg_u0 ( .ck(ispd_clk), .d(n_7135), .o(parchk_pci_cbe_en_in) );
ms00f80 output_backup_cbe_out_reg_0__u0 ( .ck(ispd_clk), .d(n_14397), .o(parchk_pci_cbe_out_in) );
ms00f80 output_backup_cbe_out_reg_1__u0 ( .ck(ispd_clk), .d(n_8531), .o(parchk_pci_cbe_out_in_1202) );
ms00f80 output_backup_cbe_out_reg_2__u0 ( .ck(ispd_clk), .d(n_14396), .o(parchk_pci_cbe_out_in_1203) );
ms00f80 output_backup_cbe_out_reg_3__u0 ( .ck(ispd_clk), .d(n_14394), .o(parchk_pci_cbe_out_in_1204) );
ms00f80 output_backup_devsel_out_reg_u0 ( .ck(ispd_clk), .d(n_14616), .o(output_backup_devsel_out_reg_Q) );
ms00f80 output_backup_frame_en_out_reg_u0 ( .ck(ispd_clk), .d(n_7210), .o(parchk_pci_frame_en_in) );
ms00f80 output_backup_frame_out_reg_u0 ( .ck(ispd_clk), .d(n_8752), .o(wbu_pciif_frame_out_in) );
ms00f80 output_backup_irdy_en_out_reg_u0 ( .ck(ispd_clk), .d(n_447), .o(parchk_pci_irdy_en_in) );
ms00f80 output_backup_irdy_out_reg_u0 ( .ck(ispd_clk), .d(n_2900), .o(out_bckp_irdy_out) );
ms00f80 output_backup_mas_ad_en_out_reg_u0 ( .ck(ispd_clk), .d(n_11450), .o(n_14905) );
ms00f80 output_backup_par_en_out_reg_u0 ( .ck(ispd_clk), .d(n_12954), .o(output_backup_par_en_out_reg_Q) );
in01s03 output_backup_par_en_out_reg_u1 ( .a(output_backup_par_en_out_reg_Q), .o(parchk_pci_par_en_in) );
ms00f80 output_backup_par_out_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15185), .o(output_backup_par_out_reg_Q) );
ms00f80 output_backup_perr_en_out_reg_u0 ( .ck(ispd_clk), .d(n_14572), .o(out_bckp_perr_en_out) );
ms00f80 output_backup_perr_out_reg_u0 ( .ck(ispd_clk), .d(n_13918), .o(output_backup_perr_out_reg_Q) );
in01s01 output_backup_perr_out_reg_u1 ( .a(output_backup_perr_out_reg_Q), .o(parchk_pci_perr_out_in) );
ms00f80 output_backup_serr_en_out_reg_u0 ( .ck(ispd_clk), .d(n_13757), .o(output_backup_serr_en_out_reg_Q) );
in01s01 output_backup_serr_en_out_reg_u1 ( .a(output_backup_serr_en_out_reg_Q), .o(parchk_pci_serr_en_in) );
ms00f80 output_backup_serr_out_reg_u0 ( .ck(ispd_clk), .d(n_13917), .o(parchk_pci_serr_out_in) );
ms00f80 output_backup_stop_out_reg_u0 ( .ck(ispd_clk), .d(n_14617), .o(output_backup_stop_out_reg_Q) );
in01s10 output_backup_stop_out_reg_u1 ( .a(output_backup_stop_out_reg_Q), .o(pciu_pciif_bckp_stop_in) );
ms00f80 output_backup_tar_ad_en_out_reg_u0 ( .ck(ispd_clk), .d(n_11448), .o(output_backup_tar_ad_en_out_reg_Q) );
in01m40 output_backup_tar_ad_en_out_reg_u1 ( .a(output_backup_tar_ad_en_out_reg_Q), .o(n_13784) );
ms00f80 output_backup_trdy_en_out_reg_u0 ( .ck(ispd_clk), .d(n_8875), .o(parchk_pci_trdy_en_in) );
ms00f80 output_backup_trdy_out_reg_u0 ( .ck(ispd_clk), .d(n_14622), .o(output_backup_trdy_out_reg_Q) );
ms00f80 parity_checker_check_for_serr_on_second_reg_u0 ( .ck(ispd_clk), .d(n_3794), .o(parity_checker_check_for_serr_on_second_reg_Q) );
in01s01 parity_checker_check_for_serr_on_second_reg_u1 ( .a(parity_checker_check_for_serr_on_second_reg_Q), .o(parity_checker_check_for_serr_on_second) );
ms00f80 parity_checker_check_perr_reg_u0 ( .ck(ispd_clk), .d(g54038_sb), .o(parity_checker_check_perr_reg_Q) );
in01s01 parity_checker_check_perr_reg_u1 ( .a(parity_checker_check_perr_reg_Q), .o(parity_checker_check_perr) );
ms00f80 parity_checker_frame_and_irdy_en_prev_prev_reg_u0 ( .ck(ispd_clk), .d(parity_checker_frame_and_irdy_en_prev), .o(parity_checker_frame_and_irdy_en_prev_prev) );
ms00f80 parity_checker_frame_and_irdy_en_prev_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15187), .o(parity_checker_frame_and_irdy_en_prev) );
ms00f80 parity_checker_frame_dec2_reg_u0 ( .ck(ispd_clk), .d(n_15302), .o(parity_checker_frame_dec2) );
ms00f80 parity_checker_master_perr_report_reg_u0 ( .ck(ispd_clk), .d(parity_checker_frame_and_irdy_en_prev_prev), .o(parity_checker_master_perr_report_reg_Q) );
in01s01 parity_checker_master_perr_report_reg_u1 ( .a(parity_checker_master_perr_report_reg_Q), .o(parity_checker_master_perr_report) );
ms00f80 parity_checker_perr_en_crit_gen_perr_en_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_14386), .o(parity_checker_pci_perr_en_reg) );
ms00f80 parity_checker_perr_sampled_reg_u0 ( .ck(ispd_clk), .d(n_14765), .o(parity_checker_perr_sampled) );
ms00f80 pci_io_mux_ad_iob0_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_13911), .o(pci_ad_o_0_) );
ms00f80 pci_io_mux_ad_iob0_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_0_) );
ms00f80 pci_io_mux_ad_iob10_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14364), .o(pci_ad_o_10_) );
ms00f80 pci_io_mux_ad_iob10_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_10_) );
ms00f80 pci_io_mux_ad_iob11_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14363), .o(pci_ad_o_11_) );
ms00f80 pci_io_mux_ad_iob11_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_11_) );
ms00f80 pci_io_mux_ad_iob12_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14362), .o(pci_ad_o_12_) );
ms00f80 pci_io_mux_ad_iob12_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_12_) );
ms00f80 pci_io_mux_ad_iob13_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14361), .o(pci_ad_o_13_) );
ms00f80 pci_io_mux_ad_iob13_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_13_) );
ms00f80 pci_io_mux_ad_iob14_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14360), .o(pci_ad_o_14_) );
ms00f80 pci_io_mux_ad_iob14_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_14_) );
ms00f80 pci_io_mux_ad_iob15_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14359), .o(pci_ad_o_15_) );
ms00f80 pci_io_mux_ad_iob15_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_15_) );
ms00f80 pci_io_mux_ad_iob16_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14358), .o(pci_ad_o_16_) );
ms00f80 pci_io_mux_ad_iob16_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_16_) );
ms00f80 pci_io_mux_ad_iob17_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14356), .o(pci_ad_o_17_) );
ms00f80 pci_io_mux_ad_iob17_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_17_) );
ms00f80 pci_io_mux_ad_iob18_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14354), .o(pci_ad_o_18_) );
ms00f80 pci_io_mux_ad_iob18_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_18_) );
ms00f80 pci_io_mux_ad_iob19_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14352), .o(pci_ad_o_19_) );
ms00f80 pci_io_mux_ad_iob19_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_19_) );
ms00f80 pci_io_mux_ad_iob1_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14086), .o(pci_ad_o_1_) );
ms00f80 pci_io_mux_ad_iob1_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_1_) );
ms00f80 pci_io_mux_ad_iob20_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14350), .o(pci_ad_o_20_) );
ms00f80 pci_io_mux_ad_iob20_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_20_) );
ms00f80 pci_io_mux_ad_iob21_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14084), .o(pci_ad_o_21_) );
ms00f80 pci_io_mux_ad_iob21_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_21_) );
ms00f80 pci_io_mux_ad_iob22_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14348), .o(pci_ad_o_22_) );
ms00f80 pci_io_mux_ad_iob22_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_22_) );
ms00f80 pci_io_mux_ad_iob23_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14342), .o(pci_ad_o_23_) );
ms00f80 pci_io_mux_ad_iob23_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_23_) );
ms00f80 pci_io_mux_ad_iob24_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14346), .o(pci_ad_o_24_) );
ms00f80 pci_io_mux_ad_iob24_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_24_) );
ms00f80 pci_io_mux_ad_iob25_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_13830), .o(pci_ad_o_25_) );
ms00f80 pci_io_mux_ad_iob25_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_25_) );
ms00f80 pci_io_mux_ad_iob26_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14077), .o(pci_ad_o_26_) );
ms00f80 pci_io_mux_ad_iob26_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_26_) );
ms00f80 pci_io_mux_ad_iob27_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14344), .o(pci_ad_o_27_) );
ms00f80 pci_io_mux_ad_iob27_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_27_) );
ms00f80 pci_io_mux_ad_iob28_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14338), .o(pci_ad_o_28_) );
ms00f80 pci_io_mux_ad_iob28_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_28_) );
ms00f80 pci_io_mux_ad_iob29_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14340), .o(pci_ad_o_29_) );
ms00f80 pci_io_mux_ad_iob29_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_29_) );
ms00f80 pci_io_mux_ad_iob2_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14336), .o(pci_ad_o_2_) );
ms00f80 pci_io_mux_ad_iob2_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_2_) );
ms00f80 pci_io_mux_ad_iob30_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14082), .o(pci_ad_o_30_) );
ms00f80 pci_io_mux_ad_iob30_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1506_n_15768), .o(pci_ad_oe_o_30_) );
ms00f80 pci_io_mux_ad_iob31_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14530), .o(pci_ad_o_31_) );
ms00f80 pci_io_mux_ad_iob31_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_31_) );
ms00f80 pci_io_mux_ad_iob3_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14334), .o(pci_ad_o_3_) );
ms00f80 pci_io_mux_ad_iob3_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_3_) );
ms00f80 pci_io_mux_ad_iob4_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14332), .o(pci_ad_o_4_) );
ms00f80 pci_io_mux_ad_iob4_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_4_) );
ms00f80 pci_io_mux_ad_iob5_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14330), .o(pci_ad_o_5_) );
ms00f80 pci_io_mux_ad_iob5_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_5_) );
ms00f80 pci_io_mux_ad_iob6_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14328), .o(pci_ad_o_6_) );
ms00f80 pci_io_mux_ad_iob6_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_6_) );
ms00f80 pci_io_mux_ad_iob7_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14326), .o(pci_ad_o_7_) );
ms00f80 pci_io_mux_ad_iob7_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_7_) );
ms00f80 pci_io_mux_ad_iob8_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14324), .o(pci_ad_o_8_) );
ms00f80 pci_io_mux_ad_iob8_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_8_) );
ms00f80 pci_io_mux_ad_iob9_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14322), .o(pci_ad_o_9_) );
ms00f80 pci_io_mux_ad_iob9_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_9_) );
ms00f80 pci_io_mux_cbe_iob0_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14393), .o(pci_cbe_o_0_) );
ms00f80 pci_io_mux_cbe_iob0_en_out_reg_u0 ( .ck(ispd_clk), .d(n_7400), .o(pci_cbe_oe_o_0_) );
ms00f80 pci_io_mux_cbe_iob1_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_8530), .o(pci_cbe_o_1_) );
ms00f80 pci_io_mux_cbe_iob1_en_out_reg_u0 ( .ck(ispd_clk), .d(n_7400), .o(pci_cbe_oe_o_1_) );
ms00f80 pci_io_mux_cbe_iob2_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14391), .o(pci_cbe_o_2_) );
ms00f80 pci_io_mux_cbe_iob2_en_out_reg_u0 ( .ck(ispd_clk), .d(n_7400), .o(pci_cbe_oe_o_2_) );
ms00f80 pci_io_mux_cbe_iob3_dat_out_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15189), .o(pci_cbe_o_3_) );
ms00f80 pci_io_mux_cbe_iob3_en_out_reg_u0 ( .ck(ispd_clk), .d(n_7400), .o(pci_cbe_oe_o_3_) );
ms00f80 pci_io_mux_devsel_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14616), .o(pci_devsel_o) );
ms00f80 pci_io_mux_devsel_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_8934), .o(pci_devsel_oe_o) );
ms00f80 pci_io_mux_frame_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_8751), .o(pci_frame_o) );
ms00f80 pci_io_mux_frame_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_7211), .o(pci_frame_oe_o) );
ms00f80 pci_io_mux_irdy_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_2900), .o(pci_irdy_o) );
ms00f80 pci_io_mux_irdy_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_333), .o(pci_irdy_oe_o) );
ms00f80 pci_io_mux_par_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15191), .o(pci_par_o) );
ms00f80 pci_io_mux_par_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_12855), .o(pci_par_oe_o) );
ms00f80 pci_io_mux_perr_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_13918), .o(pci_perr_o) );
ms00f80 pci_io_mux_perr_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_14571), .o(pci_perr_oe_o) );
ms00f80 pci_io_mux_req_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_2246), .o(pci_req_o) );
ms00f80 pci_io_mux_req_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_285), .o(pci_req_oe_o) );
ms00f80 pci_io_mux_serr_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_13917), .o(pci_serr_o) );
ms00f80 pci_io_mux_serr_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_13758), .o(pci_serr_oe_o) );
ms00f80 pci_io_mux_stop_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14617), .o(pci_stop_o) );
ms00f80 pci_io_mux_stop_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_8934), .o(pci_stop_oe_o) );
ms00f80 pci_io_mux_trdy_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14622), .o(pci_trdy_o) );
ms00f80 pci_io_mux_trdy_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_8934), .o(pci_trdy_oe_o) );
ms00f80 pci_resets_and_interrupts_inta_en_out_reg_u0 ( .ck(ispd_clk), .d(n_3315), .o(pci_inta_oe_o) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_0__u0 ( .ck(ispd_clk), .d(n_2672), .o(pci_target_unit_pcit_if_strd_addr_in) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_10__u0 ( .ck(ispd_clk), .d(n_2632), .o(pci_target_unit_pcit_if_strd_addr_in_695) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_11__u0 ( .ck(ispd_clk), .d(n_2635), .o(pci_target_unit_pcit_if_strd_addr_in_696) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_12__u0 ( .ck(ispd_clk), .d(n_2660), .o(pci_target_unit_pcit_if_strd_addr_in_697) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_13__u0 ( .ck(ispd_clk), .d(n_2658), .o(pci_target_unit_pcit_if_strd_addr_in_698) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_14__u0 ( .ck(ispd_clk), .d(n_2668), .o(pci_target_unit_pcit_if_strd_addr_in_699) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_15__u0 ( .ck(ispd_clk), .d(n_2673), .o(pci_target_unit_pcit_if_strd_addr_in_700) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_16__u0 ( .ck(ispd_clk), .d(n_2679), .o(pci_target_unit_pcit_if_strd_addr_in_701) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_17__u0 ( .ck(ispd_clk), .d(n_2636), .o(pci_target_unit_pcit_if_strd_addr_in_702) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_18__u0 ( .ck(ispd_clk), .d(n_2634), .o(pci_target_unit_pcit_if_strd_addr_in_703) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_19__u0 ( .ck(ispd_clk), .d(n_2638), .o(pci_target_unit_pcit_if_strd_addr_in_704) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_1__u0 ( .ck(ispd_clk), .d(n_2653), .o(pci_target_unit_pcit_if_strd_addr_in_686) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_20__u0 ( .ck(ispd_clk), .d(n_2646), .o(pci_target_unit_pcit_if_strd_addr_in_705) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_21__u0 ( .ck(ispd_clk), .d(n_2661), .o(pci_target_unit_pcit_if_strd_addr_in_706) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_22__u0 ( .ck(ispd_clk), .d(n_2659), .o(pci_target_unit_pcit_if_strd_addr_in_707) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_23__u0 ( .ck(ispd_clk), .d(n_2664), .o(pci_target_unit_pcit_if_strd_addr_in_708) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_24__u0 ( .ck(ispd_clk), .d(n_2665), .o(pci_target_unit_pcit_if_strd_addr_in_709) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_25__u0 ( .ck(ispd_clk), .d(n_2666), .o(pci_target_unit_pcit_if_strd_addr_in_710) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_26__u0 ( .ck(ispd_clk), .d(n_2669), .o(pci_target_unit_pcit_if_strd_addr_in_711) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_27__u0 ( .ck(ispd_clk), .d(n_2670), .o(pci_target_unit_pcit_if_strd_addr_in_712) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_28__u0 ( .ck(ispd_clk), .d(n_2674), .o(pci_target_unit_pcit_if_strd_addr_in_713) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_29__u0 ( .ck(ispd_clk), .d(n_2637), .o(pci_target_unit_pcit_if_strd_addr_in_714) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2640), .o(pci_target_unit_pcit_if_strd_addr_in_687) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_30__u0 ( .ck(ispd_clk), .d(n_2641), .o(pci_target_unit_pcit_if_strd_addr_in_715) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_31__u0 ( .ck(ispd_clk), .d(n_2656), .o(pci_target_unit_pcit_if_strd_addr_in_716) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2655), .o(pci_target_unit_pcit_if_strd_addr_in_688) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_4__u0 ( .ck(ispd_clk), .d(n_2639), .o(pci_target_unit_pcit_if_strd_addr_in_689) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_5__u0 ( .ck(ispd_clk), .d(n_2633), .o(pci_target_unit_pcit_if_strd_addr_in_690) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_6__u0 ( .ck(ispd_clk), .d(n_2645), .o(pci_target_unit_pcit_if_strd_addr_in_691) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_7__u0 ( .ck(ispd_clk), .d(n_2663), .o(pci_target_unit_pcit_if_strd_addr_in_692) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_8__u0 ( .ck(ispd_clk), .d(n_2667), .o(pci_target_unit_pcit_if_strd_addr_in_693) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_9__u0 ( .ck(ispd_clk), .d(n_2654), .o(pci_target_unit_pcit_if_strd_addr_in_694) );
ms00f80 pci_target_unit_del_sync_bc_out_reg_0__u0 ( .ck(ispd_clk), .d(n_2644), .o(pci_target_unit_pcit_if_strd_bc_in) );
ms00f80 pci_target_unit_del_sync_bc_out_reg_1__u0 ( .ck(ispd_clk), .d(n_2657), .o(pci_target_unit_pcit_if_strd_bc_in_717) );
ms00f80 pci_target_unit_del_sync_bc_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2662), .o(pci_target_unit_pcit_if_strd_bc_in_718) );
ms00f80 pci_target_unit_del_sync_bc_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2677), .o(pci_target_unit_pcit_if_strd_bc_in_719) );
ms00f80 pci_target_unit_del_sync_be_out_reg_0__u0 ( .ck(ispd_clk), .d(n_3031), .o(pci_target_unit_del_sync_be_out_reg_0__Q) );
ms00f80 pci_target_unit_del_sync_be_out_reg_1__u0 ( .ck(ispd_clk), .d(n_2652), .o(pci_target_unit_del_sync_be_out_reg_1__Q) );
ms00f80 pci_target_unit_del_sync_be_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2649), .o(pci_target_unit_del_sync_be_out_reg_2__Q) );
ms00f80 pci_target_unit_del_sync_be_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2643), .o(pci_target_unit_del_sync_be_out_reg_3__Q) );
ms00f80 pci_target_unit_del_sync_burst_out_reg_u0 ( .ck(ispd_clk), .d(n_2676), .o(pci_target_unit_wbm_sm_pci_tar_burst_ok) );
ms00f80 pci_target_unit_del_sync_comp_comp_pending_reg_u0 ( .ck(ispd_clk), .d(n_7699), .o(wbu_pci_drcomp_pending_in) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_0__u0 ( .ck(ispd_clk), .d(n_2932), .o(pci_target_unit_del_sync_comp_cycle_count_0_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_10__u0 ( .ck(ispd_clk), .d(n_3171), .o(pci_target_unit_del_sync_comp_cycle_count_10_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_11__u0 ( .ck(ispd_clk), .d(n_3355), .o(pci_target_unit_del_sync_comp_cycle_count_11_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_12__u0 ( .ck(ispd_clk), .d(n_4153), .o(pci_target_unit_del_sync_comp_cycle_count_12_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_13__u0 ( .ck(ispd_clk), .d(n_3162), .o(pci_target_unit_del_sync_comp_cycle_count_13_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_14__u0 ( .ck(ispd_clk), .d(n_3490), .o(pci_target_unit_del_sync_comp_cycle_count_14_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_15__u0 ( .ck(ispd_clk), .d(n_3497), .o(pci_target_unit_del_sync_comp_cycle_count_15_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_16__u0 ( .ck(ispd_clk), .d(n_5744), .o(pci_target_unit_del_sync_comp_cycle_count_reg_16__Q) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_1__u0 ( .ck(ispd_clk), .d(n_2938), .o(pci_target_unit_del_sync_comp_cycle_count_1_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_2__u0 ( .ck(ispd_clk), .d(n_2953), .o(pci_target_unit_del_sync_comp_cycle_count_2_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_3__u0 ( .ck(ispd_clk), .d(n_2748), .o(pci_target_unit_del_sync_comp_cycle_count_3_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_4__u0 ( .ck(ispd_clk), .d(n_2774), .o(pci_target_unit_del_sync_comp_cycle_count_4_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_5__u0 ( .ck(ispd_clk), .d(n_2937), .o(pci_target_unit_del_sync_comp_cycle_count_5_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_6__u0 ( .ck(ispd_clk), .d(n_2980), .o(pci_target_unit_del_sync_comp_cycle_count_6_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_7__u0 ( .ck(ispd_clk), .d(n_2757), .o(pci_target_unit_del_sync_comp_cycle_count_7_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_8__u0 ( .ck(ispd_clk), .d(n_3028), .o(pci_target_unit_del_sync_comp_cycle_count_8_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_9__u0 ( .ck(ispd_clk), .d(n_2952), .o(pci_target_unit_del_sync_comp_cycle_count_9_) );
ms00f80 pci_target_unit_del_sync_comp_done_reg_clr_reg_u0 ( .ck(ispd_clk), .d(n_2146), .o(pci_target_unit_del_sync_comp_done_reg_clr_reg_Q) );
in01s01 pci_target_unit_del_sync_comp_done_reg_clr_reg_u1 ( .a(pci_target_unit_del_sync_comp_done_reg_clr_reg_Q), .o(pci_target_unit_del_sync_comp_done_reg_clr) );
ms00f80 pci_target_unit_del_sync_comp_done_reg_main_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_sync_comp_done), .o(pci_target_unit_del_sync_comp_done_reg_main_reg_Q) );
in01s01 pci_target_unit_del_sync_comp_done_reg_main_reg_u1 ( .a(pci_target_unit_del_sync_comp_done_reg_main_reg_Q), .o(pci_target_unit_del_sync_comp_done_reg_main) );
ms00f80 pci_target_unit_del_sync_comp_flush_out_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_comp_cycle_count_reg_16__Q), .o(pci_target_unit_del_sync_comp_flush_out_reg_Q) );
in01s01 pci_target_unit_del_sync_comp_flush_out_reg_u1 ( .a(pci_target_unit_del_sync_comp_flush_out_reg_Q), .o(pci_target_unit_pcit_if_comp_flush_in) );
ms00f80 pci_target_unit_del_sync_comp_req_pending_reg_u0 ( .ck(ispd_clk), .d(n_7706), .o(pci_target_unit_wbm_sm_pci_tar_read_request) );
ms00f80 pci_target_unit_del_sync_comp_rty_exp_clr_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_sync_comp_rty_exp_clr), .o(pci_target_unit_del_sync_comp_rty_exp_clr_reg_Q) );
in01s01 pci_target_unit_del_sync_comp_rty_exp_clr_reg_u1 ( .a(pci_target_unit_del_sync_comp_rty_exp_clr_reg_Q), .o(pci_target_unit_del_sync_comp_rty_exp_clr) );
ms00f80 pci_target_unit_del_sync_comp_rty_exp_reg_reg_u0 ( .ck(ispd_clk), .d(n_4711), .o(pci_target_unit_del_sync_comp_rty_exp_reg) );
ms00f80 pci_target_unit_del_sync_comp_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wbu_pci_drcomp_pending_in), .o(TIMEBOOST_net_15171) );
ms00f80 pci_target_unit_del_sync_done_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_req_done_reg), .o(pci_target_unit_del_sync_sync_comp_done) );
ms00f80 pci_target_unit_del_sync_req_comp_pending_reg_u0 ( .ck(ispd_clk), .d(n_3796), .o(pci_target_unit_del_sync_req_comp_pending) );
ms00f80 pci_target_unit_del_sync_req_comp_pending_sample_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_sync_req_comp_pending), .o(pci_target_unit_del_sync_req_comp_pending_sample_reg_Q) );
in01s01 pci_target_unit_del_sync_req_comp_pending_sample_reg_u1 ( .a(pci_target_unit_del_sync_req_comp_pending_sample_reg_Q), .o(pci_target_unit_del_sync_req_comp_pending_sample) );
ms00f80 pci_target_unit_del_sync_req_done_reg_reg_u0 ( .ck(ispd_clk), .d(n_4532), .o(pci_target_unit_del_sync_req_done_reg) );
ms00f80 pci_target_unit_del_sync_req_req_pending_reg_u0 ( .ck(ispd_clk), .d(n_2445), .o(pci_target_unit_pcit_if_req_req_pending_in) );
ms00f80 pci_target_unit_del_sync_req_rty_exp_clr_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_req_rty_exp_reg), .o(pci_target_unit_del_sync_req_rty_exp_clr_reg_Q) );
in01s01 pci_target_unit_del_sync_req_rty_exp_clr_reg_u1 ( .a(pci_target_unit_del_sync_req_rty_exp_clr_reg_Q), .o(pci_target_unit_del_sync_req_rty_exp_clr) );
ms00f80 pci_target_unit_del_sync_req_rty_exp_reg_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_sync_req_rty_exp), .o(pci_target_unit_del_sync_req_rty_exp_reg) );
ms00f80 pci_target_unit_del_sync_req_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_pcit_if_req_req_pending_in), .o(pci_target_unit_del_sync_req_sync_sync_data_out_reg_0__Q) );
in01s01 pci_target_unit_del_sync_req_sync_sync_data_out_reg_0__u1 ( .a(pci_target_unit_del_sync_req_sync_sync_data_out_reg_0__Q), .o(pci_target_unit_del_sync_sync_comp_req_pending) );
ms00f80 pci_target_unit_del_sync_rty_exp_back_prop_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_738), .o(pci_target_unit_del_sync_sync_comp_rty_exp_clr) );
ms00f80 pci_target_unit_del_sync_rty_exp_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_comp_rty_exp_reg), .o(pci_target_unit_del_sync_sync_req_rty_exp) );
ms00f80 pci_target_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_42), .o(pci_target_unit_fifos_wb_clk_sync_inGreyCount) );
ms00f80 pci_target_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_inGreyCount_reg_1__Q), .o(pci_target_unit_fifos_wb_clk_sync_inGreyCount_36) );
ms00f80 pci_target_unit_fifos_inGreyCount_reg_0__u0 ( .ck(ispd_clk), .d(n_5547), .o(pci_target_unit_fifos_inGreyCount_reg_0__Q) );
in01s01 pci_target_unit_fifos_inGreyCount_reg_0__u1 ( .a(pci_target_unit_fifos_inGreyCount_reg_0__Q), .o(pci_target_unit_fifos_inGreyCount_0_) );
ms00f80 pci_target_unit_fifos_inGreyCount_reg_1__u0 ( .ck(ispd_clk), .d(n_4798), .o(pci_target_unit_fifos_inGreyCount_reg_1__Q) );
ms00f80 pci_target_unit_fifos_outGreyCount_reg_0__u0 ( .ck(ispd_clk), .d(n_13622), .o(pci_target_unit_fifos_outGreyCount_reg_0__Q) );
in01s03 pci_target_unit_fifos_outGreyCount_reg_0__u1 ( .a(pci_target_unit_fifos_outGreyCount_reg_0__Q), .o(pci_target_unit_fifos_outGreyCount_0_) );
ms00f80 pci_target_unit_fifos_outGreyCount_reg_1__u0 ( .ck(ispd_clk), .d(n_13482), .o(pci_target_unit_fifos_outGreyCount_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15193), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15195), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_100) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15197), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_101) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_39) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_40) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15199), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_1__u0 ( .ck(ispd_clk), .d(n_8854), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_2__u0 ( .ck(ispd_clk), .d(n_8855), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_2__Q) );
in01m03 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_2__u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_2__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__u0 ( .ck(ispd_clk), .d(n_8877), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_1__u0 ( .ck(ispd_clk), .d(n_8853), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_1__Q) );
in01s06 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_1__u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_1__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_1_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__u0 ( .ck(ispd_clk), .d(n_8852), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_0__Q) );
in01f20 pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_0__u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_0__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_0_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_39), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_1__Q) );
in01f20 pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_1__u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_1__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_1_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_40), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_2__Q) );
in01f40 pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_2__u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_2__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_2_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_8851), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_8850), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_8849), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(n_8848), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(n_8847), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(n_8846), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg_0__u0 ( .ck(ispd_clk), .d(n_8501), .o(pci_target_unit_fifos_pcir_whole_waddr) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg_1__u0 ( .ck(ispd_clk), .d(n_8505), .o(pci_target_unit_fifos_pcir_whole_waddr_94) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg_2__u0 ( .ck(ispd_clk), .d(n_7836), .o(n_1117) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_0_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_100), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_1_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_101), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_2_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_7830), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_7833), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_7828), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(n_8504), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(n_8502), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(n_7826), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_0__u0 ( .ck(ispd_clk), .d(n_12558), .o(pci_target_unit_pcit_if_pcir_fifo_data_in) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_10__u0 ( .ck(ispd_clk), .d(n_12557), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_775) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_11__u0 ( .ck(ispd_clk), .d(n_12556), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_776) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_12__u0 ( .ck(ispd_clk), .d(n_12555), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_777) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_13__u0 ( .ck(ispd_clk), .d(n_12554), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_778) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_14__u0 ( .ck(ispd_clk), .d(n_12553), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_779) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_15__u0 ( .ck(ispd_clk), .d(n_12771), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_780) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_16__u0 ( .ck(ispd_clk), .d(n_12552), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_781) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_17__u0 ( .ck(ispd_clk), .d(n_12551), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_782) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_18__u0 ( .ck(ispd_clk), .d(n_12550), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_783) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_19__u0 ( .ck(ispd_clk), .d(n_12549), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_784) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_1__u0 ( .ck(ispd_clk), .d(n_12548), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_766) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_20__u0 ( .ck(ispd_clk), .d(n_12547), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_785) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_21__u0 ( .ck(ispd_clk), .d(n_12546), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_786) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_22__u0 ( .ck(ispd_clk), .d(n_12545), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_787) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_23__u0 ( .ck(ispd_clk), .d(n_12544), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_788) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_24__u0 ( .ck(ispd_clk), .d(n_12543), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_789) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_25__u0 ( .ck(ispd_clk), .d(n_12770), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_790) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_26__u0 ( .ck(ispd_clk), .d(n_12542), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_791) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_27__u0 ( .ck(ispd_clk), .d(n_12541), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_792) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_28__u0 ( .ck(ispd_clk), .d(n_12540), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_793) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_29__u0 ( .ck(ispd_clk), .d(n_12539), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_794) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_2__u0 ( .ck(ispd_clk), .d(n_12538), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_767) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_30__u0 ( .ck(ispd_clk), .d(n_12537), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_795) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_31__u0 ( .ck(ispd_clk), .d(n_12536), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_796) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_37__u0 ( .ck(ispd_clk), .d(n_12535), .o(pci_target_unit_pcit_if_pcir_fifo_control_in_637) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_3__u0 ( .ck(ispd_clk), .d(n_12534), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_768) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_4__u0 ( .ck(ispd_clk), .d(n_12533), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_769) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_5__u0 ( .ck(ispd_clk), .d(n_12532), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_770) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_6__u0 ( .ck(ispd_clk), .d(n_12531), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_771) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_7__u0 ( .ck(ispd_clk), .d(n_12769), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_772) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_8__u0 ( .ck(ispd_clk), .d(n_12530), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_773) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_9__u0 ( .ck(ispd_clk), .d(n_12529), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_774) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__u0 ( .ck(ispd_clk), .d(n_7915), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__u0 ( .ck(ispd_clk), .d(n_7913), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__u0 ( .ck(ispd_clk), .d(n_7911), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__u0 ( .ck(ispd_clk), .d(n_7909), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__u0 ( .ck(ispd_clk), .d(n_7907), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__u0 ( .ck(ispd_clk), .d(n_7905), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__u0 ( .ck(ispd_clk), .d(n_7903), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__u0 ( .ck(ispd_clk), .d(n_7901), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__u0 ( .ck(ispd_clk), .d(n_7899), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__u0 ( .ck(ispd_clk), .d(n_7897), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__u0 ( .ck(ispd_clk), .d(n_7895), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__u0 ( .ck(ispd_clk), .d(n_7893), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__u0 ( .ck(ispd_clk), .d(n_7891), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__u0 ( .ck(ispd_clk), .d(n_7889), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__22__u0 ( .ck(ispd_clk), .d(n_7887), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__u0 ( .ck(ispd_clk), .d(n_7885), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__u0 ( .ck(ispd_clk), .d(n_7883), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__u0 ( .ck(ispd_clk), .d(n_7881), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__u0 ( .ck(ispd_clk), .d(n_7879), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__u0 ( .ck(ispd_clk), .d(n_7877), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__u0 ( .ck(ispd_clk), .d(n_7875), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__u0 ( .ck(ispd_clk), .d(n_7873), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__u0 ( .ck(ispd_clk), .d(n_7871), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__u0 ( .ck(ispd_clk), .d(n_7869), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__u0 ( .ck(ispd_clk), .d(n_7867), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__u0 ( .ck(ispd_clk), .d(n_7865), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__u0 ( .ck(ispd_clk), .d(n_7863), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__u0 ( .ck(ispd_clk), .d(n_7861), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__u0 ( .ck(ispd_clk), .d(n_7859), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__u0 ( .ck(ispd_clk), .d(n_7857), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__u0 ( .ck(ispd_clk), .d(n_7855), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__u0 ( .ck(ispd_clk), .d(n_7853), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__u0 ( .ck(ispd_clk), .d(n_7851), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__u0 ( .ck(ispd_clk), .d(n_7849), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__u0 ( .ck(ispd_clk), .d(n_7847), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__u0 ( .ck(ispd_clk), .d(n_7844), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__u0 ( .ck(ispd_clk), .d(n_7842), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__u0 ( .ck(ispd_clk), .d(n_7840), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__u0 ( .ck(ispd_clk), .d(n_7838), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__u0 ( .ck(ispd_clk), .d(n_8123), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__u0 ( .ck(ispd_clk), .d(n_8121), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__u0 ( .ck(ispd_clk), .d(n_8118), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__u0 ( .ck(ispd_clk), .d(n_8116), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__u0 ( .ck(ispd_clk), .d(n_8114), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__u0 ( .ck(ispd_clk), .d(n_8111), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__u0 ( .ck(ispd_clk), .d(n_8109), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__u0 ( .ck(ispd_clk), .d(n_8107), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__u0 ( .ck(ispd_clk), .d(n_8105), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__u0 ( .ck(ispd_clk), .d(n_8102), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__u0 ( .ck(ispd_clk), .d(n_8100), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__u0 ( .ck(ispd_clk), .d(n_8097), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__u0 ( .ck(ispd_clk), .d(n_8094), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__u0 ( .ck(ispd_clk), .d(n_8092), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__u0 ( .ck(ispd_clk), .d(n_8089), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__u0 ( .ck(ispd_clk), .d(n_8087), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__u0 ( .ck(ispd_clk), .d(n_8084), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__u0 ( .ck(ispd_clk), .d(n_8082), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__u0 ( .ck(ispd_clk), .d(n_8079), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__u0 ( .ck(ispd_clk), .d(n_8076), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__u0 ( .ck(ispd_clk), .d(n_8073), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__u0 ( .ck(ispd_clk), .d(n_8071), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__u0 ( .ck(ispd_clk), .d(n_8068), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__u0 ( .ck(ispd_clk), .d(n_8066), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__u0 ( .ck(ispd_clk), .d(n_8064), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__8__u0 ( .ck(ispd_clk), .d(n_8062), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__u0 ( .ck(ispd_clk), .d(n_8059), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__u0 ( .ck(ispd_clk), .d(n_8056), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__u0 ( .ck(ispd_clk), .d(n_8054), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__u0 ( .ck(ispd_clk), .d(n_8052), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__u0 ( .ck(ispd_clk), .d(n_8049), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__u0 ( .ck(ispd_clk), .d(n_8047), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__u0 ( .ck(ispd_clk), .d(n_8044), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__u0 ( .ck(ispd_clk), .d(n_8041), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__u0 ( .ck(ispd_clk), .d(n_8039), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__u0 ( .ck(ispd_clk), .d(n_8036), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__u0 ( .ck(ispd_clk), .d(n_8034), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__u0 ( .ck(ispd_clk), .d(n_8032), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__u0 ( .ck(ispd_clk), .d(n_8030), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__u0 ( .ck(ispd_clk), .d(n_8027), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__u0 ( .ck(ispd_clk), .d(n_8024), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__u0 ( .ck(ispd_clk), .d(n_8021), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__u0 ( .ck(ispd_clk), .d(n_8019), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__u0 ( .ck(ispd_clk), .d(n_8017), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__u0 ( .ck(ispd_clk), .d(n_8014), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__u0 ( .ck(ispd_clk), .d(n_8012), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__u0 ( .ck(ispd_clk), .d(n_8009), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__u0 ( .ck(ispd_clk), .d(n_8007), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__u0 ( .ck(ispd_clk), .d(n_8005), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__u0 ( .ck(ispd_clk), .d(n_8003), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__u0 ( .ck(ispd_clk), .d(n_8001), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__u0 ( .ck(ispd_clk), .d(n_7999), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__u0 ( .ck(ispd_clk), .d(n_7997), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__u0 ( .ck(ispd_clk), .d(n_7995), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__u0 ( .ck(ispd_clk), .d(n_7993), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__u0 ( .ck(ispd_clk), .d(n_7991), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__u0 ( .ck(ispd_clk), .d(n_7989), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__u0 ( .ck(ispd_clk), .d(n_7987), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__u0 ( .ck(ispd_clk), .d(n_7985), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__u0 ( .ck(ispd_clk), .d(n_7983), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__u0 ( .ck(ispd_clk), .d(n_7981), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__u0 ( .ck(ispd_clk), .d(n_7979), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__u0 ( .ck(ispd_clk), .d(n_7977), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__u0 ( .ck(ispd_clk), .d(n_7975), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__u0 ( .ck(ispd_clk), .d(n_7973), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__u0 ( .ck(ispd_clk), .d(n_7971), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__u0 ( .ck(ispd_clk), .d(n_7969), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__u0 ( .ck(ispd_clk), .d(n_7967), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__u0 ( .ck(ispd_clk), .d(n_7965), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__u0 ( .ck(ispd_clk), .d(n_7963), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__u0 ( .ck(ispd_clk), .d(n_7961), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__u0 ( .ck(ispd_clk), .d(n_7959), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__u0 ( .ck(ispd_clk), .d(n_7957), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__u0 ( .ck(ispd_clk), .d(n_7955), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__u0 ( .ck(ispd_clk), .d(n_7953), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__u0 ( .ck(ispd_clk), .d(n_7951), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__u0 ( .ck(ispd_clk), .d(n_7949), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__u0 ( .ck(ispd_clk), .d(n_7947), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__u0 ( .ck(ispd_clk), .d(n_7945), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__u0 ( .ck(ispd_clk), .d(n_7943), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__u0 ( .ck(ispd_clk), .d(n_7941), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__u0 ( .ck(ispd_clk), .d(n_7939), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__u0 ( .ck(ispd_clk), .d(n_7937), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__u0 ( .ck(ispd_clk), .d(n_7935), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__u0 ( .ck(ispd_clk), .d(n_7933), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__u0 ( .ck(ispd_clk), .d(n_7931), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__u0 ( .ck(ispd_clk), .d(n_7929), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__u0 ( .ck(ispd_clk), .d(n_7927), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__u0 ( .ck(ispd_clk), .d(n_7925), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__u0 ( .ck(ispd_clk), .d(n_7923), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__u0 ( .ck(ispd_clk), .d(n_7921), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__u0 ( .ck(ispd_clk), .d(n_7919), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__u0 ( .ck(ispd_clk), .d(n_7917), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__u0 ( .ck(ispd_clk), .d(n_8430), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__u0 ( .ck(ispd_clk), .d(n_8428), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__u0 ( .ck(ispd_clk), .d(n_8426), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__u0 ( .ck(ispd_clk), .d(n_8423), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__u0 ( .ck(ispd_clk), .d(n_8421), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__u0 ( .ck(ispd_clk), .d(n_8419), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__u0 ( .ck(ispd_clk), .d(n_8417), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__u0 ( .ck(ispd_clk), .d(n_8415), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__u0 ( .ck(ispd_clk), .d(n_8413), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__u0 ( .ck(ispd_clk), .d(n_8411), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__u0 ( .ck(ispd_clk), .d(n_8409), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__u0 ( .ck(ispd_clk), .d(n_8406), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__u0 ( .ck(ispd_clk), .d(n_8404), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__u0 ( .ck(ispd_clk), .d(n_8402), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__u0 ( .ck(ispd_clk), .d(n_8400), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__u0 ( .ck(ispd_clk), .d(n_8397), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__u0 ( .ck(ispd_clk), .d(n_8395), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__u0 ( .ck(ispd_clk), .d(n_8393), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__u0 ( .ck(ispd_clk), .d(n_8391), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__u0 ( .ck(ispd_clk), .d(n_8389), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__u0 ( .ck(ispd_clk), .d(n_8387), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__u0 ( .ck(ispd_clk), .d(n_8384), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__u0 ( .ck(ispd_clk), .d(n_8382), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__u0 ( .ck(ispd_clk), .d(n_8379), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__u0 ( .ck(ispd_clk), .d(n_8376), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__u0 ( .ck(ispd_clk), .d(n_8373), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__u0 ( .ck(ispd_clk), .d(n_8371), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__u0 ( .ck(ispd_clk), .d(n_8368), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__u0 ( .ck(ispd_clk), .d(n_8366), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__u0 ( .ck(ispd_clk), .d(n_8364), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__u0 ( .ck(ispd_clk), .d(n_8362), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__u0 ( .ck(ispd_clk), .d(n_8360), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__u0 ( .ck(ispd_clk), .d(n_8358), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__u0 ( .ck(ispd_clk), .d(n_8355), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__u0 ( .ck(ispd_clk), .d(n_8353), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__u0 ( .ck(ispd_clk), .d(n_8351), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__u0 ( .ck(ispd_clk), .d(n_8349), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__u0 ( .ck(ispd_clk), .d(n_8346), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__u0 ( .ck(ispd_clk), .d(n_8344), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__u0 ( .ck(ispd_clk), .d(n_8341), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__u0 ( .ck(ispd_clk), .d(n_8339), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__u0 ( .ck(ispd_clk), .d(n_8337), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__u0 ( .ck(ispd_clk), .d(n_8335), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__u0 ( .ck(ispd_clk), .d(n_8333), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__u0 ( .ck(ispd_clk), .d(n_8331), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__u0 ( .ck(ispd_clk), .d(n_8329), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__u0 ( .ck(ispd_clk), .d(n_8327), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__u0 ( .ck(ispd_clk), .d(n_8325), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__u0 ( .ck(ispd_clk), .d(n_8323), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__u0 ( .ck(ispd_clk), .d(n_8321), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__u0 ( .ck(ispd_clk), .d(n_8319), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__u0 ( .ck(ispd_clk), .d(n_8316), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__u0 ( .ck(ispd_clk), .d(n_8313), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__u0 ( .ck(ispd_clk), .d(n_8311), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__u0 ( .ck(ispd_clk), .d(n_8309), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__u0 ( .ck(ispd_clk), .d(n_8307), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__u0 ( .ck(ispd_clk), .d(n_8304), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__u0 ( .ck(ispd_clk), .d(n_8302), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__u0 ( .ck(ispd_clk), .d(n_8299), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__u0 ( .ck(ispd_clk), .d(n_8297), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__u0 ( .ck(ispd_clk), .d(n_8295), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__u0 ( .ck(ispd_clk), .d(n_8293), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__u0 ( .ck(ispd_clk), .d(n_8291), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__u0 ( .ck(ispd_clk), .d(n_8288), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__u0 ( .ck(ispd_clk), .d(n_8285), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__u0 ( .ck(ispd_clk), .d(n_8283), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__u0 ( .ck(ispd_clk), .d(n_8281), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__u0 ( .ck(ispd_clk), .d(n_8279), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__u0 ( .ck(ispd_clk), .d(n_8277), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__u0 ( .ck(ispd_clk), .d(n_8274), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__u0 ( .ck(ispd_clk), .d(n_8271), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__u0 ( .ck(ispd_clk), .d(n_8269), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__u0 ( .ck(ispd_clk), .d(n_8267), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__u0 ( .ck(ispd_clk), .d(n_8264), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__u0 ( .ck(ispd_clk), .d(n_8262), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__u0 ( .ck(ispd_clk), .d(n_8260), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__u0 ( .ck(ispd_clk), .d(n_8258), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__u0 ( .ck(ispd_clk), .d(n_8255), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__u0 ( .ck(ispd_clk), .d(n_8253), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__u0 ( .ck(ispd_clk), .d(n_8251), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__u0 ( .ck(ispd_clk), .d(n_8248), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__u0 ( .ck(ispd_clk), .d(n_8246), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__u0 ( .ck(ispd_clk), .d(n_8244), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__u0 ( .ck(ispd_clk), .d(n_8241), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__u0 ( .ck(ispd_clk), .d(n_8239), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__u0 ( .ck(ispd_clk), .d(n_8236), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__u0 ( .ck(ispd_clk), .d(n_8234), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__u0 ( .ck(ispd_clk), .d(n_8231), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__u0 ( .ck(ispd_clk), .d(n_8229), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__u0 ( .ck(ispd_clk), .d(n_8226), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__u0 ( .ck(ispd_clk), .d(n_8223), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__u0 ( .ck(ispd_clk), .d(n_8220), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__u0 ( .ck(ispd_clk), .d(n_8218), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__u0 ( .ck(ispd_clk), .d(n_8215), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__u0 ( .ck(ispd_clk), .d(n_8213), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__u0 ( .ck(ispd_clk), .d(n_8210), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__u0 ( .ck(ispd_clk), .d(n_8208), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__u0 ( .ck(ispd_clk), .d(n_8205), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__u0 ( .ck(ispd_clk), .d(n_8203), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__u0 ( .ck(ispd_clk), .d(n_8200), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__u0 ( .ck(ispd_clk), .d(n_8198), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__u0 ( .ck(ispd_clk), .d(n_8196), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__u0 ( .ck(ispd_clk), .d(n_8193), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__u0 ( .ck(ispd_clk), .d(n_8191), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__u0 ( .ck(ispd_clk), .d(n_8189), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__u0 ( .ck(ispd_clk), .d(n_8186), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__u0 ( .ck(ispd_clk), .d(n_8184), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__u0 ( .ck(ispd_clk), .d(n_8182), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__u0 ( .ck(ispd_clk), .d(n_8180), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__u0 ( .ck(ispd_clk), .d(n_8178), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__u0 ( .ck(ispd_clk), .d(n_8175), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__u0 ( .ck(ispd_clk), .d(n_8173), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__u0 ( .ck(ispd_clk), .d(n_8171), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__u0 ( .ck(ispd_clk), .d(n_8168), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__u0 ( .ck(ispd_clk), .d(n_8166), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__u0 ( .ck(ispd_clk), .d(n_8163), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__u0 ( .ck(ispd_clk), .d(n_8161), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__u0 ( .ck(ispd_clk), .d(n_8159), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__u0 ( .ck(ispd_clk), .d(n_8157), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__u0 ( .ck(ispd_clk), .d(n_8154), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__u0 ( .ck(ispd_clk), .d(n_8152), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__u0 ( .ck(ispd_clk), .d(n_8150), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__u0 ( .ck(ispd_clk), .d(n_8147), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__u0 ( .ck(ispd_clk), .d(n_8144), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__u0 ( .ck(ispd_clk), .d(n_8142), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__u0 ( .ck(ispd_clk), .d(n_8139), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__u0 ( .ck(ispd_clk), .d(n_8137), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__u0 ( .ck(ispd_clk), .d(n_8135), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__u0 ( .ck(ispd_clk), .d(n_8132), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__u0 ( .ck(ispd_clk), .d(n_8130), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__u0 ( .ck(ispd_clk), .d(n_8128), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__u0 ( .ck(ispd_clk), .d(n_8125), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_0__Q), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus2) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_1__Q), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_94) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_2__Q), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_95) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15201), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15203), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_74) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15205), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_75) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__u0 ( .ck(ispd_clk), .d(n_13682), .o(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__u0 ( .ck(ispd_clk), .d(n_13619), .o(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__u0 ( .ck(ispd_clk), .d(n_13618), .o(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__u0 ( .ck(ispd_clk), .d(n_16970), .o(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__u0 ( .ck(ispd_clk), .d(n_13479), .o(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__u0 ( .ck(ispd_clk), .d(n_13475), .o(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_74), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_75), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_13616), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_13614), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_13613), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_0__u0 ( .ck(ispd_clk), .d(n_13611), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_1__u0 ( .ck(ispd_clk), .d(n_13609), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_2__u0 ( .ck(ispd_clk), .d(n_13607), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_0__u0 ( .ck(ispd_clk), .d(n_13605), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_1__u0 ( .ck(ispd_clk), .d(n_13603), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_2__u0 ( .ck(ispd_clk), .d(n_13601), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(n_13599), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(n_13597), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(n_13595), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg_0__u0 ( .ck(ispd_clk), .d(n_4616), .o(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg_1__u0 ( .ck(ispd_clk), .d(n_4639), .o(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg_2__u0 ( .ck(ispd_clk), .d(n_4130), .o(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg_0__u0 ( .ck(ispd_clk), .d(n_4614), .o(pci_target_unit_fifos_pciw_whole_waddr) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg_1__u0 ( .ck(ispd_clk), .d(n_4634), .o(pci_target_unit_fifos_pciw_whole_waddr_47) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg_2__u0 ( .ck(ispd_clk), .d(n_4134), .o(n_1293) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus2), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_94), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg_2__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_95), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_4115), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_4107), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_4114), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg_0__u0 ( .ck(ispd_clk), .d(n_4113), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg_1__u0 ( .ck(ispd_clk), .d(n_4108), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg_2__u0 ( .ck(ispd_clk), .d(n_4112), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg_0__u0 ( .ck(ispd_clk), .d(n_4638), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg_1__u0 ( .ck(ispd_clk), .d(n_4138), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg_2__u0 ( .ck(ispd_clk), .d(n_4109), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(n_4636), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(n_4632), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(n_4111), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_0__u0 ( .ck(ispd_clk), .d(n_14613), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_10__u0 ( .ck(ispd_clk), .d(n_14614), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_59) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_11__u0 ( .ck(ispd_clk), .d(n_14612), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_60) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_12__u0 ( .ck(ispd_clk), .d(n_14611), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_61) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_13__u0 ( .ck(ispd_clk), .d(n_14610), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_62) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_14__u0 ( .ck(ispd_clk), .d(n_14609), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_63) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_15__u0 ( .ck(ispd_clk), .d(n_16247), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_64) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_16__u0 ( .ck(ispd_clk), .d(n_14608), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_65) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_17__u0 ( .ck(ispd_clk), .d(n_14607), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_66) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_18__u0 ( .ck(ispd_clk), .d(n_16254), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_67) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_19__u0 ( .ck(ispd_clk), .d(n_16224), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_68) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_1__u0 ( .ck(ispd_clk), .d(n_14605), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_50) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_20__u0 ( .ck(ispd_clk), .d(n_14604), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_69) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_21__u0 ( .ck(ispd_clk), .d(n_14603), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_70) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_22__u0 ( .ck(ispd_clk), .d(n_14602), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_71) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_23__u0 ( .ck(ispd_clk), .d(n_14601), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_72) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_24__u0 ( .ck(ispd_clk), .d(n_16231), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_73) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_25__u0 ( .ck(ispd_clk), .d(n_14599), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_74) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_26__u0 ( .ck(ispd_clk), .d(n_14598), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_75) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_27__u0 ( .ck(ispd_clk), .d(n_14597), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_76) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_28__u0 ( .ck(ispd_clk), .d(n_14596), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_77) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_29__u0 ( .ck(ispd_clk), .d(n_14595), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_78) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_2__u0 ( .ck(ispd_clk), .d(n_14594), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_51) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_30__u0 ( .ck(ispd_clk), .d(n_14593), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_79) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_31__u0 ( .ck(ispd_clk), .d(n_14592), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_80) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_32__u0 ( .ck(ispd_clk), .d(n_14591), .o(pci_target_unit_wbm_sm_pciw_fifo_cbe_in) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_33__u0 ( .ck(ispd_clk), .d(n_14590), .o(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_81) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_34__u0 ( .ck(ispd_clk), .d(n_14589), .o(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_82) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_35__u0 ( .ck(ispd_clk), .d(n_14588), .o(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_83) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_36__u0 ( .ck(ispd_clk), .d(n_16213), .o(pci_target_unit_wbm_sm_pciw_fifo_control_in) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_37__u0 ( .ck(ispd_clk), .d(n_14585), .o(pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_37__Q) );
in01m03 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_37__u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_37__Q), .o(pci_target_unit_wbm_sm_pciw_fifo_control_in_84) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_38__u0 ( .ck(ispd_clk), .d(n_16173), .o(pci_target_unit_wbm_sm_pciw_fifo_control_in_85) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_39__u0 ( .ck(ispd_clk), .d(n_14583), .o(pci_target_unit_wbm_sm_pciw_fifo_control_in_86) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_3__u0 ( .ck(ispd_clk), .d(n_14582), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_52) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_4__u0 ( .ck(ispd_clk), .d(n_16240), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_53) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_5__u0 ( .ck(ispd_clk), .d(n_14580), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_54) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_6__u0 ( .ck(ispd_clk), .d(n_14579), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_55) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_7__u0 ( .ck(ispd_clk), .d(n_16261), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_56) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_8__u0 ( .ck(ispd_clk), .d(n_14578), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_57) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_9__u0 ( .ck(ispd_clk), .d(n_14577), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_58) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__u0 ( .ck(ispd_clk), .d(n_6963), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__u0 ( .ck(ispd_clk), .d(n_5225), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__u0 ( .ck(ispd_clk), .d(n_5223), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__12__u0 ( .ck(ispd_clk), .d(n_5221), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__u0 ( .ck(ispd_clk), .d(n_5218), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__u0 ( .ck(ispd_clk), .d(n_5216), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__15__u0 ( .ck(ispd_clk), .d(n_5214), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__u0 ( .ck(ispd_clk), .d(n_5212), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__u0 ( .ck(ispd_clk), .d(n_5207), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__18__u0 ( .ck(ispd_clk), .d(n_5203), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__u0 ( .ck(ispd_clk), .d(n_5200), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__1__u0 ( .ck(ispd_clk), .d(n_6961), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__u0 ( .ck(ispd_clk), .d(n_5198), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__21__u0 ( .ck(ispd_clk), .d(n_5196), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__u0 ( .ck(ispd_clk), .d(n_5194), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__u0 ( .ck(ispd_clk), .d(n_5192), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__u0 ( .ck(ispd_clk), .d(n_5190), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__u0 ( .ck(ispd_clk), .d(n_5188), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__u0 ( .ck(ispd_clk), .d(n_5185), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__u0 ( .ck(ispd_clk), .d(n_5183), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__u0 ( .ck(ispd_clk), .d(n_5181), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__u0 ( .ck(ispd_clk), .d(n_5179), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__u0 ( .ck(ispd_clk), .d(n_4963), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__u0 ( .ck(ispd_clk), .d(n_5176), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__u0 ( .ck(ispd_clk), .d(n_5174), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__u0 ( .ck(ispd_clk), .d(n_7125), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__u0 ( .ck(ispd_clk), .d(n_5170), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__u0 ( .ck(ispd_clk), .d(n_5168), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__u0 ( .ck(ispd_clk), .d(n_5166), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__36__u0 ( .ck(ispd_clk), .d(n_7123), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__36__Q) );
in01s01 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__36__u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__36__Q), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_0__153) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__u0 ( .ck(ispd_clk), .d(n_7681), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__u0 ( .ck(ispd_clk), .d(n_4926), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__u0 ( .ck(ispd_clk), .d(n_4605), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__u0 ( .ck(ispd_clk), .d(n_5163), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__u0 ( .ck(ispd_clk), .d(n_5161), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__u0 ( .ck(ispd_clk), .d(n_5158), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__6__u0 ( .ck(ispd_clk), .d(n_5156), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__u0 ( .ck(ispd_clk), .d(n_5153), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__u0 ( .ck(ispd_clk), .d(n_5151), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__u0 ( .ck(ispd_clk), .d(n_5146), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__u0 ( .ck(ispd_clk), .d(n_6956), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__u0 ( .ck(ispd_clk), .d(n_5140), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__u0 ( .ck(ispd_clk), .d(n_5138), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__12__u0 ( .ck(ispd_clk), .d(n_4978), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__u0 ( .ck(ispd_clk), .d(n_5136), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__14__u0 ( .ck(ispd_clk), .d(n_5134), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__15__u0 ( .ck(ispd_clk), .d(n_5132), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__16__u0 ( .ck(ispd_clk), .d(n_4959), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__u0 ( .ck(ispd_clk), .d(n_5130), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__18__u0 ( .ck(ispd_clk), .d(n_5128), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__u0 ( .ck(ispd_clk), .d(n_5126), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__u0 ( .ck(ispd_clk), .d(n_6953), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__u0 ( .ck(ispd_clk), .d(n_5124), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__21__u0 ( .ck(ispd_clk), .d(n_5120), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__u0 ( .ck(ispd_clk), .d(n_5118), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__u0 ( .ck(ispd_clk), .d(n_5116), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__u0 ( .ck(ispd_clk), .d(n_5114), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__u0 ( .ck(ispd_clk), .d(n_5112), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__u0 ( .ck(ispd_clk), .d(n_5110), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__u0 ( .ck(ispd_clk), .d(n_5108), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__u0 ( .ck(ispd_clk), .d(n_5106), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__u0 ( .ck(ispd_clk), .d(n_5104), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__u0 ( .ck(ispd_clk), .d(n_5102), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__u0 ( .ck(ispd_clk), .d(n_5100), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__u0 ( .ck(ispd_clk), .d(n_5098), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__u0 ( .ck(ispd_clk), .d(n_7121), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__u0 ( .ck(ispd_clk), .d(n_5096), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__u0 ( .ck(ispd_clk), .d(n_5094), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__u0 ( .ck(ispd_clk), .d(n_5092), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__36__u0 ( .ck(ispd_clk), .d(n_7119), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__36__Q) );
in01s01 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__36__u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__36__Q), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_1__192) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__u0 ( .ck(ispd_clk), .d(n_7679), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__u0 ( .ck(ispd_clk), .d(n_4924), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__u0 ( .ck(ispd_clk), .d(n_4603), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__u0 ( .ck(ispd_clk), .d(n_5088), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__u0 ( .ck(ispd_clk), .d(n_5086), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__u0 ( .ck(ispd_clk), .d(n_5084), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__u0 ( .ck(ispd_clk), .d(n_5082), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__u0 ( .ck(ispd_clk), .d(n_5080), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__u0 ( .ck(ispd_clk), .d(n_5078), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__u0 ( .ck(ispd_clk), .d(n_5076), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__u0 ( .ck(ispd_clk), .d(n_6951), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__u0 ( .ck(ispd_clk), .d(n_5074), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__u0 ( .ck(ispd_clk), .d(n_5071), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__12__u0 ( .ck(ispd_clk), .d(n_5068), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__13__u0 ( .ck(ispd_clk), .d(n_5064), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__u0 ( .ck(ispd_clk), .d(n_5060), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__u0 ( .ck(ispd_clk), .d(n_5058), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__16__u0 ( .ck(ispd_clk), .d(n_5056), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__u0 ( .ck(ispd_clk), .d(n_5054), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__u0 ( .ck(ispd_clk), .d(n_5052), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__u0 ( .ck(ispd_clk), .d(n_5050), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__u0 ( .ck(ispd_clk), .d(n_6948), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__u0 ( .ck(ispd_clk), .d(n_5048), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__21__u0 ( .ck(ispd_clk), .d(n_5046), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__u0 ( .ck(ispd_clk), .d(n_5044), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__u0 ( .ck(ispd_clk), .d(n_5042), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__u0 ( .ck(ispd_clk), .d(n_5040), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__u0 ( .ck(ispd_clk), .d(n_5038), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__u0 ( .ck(ispd_clk), .d(n_5036), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__u0 ( .ck(ispd_clk), .d(n_5033), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__28__u0 ( .ck(ispd_clk), .d(n_5031), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__u0 ( .ck(ispd_clk), .d(n_5029), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__u0 ( .ck(ispd_clk), .d(n_5027), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__u0 ( .ck(ispd_clk), .d(n_5025), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__u0 ( .ck(ispd_clk), .d(n_5023), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__u0 ( .ck(ispd_clk), .d(n_7117), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__u0 ( .ck(ispd_clk), .d(n_5021), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__u0 ( .ck(ispd_clk), .d(n_5018), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__u0 ( .ck(ispd_clk), .d(n_5016), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__36__u0 ( .ck(ispd_clk), .d(n_7126), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__36__Q) );
in01s01 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__36__u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__36__Q), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_2__231) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__u0 ( .ck(ispd_clk), .d(n_7683), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__u0 ( .ck(ispd_clk), .d(n_4922), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__u0 ( .ck(ispd_clk), .d(n_4607), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__u0 ( .ck(ispd_clk), .d(n_5066), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__u0 ( .ck(ispd_clk), .d(n_5205), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__u0 ( .ck(ispd_clk), .d(n_4957), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__u0 ( .ck(ispd_clk), .d(n_5014), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__u0 ( .ck(ispd_clk), .d(n_4961), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__u0 ( .ck(ispd_clk), .d(n_5012), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__u0 ( .ck(ispd_clk), .d(n_5062), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__u0 ( .ck(ispd_clk), .d(n_6946), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__u0 ( .ck(ispd_clk), .d(n_5009), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__u0 ( .ck(ispd_clk), .d(n_5149), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__12__u0 ( .ck(ispd_clk), .d(n_5090), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__13__u0 ( .ck(ispd_clk), .d(n_5006), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__u0 ( .ck(ispd_clk), .d(n_5003), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__u0 ( .ck(ispd_clk), .d(n_5122), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__16__u0 ( .ck(ispd_clk), .d(n_5001), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__u0 ( .ck(ispd_clk), .d(n_5143), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__u0 ( .ck(ispd_clk), .d(n_4999), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__u0 ( .ck(ispd_clk), .d(n_5172), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__u0 ( .ck(ispd_clk), .d(n_6958), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__u0 ( .ck(ispd_clk), .d(n_4996), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__21__u0 ( .ck(ispd_clk), .d(n_4993), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__u0 ( .ck(ispd_clk), .d(n_5210), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__u0 ( .ck(ispd_clk), .d(n_4991), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__u0 ( .ck(ispd_clk), .d(n_4988), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__u0 ( .ck(ispd_clk), .d(n_4986), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__u0 ( .ck(ispd_clk), .d(n_5227), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__u0 ( .ck(ispd_clk), .d(n_4984), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__28__u0 ( .ck(ispd_clk), .d(n_4941), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__u0 ( .ck(ispd_clk), .d(n_4982), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__u0 ( .ck(ispd_clk), .d(n_4943), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__u0 ( .ck(ispd_clk), .d(n_4980), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__u0 ( .ck(ispd_clk), .d(n_4945), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__u0 ( .ck(ispd_clk), .d(n_7112), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__u0 ( .ck(ispd_clk), .d(n_4949), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__u0 ( .ck(ispd_clk), .d(n_4955), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__u0 ( .ck(ispd_clk), .d(n_4953), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__36__u0 ( .ck(ispd_clk), .d(n_7122), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__36__Q) );
in01s01 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__36__u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__36__Q), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_3__270) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__u0 ( .ck(ispd_clk), .d(n_7677), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__u0 ( .ck(ispd_clk), .d(n_4920), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__u0 ( .ck(ispd_clk), .d(n_4601), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__u0 ( .ck(ispd_clk), .d(n_4975), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__u0 ( .ck(ispd_clk), .d(n_4947), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__u0 ( .ck(ispd_clk), .d(n_4973), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__u0 ( .ck(ispd_clk), .d(n_4970), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__u0 ( .ck(ispd_clk), .d(n_4968), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__u0 ( .ck(ispd_clk), .d(n_4951), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__u0 ( .ck(ispd_clk), .d(n_4965), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__u0 ( .ck(ispd_clk), .d(n_6977), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__u0 ( .ck(ispd_clk), .d(n_5414), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__u0 ( .ck(ispd_clk), .d(n_5308), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__u0 ( .ck(ispd_clk), .d(n_5361), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__13__u0 ( .ck(ispd_clk), .d(n_5363), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__14__u0 ( .ck(ispd_clk), .d(n_5366), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__u0 ( .ck(ispd_clk), .d(n_5371), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__16__u0 ( .ck(ispd_clk), .d(n_5380), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__u0 ( .ck(ispd_clk), .d(n_5386), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__u0 ( .ck(ispd_clk), .d(n_5388), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__u0 ( .ck(ispd_clk), .d(n_5409), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__u0 ( .ck(ispd_clk), .d(n_6975), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__u0 ( .ck(ispd_clk), .d(n_5290), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__u0 ( .ck(ispd_clk), .d(n_5303), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__u0 ( .ck(ispd_clk), .d(n_5300), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__u0 ( .ck(ispd_clk), .d(n_5406), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__u0 ( .ck(ispd_clk), .d(n_5404), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__u0 ( .ck(ispd_clk), .d(n_5318), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__u0 ( .ck(ispd_clk), .d(n_5402), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__u0 ( .ck(ispd_clk), .d(n_5337), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__u0 ( .ck(ispd_clk), .d(n_5399), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__u0 ( .ck(ispd_clk), .d(n_5354), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__u0 ( .ck(ispd_clk), .d(n_5418), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__u0 ( .ck(ispd_clk), .d(n_5421), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__u0 ( .ck(ispd_clk), .d(n_5396), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__u0 ( .ck(ispd_clk), .d(n_7128), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__u0 ( .ck(ispd_clk), .d(n_5393), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__u0 ( .ck(ispd_clk), .d(n_5391), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__u0 ( .ck(ispd_clk), .d(n_5305), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__u0 ( .ck(ispd_clk), .d(n_6115), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__u0 ( .ck(ispd_clk), .d(n_7692), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__u0 ( .ck(ispd_clk), .d(n_4928), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__u0 ( .ck(ispd_clk), .d(n_4623), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__u0 ( .ck(ispd_clk), .d(n_5323), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__u0 ( .ck(ispd_clk), .d(n_5332), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__u0 ( .ck(ispd_clk), .d(n_5315), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__u0 ( .ck(ispd_clk), .d(n_5412), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__u0 ( .ck(ispd_clk), .d(n_5267), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__u0 ( .ck(ispd_clk), .d(n_5416), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__u0 ( .ck(ispd_clk), .d(n_5448), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__u0 ( .ck(ispd_clk), .d(n_6971), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__u0 ( .ck(ispd_clk), .d(n_5383), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__u0 ( .ck(ispd_clk), .d(n_5265), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__u0 ( .ck(ispd_clk), .d(n_5378), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__13__u0 ( .ck(ispd_clk), .d(n_5275), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__u0 ( .ck(ispd_clk), .d(n_5376), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__15__u0 ( .ck(ispd_clk), .d(n_5281), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__16__u0 ( .ck(ispd_clk), .d(n_5288), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__u0 ( .ck(ispd_clk), .d(n_5296), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__u0 ( .ck(ispd_clk), .d(n_5373), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__u0 ( .ck(ispd_clk), .d(n_5298), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__u0 ( .ck(ispd_clk), .d(n_6967), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__u0 ( .ck(ispd_clk), .d(n_5237), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__u0 ( .ck(ispd_clk), .d(n_5368), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__u0 ( .ck(ispd_clk), .d(n_5244), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__u0 ( .ck(ispd_clk), .d(n_5255), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__u0 ( .ck(ispd_clk), .d(n_5258), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__u0 ( .ck(ispd_clk), .d(n_5424), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__u0 ( .ck(ispd_clk), .d(n_5429), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__u0 ( .ck(ispd_clk), .d(n_5433), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__u0 ( .ck(ispd_clk), .d(n_5441), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__u0 ( .ck(ispd_clk), .d(n_5450), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__u0 ( .ck(ispd_clk), .d(n_5458), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__u0 ( .ck(ispd_clk), .d(n_5461), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__u0 ( .ck(ispd_clk), .d(n_5463), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__u0 ( .ck(ispd_clk), .d(n_7134), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__u0 ( .ck(ispd_clk), .d(n_5478), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__u0 ( .ck(ispd_clk), .d(n_5481), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__u0 ( .ck(ispd_clk), .d(n_5491), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__u0 ( .ck(ispd_clk), .d(n_6132), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__u0 ( .ck(ispd_clk), .d(n_7689), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__u0 ( .ck(ispd_clk), .d(n_4932), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__u0 ( .ck(ispd_clk), .d(n_4627), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__u0 ( .ck(ispd_clk), .d(n_5493), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__u0 ( .ck(ispd_clk), .d(n_5497), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__u0 ( .ck(ispd_clk), .d(n_5501), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__u0 ( .ck(ispd_clk), .d(n_5505), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__u0 ( .ck(ispd_clk), .d(n_5358), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__u0 ( .ck(ispd_clk), .d(n_5509), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__u0 ( .ck(ispd_clk), .d(n_5511), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__u0 ( .ck(ispd_clk), .d(n_6980), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__u0 ( .ck(ispd_clk), .d(n_5470), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__u0 ( .ck(ispd_clk), .d(n_5356), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__12__u0 ( .ck(ispd_clk), .d(n_5539), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__u0 ( .ck(ispd_clk), .d(n_5534), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__14__u0 ( .ck(ispd_clk), .d(n_5248), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__u0 ( .ck(ispd_clk), .d(n_5351), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__16__u0 ( .ck(ispd_clk), .d(n_5531), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__u0 ( .ck(ispd_clk), .d(n_5349), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__u0 ( .ck(ispd_clk), .d(n_5483), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__u0 ( .ck(ispd_clk), .d(n_5347), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__u0 ( .ck(ispd_clk), .d(n_5716), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__u0 ( .ck(ispd_clk), .d(n_5345), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__u0 ( .ck(ispd_clk), .d(n_5521), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__u0 ( .ck(ispd_clk), .d(n_5342), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__u0 ( .ck(ispd_clk), .d(n_5528), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__u0 ( .ck(ispd_clk), .d(n_5499), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__u0 ( .ck(ispd_clk), .d(n_5260), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__u0 ( .ck(ispd_clk), .d(n_5339), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__u0 ( .ck(ispd_clk), .d(n_5240), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__28__u0 ( .ck(ispd_clk), .d(n_5242), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__u0 ( .ck(ispd_clk), .d(n_5253), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__u0 ( .ck(ispd_clk), .d(n_5427), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__u0 ( .ck(ispd_clk), .d(n_5446), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__u0 ( .ck(ispd_clk), .d(n_5467), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__u0 ( .ck(ispd_clk), .d(n_7130), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__u0 ( .ck(ispd_clk), .d(n_5335), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__u0 ( .ck(ispd_clk), .d(n_5537), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__u0 ( .ck(ispd_clk), .d(n_5489), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__u0 ( .ck(ispd_clk), .d(n_6135), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__u0 ( .ck(ispd_clk), .d(n_7694), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__u0 ( .ck(ispd_clk), .d(n_4930), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__u0 ( .ck(ispd_clk), .d(n_4625), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__u0 ( .ck(ispd_clk), .d(n_5503), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__u0 ( .ck(ispd_clk), .d(n_5330), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__u0 ( .ck(ispd_clk), .d(n_5517), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__u0 ( .ck(ispd_clk), .d(n_5513), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__u0 ( .ck(ispd_clk), .d(n_5523), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__u0 ( .ck(ispd_clk), .d(n_5327), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__u0 ( .ck(ispd_clk), .d(n_5543), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__u0 ( .ck(ispd_clk), .d(n_6969), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__u0 ( .ck(ispd_clk), .d(n_5277), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__u0 ( .ck(ispd_clk), .d(n_5285), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__u0 ( .ck(ispd_clk), .d(n_5325), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__u0 ( .ck(ispd_clk), .d(n_5438), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__14__u0 ( .ck(ispd_clk), .d(n_5431), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__u0 ( .ck(ispd_clk), .d(n_5454), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__16__u0 ( .ck(ispd_clk), .d(n_5320), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__u0 ( .ck(ispd_clk), .d(n_5272), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__u0 ( .ck(ispd_clk), .d(n_5293), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__u0 ( .ck(ispd_clk), .d(n_5235), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__u0 ( .ck(ispd_clk), .d(n_6973), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__u0 ( .ck(ispd_clk), .d(n_5246), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__u0 ( .ck(ispd_clk), .d(n_5486), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__22__u0 ( .ck(ispd_clk), .d(n_5495), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__u0 ( .ck(ispd_clk), .d(n_5313), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__u0 ( .ck(ispd_clk), .d(n_5519), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__u0 ( .ck(ispd_clk), .d(n_5526), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__u0 ( .ck(ispd_clk), .d(n_5435), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__u0 ( .ck(ispd_clk), .d(n_5452), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__28__u0 ( .ck(ispd_clk), .d(n_5311), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__u0 ( .ck(ispd_clk), .d(n_5456), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__u0 ( .ck(ispd_clk), .d(n_5507), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__u0 ( .ck(ispd_clk), .d(n_5476), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__u0 ( .ck(ispd_clk), .d(n_5541), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__u0 ( .ck(ispd_clk), .d(n_7132), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__u0 ( .ck(ispd_clk), .d(n_5444), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__u0 ( .ck(ispd_clk), .d(n_5465), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__u0 ( .ck(ispd_clk), .d(n_5515), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__u0 ( .ck(ispd_clk), .d(n_6125), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__u0 ( .ck(ispd_clk), .d(n_7687), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__u0 ( .ck(ispd_clk), .d(n_4934), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__u0 ( .ck(ispd_clk), .d(n_4621), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__u0 ( .ck(ispd_clk), .d(n_5251), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__u0 ( .ck(ispd_clk), .d(n_5472), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__u0 ( .ck(ispd_clk), .d(n_5263), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__u0 ( .ck(ispd_clk), .d(n_5474), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__u0 ( .ck(ispd_clk), .d(n_5269), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__u0 ( .ck(ispd_clk), .d(n_5279), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__u0 ( .ck(ispd_clk), .d(n_5283), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_inTransactionCount_reg_0__u0 ( .ck(ispd_clk), .d(n_4797), .o(pci_target_unit_fifos_pciw_inTransactionCount_0_) );
ms00f80 pci_target_unit_fifos_pciw_inTransactionCount_reg_1__u0 ( .ck(ispd_clk), .d(n_5548), .o(pci_target_unit_fifos_pciw_inTransactionCount_reg_1__Q) );
in01s01 pci_target_unit_fifos_pciw_inTransactionCount_reg_1__u1 ( .a(pci_target_unit_fifos_pciw_inTransactionCount_reg_1__Q), .o(pci_target_unit_fifos_pciw_inTransactionCount_1_) );
ms00f80 pci_target_unit_fifos_pciw_outTransactionCount_reg_0__u0 ( .ck(ispd_clk), .d(n_13483), .o(pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pciw_outTransactionCount_reg_1__u0 ( .ck(ispd_clk), .d(n_13623), .o(pci_target_unit_fifos_pciw_outTransactionCount_reg_1__Q) );
in01s01 pci_target_unit_fifos_pciw_outTransactionCount_reg_1__u1 ( .a(pci_target_unit_fifos_pciw_outTransactionCount_reg_1__Q), .o(pci_target_unit_fifos_pciw_outTransactionCount_1_) );
ms00f80 pci_target_unit_fifos_wb_clk_inGreyCount_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_wb_clk_sync_inGreyCount), .o(pci_target_unit_fifos_wb_clk_inGreyCount_0_) );
ms00f80 pci_target_unit_fifos_wb_clk_inGreyCount_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_wb_clk_sync_inGreyCount_36), .o(pci_target_unit_fifos_wb_clk_inGreyCount_1_) );
ms00f80 pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg_u0 ( .ck(ispd_clk), .d(n_4667), .o(pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg_Q) );
in01s06 pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg_u1 ( .a(pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg_Q), .o(pci_target_unit_fifos_pcir_flush_in) );
ms00f80 pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg_u0 ( .ck(ispd_clk), .d(n_12170), .o(pci_target_unit_pci_target_if_keep_desconnect_wo_data_set) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_0__u0 ( .ck(ispd_clk), .d(n_2603), .o(pci_target_unit_pci_target_if_norm_address_reg_0__Q) );
in01s01 pci_target_unit_pci_target_if_norm_address_reg_0__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_0__Q), .o(pci_target_unit_del_sync_addr_in) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_10__u0 ( .ck(ispd_clk), .d(n_2592), .o(pci_target_unit_del_sync_addr_in_213) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_11__u0 ( .ck(ispd_clk), .d(n_2595), .o(pci_target_unit_del_sync_addr_in_214) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_12__u0 ( .ck(ispd_clk), .d(n_2576), .o(pci_target_unit_del_sync_addr_in_215) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_13__u0 ( .ck(ispd_clk), .d(n_2593), .o(pci_target_unit_del_sync_addr_in_216) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_14__u0 ( .ck(ispd_clk), .d(n_2573), .o(pci_target_unit_del_sync_addr_in_217) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_15__u0 ( .ck(ispd_clk), .d(n_2574), .o(pci_target_unit_del_sync_addr_in_218) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_16__u0 ( .ck(ispd_clk), .d(n_2577), .o(pci_target_unit_del_sync_addr_in_219) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_17__u0 ( .ck(ispd_clk), .d(n_2570), .o(pci_target_unit_del_sync_addr_in_220) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_18__u0 ( .ck(ispd_clk), .d(n_2594), .o(pci_target_unit_del_sync_addr_in_221) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_19__u0 ( .ck(ispd_clk), .d(n_2588), .o(pci_target_unit_del_sync_addr_in_222) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_1__u0 ( .ck(ispd_clk), .d(n_2794), .o(pci_target_unit_pci_target_if_norm_address_reg_1__Q) );
in01s01 pci_target_unit_pci_target_if_norm_address_reg_1__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_1__Q), .o(pci_target_unit_del_sync_addr_in_204) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_20__u0 ( .ck(ispd_clk), .d(n_2571), .o(pci_target_unit_del_sync_addr_in_223) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_21__u0 ( .ck(ispd_clk), .d(n_2581), .o(pci_target_unit_del_sync_addr_in_224) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_22__u0 ( .ck(ispd_clk), .d(n_2590), .o(pci_target_unit_del_sync_addr_in_225) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_23__u0 ( .ck(ispd_clk), .d(n_2482), .o(pci_target_unit_del_sync_addr_in_226) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_24__u0 ( .ck(ispd_clk), .d(n_2572), .o(pci_target_unit_del_sync_addr_in_227) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_25__u0 ( .ck(ispd_clk), .d(n_2582), .o(pci_target_unit_del_sync_addr_in_228) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_26__u0 ( .ck(ispd_clk), .d(n_2583), .o(pci_target_unit_del_sync_addr_in_229) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_27__u0 ( .ck(ispd_clk), .d(n_2584), .o(pci_target_unit_del_sync_addr_in_230) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_28__u0 ( .ck(ispd_clk), .d(n_2585), .o(pci_target_unit_del_sync_addr_in_231) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_29__u0 ( .ck(ispd_clk), .d(n_2569), .o(pci_target_unit_del_sync_addr_in_232) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_2__u0 ( .ck(ispd_clk), .d(n_2792), .o(pci_target_unit_pci_target_if_norm_address_reg_2__Q) );
in01s01 pci_target_unit_pci_target_if_norm_address_reg_2__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_2__Q), .o(pci_target_unit_del_sync_addr_in_205) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_30__u0 ( .ck(ispd_clk), .d(n_2587), .o(pci_target_unit_del_sync_addr_in_233) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_31__u0 ( .ck(ispd_clk), .d(n_2586), .o(pci_target_unit_del_sync_addr_in_234) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_3__u0 ( .ck(ispd_clk), .d(n_2789), .o(pci_target_unit_pci_target_if_norm_address_reg_3__Q) );
in01s01 pci_target_unit_pci_target_if_norm_address_reg_3__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_3__Q), .o(pci_target_unit_del_sync_addr_in_206) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_4__u0 ( .ck(ispd_clk), .d(n_2734), .o(pci_target_unit_pci_target_if_norm_address_reg_4__Q) );
in01s01 pci_target_unit_pci_target_if_norm_address_reg_4__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_4__Q), .o(pci_target_unit_del_sync_addr_in_207) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_5__u0 ( .ck(ispd_clk), .d(n_2605), .o(pci_target_unit_pci_target_if_norm_address_reg_5__Q) );
in01s01 pci_target_unit_pci_target_if_norm_address_reg_5__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_5__Q), .o(pci_target_unit_del_sync_addr_in_208) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_6__u0 ( .ck(ispd_clk), .d(n_2787), .o(pci_target_unit_pci_target_if_norm_address_reg_6__Q) );
in01s01 pci_target_unit_pci_target_if_norm_address_reg_6__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_6__Q), .o(pci_target_unit_del_sync_addr_in_209) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_7__u0 ( .ck(ispd_clk), .d(n_2608), .o(pci_target_unit_pci_target_if_norm_address_reg_7__Q) );
in01s01 pci_target_unit_pci_target_if_norm_address_reg_7__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_7__Q), .o(pci_target_unit_del_sync_addr_in_210) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_8__u0 ( .ck(ispd_clk), .d(n_2611), .o(pci_target_unit_pci_target_if_norm_address_reg_8__Q) );
in01s01 pci_target_unit_pci_target_if_norm_address_reg_8__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_8__Q), .o(pci_target_unit_del_sync_addr_in_211) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_9__u0 ( .ck(ispd_clk), .d(n_2613), .o(pci_target_unit_pci_target_if_norm_address_reg_9__Q) );
in01s01 pci_target_unit_pci_target_if_norm_address_reg_9__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_9__Q), .o(pci_target_unit_del_sync_addr_in_212) );
ms00f80 pci_target_unit_pci_target_if_norm_bc_reg_0__u0 ( .ck(ispd_clk), .d(n_3220), .o(pci_target_unit_del_sync_bc_in) );
ms00f80 pci_target_unit_pci_target_if_norm_bc_reg_1__u0 ( .ck(ispd_clk), .d(n_2793), .o(pci_target_unit_del_sync_bc_in_201) );
ms00f80 pci_target_unit_pci_target_if_norm_bc_reg_2__u0 ( .ck(ispd_clk), .d(n_2575), .o(pci_target_unit_del_sync_bc_in_202) );
ms00f80 pci_target_unit_pci_target_if_norm_bc_reg_3__u0 ( .ck(ispd_clk), .d(n_2579), .o(pci_target_unit_del_sync_bc_in_203) );
ms00f80 pci_target_unit_pci_target_if_norm_prf_en_reg_u0 ( .ck(ispd_clk), .d(n_8659), .o(pci_target_unit_pci_target_if_norm_prf_en) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_reg_1__u0 ( .ck(ispd_clk), .d(n_13146), .o(pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_77) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_0__u0 ( .ck(ispd_clk), .d(n_12980), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_0__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_10__u0 ( .ck(ispd_clk), .d(n_12978), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_10__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_11__u0 ( .ck(ispd_clk), .d(n_12976), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_11__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_12__u0 ( .ck(ispd_clk), .d(n_12974), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_12__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_13__u0 ( .ck(ispd_clk), .d(n_12972), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_13__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_14__u0 ( .ck(ispd_clk), .d(n_12970), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_14__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_15__u0 ( .ck(ispd_clk), .d(n_13097), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_15__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_16__u0 ( .ck(ispd_clk), .d(n_12968), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_16__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_17__u0 ( .ck(ispd_clk), .d(n_12966), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_17__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_18__u0 ( .ck(ispd_clk), .d(n_13095), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_18__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_19__u0 ( .ck(ispd_clk), .d(n_13094), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_19__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_1__u0 ( .ck(ispd_clk), .d(n_13093), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_1__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_20__u0 ( .ck(ispd_clk), .d(n_13091), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_20__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_21__u0 ( .ck(ispd_clk), .d(n_13090), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_21__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_22__u0 ( .ck(ispd_clk), .d(n_13089), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_22__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_23__u0 ( .ck(ispd_clk), .d(n_13088), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_23__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_24__u0 ( .ck(ispd_clk), .d(n_13087), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_24__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_25__u0 ( .ck(ispd_clk), .d(n_13125), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_25__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_26__u0 ( .ck(ispd_clk), .d(n_13086), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_26__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_27__u0 ( .ck(ispd_clk), .d(n_13085), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_27__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_28__u0 ( .ck(ispd_clk), .d(n_13084), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_28__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_29__u0 ( .ck(ispd_clk), .d(n_13083), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_29__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_2__u0 ( .ck(ispd_clk), .d(n_13082), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_2__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_30__u0 ( .ck(ispd_clk), .d(n_13081), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_30__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_31__u0 ( .ck(ispd_clk), .d(n_13080), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_31__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_3__u0 ( .ck(ispd_clk), .d(n_13079), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_3__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_4__u0 ( .ck(ispd_clk), .d(n_13078), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_4__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_5__u0 ( .ck(ispd_clk), .d(n_13077), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_5__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_6__u0 ( .ck(ispd_clk), .d(n_13076), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_6__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_7__u0 ( .ck(ispd_clk), .d(n_13123), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_7__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_8__u0 ( .ck(ispd_clk), .d(n_13075), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_8__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_9__u0 ( .ck(ispd_clk), .d(n_13074), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_9__Q) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_2776), .o(pci_target_unit_fifos_pciw_addr_data_in) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_10__u0 ( .ck(ispd_clk), .d(n_2519), .o(pci_target_unit_fifos_pciw_addr_data_in_130) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_11__u0 ( .ck(ispd_clk), .d(n_2517), .o(pci_target_unit_fifos_pciw_addr_data_in_131) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_12__u0 ( .ck(ispd_clk), .d(n_2546), .o(pci_target_unit_fifos_pciw_addr_data_in_132) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_13__u0 ( .ck(ispd_clk), .d(n_2534), .o(pci_target_unit_fifos_pciw_addr_data_in_133) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_14__u0 ( .ck(ispd_clk), .d(n_2496), .o(pci_target_unit_fifos_pciw_addr_data_in_134) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_15__u0 ( .ck(ispd_clk), .d(n_2498), .o(pci_target_unit_fifos_pciw_addr_data_in_135) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_16__u0 ( .ck(ispd_clk), .d(n_2537), .o(pci_target_unit_fifos_pciw_addr_data_in_136) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_17__u0 ( .ck(ispd_clk), .d(n_2536), .o(pci_target_unit_fifos_pciw_addr_data_in_137) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_18__u0 ( .ck(ispd_clk), .d(n_2530), .o(pci_target_unit_fifos_pciw_addr_data_in_138) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_19__u0 ( .ck(ispd_clk), .d(n_2528), .o(pci_target_unit_fifos_pciw_addr_data_in_139) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_1__u0 ( .ck(ispd_clk), .d(n_2973), .o(pci_target_unit_fifos_pciw_addr_data_in_121) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_20__u0 ( .ck(ispd_clk), .d(n_2540), .o(pci_target_unit_fifos_pciw_addr_data_in_140) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_21__u0 ( .ck(ispd_clk), .d(n_2531), .o(pci_target_unit_fifos_pciw_addr_data_in_141) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_22__u0 ( .ck(ispd_clk), .d(n_2514), .o(pci_target_unit_fifos_pciw_addr_data_in_142) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_23__u0 ( .ck(ispd_clk), .d(n_2539), .o(pci_target_unit_fifos_pciw_addr_data_in_143) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_24__u0 ( .ck(ispd_clk), .d(n_2502), .o(pci_target_unit_fifos_pciw_addr_data_in_144) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_25__u0 ( .ck(ispd_clk), .d(n_2522), .o(pci_target_unit_fifos_pciw_addr_data_in_145) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_26__u0 ( .ck(ispd_clk), .d(n_2533), .o(pci_target_unit_fifos_pciw_addr_data_in_146) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_27__u0 ( .ck(ispd_clk), .d(n_2543), .o(pci_target_unit_fifos_pciw_addr_data_in_147) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_28__u0 ( .ck(ispd_clk), .d(n_2518), .o(pci_target_unit_fifos_pciw_addr_data_in_148) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_29__u0 ( .ck(ispd_clk), .d(n_2505), .o(pci_target_unit_fifos_pciw_addr_data_in_149) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2516), .o(pci_target_unit_fifos_pciw_addr_data_in_122) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_30__u0 ( .ck(ispd_clk), .d(n_2510), .o(pci_target_unit_fifos_pciw_addr_data_in_150) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_31__u0 ( .ck(ispd_clk), .d(n_2497), .o(pci_target_unit_fifos_pciw_addr_data_in_151) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2500), .o(pci_target_unit_fifos_pciw_addr_data_in_123) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_4__u0 ( .ck(ispd_clk), .d(n_2527), .o(pci_target_unit_fifos_pciw_addr_data_in_124) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_5__u0 ( .ck(ispd_clk), .d(n_2545), .o(pci_target_unit_fifos_pciw_addr_data_in_125) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_6__u0 ( .ck(ispd_clk), .d(n_2513), .o(pci_target_unit_fifos_pciw_addr_data_in_126) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_7__u0 ( .ck(ispd_clk), .d(n_2542), .o(pci_target_unit_fifos_pciw_addr_data_in_127) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_8__u0 ( .ck(ispd_clk), .d(n_2508), .o(pci_target_unit_fifos_pciw_addr_data_in_128) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_9__u0 ( .ck(ispd_clk), .d(n_2504), .o(pci_target_unit_fifos_pciw_addr_data_in_129) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg_0__u0 ( .ck(ispd_clk), .d(n_3000), .o(pci_target_unit_fifos_pciw_cbe_in) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg_1__u0 ( .ck(ispd_clk), .d(n_2501), .o(pci_target_unit_fifos_pciw_cbe_in_152) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2524), .o(pci_target_unit_fifos_pciw_cbe_in_153) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2521), .o(pci_target_unit_fifos_pciw_cbe_in_154) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_0__u0 ( .ck(ispd_clk), .d(FE_OFN793_n_2547), .o(pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_0__Q) );
in01s01 pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_0__u1 ( .a(pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_0__Q), .o(pci_target_unit_fifos_pciw_control_in) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_1__u0 ( .ck(ispd_clk), .d(n_4142), .o(pci_target_unit_fifos_pciw_control_in_155) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2729), .o(pci_target_unit_fifos_pciw_control_in_156) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2031), .o(pci_target_unit_fifos_pciw_control_in_157) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_wenable_out_reg_u0 ( .ck(ispd_clk), .d(n_8566), .o(pci_target_unit_fifos_pciw_wenable_in) );
ms00f80 pci_target_unit_pci_target_if_same_read_reg_reg_u0 ( .ck(ispd_clk), .d(n_5640), .o(pci_target_unit_pci_target_if_same_read_reg) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_0__u0 ( .ck(ispd_clk), .d(n_2602), .o(conf_w_addr_in) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_1__u0 ( .ck(ispd_clk), .d(n_2780), .o(conf_w_addr_in_931) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_2__u0 ( .ck(ispd_clk), .d(n_4214), .o(conf_w_addr_in_932) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_3__u0 ( .ck(ispd_clk), .d(n_3216), .o(conf_w_addr_in_933) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_4__u0 ( .ck(ispd_clk), .d(n_2781), .o(n_2078) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_5__u0 ( .ck(ispd_clk), .d(n_2782), .o(conf_w_addr_in_935) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_6__u0 ( .ck(ispd_clk), .d(n_2784), .o(n_15998) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_7__u0 ( .ck(ispd_clk), .d(n_2745), .o(conf_w_addr_in_937) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_8__u0 ( .ck(ispd_clk), .d(n_2786), .o(conf_w_addr_in_938) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_9__u0 ( .ck(ispd_clk), .d(n_2785), .o(conf_w_addr_in_939) );
ms00f80 pci_target_unit_pci_target_if_target_rd_reg_u0 ( .ck(ispd_clk), .d(n_3380), .o(pci_target_unit_pci_target_if_target_rd_completed) );
ms00f80 pci_target_unit_pci_target_sm_backoff_reg_u0 ( .ck(ispd_clk), .d(n_14630), .o(pci_target_unit_pci_target_sm_backoff) );
ms00f80 pci_target_unit_pci_target_sm_bckp_trdy_reg_reg_u0 ( .ck(ispd_clk), .d(output_backup_trdy_out_reg_Q), .o(pci_target_unit_pci_target_sm_bckp_trdy_reg_reg_Q) );
in01f20 pci_target_unit_pci_target_sm_bckp_trdy_reg_reg_u1 ( .a(pci_target_unit_pci_target_sm_bckp_trdy_reg_reg_Q), .o(n_2597) );
ms00f80 pci_target_unit_pci_target_sm_c_state_reg_0__u0 ( .ck(ispd_clk), .d(n_9180), .o(n_1628) );
ms00f80 pci_target_unit_pci_target_sm_c_state_reg_1__u0 ( .ck(ispd_clk), .d(n_9179), .o(pci_target_unit_pci_target_sm_n_2) );
ms00f80 pci_target_unit_pci_target_sm_c_state_reg_2__u0 ( .ck(ispd_clk), .d(n_9176), .o(pci_target_unit_pci_target_sm_n_3) );
ms00f80 pci_target_unit_pci_target_sm_cnf_progress_reg_u0 ( .ck(ispd_clk), .d(n_2946), .o(pci_target_unit_pci_target_sm_cnf_progress) );
ms00f80 pci_target_unit_pci_target_sm_master_will_request_read_reg_u0 ( .ck(ispd_clk), .d(n_8528), .o(pci_target_unit_pci_target_sm_master_will_request_read) );
ms00f80 pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg_u0 ( .ck(ispd_clk), .d(n_8574), .o(n_2314) );
ms00f80 pci_target_unit_pci_target_sm_previous_frame_reg_u0 ( .ck(ispd_clk), .d(n_15302), .o(pci_target_unit_pci_target_sm_previous_frame) );
ms00f80 pci_target_unit_pci_target_sm_rd_from_fifo_reg_u0 ( .ck(ispd_clk), .d(n_3364), .o(pci_target_unit_pci_target_sm_rd_from_fifo) );
ms00f80 pci_target_unit_pci_target_sm_rd_progress_reg_u0 ( .ck(ispd_clk), .d(n_8688), .o(pci_target_unit_pci_target_sm_rd_progress) );
ms00f80 pci_target_unit_pci_target_sm_rd_request_reg_u0 ( .ck(ispd_clk), .d(n_8687), .o(pci_target_unit_pci_target_sm_rd_request_reg_Q) );
in01s01 pci_target_unit_pci_target_sm_rd_request_reg_u1 ( .a(pci_target_unit_pci_target_sm_rd_request_reg_Q), .o(pci_target_unit_pci_target_sm_rd_request) );
ms00f80 pci_target_unit_pci_target_sm_read_completed_reg_reg_u0 ( .ck(ispd_clk), .d(n_2337), .o(pci_target_unit_pci_target_sm_read_completed_reg_reg_Q) );
in01f10 pci_target_unit_pci_target_sm_read_completed_reg_reg_u1 ( .a(pci_target_unit_pci_target_sm_read_completed_reg_reg_Q), .o(pci_target_unit_pci_target_sm_read_completed_reg) );
ms00f80 pci_target_unit_pci_target_sm_rw_cbe0_reg_u0 ( .ck(ispd_clk), .d(n_3219), .o(n_978) );
ms00f80 pci_target_unit_pci_target_sm_same_read_reg_reg_u0 ( .ck(ispd_clk), .d(n_4895), .o(pci_target_unit_pci_target_sm_same_read_reg) );
ms00f80 pci_target_unit_pci_target_sm_state_backoff_reg_reg_u0 ( .ck(ispd_clk), .d(n_2140), .o(pci_target_unit_pci_target_sm_state_backoff_reg_reg_Q) );
ms00f80 pci_target_unit_pci_target_sm_state_transfere_reg_reg_u0 ( .ck(ispd_clk), .d(n_13817), .o(pci_target_unit_pci_target_sm_state_transfere_reg_reg_Q) );
in01s10 pci_target_unit_pci_target_sm_state_transfere_reg_reg_u1 ( .a(pci_target_unit_pci_target_sm_state_transfere_reg_reg_Q), .o(pci_target_unit_pci_target_sm_state_transfere_reg) );
ms00f80 pci_target_unit_pci_target_sm_wr_progress_reg_u0 ( .ck(ispd_clk), .d(n_8573), .o(pci_target_unit_pci_target_sm_wr_progress) );
ms00f80 pci_target_unit_pci_target_sm_wr_to_fifo_reg_u0 ( .ck(ispd_clk), .d(n_3499), .o(pci_target_unit_pci_target_sm_wr_to_fifo) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_0__u0 ( .ck(ispd_clk), .d(n_14804), .o(wbm_adr_o_0_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_10__u0 ( .ck(ispd_clk), .d(n_14813), .o(wbm_adr_o_10_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_11__u0 ( .ck(ispd_clk), .d(n_14812), .o(wbm_adr_o_11_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_12__u0 ( .ck(ispd_clk), .d(n_14811), .o(wbm_adr_o_12_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_13__u0 ( .ck(ispd_clk), .d(n_14810), .o(wbm_adr_o_13_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_14__u0 ( .ck(ispd_clk), .d(n_14847), .o(wbm_adr_o_14_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_15__u0 ( .ck(ispd_clk), .d(n_14808), .o(wbm_adr_o_15_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_16__u0 ( .ck(ispd_clk), .d(n_14848), .o(wbm_adr_o_16_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_17__u0 ( .ck(ispd_clk), .d(n_14828), .o(wbm_adr_o_17_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_18__u0 ( .ck(ispd_clk), .d(n_14803), .o(wbm_adr_o_18_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_19__u0 ( .ck(ispd_clk), .d(n_14826), .o(wbm_adr_o_19_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_1__u0 ( .ck(ispd_clk), .d(n_14805), .o(wbm_adr_o_1_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_20__u0 ( .ck(ispd_clk), .d(n_14825), .o(wbm_adr_o_20_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_21__u0 ( .ck(ispd_clk), .d(n_14818), .o(wbm_adr_o_21_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_22__u0 ( .ck(ispd_clk), .d(n_14824), .o(wbm_adr_o_22_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_23__u0 ( .ck(ispd_clk), .d(n_14846), .o(wbm_adr_o_23_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_24__u0 ( .ck(ispd_clk), .d(n_14822), .o(wbm_adr_o_24_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_25__u0 ( .ck(ispd_clk), .d(n_14821), .o(wbm_adr_o_25_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_26__u0 ( .ck(ispd_clk), .d(n_14845), .o(wbm_adr_o_26_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_27__u0 ( .ck(ispd_clk), .d(n_14819), .o(wbm_adr_o_27_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_28__u0 ( .ck(ispd_clk), .d(n_14815), .o(wbm_adr_o_28_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_29__u0 ( .ck(ispd_clk), .d(n_14817), .o(wbm_adr_o_29_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_2__u0 ( .ck(ispd_clk), .d(n_14844), .o(wbm_adr_o_2_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_30__u0 ( .ck(ispd_clk), .d(n_14816), .o(wbm_adr_o_30_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_31__u0 ( .ck(ispd_clk), .d(n_14814), .o(wbm_adr_o_31_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_3__u0 ( .ck(ispd_clk), .d(n_14842), .o(wbm_adr_o_3_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_4__u0 ( .ck(ispd_clk), .d(n_14841), .o(wbm_adr_o_4_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_5__u0 ( .ck(ispd_clk), .d(n_14840), .o(wbm_adr_o_5_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_6__u0 ( .ck(ispd_clk), .d(n_14838), .o(wbm_adr_o_6_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_7__u0 ( .ck(ispd_clk), .d(n_14807), .o(wbm_adr_o_7_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_8__u0 ( .ck(ispd_clk), .d(n_14836), .o(wbm_adr_o_8_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_9__u0 ( .ck(ispd_clk), .d(n_14834), .o(wbm_adr_o_9_) );
ms00f80 pci_target_unit_wishbone_master_addr_into_cnt_reg_reg_u0 ( .ck(ispd_clk), .d(n_8757), .o(pci_target_unit_wishbone_master_addr_into_cnt_reg) );
ms00f80 pci_target_unit_wishbone_master_bc_register_reg_0__u0 ( .ck(ispd_clk), .d(n_14687), .o(pci_target_unit_wishbone_master_bc_register_reg_0__Q) );
ms00f80 pci_target_unit_wishbone_master_bc_register_reg_1__u0 ( .ck(ispd_clk), .d(n_14686), .o(pci_target_unit_wishbone_master_bc_register_reg_1__Q) );
ms00f80 pci_target_unit_wishbone_master_bc_register_reg_2__u0 ( .ck(ispd_clk), .d(n_14685), .o(pci_target_unit_wishbone_master_bc_register_reg_2__Q) );
ms00f80 pci_target_unit_wishbone_master_bc_register_reg_3__u0 ( .ck(ispd_clk), .d(n_14683), .o(pci_target_unit_wishbone_master_bc_register_reg_3__Q) );
ms00f80 pci_target_unit_wishbone_master_burst_chopped_delayed_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_wishbone_master_burst_chopped), .o(pci_target_unit_wishbone_master_burst_chopped_delayed_reg_Q) );
in01f20 pci_target_unit_wishbone_master_burst_chopped_delayed_reg_u1 ( .a(pci_target_unit_wishbone_master_burst_chopped_delayed_reg_Q), .o(pci_target_unit_wishbone_master_burst_chopped_delayed) );
ms00f80 pci_target_unit_wishbone_master_burst_chopped_reg_u0 ( .ck(ispd_clk), .d(n_14694), .o(pci_target_unit_wishbone_master_burst_chopped) );
ms00f80 pci_target_unit_wishbone_master_c_state_reg_0__u0 ( .ck(ispd_clk), .d(n_16167), .o(pci_target_unit_wishbone_master_c_state_0_) );
ms00f80 pci_target_unit_wishbone_master_c_state_reg_1__u0 ( .ck(ispd_clk), .d(n_8452), .o(pci_target_unit_wishbone_master_c_state_1_) );
ms00f80 pci_target_unit_wishbone_master_c_state_reg_2__u0 ( .ck(ispd_clk), .d(n_15188), .o(pci_target_unit_wishbone_master_c_state_2_) );
ms00f80 pci_target_unit_wishbone_master_first_data_is_burst_reg_reg_u0 ( .ck(ispd_clk), .d(n_10787), .o(pci_target_unit_wishbone_master_first_data_is_burst_reg) );
ms00f80 pci_target_unit_wishbone_master_first_wb_data_access_reg_u0 ( .ck(ispd_clk), .d(n_13789), .o(pci_target_unit_wishbone_master_first_wb_data_access) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_control_out_reg_1__u0 ( .ck(ispd_clk), .d(n_3223), .o(pci_target_unit_fifos_pcir_control_in_192) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_0__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15207), .o(pci_target_unit_fifos_pcir_data_in) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_10__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15209), .o(pci_target_unit_fifos_pcir_data_in_167) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_11__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15211), .o(pci_target_unit_fifos_pcir_data_in_168) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_12__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15213), .o(pci_target_unit_fifos_pcir_data_in_169) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_13__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15215), .o(pci_target_unit_fifos_pcir_data_in_170) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_14__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15217), .o(pci_target_unit_fifos_pcir_data_in_171) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_15__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15219), .o(pci_target_unit_fifos_pcir_data_in_172) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_16__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15221), .o(pci_target_unit_fifos_pcir_data_in_173) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_17__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15223), .o(pci_target_unit_fifos_pcir_data_in_174) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_18__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15225), .o(pci_target_unit_fifos_pcir_data_in_175) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_19__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15227), .o(pci_target_unit_fifos_pcir_data_in_176) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_1__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15229), .o(pci_target_unit_fifos_pcir_data_in_158) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_20__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15231), .o(pci_target_unit_fifos_pcir_data_in_177) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_21__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15233), .o(pci_target_unit_fifos_pcir_data_in_178) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_22__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15235), .o(pci_target_unit_fifos_pcir_data_in_179) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_23__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15237), .o(pci_target_unit_fifos_pcir_data_in_180) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_24__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15239), .o(pci_target_unit_fifos_pcir_data_in_181) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_25__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15241), .o(pci_target_unit_fifos_pcir_data_in_182) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_26__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15243), .o(pci_target_unit_fifos_pcir_data_in_183) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_27__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15245), .o(pci_target_unit_fifos_pcir_data_in_184) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_28__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15247), .o(pci_target_unit_fifos_pcir_data_in_185) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_29__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15249), .o(pci_target_unit_fifos_pcir_data_in_186) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_2__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15251), .o(pci_target_unit_fifos_pcir_data_in_159) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_30__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15253), .o(pci_target_unit_fifos_pcir_data_in_187) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_31__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15255), .o(pci_target_unit_fifos_pcir_data_in_188) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_3__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15257), .o(pci_target_unit_fifos_pcir_data_in_160) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_4__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15259), .o(pci_target_unit_fifos_pcir_data_in_161) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_5__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15261), .o(pci_target_unit_fifos_pcir_data_in_162) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_6__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15263), .o(pci_target_unit_fifos_pcir_data_in_163) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_7__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15265), .o(pci_target_unit_fifos_pcir_data_in_164) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_8__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15267), .o(pci_target_unit_fifos_pcir_data_in_165) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_9__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_15269), .o(pci_target_unit_fifos_pcir_data_in_166) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_wenable_out_reg_u0 ( .ck(ispd_clk), .d(n_3224), .o(pci_target_unit_fifos_pcir_wenable_in) );
ms00f80 pci_target_unit_wishbone_master_read_bound_reg_u0 ( .ck(ispd_clk), .d(n_7401), .o(pci_target_unit_wishbone_master_read_bound) );
ms00f80 pci_target_unit_wishbone_master_read_count_reg_0__u0 ( .ck(ispd_clk), .d(n_7575), .o(pci_target_unit_wishbone_master_read_count_0_) );
ms00f80 pci_target_unit_wishbone_master_read_count_reg_1__u0 ( .ck(ispd_clk), .d(n_7609), .o(pci_target_unit_wishbone_master_read_count_1_) );
ms00f80 pci_target_unit_wishbone_master_read_count_reg_2__u0 ( .ck(ispd_clk), .d(n_7791), .o(pci_target_unit_wishbone_master_read_count_reg_2__Q) );
ms00f80 pci_target_unit_wishbone_master_reset_rty_cnt_reg_u0 ( .ck(ispd_clk), .d(n_8494), .o(pci_target_unit_wishbone_master_reset_rty_cnt_reg_Q) );
in01s01 pci_target_unit_wishbone_master_reset_rty_cnt_reg_u1 ( .a(pci_target_unit_wishbone_master_reset_rty_cnt_reg_Q), .o(pci_target_unit_wishbone_master_reset_rty_cnt) );
ms00f80 pci_target_unit_wishbone_master_retried_reg_u0 ( .ck(ispd_clk), .d(n_3268), .o(pci_target_unit_wishbone_master_retried) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_0__u0 ( .ck(ispd_clk), .d(n_8818), .o(pci_target_unit_wishbone_master_rty_counter_0_) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_1__u0 ( .ck(ispd_clk), .d(n_8721), .o(pci_target_unit_wishbone_master_rty_counter_1_) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_2__u0 ( .ck(ispd_clk), .d(n_8726), .o(n_1263) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_3__u0 ( .ck(ispd_clk), .d(n_8725), .o(pci_target_unit_wishbone_master_rty_counter_3_) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_4__u0 ( .ck(ispd_clk), .d(n_8724), .o(pci_target_unit_wishbone_master_rty_counter_4_) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_5__u0 ( .ck(ispd_clk), .d(n_8734), .o(pci_target_unit_wishbone_master_rty_counter_5_) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_6__u0 ( .ck(ispd_clk), .d(n_8733), .o(pci_target_unit_wishbone_master_rty_counter_6_) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_7__u0 ( .ck(ispd_clk), .d(n_8731), .o(pci_target_unit_wishbone_master_rty_counter_7_) );
ms00f80 pci_target_unit_wishbone_master_w_attempt_reg_u0 ( .ck(ispd_clk), .d(n_8565), .o(n_16501) );
ms00f80 pci_target_unit_wishbone_master_wb_cti_o_reg_0__u0 ( .ck(ispd_clk), .d(n_14904), .o(wbm_cti_o_0_) );
ms00f80 pci_target_unit_wishbone_master_wb_cti_o_reg_1__u0 ( .ck(ispd_clk), .d(n_14629), .o(wbm_cti_o_1_) );
ms00f80 pci_target_unit_wishbone_master_wb_cti_o_reg_2__u0 ( .ck(ispd_clk), .d(n_14903), .o(wbm_cti_o_2_) );
ms00f80 pci_target_unit_wishbone_master_wb_cyc_o_reg_u0 ( .ck(ispd_clk), .d(n_13624), .o(pci_target_unit_wishbone_master_wb_cyc_o_reg_Q) );
in01s10 pci_target_unit_wishbone_master_wb_cyc_o_reg_u1 ( .a(pci_target_unit_wishbone_master_wb_cyc_o_reg_Q), .o(wbm_cyc_o_1378) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_0__u0 ( .ck(ispd_clk), .d(n_14887), .o(wbm_dat_o_0_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_10__u0 ( .ck(ispd_clk), .d(n_15197), .o(wbm_dat_o_10_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_11__u0 ( .ck(ispd_clk), .d(n_14885), .o(wbm_dat_o_11_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_12__u0 ( .ck(ispd_clk), .d(n_14884), .o(wbm_dat_o_12_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_13__u0 ( .ck(ispd_clk), .d(n_14883), .o(wbm_dat_o_13_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_14__u0 ( .ck(ispd_clk), .d(n_14881), .o(wbm_dat_o_14_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_15__u0 ( .ck(ispd_clk), .d(n_14851), .o(wbm_dat_o_15_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_16__u0 ( .ck(ispd_clk), .d(n_14879), .o(wbm_dat_o_16_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_17__u0 ( .ck(ispd_clk), .d(n_14880), .o(wbm_dat_o_17_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_18__u0 ( .ck(ispd_clk), .d(n_14850), .o(wbm_dat_o_18_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_19__u0 ( .ck(ispd_clk), .d(n_14877), .o(wbm_dat_o_19_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_1__u0 ( .ck(ispd_clk), .d(n_14875), .o(wbm_dat_o_1_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_20__u0 ( .ck(ispd_clk), .d(n_14873), .o(wbm_dat_o_20_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_21__u0 ( .ck(ispd_clk), .d(n_14871), .o(wbm_dat_o_21_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_22__u0 ( .ck(ispd_clk), .d(n_16304), .o(wbm_dat_o_22_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_23__u0 ( .ck(ispd_clk), .d(n_14869), .o(wbm_dat_o_23_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_24__u0 ( .ck(ispd_clk), .d(n_14867), .o(wbm_dat_o_24_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_25__u0 ( .ck(ispd_clk), .d(n_14866), .o(wbm_dat_o_25_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_26__u0 ( .ck(ispd_clk), .d(n_14865), .o(wbm_dat_o_26_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_27__u0 ( .ck(ispd_clk), .d(n_14863), .o(wbm_dat_o_27_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_28__u0 ( .ck(ispd_clk), .d(n_14864), .o(wbm_dat_o_28_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_29__u0 ( .ck(ispd_clk), .d(n_14862), .o(wbm_dat_o_29_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_2__u0 ( .ck(ispd_clk), .d(n_14861), .o(wbm_dat_o_2_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_30__u0 ( .ck(ispd_clk), .d(n_14860), .o(wbm_dat_o_30_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_31__u0 ( .ck(ispd_clk), .d(n_14856), .o(wbm_dat_o_31_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_3__u0 ( .ck(ispd_clk), .d(n_14859), .o(wbm_dat_o_3_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_4__u0 ( .ck(ispd_clk), .d(n_14858), .o(wbm_dat_o_4_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_5__u0 ( .ck(ispd_clk), .d(n_14855), .o(wbm_dat_o_5_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_6__u0 ( .ck(ispd_clk), .d(n_14854), .o(wbm_dat_o_6_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_7__u0 ( .ck(ispd_clk), .d(n_14849), .o(wbm_dat_o_7_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_8__u0 ( .ck(ispd_clk), .d(n_14853), .o(wbm_dat_o_8_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_9__u0 ( .ck(ispd_clk), .d(n_14852), .o(wbm_dat_o_9_) );
ms00f80 pci_target_unit_wishbone_master_wb_read_done_out_reg_u0 ( .ck(ispd_clk), .d(n_4896), .o(pci_target_unit_del_sync_comp_in) );
ms00f80 pci_target_unit_wishbone_master_wb_sel_o_reg_0__u0 ( .ck(ispd_clk), .d(n_14897), .o(wbm_sel_o_0_) );
ms00f80 pci_target_unit_wishbone_master_wb_sel_o_reg_1__u0 ( .ck(ispd_clk), .d(n_14894), .o(wbm_sel_o_1_) );
ms00f80 pci_target_unit_wishbone_master_wb_sel_o_reg_2__u0 ( .ck(ispd_clk), .d(n_14896), .o(wbm_sel_o_2_) );
ms00f80 pci_target_unit_wishbone_master_wb_sel_o_reg_3__u0 ( .ck(ispd_clk), .d(n_14893), .o(wbm_sel_o_3_) );
ms00f80 pci_target_unit_wishbone_master_wb_stb_o_reg_u0 ( .ck(ispd_clk), .d(n_13624), .o(wbm_stb_o) );
ms00f80 pci_target_unit_wishbone_master_wb_we_o_reg_u0 ( .ck(ispd_clk), .d(n_13481), .o(wbm_we_o) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_0__u0 ( .ck(ispd_clk), .d(n_9402), .o(wishbone_slave_unit_del_sync_addr_out_reg_0__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_10__u0 ( .ck(ispd_clk), .d(n_9400), .o(wishbone_slave_unit_del_sync_addr_out_reg_10__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_11__u0 ( .ck(ispd_clk), .d(n_9398), .o(wishbone_slave_unit_del_sync_addr_out_reg_11__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_12__u0 ( .ck(ispd_clk), .d(n_8989), .o(wishbone_slave_unit_del_sync_addr_out_reg_12__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_13__u0 ( .ck(ispd_clk), .d(n_9396), .o(wishbone_slave_unit_del_sync_addr_out_reg_13__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_14__u0 ( .ck(ispd_clk), .d(n_8986), .o(wishbone_slave_unit_del_sync_addr_out_reg_14__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_15__u0 ( .ck(ispd_clk), .d(n_9393), .o(wishbone_slave_unit_del_sync_addr_out_reg_15__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_16__u0 ( .ck(ispd_clk), .d(n_9391), .o(wishbone_slave_unit_del_sync_addr_out_reg_16__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_17__u0 ( .ck(ispd_clk), .d(n_9389), .o(wishbone_slave_unit_del_sync_addr_out_reg_17__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_18__u0 ( .ck(ispd_clk), .d(n_9387), .o(wishbone_slave_unit_del_sync_addr_out_reg_18__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_19__u0 ( .ck(ispd_clk), .d(n_9385), .o(wishbone_slave_unit_del_sync_addr_out_reg_19__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_1__u0 ( .ck(ispd_clk), .d(n_9383), .o(wishbone_slave_unit_del_sync_addr_out_reg_1__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_20__u0 ( .ck(ispd_clk), .d(n_9381), .o(wishbone_slave_unit_del_sync_addr_out_reg_20__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_21__u0 ( .ck(ispd_clk), .d(n_9379), .o(wishbone_slave_unit_del_sync_addr_out_reg_21__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_22__u0 ( .ck(ispd_clk), .d(n_8983), .o(wishbone_slave_unit_del_sync_addr_out_reg_22__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_23__u0 ( .ck(ispd_clk), .d(n_9377), .o(wishbone_slave_unit_del_sync_addr_out_reg_23__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_24__u0 ( .ck(ispd_clk), .d(n_9374), .o(wishbone_slave_unit_del_sync_addr_out_reg_24__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_25__u0 ( .ck(ispd_clk), .d(n_8981), .o(wishbone_slave_unit_del_sync_addr_out_reg_25__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_26__u0 ( .ck(ispd_clk), .d(n_9371), .o(wishbone_slave_unit_del_sync_addr_out_reg_26__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_27__u0 ( .ck(ispd_clk), .d(n_9368), .o(wishbone_slave_unit_del_sync_addr_out_reg_27__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_28__u0 ( .ck(ispd_clk), .d(n_9366), .o(wishbone_slave_unit_del_sync_addr_out_reg_28__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_29__u0 ( .ck(ispd_clk), .d(n_9363), .o(wishbone_slave_unit_del_sync_addr_out_reg_29__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_2__u0 ( .ck(ispd_clk), .d(n_8979), .o(wishbone_slave_unit_del_sync_addr_out_reg_2__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_30__u0 ( .ck(ispd_clk), .d(n_9361), .o(wishbone_slave_unit_del_sync_addr_out_reg_30__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_31__u0 ( .ck(ispd_clk), .d(n_9358), .o(wishbone_slave_unit_del_sync_addr_out_reg_31__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_3__u0 ( .ck(ispd_clk), .d(n_9355), .o(wishbone_slave_unit_del_sync_addr_out_reg_3__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_4__u0 ( .ck(ispd_clk), .d(n_8977), .o(wishbone_slave_unit_del_sync_addr_out_reg_4__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_5__u0 ( .ck(ispd_clk), .d(n_8975), .o(wishbone_slave_unit_del_sync_addr_out_reg_5__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_6__u0 ( .ck(ispd_clk), .d(n_8973), .o(wishbone_slave_unit_del_sync_addr_out_reg_6__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_7__u0 ( .ck(ispd_clk), .d(n_9353), .o(wishbone_slave_unit_del_sync_addr_out_reg_7__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_8__u0 ( .ck(ispd_clk), .d(n_9350), .o(wishbone_slave_unit_del_sync_addr_out_reg_8__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_9__u0 ( .ck(ispd_clk), .d(n_9348), .o(wishbone_slave_unit_del_sync_addr_out_reg_9__Q) );
ms00f80 wishbone_slave_unit_del_sync_bc_out_reg_0__u0 ( .ck(ispd_clk), .d(n_8598), .o(wishbone_slave_unit_del_sync_bc_out_reg_0__Q) );
in01s02 wishbone_slave_unit_del_sync_bc_out_reg_0__u1 ( .a(wishbone_slave_unit_del_sync_bc_out_reg_0__Q), .o(wishbone_slave_unit_pcim_if_del_bc_in) );
ms00f80 wishbone_slave_unit_del_sync_bc_out_reg_1__u0 ( .ck(ispd_clk), .d(n_8677), .o(wishbone_slave_unit_del_sync_bc_out_reg_1__Q) );
ms00f80 wishbone_slave_unit_del_sync_bc_out_reg_2__u0 ( .ck(ispd_clk), .d(n_8723), .o(wishbone_slave_unit_del_sync_bc_out_reg_2__Q) );
in01s01 wishbone_slave_unit_del_sync_bc_out_reg_2__u1 ( .a(wishbone_slave_unit_del_sync_bc_out_reg_2__Q), .o(wishbone_slave_unit_pcim_if_del_bc_in_382) );
ms00f80 wishbone_slave_unit_del_sync_bc_out_reg_3__u0 ( .ck(ispd_clk), .d(n_8796), .o(wishbone_slave_unit_del_sync_bc_out_reg_3__Q) );
in01s01 wishbone_slave_unit_del_sync_bc_out_reg_3__u1 ( .a(wishbone_slave_unit_del_sync_bc_out_reg_3__Q), .o(wishbone_slave_unit_pcim_if_del_bc_in_383) );
ms00f80 wishbone_slave_unit_del_sync_be_out_reg_0__u0 ( .ck(ispd_clk), .d(n_8676), .o(wishbone_slave_unit_fifos_wbr_be_in) );
ms00f80 wishbone_slave_unit_del_sync_be_out_reg_1__u0 ( .ck(ispd_clk), .d(n_8675), .o(wishbone_slave_unit_fifos_wbr_be_in_264) );
ms00f80 wishbone_slave_unit_del_sync_be_out_reg_2__u0 ( .ck(ispd_clk), .d(n_8674), .o(wishbone_slave_unit_fifos_wbr_be_in_265) );
ms00f80 wishbone_slave_unit_del_sync_be_out_reg_3__u0 ( .ck(ispd_clk), .d(n_8673), .o(wishbone_slave_unit_fifos_wbr_be_in_266) );
ms00f80 wishbone_slave_unit_del_sync_burst_out_reg_u0 ( .ck(ispd_clk), .d(n_8843), .o(wishbone_slave_unit_pcim_if_del_burst_in) );
ms00f80 wishbone_slave_unit_del_sync_comp_comp_pending_reg_u0 ( .ck(ispd_clk), .d(n_8496), .o(wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_0__u0 ( .ck(ispd_clk), .d(n_8652), .o(wishbone_slave_unit_del_sync_comp_cycle_count_0_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_10__u0 ( .ck(ispd_clk), .d(n_8656), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_10__Q) );
in01s06 wishbone_slave_unit_del_sync_comp_cycle_count_reg_10__u1 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_10__Q), .o(wishbone_slave_unit_del_sync_comp_cycle_count_10_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_11__u0 ( .ck(ispd_clk), .d(n_8651), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_11__Q) );
in01m01 wishbone_slave_unit_del_sync_comp_cycle_count_reg_11__u1 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_11__Q), .o(wishbone_slave_unit_del_sync_comp_cycle_count_11_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_12__u0 ( .ck(ispd_clk), .d(n_8662), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_12__Q) );
in01s01 wishbone_slave_unit_del_sync_comp_cycle_count_reg_12__u1 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_12__Q), .o(wishbone_slave_unit_del_sync_comp_cycle_count_12_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__u0 ( .ck(ispd_clk), .d(n_8650), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__u0 ( .ck(ispd_clk), .d(n_8649), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__u0 ( .ck(ispd_clk), .d(n_8648), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__Q) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__u0 ( .ck(ispd_clk), .d(n_8579), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_1__u0 ( .ck(ispd_clk), .d(n_8658), .o(wishbone_slave_unit_del_sync_comp_cycle_count_1_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_2__u0 ( .ck(ispd_clk), .d(n_8647), .o(wishbone_slave_unit_del_sync_comp_cycle_count_2_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_3__u0 ( .ck(ispd_clk), .d(n_8646), .o(wishbone_slave_unit_del_sync_comp_cycle_count_3_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_4__u0 ( .ck(ispd_clk), .d(n_8645), .o(wishbone_slave_unit_del_sync_comp_cycle_count_4_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_5__u0 ( .ck(ispd_clk), .d(n_8644), .o(wishbone_slave_unit_del_sync_comp_cycle_count_5_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_6__u0 ( .ck(ispd_clk), .d(n_8643), .o(wishbone_slave_unit_del_sync_comp_cycle_count_6_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_7__u0 ( .ck(ispd_clk), .d(n_8642), .o(wishbone_slave_unit_del_sync_comp_cycle_count_7_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_8__u0 ( .ck(ispd_clk), .d(n_8661), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_8__Q) );
in01s06 wishbone_slave_unit_del_sync_comp_cycle_count_reg_8__u1 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_8__Q), .o(wishbone_slave_unit_del_sync_comp_cycle_count_8_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_9__u0 ( .ck(ispd_clk), .d(n_8655), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_9__Q) );
in01s06 wishbone_slave_unit_del_sync_comp_cycle_count_reg_9__u1 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_9__Q), .o(wishbone_slave_unit_del_sync_comp_cycle_count_9_) );
ms00f80 wishbone_slave_unit_del_sync_comp_done_reg_clr_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_comp_done_reg_main), .o(wishbone_slave_unit_del_sync_comp_done_reg_clr_reg_Q) );
in01s01 wishbone_slave_unit_del_sync_comp_done_reg_clr_reg_u1 ( .a(wishbone_slave_unit_del_sync_comp_done_reg_clr_reg_Q), .o(wishbone_slave_unit_del_sync_comp_done_reg_clr) );
ms00f80 wishbone_slave_unit_del_sync_comp_done_reg_main_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_sync_comp_done), .o(wishbone_slave_unit_del_sync_comp_done_reg_main) );
ms00f80 wishbone_slave_unit_del_sync_comp_flush_out_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q), .o(wishbone_slave_unit_del_sync_comp_flush_out) );
ms00f80 wishbone_slave_unit_del_sync_comp_req_pending_reg_u0 ( .ck(ispd_clk), .d(n_7716), .o(wishbone_slave_unit_del_sync_comp_req_pending_reg_Q) );
in01s06 wishbone_slave_unit_del_sync_comp_req_pending_reg_u1 ( .a(wishbone_slave_unit_del_sync_comp_req_pending_reg_Q), .o(wishbone_slave_unit_pcim_if_del_req_in) );
ms00f80 wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_sync_comp_rty_exp_clr), .o(wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg_Q) );
in01s01 wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg_u1 ( .a(wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg_Q), .o(wishbone_slave_unit_del_sync_comp_rty_exp_clr) );
ms00f80 wishbone_slave_unit_del_sync_comp_rty_exp_reg_reg_u0 ( .ck(ispd_clk), .d(n_4140), .o(wishbone_slave_unit_del_sync_comp_rty_exp_reg) );
ms00f80 wishbone_slave_unit_del_sync_comp_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q), .o(TIMEBOOST_net_15173) );
ms00f80 wishbone_slave_unit_del_sync_done_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_325), .o(wishbone_slave_unit_del_sync_sync_comp_done) );
ms00f80 wishbone_slave_unit_del_sync_req_comp_pending_reg_u0 ( .ck(ispd_clk), .d(n_14621), .o(wishbone_slave_unit_del_sync_req_comp_pending) );
ms00f80 wishbone_slave_unit_del_sync_req_comp_pending_sample_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_sync_req_comp_pending), .o(wishbone_slave_unit_del_sync_req_comp_pending_sample_reg_Q) );
in01s01 wishbone_slave_unit_del_sync_req_comp_pending_sample_reg_u1 ( .a(wishbone_slave_unit_del_sync_req_comp_pending_sample_reg_Q), .o(wishbone_slave_unit_del_sync_req_comp_pending_sample) );
ms00f80 wishbone_slave_unit_del_sync_req_done_reg_reg_u0 ( .ck(ispd_clk), .d(n_14623), .o(wishbone_slave_unit_del_sync_req_done_reg_reg_Q) );
in01s01 wishbone_slave_unit_del_sync_req_done_reg_reg_u1 ( .a(wishbone_slave_unit_del_sync_req_done_reg_reg_Q), .o(wishbone_slave_unit_del_sync_req_done_reg) );
ms00f80 wishbone_slave_unit_del_sync_req_req_pending_reg_u0 ( .ck(ispd_clk), .d(n_8495), .o(wishbone_slave_unit_wbs_sm_del_req_pending_in) );
ms00f80 wishbone_slave_unit_del_sync_req_rty_exp_clr_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_req_rty_exp_reg), .o(wishbone_slave_unit_del_sync_req_rty_exp_clr_reg_Q) );
in01s01 wishbone_slave_unit_del_sync_req_rty_exp_clr_reg_u1 ( .a(wishbone_slave_unit_del_sync_req_rty_exp_clr_reg_Q), .o(wishbone_slave_unit_del_sync_req_rty_exp_clr) );
ms00f80 wishbone_slave_unit_del_sync_req_rty_exp_reg_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_sync_req_rty_exp), .o(wishbone_slave_unit_del_sync_req_rty_exp_reg) );
ms00f80 wishbone_slave_unit_del_sync_req_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_wbs_sm_del_req_pending_in), .o(wishbone_slave_unit_del_sync_sync_comp_req_pending) );
ms00f80 wishbone_slave_unit_del_sync_rty_exp_back_prop_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_2386), .o(wishbone_slave_unit_del_sync_sync_comp_rty_exp_clr) );
ms00f80 wishbone_slave_unit_del_sync_rty_exp_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_comp_rty_exp_reg), .o(wishbone_slave_unit_del_sync_sync_req_rty_exp) );
ms00f80 wishbone_slave_unit_del_sync_we_out_reg_u0 ( .ck(ispd_clk), .d(n_8672), .o(wishbone_slave_unit_del_sync_we_out_reg_Q) );
in01s10 wishbone_slave_unit_del_sync_we_out_reg_u1 ( .a(wishbone_slave_unit_del_sync_we_out_reg_Q), .o(wishbone_slave_unit_pcim_if_del_we_in) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_70), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_70) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_10__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_80), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_80) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_11__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_81), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_81) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_12__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_82), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_82) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_13__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_83), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_83) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_14__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_84), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_84) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_15__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_85), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_85) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_16__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_86), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_86) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_17__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_87), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_87) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_18__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_88), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_88) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_19__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_89), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_89) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_71), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_71) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_20__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_90), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_90) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_21__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_91), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_91) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_22__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_92), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_92) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_23__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_93), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_93) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_24__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_94), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_94) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_25__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_95), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_95) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_26__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_96), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_96) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_27__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_97), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_97) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_28__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_98), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_98) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_29__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_99), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_99) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_72), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_72) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_30__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_100), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_100) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_31__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_101), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_101) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_73), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_73) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_4__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_74), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_74) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_5__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_75), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_75) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_6__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_76), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_76) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_7__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_77), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_77) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_8__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_78), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_78) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_9__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_79), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_79) );
ms00f80 wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_22), .o(wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount) );
ms00f80 wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_inGreyCount_reg_1__Q), .o(wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_49) );
ms00f80 wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_inGreyCount_reg_2__Q), .o(wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_50) );
ms00f80 wishbone_slave_unit_fifos_inGreyCount_reg_0__u0 ( .ck(ispd_clk), .d(n_9145), .o(wishbone_slave_unit_fifos_inGreyCount_reg_0__Q) );
in01s01 wishbone_slave_unit_fifos_inGreyCount_reg_0__u1 ( .a(wishbone_slave_unit_fifos_inGreyCount_reg_0__Q), .o(wishbone_slave_unit_fifos_inGreyCount_0_) );
ms00f80 wishbone_slave_unit_fifos_inGreyCount_reg_1__u0 ( .ck(ispd_clk), .d(n_8920), .o(wishbone_slave_unit_fifos_inGreyCount_reg_1__Q) );
ms00f80 wishbone_slave_unit_fifos_inGreyCount_reg_2__u0 ( .ck(ispd_clk), .d(n_8919), .o(wishbone_slave_unit_fifos_inGreyCount_reg_2__Q) );
ms00f80 wishbone_slave_unit_fifos_outGreyCount_reg_0__u0 ( .ck(ispd_clk), .d(n_8717), .o(wishbone_slave_unit_fifos_outGreyCount_0_) );
ms00f80 wishbone_slave_unit_fifos_outGreyCount_reg_1__u0 ( .ck(ispd_clk), .d(n_8589), .o(wishbone_slave_unit_fifos_outGreyCount_1_) );
ms00f80 wishbone_slave_unit_fifos_outGreyCount_reg_2__u0 ( .ck(ispd_clk), .d(n_8585), .o(wishbone_slave_unit_fifos_outGreyCount_2_) );
ms00f80 wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount), .o(wishbone_slave_unit_fifos_pci_clk_inGreyCount_0_) );
ms00f80 wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_49), .o(wishbone_slave_unit_fifos_pci_clk_inGreyCount_1_) );
ms00f80 wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_50), .o(wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_2__Q) );
in01f20 wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_2__u1 ( .a(wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_2__Q), .o(wishbone_slave_unit_fifos_pci_clk_inGreyCount_2_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_276), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_45) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_46) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_47) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_0__u0 ( .ck(ispd_clk), .d(n_9942), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_0__Q) );
in01s20 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_0__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_1__u0 ( .ck(ispd_clk), .d(n_9238), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_1__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_1__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_1__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_1_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_2__u0 ( .ck(ispd_clk), .d(n_9239), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_2__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_2__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_2__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_3__u0 ( .ck(ispd_clk), .d(n_9241), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_3__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_3__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_3__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_3_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_0__u0 ( .ck(ispd_clk), .d(n_9947), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_0__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_0__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_0__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_0_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_1__u0 ( .ck(ispd_clk), .d(n_9932), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_1__Q) );
in01m06 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_1__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_1__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_1_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_2__u0 ( .ck(ispd_clk), .d(n_9931), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_2__Q) );
in01s20 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_2__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_2__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__u0 ( .ck(ispd_clk), .d(n_9154), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_0__Q) );
in01f40 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_0__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_0__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_0_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_45), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_1__Q) );
in01f40 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_1__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_1__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_1_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_46), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_2__Q) );
in01f40 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_2__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_2__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_2_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_47), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_3__Q) );
in01f40 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_3__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_3__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_3_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_9237), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_0_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_9236), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_1_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_9235), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_2_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg_3__u0 ( .ck(ispd_clk), .d(n_9234), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_3_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg_0__u0 ( .ck(ispd_clk), .d(n_6112), .o(wishbone_slave_unit_fifos_wbr_whole_waddr) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg_1__u0 ( .ck(ispd_clk), .d(n_7393), .o(wishbone_slave_unit_fifos_wbr_whole_waddr_104) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg_2__u0 ( .ck(ispd_clk), .d(n_5770), .o(wishbone_slave_unit_fifos_wbr_whole_waddr_105) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg_3__u0 ( .ck(ispd_clk), .d(n_6138), .o(wishbone_slave_unit_fifos_wbr_whole_waddr_106) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_7137), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_0__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_0__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_0__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_0_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_6937), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_5768), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__u0 ( .ck(ispd_clk), .d(n_5766), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_0__u0 ( .ck(ispd_clk), .d(n_13131), .o(wbs_wbb3_2_wbb2_dat_o_i) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_10__u0 ( .ck(ispd_clk), .d(n_13401), .o(wbs_wbb3_2_wbb2_dat_o_i_109) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_11__u0 ( .ck(ispd_clk), .d(n_13400), .o(wbs_wbb3_2_wbb2_dat_o_i_110) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_12__u0 ( .ck(ispd_clk), .d(n_13130), .o(wbs_wbb3_2_wbb2_dat_o_i_111) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_13__u0 ( .ck(ispd_clk), .d(n_13129), .o(wbs_wbb3_2_wbb2_dat_o_i_112) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_14__u0 ( .ck(ispd_clk), .d(n_13128), .o(wbs_wbb3_2_wbb2_dat_o_i_113) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_15__u0 ( .ck(ispd_clk), .d(n_13318), .o(wbs_wbb3_2_wbb2_dat_o_i_114) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_16__u0 ( .ck(ispd_clk), .d(n_13399), .o(wbs_wbb3_2_wbb2_dat_o_i_115) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_17__u0 ( .ck(ispd_clk), .d(n_13144), .o(wbs_wbb3_2_wbb2_dat_o_i_116) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_18__u0 ( .ck(ispd_clk), .d(n_13409), .o(wbs_wbb3_2_wbb2_dat_o_i_117) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_19__u0 ( .ck(ispd_clk), .d(n_13408), .o(wbs_wbb3_2_wbb2_dat_o_i_118) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_1__u0 ( .ck(ispd_clk), .d(n_13407), .o(wbs_wbb3_2_wbb2_dat_o_i_100) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_20__u0 ( .ck(ispd_clk), .d(n_13143), .o(wbs_wbb3_2_wbb2_dat_o_i_119) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_21__u0 ( .ck(ispd_clk), .d(n_13406), .o(wbs_wbb3_2_wbb2_dat_o_i_120) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_22__u0 ( .ck(ispd_clk), .d(n_13405), .o(wbs_wbb3_2_wbb2_dat_o_i_121) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_23__u0 ( .ck(ispd_clk), .d(n_13142), .o(wbs_wbb3_2_wbb2_dat_o_i_122) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_24__u0 ( .ck(ispd_clk), .d(n_13323), .o(wbs_wbb3_2_wbb2_dat_o_i_123) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_25__u0 ( .ck(ispd_clk), .d(n_15942), .o(wbs_wbb3_2_wbb2_dat_o_i_124) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_26__u0 ( .ck(ispd_clk), .d(n_13141), .o(wbs_wbb3_2_wbb2_dat_o_i_125) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_27__u0 ( .ck(ispd_clk), .d(n_13321), .o(wbs_wbb3_2_wbb2_dat_o_i_126) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_28__u0 ( .ck(ispd_clk), .d(n_13140), .o(wbs_wbb3_2_wbb2_dat_o_i_127) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_29__u0 ( .ck(ispd_clk), .d(n_13139), .o(wbs_wbb3_2_wbb2_dat_o_i_128) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_2__u0 ( .ck(ispd_clk), .d(n_13320), .o(wbs_wbb3_2_wbb2_dat_o_i_101) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_30__u0 ( .ck(ispd_clk), .d(n_13404), .o(wbs_wbb3_2_wbb2_dat_o_i_129) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_31__u0 ( .ck(ispd_clk), .d(n_13138), .o(wbs_wbb3_2_wbb2_dat_o_i_130) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_36__u0 ( .ck(ispd_clk), .d(n_13319), .o(wishbone_slave_unit_wbs_sm_wbr_control_in) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_37__u0 ( .ck(ispd_clk), .d(n_13137), .o(wishbone_slave_unit_wbs_sm_wbr_control_in_190) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_3__u0 ( .ck(ispd_clk), .d(n_13136), .o(wbs_wbb3_2_wbb2_dat_o_i_102) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_4__u0 ( .ck(ispd_clk), .d(n_13135), .o(wbs_wbb3_2_wbb2_dat_o_i_103) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_5__u0 ( .ck(ispd_clk), .d(n_13403), .o(wbs_wbb3_2_wbb2_dat_o_i_104) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_6__u0 ( .ck(ispd_clk), .d(n_13402), .o(wbs_wbb3_2_wbb2_dat_o_i_105) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_7__u0 ( .ck(ispd_clk), .d(n_13134), .o(wbs_wbb3_2_wbb2_dat_o_i_106) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_8__u0 ( .ck(ispd_clk), .d(n_13133), .o(wbs_wbb3_2_wbb2_dat_o_i_107) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_9__u0 ( .ck(ispd_clk), .d(n_13132), .o(wbs_wbb3_2_wbb2_dat_o_i_108) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__u0 ( .ck(ispd_clk), .d(n_6926), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__u0 ( .ck(ispd_clk), .d(n_6924), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__u0 ( .ck(ispd_clk), .d(n_6922), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__12__u0 ( .ck(ispd_clk), .d(n_6920), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__12__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__12__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__12__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__51) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__u0 ( .ck(ispd_clk), .d(n_6919), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__u0 ( .ck(ispd_clk), .d(n_6917), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__15__u0 ( .ck(ispd_clk), .d(n_6915), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__u0 ( .ck(ispd_clk), .d(n_6913), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__17__u0 ( .ck(ispd_clk), .d(n_6911), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__17__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__17__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__17__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__56) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__u0 ( .ck(ispd_clk), .d(n_6910), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__u0 ( .ck(ispd_clk), .d(n_6908), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__1__u0 ( .ck(ispd_clk), .d(n_6905), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__20__u0 ( .ck(ispd_clk), .d(n_6903), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__20__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__20__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__20__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__59) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__u0 ( .ck(ispd_clk), .d(n_6902), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__u0 ( .ck(ispd_clk), .d(n_6900), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__23__u0 ( .ck(ispd_clk), .d(n_6898), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__23__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__23__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__23__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__62) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__u0 ( .ck(ispd_clk), .d(n_6897), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__u0 ( .ck(ispd_clk), .d(n_6895), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__u0 ( .ck(ispd_clk), .d(n_6892), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__u0 ( .ck(ispd_clk), .d(n_6889), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__28__u0 ( .ck(ispd_clk), .d(n_6887), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__28__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__28__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__28__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__67) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__u0 ( .ck(ispd_clk), .d(n_6885), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__u0 ( .ck(ispd_clk), .d(n_6883), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__30__u0 ( .ck(ispd_clk), .d(n_6878), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__31__u0 ( .ck(ispd_clk), .d(n_6876), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__31__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__31__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__31__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__70) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__u0 ( .ck(ispd_clk), .d(n_6097), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__u0 ( .ck(ispd_clk), .d(n_7392), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__u0 ( .ck(ispd_clk), .d(n_6875), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__4__u0 ( .ck(ispd_clk), .d(n_6872), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__4__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__4__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__4__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__43) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__5__u0 ( .ck(ispd_clk), .d(n_6140), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__u0 ( .ck(ispd_clk), .d(n_6871), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__7__u0 ( .ck(ispd_clk), .d(n_6869), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__7__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__7__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__7__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__46) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__8__u0 ( .ck(ispd_clk), .d(n_6868), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__8__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__8__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__8__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__47) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__u0 ( .ck(ispd_clk), .d(n_6867), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__u0 ( .ck(ispd_clk), .d(n_6865), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__u0 ( .ck(ispd_clk), .d(n_6932), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__u0 ( .ck(ispd_clk), .d(n_6863), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__u0 ( .ck(ispd_clk), .d(n_6861), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__13__u0 ( .ck(ispd_clk), .d(n_6859), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__14__u0 ( .ck(ispd_clk), .d(n_6857), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__u0 ( .ck(ispd_clk), .d(n_6855), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__u0 ( .ck(ispd_clk), .d(n_6853), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__17__u0 ( .ck(ispd_clk), .d(n_6851), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__u0 ( .ck(ispd_clk), .d(n_6934), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__u0 ( .ck(ispd_clk), .d(n_6849), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__1__u0 ( .ck(ispd_clk), .d(n_6847), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__20__u0 ( .ck(ispd_clk), .d(n_6845), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__u0 ( .ck(ispd_clk), .d(n_6709), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__u0 ( .ck(ispd_clk), .d(n_6842), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__u0 ( .ck(ispd_clk), .d(n_6840), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__u0 ( .ck(ispd_clk), .d(n_6837), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__u0 ( .ck(ispd_clk), .d(n_6835), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__u0 ( .ck(ispd_clk), .d(n_6833), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__u0 ( .ck(ispd_clk), .d(n_6747), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__u0 ( .ck(ispd_clk), .d(n_6830), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__u0 ( .ck(ispd_clk), .d(n_6828), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__u0 ( .ck(ispd_clk), .d(n_6826), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__u0 ( .ck(ispd_clk), .d(n_6824), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__31__u0 ( .ck(ispd_clk), .d(n_6821), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__u0 ( .ck(ispd_clk), .d(n_6129), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__u0 ( .ck(ispd_clk), .d(n_7390), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__u0 ( .ck(ispd_clk), .d(n_6819), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__u0 ( .ck(ispd_clk), .d(n_6816), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__u0 ( .ck(ispd_clk), .d(n_6880), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__u0 ( .ck(ispd_clk), .d(n_6814), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__u0 ( .ck(ispd_clk), .d(n_6812), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__u0 ( .ck(ispd_clk), .d(n_6809), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__u0 ( .ck(ispd_clk), .d(n_6150), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__u0 ( .ck(ispd_clk), .d(n_6095), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__u0 ( .ck(ispd_clk), .d(n_5812), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__u0 ( .ck(ispd_clk), .d(n_6093), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__u0 ( .ck(ispd_clk), .d(n_6091), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__u0 ( .ck(ispd_clk), .d(n_5816), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__u0 ( .ck(ispd_clk), .d(n_6089), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__u0 ( .ck(ispd_clk), .d(n_6099), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__u0 ( .ck(ispd_clk), .d(n_6087), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__u0 ( .ck(ispd_clk), .d(n_6085), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__u0 ( .ck(ispd_clk), .d(n_6103), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__u0 ( .ck(ispd_clk), .d(n_6083), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__u0 ( .ck(ispd_clk), .d(n_6107), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__u0 ( .ck(ispd_clk), .d(n_6081), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__u0 ( .ck(ispd_clk), .d(n_5840), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__u0 ( .ck(ispd_clk), .d(n_5848), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__u0 ( .ck(ispd_clk), .d(n_6079), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__u0 ( .ck(ispd_clk), .d(n_6077), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__u0 ( .ck(ispd_clk), .d(n_6111), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__26__u0 ( .ck(ispd_clk), .d(n_6075), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__u0 ( .ck(ispd_clk), .d(n_5810), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__u0 ( .ck(ispd_clk), .d(n_5806), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__u0 ( .ck(ispd_clk), .d(n_5822), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__u0 ( .ck(ispd_clk), .d(n_6073), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__u0 ( .ck(ispd_clk), .d(n_5792), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__u0 ( .ck(ispd_clk), .d(n_6071), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__u0 ( .ck(ispd_clk), .d(n_5790), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__37__u0 ( .ck(ispd_clk), .d(n_7388), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__37__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__37__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__37__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_11__466) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__u0 ( .ck(ispd_clk), .d(n_5981), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__u0 ( .ck(ispd_clk), .d(n_6069), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__u0 ( .ck(ispd_clk), .d(n_6109), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__u0 ( .ck(ispd_clk), .d(n_6067), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__u0 ( .ck(ispd_clk), .d(n_6065), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__u0 ( .ck(ispd_clk), .d(n_6063), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__u0 ( .ck(ispd_clk), .d(n_6101), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__u0 ( .ck(ispd_clk), .d(n_6806), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__u0 ( .ck(ispd_clk), .d(n_6804), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__u0 ( .ck(ispd_clk), .d(n_6801), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__u0 ( .ck(ispd_clk), .d(n_6799), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__u0 ( .ck(ispd_clk), .d(n_6797), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__u0 ( .ck(ispd_clk), .d(n_6795), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__u0 ( .ck(ispd_clk), .d(n_6156), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__16__u0 ( .ck(ispd_clk), .d(n_6793), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__16__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__16__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__16__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__484) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__u0 ( .ck(ispd_clk), .d(n_6158), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__u0 ( .ck(ispd_clk), .d(n_6791), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__19__u0 ( .ck(ispd_clk), .d(n_6789), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__19__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__19__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__19__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__487) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__u0 ( .ck(ispd_clk), .d(n_6788), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__u0 ( .ck(ispd_clk), .d(n_6785), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__u0 ( .ck(ispd_clk), .d(n_6783), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__u0 ( .ck(ispd_clk), .d(n_6781), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__23__u0 ( .ck(ispd_clk), .d(n_6778), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__u0 ( .ck(ispd_clk), .d(n_6776), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__25__u0 ( .ck(ispd_clk), .d(n_6774), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__u0 ( .ck(ispd_clk), .d(n_6929), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__u0 ( .ck(ispd_clk), .d(n_6772), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__28__u0 ( .ck(ispd_clk), .d(n_6770), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__u0 ( .ck(ispd_clk), .d(n_6768), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__u0 ( .ck(ispd_clk), .d(n_6766), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__u0 ( .ck(ispd_clk), .d(n_6763), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__u0 ( .ck(ispd_clk), .d(n_6761), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__u0 ( .ck(ispd_clk), .d(n_6127), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__u0 ( .ck(ispd_clk), .d(n_7366), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__u0 ( .ck(ispd_clk), .d(n_6759), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__u0 ( .ck(ispd_clk), .d(n_6757), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__u0 ( .ck(ispd_clk), .d(n_6754), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__u0 ( .ck(ispd_clk), .d(n_6514), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__u0 ( .ck(ispd_clk), .d(n_6752), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__u0 ( .ck(ispd_clk), .d(n_6745), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__u0 ( .ck(ispd_clk), .d(n_6749), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__0__u0 ( .ck(ispd_clk), .d(n_6061), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__0__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__0__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__0__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__u0 ( .ck(ispd_clk), .d(n_6060), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__u0 ( .ck(ispd_clk), .d(n_6058), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__u0 ( .ck(ispd_clk), .d(n_6056), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__u0 ( .ck(ispd_clk), .d(n_5772), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__u0 ( .ck(ispd_clk), .d(n_5774), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__15__u0 ( .ck(ispd_clk), .d(n_6054), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__15__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__15__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__15__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__522) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__u0 ( .ck(ispd_clk), .d(n_5804), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__u0 ( .ck(ispd_clk), .d(n_6053), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__u0 ( .ck(ispd_clk), .d(n_5838), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__u0 ( .ck(ispd_clk), .d(n_6051), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__u0 ( .ck(ispd_clk), .d(n_5844), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__u0 ( .ck(ispd_clk), .d(n_6049), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__u0 ( .ck(ispd_clk), .d(n_6047), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__u0 ( .ck(ispd_clk), .d(n_5854), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__u0 ( .ck(ispd_clk), .d(n_5858), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__24__u0 ( .ck(ispd_clk), .d(n_5967), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__24__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__24__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__24__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__531) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__25__u0 ( .ck(ispd_clk), .d(n_5850), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__25__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__25__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__25__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__532) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__u0 ( .ck(ispd_clk), .d(n_6045), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__u0 ( .ck(ispd_clk), .d(n_5794), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__u0 ( .ck(ispd_clk), .d(n_6043), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__29__u0 ( .ck(ispd_clk), .d(n_6041), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__29__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__29__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__29__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__536) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__2__u0 ( .ck(ispd_clk), .d(n_6040), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__2__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__2__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__2__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__509) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__u0 ( .ck(ispd_clk), .d(n_5936), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__31__u0 ( .ck(ispd_clk), .d(n_6039), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__u0 ( .ck(ispd_clk), .d(n_5800), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__37__u0 ( .ck(ispd_clk), .d(n_7387), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__37__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__37__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__37__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__544) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__u0 ( .ck(ispd_clk), .d(n_5870), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__u0 ( .ck(ispd_clk), .d(n_6037), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__u0 ( .ck(ispd_clk), .d(n_5776), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__u0 ( .ck(ispd_clk), .d(n_6035), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__u0 ( .ck(ispd_clk), .d(n_5814), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__u0 ( .ck(ispd_clk), .d(n_6033), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__u0 ( .ck(ispd_clk), .d(n_5833), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__u0 ( .ck(ispd_clk), .d(n_6031), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__u0 ( .ck(ispd_clk), .d(n_6029), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__u0 ( .ck(ispd_clk), .d(n_5862), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__u0 ( .ck(ispd_clk), .d(n_6027), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__u0 ( .ck(ispd_clk), .d(n_6025), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__u0 ( .ck(ispd_clk), .d(n_6023), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__u0 ( .ck(ispd_clk), .d(n_5796), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__u0 ( .ck(ispd_clk), .d(n_6021), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__u0 ( .ck(ispd_clk), .d(n_6019), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__u0 ( .ck(ispd_clk), .d(n_6017), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__u0 ( .ck(ispd_clk), .d(n_6015), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__u0 ( .ck(ispd_clk), .d(n_6013), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__u0 ( .ck(ispd_clk), .d(n_6105), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__u0 ( .ck(ispd_clk), .d(n_6011), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__u0 ( .ck(ispd_clk), .d(n_6009), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__u0 ( .ck(ispd_clk), .d(n_6007), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__u0 ( .ck(ispd_clk), .d(n_5830), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__u0 ( .ck(ispd_clk), .d(n_6005), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__u0 ( .ck(ispd_clk), .d(n_6003), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__u0 ( .ck(ispd_clk), .d(n_6001), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__u0 ( .ck(ispd_clk), .d(n_5798), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__u0 ( .ck(ispd_clk), .d(n_5999), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__u0 ( .ck(ispd_clk), .d(n_5997), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__u0 ( .ck(ispd_clk), .d(n_5995), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__u0 ( .ck(ispd_clk), .d(n_5993), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__u0 ( .ck(ispd_clk), .d(n_5991), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__37__u0 ( .ck(ispd_clk), .d(n_7364), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__37__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__37__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__37__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_14__583) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__u0 ( .ck(ispd_clk), .d(n_5989), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__u0 ( .ck(ispd_clk), .d(n_5987), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__u0 ( .ck(ispd_clk), .d(n_5985), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__u0 ( .ck(ispd_clk), .d(n_5827), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__u0 ( .ck(ispd_clk), .d(n_5983), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__u0 ( .ck(ispd_clk), .d(n_5868), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__u0 ( .ck(ispd_clk), .d(n_5979), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__u0 ( .ck(ispd_clk), .d(n_5856), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__u0 ( .ck(ispd_clk), .d(n_5842), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__u0 ( .ck(ispd_clk), .d(n_5977), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__u0 ( .ck(ispd_clk), .d(n_5975), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__u0 ( .ck(ispd_clk), .d(n_5973), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__u0 ( .ck(ispd_clk), .d(n_5864), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__u0 ( .ck(ispd_clk), .d(n_5971), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__u0 ( .ck(ispd_clk), .d(n_5824), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__u0 ( .ck(ispd_clk), .d(n_5969), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__u0 ( .ck(ispd_clk), .d(n_5866), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__u0 ( .ck(ispd_clk), .d(n_5966), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__u0 ( .ck(ispd_clk), .d(n_5964), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__u0 ( .ck(ispd_clk), .d(n_5962), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__u0 ( .ck(ispd_clk), .d(n_5782), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__u0 ( .ck(ispd_clk), .d(n_5960), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__u0 ( .ck(ispd_clk), .d(n_5784), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__u0 ( .ck(ispd_clk), .d(n_5958), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__u0 ( .ck(ispd_clk), .d(n_5786), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__u0 ( .ck(ispd_clk), .d(n_5956), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__u0 ( .ck(ispd_clk), .d(n_5954), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__u0 ( .ck(ispd_clk), .d(n_5952), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__u0 ( .ck(ispd_clk), .d(n_5788), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__u0 ( .ck(ispd_clk), .d(n_5950), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__u0 ( .ck(ispd_clk), .d(n_5802), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__31__u0 ( .ck(ispd_clk), .d(n_5948), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__u0 ( .ck(ispd_clk), .d(n_5808), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__37__u0 ( .ck(ispd_clk), .d(n_7386), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__37__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__37__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__37__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_15__622) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__u0 ( .ck(ispd_clk), .d(n_5819), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__u0 ( .ck(ispd_clk), .d(n_5946), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__u0 ( .ck(ispd_clk), .d(n_5860), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__u0 ( .ck(ispd_clk), .d(n_5780), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__u0 ( .ck(ispd_clk), .d(n_5778), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__u0 ( .ck(ispd_clk), .d(n_5944), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__u0 ( .ck(ispd_clk), .d(n_5942), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__u0 ( .ck(ispd_clk), .d(n_6743), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__u0 ( .ck(ispd_clk), .d(n_6741), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__u0 ( .ck(ispd_clk), .d(n_6738), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__u0 ( .ck(ispd_clk), .d(n_6735), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__u0 ( .ck(ispd_clk), .d(n_6733), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__u0 ( .ck(ispd_clk), .d(n_6731), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__u0 ( .ck(ispd_clk), .d(n_6729), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__u0 ( .ck(ispd_clk), .d(n_6726), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__u0 ( .ck(ispd_clk), .d(n_6724), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__u0 ( .ck(ispd_clk), .d(n_6162), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__u0 ( .ck(ispd_clk), .d(n_6722), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__u0 ( .ck(ispd_clk), .d(n_6720), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__u0 ( .ck(ispd_clk), .d(n_6718), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__u0 ( .ck(ispd_clk), .d(n_6716), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__u0 ( .ck(ispd_clk), .d(n_6142), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__23__u0 ( .ck(ispd_clk), .d(n_6714), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__u0 ( .ck(ispd_clk), .d(n_6152), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__u0 ( .ck(ispd_clk), .d(n_6712), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__u0 ( .ck(ispd_clk), .d(n_6154), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__u0 ( .ck(ispd_clk), .d(n_6707), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__u0 ( .ck(ispd_clk), .d(n_6705), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__u0 ( .ck(ispd_clk), .d(n_6144), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__u0 ( .ck(ispd_clk), .d(n_6146), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__u0 ( .ck(ispd_clk), .d(n_6703), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__u0 ( .ck(ispd_clk), .d(n_6148), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__u0 ( .ck(ispd_clk), .d(n_5836), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__u0 ( .ck(ispd_clk), .d(n_7385), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__u0 ( .ck(ispd_clk), .d(n_6701), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__u0 ( .ck(ispd_clk), .d(n_6699), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__u0 ( .ck(ispd_clk), .d(n_6171), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__u0 ( .ck(ispd_clk), .d(n_6697), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__u0 ( .ck(ispd_clk), .d(n_6695), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__u0 ( .ck(ispd_clk), .d(n_6693), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__u0 ( .ck(ispd_clk), .d(n_6691), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__u0 ( .ck(ispd_clk), .d(n_6689), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__u0 ( .ck(ispd_clk), .d(n_6686), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__u0 ( .ck(ispd_clk), .d(n_6684), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__u0 ( .ck(ispd_clk), .d(n_6682), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__u0 ( .ck(ispd_clk), .d(n_6680), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__u0 ( .ck(ispd_clk), .d(n_6678), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__u0 ( .ck(ispd_clk), .d(n_6676), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__u0 ( .ck(ispd_clk), .d(n_6674), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__u0 ( .ck(ispd_clk), .d(n_6672), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__u0 ( .ck(ispd_clk), .d(n_6670), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__u0 ( .ck(ispd_clk), .d(n_6668), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__u0 ( .ck(ispd_clk), .d(n_6665), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__u0 ( .ck(ispd_clk), .d(n_6662), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__u0 ( .ck(ispd_clk), .d(n_6659), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__u0 ( .ck(ispd_clk), .d(n_6657), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__u0 ( .ck(ispd_clk), .d(n_6654), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__u0 ( .ck(ispd_clk), .d(n_6651), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__u0 ( .ck(ispd_clk), .d(n_6649), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__u0 ( .ck(ispd_clk), .d(n_6647), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__u0 ( .ck(ispd_clk), .d(n_6644), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__28__u0 ( .ck(ispd_clk), .d(n_6641), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__u0 ( .ck(ispd_clk), .d(n_6639), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__u0 ( .ck(ispd_clk), .d(n_6636), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__u0 ( .ck(ispd_clk), .d(n_6634), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__u0 ( .ck(ispd_clk), .d(n_6631), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__u0 ( .ck(ispd_clk), .d(n_5940), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__u0 ( .ck(ispd_clk), .d(n_7383), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__u0 ( .ck(ispd_clk), .d(n_6629), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__u0 ( .ck(ispd_clk), .d(n_6626), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__u0 ( .ck(ispd_clk), .d(n_6623), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__6__u0 ( .ck(ispd_clk), .d(n_6621), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__6__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__6__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__6__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_2__6) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__u0 ( .ck(ispd_clk), .d(n_6620), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__8__u0 ( .ck(ispd_clk), .d(n_6617), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__u0 ( .ck(ispd_clk), .d(n_6615), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__u0 ( .ck(ispd_clk), .d(n_6613), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__u0 ( .ck(ispd_clk), .d(n_6610), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__u0 ( .ck(ispd_clk), .d(n_6607), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__u0 ( .ck(ispd_clk), .d(n_6605), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__u0 ( .ck(ispd_clk), .d(n_6603), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__14__u0 ( .ck(ispd_clk), .d(n_6601), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__u0 ( .ck(ispd_clk), .d(n_6598), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__u0 ( .ck(ispd_clk), .d(n_6596), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__u0 ( .ck(ispd_clk), .d(n_6594), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__u0 ( .ck(ispd_clk), .d(n_6592), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__u0 ( .ck(ispd_clk), .d(n_6589), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__u0 ( .ck(ispd_clk), .d(n_6587), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__u0 ( .ck(ispd_clk), .d(n_6585), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__21__u0 ( .ck(ispd_clk), .d(n_6582), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__21__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__21__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__21__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__177) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__22__u0 ( .ck(ispd_clk), .d(n_6580), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__22__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__22__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__22__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__178) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__u0 ( .ck(ispd_clk), .d(n_6578), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__u0 ( .ck(ispd_clk), .d(n_6575), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__u0 ( .ck(ispd_clk), .d(n_6572), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__26__u0 ( .ck(ispd_clk), .d(n_6569), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__27__u0 ( .ck(ispd_clk), .d(n_6567), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__27__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__27__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__27__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__183) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__u0 ( .ck(ispd_clk), .d(n_6566), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__u0 ( .ck(ispd_clk), .d(n_6563), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__u0 ( .ck(ispd_clk), .d(n_6561), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__u0 ( .ck(ispd_clk), .d(n_6558), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__u0 ( .ck(ispd_clk), .d(n_6556), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__u0 ( .ck(ispd_clk), .d(n_6123), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__u0 ( .ck(ispd_clk), .d(n_7381), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__u0 ( .ck(ispd_clk), .d(n_6553), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__u0 ( .ck(ispd_clk), .d(n_6550), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__u0 ( .ck(ispd_clk), .d(n_6548), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__u0 ( .ck(ispd_clk), .d(n_6546), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__u0 ( .ck(ispd_clk), .d(n_6543), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__8__u0 ( .ck(ispd_clk), .d(n_6541), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__u0 ( .ck(ispd_clk), .d(n_6538), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__0__u0 ( .ck(ispd_clk), .d(n_6536), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__u0 ( .ck(ispd_clk), .d(n_6534), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__u0 ( .ck(ispd_clk), .d(n_6532), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__u0 ( .ck(ispd_clk), .d(n_6530), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__u0 ( .ck(ispd_clk), .d(n_6528), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__u0 ( .ck(ispd_clk), .d(n_6526), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__15__u0 ( .ck(ispd_clk), .d(n_6523), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__u0 ( .ck(ispd_clk), .d(n_6521), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__u0 ( .ck(ispd_clk), .d(n_6518), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__u0 ( .ck(ispd_clk), .d(n_6516), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__u0 ( .ck(ispd_clk), .d(n_6166), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__u0 ( .ck(ispd_clk), .d(n_6512), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__u0 ( .ck(ispd_clk), .d(n_6509), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__u0 ( .ck(ispd_clk), .d(n_6168), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__22__u0 ( .ck(ispd_clk), .d(n_6506), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__u0 ( .ck(ispd_clk), .d(n_6504), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__u0 ( .ck(ispd_clk), .d(n_6501), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__u0 ( .ck(ispd_clk), .d(n_6498), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__u0 ( .ck(ispd_clk), .d(n_6495), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__u0 ( .ck(ispd_clk), .d(n_6493), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__u0 ( .ck(ispd_clk), .d(n_6490), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__u0 ( .ck(ispd_clk), .d(n_6488), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__u0 ( .ck(ispd_clk), .d(n_6485), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__u0 ( .ck(ispd_clk), .d(n_6483), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__u0 ( .ck(ispd_clk), .d(n_6480), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__u0 ( .ck(ispd_clk), .d(n_5938), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__u0 ( .ck(ispd_clk), .d(n_7379), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__u0 ( .ck(ispd_clk), .d(n_6477), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__u0 ( .ck(ispd_clk), .d(n_6475), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__u0 ( .ck(ispd_clk), .d(n_6473), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__u0 ( .ck(ispd_clk), .d(n_6470), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__u0 ( .ck(ispd_clk), .d(n_6468), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__u0 ( .ck(ispd_clk), .d(n_6465), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__u0 ( .ck(ispd_clk), .d(n_6463), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__u0 ( .ck(ispd_clk), .d(n_6461), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__u0 ( .ck(ispd_clk), .d(n_6458), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__u0 ( .ck(ispd_clk), .d(n_6160), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__u0 ( .ck(ispd_clk), .d(n_6456), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__u0 ( .ck(ispd_clk), .d(n_6453), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__14__u0 ( .ck(ispd_clk), .d(n_6451), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__u0 ( .ck(ispd_clk), .d(n_6448), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__u0 ( .ck(ispd_clk), .d(n_6446), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__u0 ( .ck(ispd_clk), .d(n_6443), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__u0 ( .ck(ispd_clk), .d(n_6440), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__u0 ( .ck(ispd_clk), .d(n_6438), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__u0 ( .ck(ispd_clk), .d(n_6435), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__u0 ( .ck(ispd_clk), .d(n_6433), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__u0 ( .ck(ispd_clk), .d(n_6430), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__u0 ( .ck(ispd_clk), .d(n_6427), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__u0 ( .ck(ispd_clk), .d(n_6425), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__u0 ( .ck(ispd_clk), .d(n_6423), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__u0 ( .ck(ispd_clk), .d(n_6420), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__26__u0 ( .ck(ispd_clk), .d(n_6417), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__u0 ( .ck(ispd_clk), .d(n_6415), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__u0 ( .ck(ispd_clk), .d(n_6413), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__u0 ( .ck(ispd_clk), .d(n_6410), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__u0 ( .ck(ispd_clk), .d(n_6407), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__u0 ( .ck(ispd_clk), .d(n_6405), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__u0 ( .ck(ispd_clk), .d(n_6402), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__u0 ( .ck(ispd_clk), .d(n_6121), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__u0 ( .ck(ispd_clk), .d(n_7377), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__u0 ( .ck(ispd_clk), .d(n_6400), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__u0 ( .ck(ispd_clk), .d(n_6398), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__u0 ( .ck(ispd_clk), .d(n_6395), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__u0 ( .ck(ispd_clk), .d(n_6393), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__u0 ( .ck(ispd_clk), .d(n_6390), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__u0 ( .ck(ispd_clk), .d(n_6388), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__u0 ( .ck(ispd_clk), .d(n_6386), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__u0 ( .ck(ispd_clk), .d(n_6384), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__u0 ( .ck(ispd_clk), .d(n_6382), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__u0 ( .ck(ispd_clk), .d(n_6379), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__u0 ( .ck(ispd_clk), .d(n_6376), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__13__u0 ( .ck(ispd_clk), .d(n_6374), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__13__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__13__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__13__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__247) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__14__u0 ( .ck(ispd_clk), .d(n_6373), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__14__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__14__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__14__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__248) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__15__u0 ( .ck(ispd_clk), .d(n_6372), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__15__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__15__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__15__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__249) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__u0 ( .ck(ispd_clk), .d(n_6371), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__u0 ( .ck(ispd_clk), .d(n_6369), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__u0 ( .ck(ispd_clk), .d(n_6366), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__u0 ( .ck(ispd_clk), .d(n_6364), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__u0 ( .ck(ispd_clk), .d(n_6361), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__20__u0 ( .ck(ispd_clk), .d(n_6358), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__u0 ( .ck(ispd_clk), .d(n_6355), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__22__u0 ( .ck(ispd_clk), .d(n_6353), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__u0 ( .ck(ispd_clk), .d(n_6350), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__24__u0 ( .ck(ispd_clk), .d(n_6348), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__24__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__24__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__24__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__258) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__u0 ( .ck(ispd_clk), .d(n_6347), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__26__u0 ( .ck(ispd_clk), .d(n_6345), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__26__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__26__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__26__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__260) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__u0 ( .ck(ispd_clk), .d(n_6344), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__u0 ( .ck(ispd_clk), .d(n_6342), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__u0 ( .ck(ispd_clk), .d(n_6340), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__2__u0 ( .ck(ispd_clk), .d(n_6338), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__2__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__2__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__2__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__236) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__u0 ( .ck(ispd_clk), .d(n_6337), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__31__u0 ( .ck(ispd_clk), .d(n_6335), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__31__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__31__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__31__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__265) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__u0 ( .ck(ispd_clk), .d(n_6119), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__37__u0 ( .ck(ispd_clk), .d(n_7375), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__37__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__37__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__37__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__271) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__3__u0 ( .ck(ispd_clk), .d(n_6334), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__3__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__3__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__3__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__237) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__4__u0 ( .ck(ispd_clk), .d(n_6333), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__4__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__4__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__4__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__238) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__u0 ( .ck(ispd_clk), .d(n_6331), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__u0 ( .ck(ispd_clk), .d(n_6329), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__u0 ( .ck(ispd_clk), .d(n_6327), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__u0 ( .ck(ispd_clk), .d(n_6325), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__9__u0 ( .ck(ispd_clk), .d(n_6323), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__9__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__9__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__9__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__243) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__u0 ( .ck(ispd_clk), .d(n_5846), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__u0 ( .ck(ispd_clk), .d(n_5934), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__u0 ( .ck(ispd_clk), .d(n_5932), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__u0 ( .ck(ispd_clk), .d(n_5930), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__u0 ( .ck(ispd_clk), .d(n_5928), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__14__u0 ( .ck(ispd_clk), .d(n_5926), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__u0 ( .ck(ispd_clk), .d(n_5924), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__u0 ( .ck(ispd_clk), .d(n_5922), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__u0 ( .ck(ispd_clk), .d(n_5920), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__18__u0 ( .ck(ispd_clk), .d(n_5918), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__u0 ( .ck(ispd_clk), .d(n_5916), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__1__u0 ( .ck(ispd_clk), .d(n_5914), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__20__u0 ( .ck(ispd_clk), .d(n_5912), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__u0 ( .ck(ispd_clk), .d(n_5910), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__22__u0 ( .ck(ispd_clk), .d(n_5908), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__u0 ( .ck(ispd_clk), .d(n_5906), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__u0 ( .ck(ispd_clk), .d(n_5852), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__u0 ( .ck(ispd_clk), .d(n_5904), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__u0 ( .ck(ispd_clk), .d(n_5902), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__u0 ( .ck(ispd_clk), .d(n_5900), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__u0 ( .ck(ispd_clk), .d(n_5898), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__u0 ( .ck(ispd_clk), .d(n_5896), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__u0 ( .ck(ispd_clk), .d(n_5894), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__30__u0 ( .ck(ispd_clk), .d(n_5892), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__31__u0 ( .ck(ispd_clk), .d(n_5890), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__u0 ( .ck(ispd_clk), .d(n_5888), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__37__u0 ( .ck(ispd_clk), .d(n_7374), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__37__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__37__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__37__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_7__310) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__u0 ( .ck(ispd_clk), .d(n_5886), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__u0 ( .ck(ispd_clk), .d(n_5884), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__u0 ( .ck(ispd_clk), .d(n_5882), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__u0 ( .ck(ispd_clk), .d(n_5880), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__u0 ( .ck(ispd_clk), .d(n_5878), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__u0 ( .ck(ispd_clk), .d(n_5876), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__u0 ( .ck(ispd_clk), .d(n_5874), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__u0 ( .ck(ispd_clk), .d(n_6321), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__u0 ( .ck(ispd_clk), .d(n_6318), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__u0 ( .ck(ispd_clk), .d(n_6315), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__u0 ( .ck(ispd_clk), .d(n_6313), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__u0 ( .ck(ispd_clk), .d(n_6311), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__u0 ( .ck(ispd_clk), .d(n_6308), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__u0 ( .ck(ispd_clk), .d(n_6305), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__u0 ( .ck(ispd_clk), .d(n_6303), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__u0 ( .ck(ispd_clk), .d(n_6301), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__18__u0 ( .ck(ispd_clk), .d(n_6298), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__18__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__18__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__18__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__330) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__u0 ( .ck(ispd_clk), .d(n_6297), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__u0 ( .ck(ispd_clk), .d(n_6295), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__u0 ( .ck(ispd_clk), .d(n_6292), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__u0 ( .ck(ispd_clk), .d(n_6289), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__u0 ( .ck(ispd_clk), .d(n_6286), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__u0 ( .ck(ispd_clk), .d(n_6284), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__u0 ( .ck(ispd_clk), .d(n_6281), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__u0 ( .ck(ispd_clk), .d(n_6278), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__26__u0 ( .ck(ispd_clk), .d(n_6164), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__u0 ( .ck(ispd_clk), .d(n_6276), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__u0 ( .ck(ispd_clk), .d(n_6273), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__u0 ( .ck(ispd_clk), .d(n_6271), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__u0 ( .ck(ispd_clk), .d(n_6268), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__30__u0 ( .ck(ispd_clk), .d(n_6266), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__30__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__30__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__30__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__342) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__u0 ( .ck(ispd_clk), .d(n_6264), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__u0 ( .ck(ispd_clk), .d(n_5872), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__u0 ( .ck(ispd_clk), .d(n_7371), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__u0 ( .ck(ispd_clk), .d(n_6261), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__u0 ( .ck(ispd_clk), .d(n_6259), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__u0 ( .ck(ispd_clk), .d(n_6257), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__u0 ( .ck(ispd_clk), .d(n_6254), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__u0 ( .ck(ispd_clk), .d(n_6252), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__u0 ( .ck(ispd_clk), .d(n_6249), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__u0 ( .ck(ispd_clk), .d(n_6246), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__u0 ( .ck(ispd_clk), .d(n_6243), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__u0 ( .ck(ispd_clk), .d(n_6240), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__u0 ( .ck(ispd_clk), .d(n_6238), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__12__u0 ( .ck(ispd_clk), .d(n_6235), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__12__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__12__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__12__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__363) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__u0 ( .ck(ispd_clk), .d(n_6234), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__u0 ( .ck(ispd_clk), .d(n_6231), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__365) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__u0 ( .ck(ispd_clk), .d(n_6230), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__u0 ( .ck(ispd_clk), .d(n_6228), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__u0 ( .ck(ispd_clk), .d(n_6226), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__u0 ( .ck(ispd_clk), .d(n_6223), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__u0 ( .ck(ispd_clk), .d(n_6221), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__1__u0 ( .ck(ispd_clk), .d(n_6216), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__20__u0 ( .ck(ispd_clk), .d(n_6213), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__u0 ( .ck(ispd_clk), .d(n_6211), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__u0 ( .ck(ispd_clk), .d(n_6208), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__23__u0 ( .ck(ispd_clk), .d(n_6206), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__23__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__23__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__23__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__374) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__u0 ( .ck(ispd_clk), .d(n_6204), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__25__u0 ( .ck(ispd_clk), .d(n_6201), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__25__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__25__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__25__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__376) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__26__u0 ( .ck(ispd_clk), .d(n_6200), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__26__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__26__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__26__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__377) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__u0 ( .ck(ispd_clk), .d(n_6199), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__28__u0 ( .ck(ispd_clk), .d(n_6196), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__28__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__28__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__28__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__379) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__29__u0 ( .ck(ispd_clk), .d(n_6195), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__29__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__29__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__29__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__380) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__u0 ( .ck(ispd_clk), .d(n_6193), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__u0 ( .ck(ispd_clk), .d(n_6191), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__31__u0 ( .ck(ispd_clk), .d(n_6189), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__u0 ( .ck(ispd_clk), .d(n_6117), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__u0 ( .ck(ispd_clk), .d(n_7368), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__u0 ( .ck(ispd_clk), .d(n_6186), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__u0 ( .ck(ispd_clk), .d(n_6184), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__u0 ( .ck(ispd_clk), .d(n_6181), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__u0 ( .ck(ispd_clk), .d(n_6179), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__7__u0 ( .ck(ispd_clk), .d(n_6177), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__7__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__7__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__7__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__358) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__8__u0 ( .ck(ispd_clk), .d(n_6175), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__8__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__8__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__8__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__359) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__9__u0 ( .ck(ispd_clk), .d(n_6173), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__9__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__9__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__9__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__360) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_0__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus1) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_1__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_93) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_2__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_94) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_3__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_95) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_70) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_71) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_72) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg_0__u0 ( .ck(ispd_clk), .d(n_8765), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg_1__u0 ( .ck(ispd_clk), .d(n_8713), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg_2__u0 ( .ck(ispd_clk), .d(n_8716), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg_3__u0 ( .ck(ispd_clk), .d(n_8714), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg_0__u0 ( .ck(ispd_clk), .d(n_8745), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg_1__u0 ( .ck(ispd_clk), .d(n_8784), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg_2__u0 ( .ck(ispd_clk), .d(n_8712), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg_3__u0 ( .ck(ispd_clk), .d(n_8711), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_70), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_71), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_72), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_8709), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_8708), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_8707), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_3__u0 ( .ck(ispd_clk), .d(n_8705), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_0__u0 ( .ck(ispd_clk), .d(n_8703), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_1__u0 ( .ck(ispd_clk), .d(n_8701), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_2__u0 ( .ck(ispd_clk), .d(n_8699), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_3__u0 ( .ck(ispd_clk), .d(n_8697), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(n_8695), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(n_8694), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(n_8693), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg_3__u0 ( .ck(ispd_clk), .d(n_8692), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg_0__u0 ( .ck(ispd_clk), .d(n_9340), .o(wishbone_slave_unit_fifos_wbw_whole_waddr) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg_1__u0 ( .ck(ispd_clk), .d(n_9343), .o(wishbone_slave_unit_fifos_wbw_whole_waddr_55) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg_2__u0 ( .ck(ispd_clk), .d(n_9194), .o(wishbone_slave_unit_fifos_wbw_whole_waddr_56) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg_3__u0 ( .ck(ispd_clk), .d(n_9189), .o(wishbone_slave_unit_fifos_wbw_whole_waddr_57) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus1), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_93), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_94), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_95), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_9187), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_9185), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_9184), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg_3__u0 ( .ck(ispd_clk), .d(n_9183), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(n_9342), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(n_9192), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(n_9182), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg_3__u0 ( .ck(ispd_clk), .d(n_9181), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_0__u0 ( .ck(ispd_clk), .d(n_12853), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_10__u0 ( .ck(ispd_clk), .d(n_12852), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_393) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_11__u0 ( .ck(ispd_clk), .d(n_12851), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_394) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_12__u0 ( .ck(ispd_clk), .d(n_12850), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_395) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_13__u0 ( .ck(ispd_clk), .d(n_12849), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_396) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_14__u0 ( .ck(ispd_clk), .d(n_12848), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_397) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_15__u0 ( .ck(ispd_clk), .d(n_12847), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_398) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_16__u0 ( .ck(ispd_clk), .d(n_12846), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_399) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_17__u0 ( .ck(ispd_clk), .d(n_12845), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_400) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_18__u0 ( .ck(ispd_clk), .d(n_15565), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_401) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_19__u0 ( .ck(ispd_clk), .d(n_12843), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_402) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_1__u0 ( .ck(ispd_clk), .d(n_12842), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_384) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_20__u0 ( .ck(ispd_clk), .d(n_12841), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_403) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_21__u0 ( .ck(ispd_clk), .d(n_12775), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_404) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_22__u0 ( .ck(ispd_clk), .d(n_12840), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_405) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_23__u0 ( .ck(ispd_clk), .d(n_12839), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_406) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_24__u0 ( .ck(ispd_clk), .d(n_15540), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_407) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_25__u0 ( .ck(ispd_clk), .d(n_12774), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_408) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_26__u0 ( .ck(ispd_clk), .d(n_12951), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_409) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_27__u0 ( .ck(ispd_clk), .d(n_12837), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_410) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_28__u0 ( .ck(ispd_clk), .d(n_12836), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_411) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_29__u0 ( .ck(ispd_clk), .d(n_12835), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_412) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_2__u0 ( .ck(ispd_clk), .d(n_12834), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_385) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_30__u0 ( .ck(ispd_clk), .d(n_12773), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_413) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_31__u0 ( .ck(ispd_clk), .d(n_12833), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_414) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_32__u0 ( .ck(ispd_clk), .d(n_12832), .o(wishbone_slave_unit_pcim_if_wbw_cbe_in) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__u0 ( .ck(ispd_clk), .d(n_12831), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_34__u0 ( .ck(ispd_clk), .d(n_12830), .o(wishbone_slave_unit_pcim_if_wbw_cbe_in_416) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_35__u0 ( .ck(ispd_clk), .d(n_12829), .o(wishbone_slave_unit_pcim_if_wbw_cbe_in_417) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__u0 ( .ck(ispd_clk), .d(n_12828), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_3__u0 ( .ck(ispd_clk), .d(n_12827), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_386) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_4__u0 ( .ck(ispd_clk), .d(n_12826), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_387) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_5__u0 ( .ck(ispd_clk), .d(n_12825), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_388) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_6__u0 ( .ck(ispd_clk), .d(n_12824), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_389) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_7__u0 ( .ck(ispd_clk), .d(n_12823), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_390) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_8__u0 ( .ck(ispd_clk), .d(n_12822), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_391) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_9__u0 ( .ck(ispd_clk), .d(n_12821), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_392) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__u0 ( .ck(ispd_clk), .d(n_11513), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__u0 ( .ck(ispd_clk), .d(n_11512), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__u0 ( .ck(ispd_clk), .d(n_11510), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__u0 ( .ck(ispd_clk), .d(n_10424), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__u0 ( .ck(ispd_clk), .d(n_11509), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__u0 ( .ck(ispd_clk), .d(n_10423), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__u0 ( .ck(ispd_clk), .d(n_11507), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__u0 ( .ck(ispd_clk), .d(n_11505), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__u0 ( .ck(ispd_clk), .d(n_11503), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__u0 ( .ck(ispd_clk), .d(n_11502), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__u0 ( .ck(ispd_clk), .d(n_11500), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__u0 ( .ck(ispd_clk), .d(n_11499), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__u0 ( .ck(ispd_clk), .d(n_11497), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__u0 ( .ck(ispd_clk), .d(n_11496), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__u0 ( .ck(ispd_clk), .d(n_10421), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__u0 ( .ck(ispd_clk), .d(n_11495), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__u0 ( .ck(ispd_clk), .d(n_11493), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__u0 ( .ck(ispd_clk), .d(n_10419), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__u0 ( .ck(ispd_clk), .d(n_11492), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__u0 ( .ck(ispd_clk), .d(n_11490), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__u0 ( .ck(ispd_clk), .d(n_11489), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__u0 ( .ck(ispd_clk), .d(n_11487), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__u0 ( .ck(ispd_clk), .d(n_10418), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__u0 ( .ck(ispd_clk), .d(n_11485), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__u0 ( .ck(ispd_clk), .d(n_11484), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__u0 ( .ck(ispd_clk), .d(n_10829), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__u0 ( .ck(ispd_clk), .d(n_10828), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__u0 ( .ck(ispd_clk), .d(n_10366), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__u0 ( .ck(ispd_clk), .d(n_11710), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__u0 ( .ck(ispd_clk), .d(n_8959), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__u0 ( .ck(ispd_clk), .d(n_11483), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__u0 ( .ck(ispd_clk), .d(n_10417), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__u0 ( .ck(ispd_clk), .d(n_10416), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__u0 ( .ck(ispd_clk), .d(n_10414), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__u0 ( .ck(ispd_clk), .d(n_11482), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__u0 ( .ck(ispd_clk), .d(n_11480), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__u0 ( .ck(ispd_clk), .d(n_11479), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__u0 ( .ck(ispd_clk), .d(n_11698), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__u0 ( .ck(ispd_clk), .d(n_11697), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__u0 ( .ck(ispd_clk), .d(n_11696), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__u0 ( .ck(ispd_clk), .d(n_10515), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__u0 ( .ck(ispd_clk), .d(n_11695), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__u0 ( .ck(ispd_clk), .d(n_10513), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__u0 ( .ck(ispd_clk), .d(n_11694), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__u0 ( .ck(ispd_clk), .d(n_11693), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__u0 ( .ck(ispd_clk), .d(n_11692), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__u0 ( .ck(ispd_clk), .d(n_11691), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__u0 ( .ck(ispd_clk), .d(n_11690), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__u0 ( .ck(ispd_clk), .d(n_11689), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__u0 ( .ck(ispd_clk), .d(n_11688), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__u0 ( .ck(ispd_clk), .d(n_11687), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__u0 ( .ck(ispd_clk), .d(n_10511), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__u0 ( .ck(ispd_clk), .d(n_11686), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__u0 ( .ck(ispd_clk), .d(n_11685), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__u0 ( .ck(ispd_clk), .d(n_10509), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__u0 ( .ck(ispd_clk), .d(n_11684), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__u0 ( .ck(ispd_clk), .d(n_11683), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__u0 ( .ck(ispd_clk), .d(n_11682), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__u0 ( .ck(ispd_clk), .d(n_11681), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__u0 ( .ck(ispd_clk), .d(n_10508), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__u0 ( .ck(ispd_clk), .d(n_11680), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__u0 ( .ck(ispd_clk), .d(n_11679), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__u0 ( .ck(ispd_clk), .d(n_10848), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__u0 ( .ck(ispd_clk), .d(n_10847), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__u0 ( .ck(ispd_clk), .d(n_10506), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__u0 ( .ck(ispd_clk), .d(n_11708), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__u0 ( .ck(ispd_clk), .d(n_8916), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__u0 ( .ck(ispd_clk), .d(n_11677), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__u0 ( .ck(ispd_clk), .d(n_10503), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__u0 ( .ck(ispd_clk), .d(n_10501), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__u0 ( .ck(ispd_clk), .d(n_10499), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__u0 ( .ck(ispd_clk), .d(n_11676), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__8__u0 ( .ck(ispd_clk), .d(n_11675), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__u0 ( .ck(ispd_clk), .d(n_11674), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__u0 ( .ck(ispd_clk), .d(n_11336), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__u0 ( .ck(ispd_clk), .d(n_11334), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__u0 ( .ck(ispd_clk), .d(n_11332), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__u0 ( .ck(ispd_clk), .d(n_10365), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__u0 ( .ck(ispd_clk), .d(n_11330), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__u0 ( .ck(ispd_clk), .d(n_10363), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__u0 ( .ck(ispd_clk), .d(n_11328), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__u0 ( .ck(ispd_clk), .d(n_11327), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__u0 ( .ck(ispd_clk), .d(n_11324), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__u0 ( .ck(ispd_clk), .d(n_11326), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__u0 ( .ck(ispd_clk), .d(n_11322), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__u0 ( .ck(ispd_clk), .d(n_11320), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__u0 ( .ck(ispd_clk), .d(n_11318), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__u0 ( .ck(ispd_clk), .d(n_11316), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__u0 ( .ck(ispd_clk), .d(n_10362), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__u0 ( .ck(ispd_clk), .d(n_11314), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__u0 ( .ck(ispd_clk), .d(n_11311), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__u0 ( .ck(ispd_clk), .d(n_10361), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__u0 ( .ck(ispd_clk), .d(n_11309), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__u0 ( .ck(ispd_clk), .d(n_11307), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__u0 ( .ck(ispd_clk), .d(n_11306), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__u0 ( .ck(ispd_clk), .d(n_11305), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__u0 ( .ck(ispd_clk), .d(n_10359), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__u0 ( .ck(ispd_clk), .d(n_11303), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__u0 ( .ck(ispd_clk), .d(n_11302), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__u0 ( .ck(ispd_clk), .d(n_10823), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__u0 ( .ck(ispd_clk), .d(n_10821), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__u0 ( .ck(ispd_clk), .d(n_10357), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__u0 ( .ck(ispd_clk), .d(n_11300), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__36__u0 ( .ck(ispd_clk), .d(n_8955), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__36__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__36__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__36__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_11__465) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__u0 ( .ck(ispd_clk), .d(n_11297), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__u0 ( .ck(ispd_clk), .d(n_10355), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__u0 ( .ck(ispd_clk), .d(n_10353), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__u0 ( .ck(ispd_clk), .d(n_10351), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__u0 ( .ck(ispd_clk), .d(n_11295), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__u0 ( .ck(ispd_clk), .d(n_11293), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__u0 ( .ck(ispd_clk), .d(n_11290), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__u0 ( .ck(ispd_clk), .d(n_11672), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__u0 ( .ck(ispd_clk), .d(n_11671), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__u0 ( .ck(ispd_clk), .d(n_11670), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__u0 ( .ck(ispd_clk), .d(n_10497), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__u0 ( .ck(ispd_clk), .d(n_11669), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__u0 ( .ck(ispd_clk), .d(n_10495), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__u0 ( .ck(ispd_clk), .d(n_11668), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__u0 ( .ck(ispd_clk), .d(n_11667), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__u0 ( .ck(ispd_clk), .d(n_11666), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__u0 ( .ck(ispd_clk), .d(n_11665), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__u0 ( .ck(ispd_clk), .d(n_11663), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__u0 ( .ck(ispd_clk), .d(n_11662), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__u0 ( .ck(ispd_clk), .d(n_11660), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__u0 ( .ck(ispd_clk), .d(n_11661), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__u0 ( .ck(ispd_clk), .d(n_10493), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__u0 ( .ck(ispd_clk), .d(n_11659), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__u0 ( .ck(ispd_clk), .d(n_11657), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__u0 ( .ck(ispd_clk), .d(n_10491), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__u0 ( .ck(ispd_clk), .d(n_11655), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__u0 ( .ck(ispd_clk), .d(n_11653), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__u0 ( .ck(ispd_clk), .d(n_11652), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__u0 ( .ck(ispd_clk), .d(n_11651), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__u0 ( .ck(ispd_clk), .d(n_10489), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__u0 ( .ck(ispd_clk), .d(n_11650), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__u0 ( .ck(ispd_clk), .d(n_11648), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__u0 ( .ck(ispd_clk), .d(n_10845), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__u0 ( .ck(ispd_clk), .d(n_10843), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__u0 ( .ck(ispd_clk), .d(n_10487), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__u0 ( .ck(ispd_clk), .d(n_11707), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__u0 ( .ck(ispd_clk), .d(n_8914), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__u0 ( .ck(ispd_clk), .d(n_11647), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__u0 ( .ck(ispd_clk), .d(n_10485), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__u0 ( .ck(ispd_clk), .d(n_10483), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__u0 ( .ck(ispd_clk), .d(n_10481), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__u0 ( .ck(ispd_clk), .d(n_11645), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__u0 ( .ck(ispd_clk), .d(n_11644), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__u0 ( .ck(ispd_clk), .d(n_11642), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__u0 ( .ck(ispd_clk), .d(n_11289), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__10__u0 ( .ck(ispd_clk), .d(n_11287), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__u0 ( .ck(ispd_clk), .d(n_11286), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__u0 ( .ck(ispd_clk), .d(n_10349), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__u0 ( .ck(ispd_clk), .d(n_11285), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__u0 ( .ck(ispd_clk), .d(n_10348), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__u0 ( .ck(ispd_clk), .d(n_11284), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__u0 ( .ck(ispd_clk), .d(n_11283), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__u0 ( .ck(ispd_clk), .d(n_11282), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__u0 ( .ck(ispd_clk), .d(n_11281), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__u0 ( .ck(ispd_clk), .d(n_11280), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__u0 ( .ck(ispd_clk), .d(n_11279), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__u0 ( .ck(ispd_clk), .d(n_11277), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__u0 ( .ck(ispd_clk), .d(n_11276), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__22__u0 ( .ck(ispd_clk), .d(n_10346), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__u0 ( .ck(ispd_clk), .d(n_11274), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__u0 ( .ck(ispd_clk), .d(n_11273), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__u0 ( .ck(ispd_clk), .d(n_10344), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__u0 ( .ck(ispd_clk), .d(n_11271), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__u0 ( .ck(ispd_clk), .d(n_11270), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__u0 ( .ck(ispd_clk), .d(n_11268), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__u0 ( .ck(ispd_clk), .d(n_11266), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__u0 ( .ck(ispd_clk), .d(n_10343), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__u0 ( .ck(ispd_clk), .d(n_11265), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__u0 ( .ck(ispd_clk), .d(n_11264), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__u0 ( .ck(ispd_clk), .d(n_10820), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__u0 ( .ck(ispd_clk), .d(n_10819), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__u0 ( .ck(ispd_clk), .d(n_10342), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__u0 ( .ck(ispd_clk), .d(n_11262), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__36__u0 ( .ck(ispd_clk), .d(n_8900), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__36__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__36__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__36__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_13__543) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__u0 ( .ck(ispd_clk), .d(n_11261), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__u0 ( .ck(ispd_clk), .d(n_10340), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__u0 ( .ck(ispd_clk), .d(n_10338), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__u0 ( .ck(ispd_clk), .d(n_10336), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__u0 ( .ck(ispd_clk), .d(n_11260), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__u0 ( .ck(ispd_clk), .d(n_11259), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__u0 ( .ck(ispd_clk), .d(n_11258), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__u0 ( .ck(ispd_clk), .d(n_11256), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__u0 ( .ck(ispd_clk), .d(n_11255), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__u0 ( .ck(ispd_clk), .d(n_11254), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__u0 ( .ck(ispd_clk), .d(n_10334), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__u0 ( .ck(ispd_clk), .d(n_11252), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__u0 ( .ck(ispd_clk), .d(n_10332), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__u0 ( .ck(ispd_clk), .d(n_11251), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__u0 ( .ck(ispd_clk), .d(n_11250), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__u0 ( .ck(ispd_clk), .d(n_11249), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__u0 ( .ck(ispd_clk), .d(n_11247), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__u0 ( .ck(ispd_clk), .d(n_11246), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__u0 ( .ck(ispd_clk), .d(n_11245), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__u0 ( .ck(ispd_clk), .d(n_11244), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__u0 ( .ck(ispd_clk), .d(n_11243), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__u0 ( .ck(ispd_clk), .d(n_10331), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__u0 ( .ck(ispd_clk), .d(n_11242), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__u0 ( .ck(ispd_clk), .d(n_11241), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__u0 ( .ck(ispd_clk), .d(n_10329), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__u0 ( .ck(ispd_clk), .d(n_11240), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__u0 ( .ck(ispd_clk), .d(n_11239), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__u0 ( .ck(ispd_clk), .d(n_11238), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__u0 ( .ck(ispd_clk), .d(n_11236), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__u0 ( .ck(ispd_clk), .d(n_10327), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__u0 ( .ck(ispd_clk), .d(n_11235), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__u0 ( .ck(ispd_clk), .d(n_11234), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__u0 ( .ck(ispd_clk), .d(n_10817), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__u0 ( .ck(ispd_clk), .d(n_10815), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__u0 ( .ck(ispd_clk), .d(n_10325), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__u0 ( .ck(ispd_clk), .d(n_11232), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__36__u0 ( .ck(ispd_clk), .d(n_8899), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__36__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__36__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__36__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_14__582) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__u0 ( .ck(ispd_clk), .d(n_11230), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__u0 ( .ck(ispd_clk), .d(n_10323), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__u0 ( .ck(ispd_clk), .d(n_10321), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__u0 ( .ck(ispd_clk), .d(n_10319), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__u0 ( .ck(ispd_clk), .d(n_11229), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__u0 ( .ck(ispd_clk), .d(n_11228), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__u0 ( .ck(ispd_clk), .d(n_11226), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__u0 ( .ck(ispd_clk), .d(n_11224), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__u0 ( .ck(ispd_clk), .d(n_11223), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__u0 ( .ck(ispd_clk), .d(n_11222), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__u0 ( .ck(ispd_clk), .d(n_10317), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__u0 ( .ck(ispd_clk), .d(n_11220), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__u0 ( .ck(ispd_clk), .d(n_10316), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__u0 ( .ck(ispd_clk), .d(n_11219), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__u0 ( .ck(ispd_clk), .d(n_11218), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__u0 ( .ck(ispd_clk), .d(n_11217), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__u0 ( .ck(ispd_clk), .d(n_11216), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__u0 ( .ck(ispd_clk), .d(n_11215), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__u0 ( .ck(ispd_clk), .d(n_11214), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__u0 ( .ck(ispd_clk), .d(n_11213), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__u0 ( .ck(ispd_clk), .d(n_11212), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__22__u0 ( .ck(ispd_clk), .d(n_10314), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__u0 ( .ck(ispd_clk), .d(n_11211), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__u0 ( .ck(ispd_clk), .d(n_11209), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__u0 ( .ck(ispd_clk), .d(n_10312), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__u0 ( .ck(ispd_clk), .d(n_11208), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__u0 ( .ck(ispd_clk), .d(n_11207), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__u0 ( .ck(ispd_clk), .d(n_11206), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__u0 ( .ck(ispd_clk), .d(n_11205), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__u0 ( .ck(ispd_clk), .d(n_10311), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__u0 ( .ck(ispd_clk), .d(n_11203), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__u0 ( .ck(ispd_clk), .d(n_11202), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__u0 ( .ck(ispd_clk), .d(n_10813), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__u0 ( .ck(ispd_clk), .d(n_10812), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__u0 ( .ck(ispd_clk), .d(n_10310), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__u0 ( .ck(ispd_clk), .d(n_11200), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__36__u0 ( .ck(ispd_clk), .d(n_8898), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__36__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__36__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__36__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_15__621) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__u0 ( .ck(ispd_clk), .d(n_11198), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__u0 ( .ck(ispd_clk), .d(n_10308), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__u0 ( .ck(ispd_clk), .d(n_10306), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__u0 ( .ck(ispd_clk), .d(n_10304), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__u0 ( .ck(ispd_clk), .d(n_11196), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__8__u0 ( .ck(ispd_clk), .d(n_11194), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__u0 ( .ck(ispd_clk), .d(n_11193), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__u0 ( .ck(ispd_clk), .d(n_11478), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__u0 ( .ck(ispd_clk), .d(n_11477), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__u0 ( .ck(ispd_clk), .d(n_11476), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__u0 ( .ck(ispd_clk), .d(n_10413), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__u0 ( .ck(ispd_clk), .d(n_11474), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__u0 ( .ck(ispd_clk), .d(n_10412), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__u0 ( .ck(ispd_clk), .d(n_11473), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__u0 ( .ck(ispd_clk), .d(n_11472), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__u0 ( .ck(ispd_clk), .d(n_11470), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__u0 ( .ck(ispd_clk), .d(n_11468), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__u0 ( .ck(ispd_clk), .d(n_11467), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__u0 ( .ck(ispd_clk), .d(n_11466), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__u0 ( .ck(ispd_clk), .d(n_11464), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__u0 ( .ck(ispd_clk), .d(n_11463), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__u0 ( .ck(ispd_clk), .d(n_10411), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__u0 ( .ck(ispd_clk), .d(n_11462), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__u0 ( .ck(ispd_clk), .d(n_11460), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__u0 ( .ck(ispd_clk), .d(n_10410), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__u0 ( .ck(ispd_clk), .d(n_11458), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__u0 ( .ck(ispd_clk), .d(n_11457), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__u0 ( .ck(ispd_clk), .d(n_11456), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__29__u0 ( .ck(ispd_clk), .d(n_11454), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__u0 ( .ck(ispd_clk), .d(n_10408), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__u0 ( .ck(ispd_clk), .d(n_11451), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__u0 ( .ck(ispd_clk), .d(n_11452), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__u0 ( .ck(ispd_clk), .d(n_10810), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__u0 ( .ck(ispd_clk), .d(n_10807), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__u0 ( .ck(ispd_clk), .d(n_10302), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__u0 ( .ck(ispd_clk), .d(n_11706), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__u0 ( .ck(ispd_clk), .d(n_8912), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__u0 ( .ck(ispd_clk), .d(n_11449), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__u0 ( .ck(ispd_clk), .d(n_10407), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__u0 ( .ck(ispd_clk), .d(n_10405), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__u0 ( .ck(ispd_clk), .d(n_10404), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__u0 ( .ck(ispd_clk), .d(n_11446), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__u0 ( .ck(ispd_clk), .d(n_11445), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__u0 ( .ck(ispd_clk), .d(n_11443), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__u0 ( .ck(ispd_clk), .d(n_11442), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__u0 ( .ck(ispd_clk), .d(n_11441), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__u0 ( .ck(ispd_clk), .d(n_11440), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__u0 ( .ck(ispd_clk), .d(n_10402), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__u0 ( .ck(ispd_clk), .d(n_11438), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__u0 ( .ck(ispd_clk), .d(n_10401), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__u0 ( .ck(ispd_clk), .d(n_11437), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__u0 ( .ck(ispd_clk), .d(n_11436), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__u0 ( .ck(ispd_clk), .d(n_11435), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__u0 ( .ck(ispd_clk), .d(n_11431), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__u0 ( .ck(ispd_clk), .d(n_11434), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__u0 ( .ck(ispd_clk), .d(n_11433), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__u0 ( .ck(ispd_clk), .d(n_11432), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__u0 ( .ck(ispd_clk), .d(n_11429), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__u0 ( .ck(ispd_clk), .d(n_10400), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__u0 ( .ck(ispd_clk), .d(n_11427), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__u0 ( .ck(ispd_clk), .d(n_11425), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__u0 ( .ck(ispd_clk), .d(n_10399), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__u0 ( .ck(ispd_clk), .d(n_11424), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__u0 ( .ck(ispd_clk), .d(n_11423), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__u0 ( .ck(ispd_clk), .d(n_11421), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__u0 ( .ck(ispd_clk), .d(n_11420), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__u0 ( .ck(ispd_clk), .d(n_10397), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__u0 ( .ck(ispd_clk), .d(n_11419), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__u0 ( .ck(ispd_clk), .d(n_11418), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__u0 ( .ck(ispd_clk), .d(n_10806), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__u0 ( .ck(ispd_clk), .d(n_10804), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__u0 ( .ck(ispd_clk), .d(n_10300), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__u0 ( .ck(ispd_clk), .d(n_11705), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__u0 ( .ck(ispd_clk), .d(n_8910), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__u0 ( .ck(ispd_clk), .d(n_11417), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__u0 ( .ck(ispd_clk), .d(n_10396), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__u0 ( .ck(ispd_clk), .d(n_10394), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__u0 ( .ck(ispd_clk), .d(n_10393), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__u0 ( .ck(ispd_clk), .d(n_11415), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__u0 ( .ck(ispd_clk), .d(n_11414), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__u0 ( .ck(ispd_clk), .d(n_11413), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__u0 ( .ck(ispd_clk), .d(n_11641), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__u0 ( .ck(ispd_clk), .d(n_11640), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__u0 ( .ck(ispd_clk), .d(n_11639), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__u0 ( .ck(ispd_clk), .d(n_10479), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__u0 ( .ck(ispd_clk), .d(n_11638), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__u0 ( .ck(ispd_clk), .d(n_10478), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__u0 ( .ck(ispd_clk), .d(n_11637), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__u0 ( .ck(ispd_clk), .d(n_11635), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__u0 ( .ck(ispd_clk), .d(n_11634), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__u0 ( .ck(ispd_clk), .d(n_11631), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__u0 ( .ck(ispd_clk), .d(n_11633), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__u0 ( .ck(ispd_clk), .d(n_11632), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__u0 ( .ck(ispd_clk), .d(n_11630), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__u0 ( .ck(ispd_clk), .d(n_11628), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__u0 ( .ck(ispd_clk), .d(n_10477), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__u0 ( .ck(ispd_clk), .d(n_11626), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__u0 ( .ck(ispd_clk), .d(n_11625), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__u0 ( .ck(ispd_clk), .d(n_10476), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__u0 ( .ck(ispd_clk), .d(n_11624), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__u0 ( .ck(ispd_clk), .d(n_11623), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__u0 ( .ck(ispd_clk), .d(n_11622), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__u0 ( .ck(ispd_clk), .d(n_11620), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__u0 ( .ck(ispd_clk), .d(n_10474), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__u0 ( .ck(ispd_clk), .d(n_11618), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__u0 ( .ck(ispd_clk), .d(n_11617), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__u0 ( .ck(ispd_clk), .d(n_10841), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__u0 ( .ck(ispd_clk), .d(n_10839), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__u0 ( .ck(ispd_clk), .d(n_10473), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__u0 ( .ck(ispd_clk), .d(n_11712), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__u0 ( .ck(ispd_clk), .d(n_8908), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__u0 ( .ck(ispd_clk), .d(n_11616), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__u0 ( .ck(ispd_clk), .d(n_10469), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__u0 ( .ck(ispd_clk), .d(n_10470), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__u0 ( .ck(ispd_clk), .d(n_10467), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__u0 ( .ck(ispd_clk), .d(n_11614), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__u0 ( .ck(ispd_clk), .d(n_11613), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__u0 ( .ck(ispd_clk), .d(n_11611), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__u0 ( .ck(ispd_clk), .d(n_11411), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__u0 ( .ck(ispd_clk), .d(n_11410), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__u0 ( .ck(ispd_clk), .d(n_11408), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__u0 ( .ck(ispd_clk), .d(n_10391), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__u0 ( .ck(ispd_clk), .d(n_11406), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__u0 ( .ck(ispd_clk), .d(n_10390), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__u0 ( .ck(ispd_clk), .d(n_11405), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__u0 ( .ck(ispd_clk), .d(n_11403), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__u0 ( .ck(ispd_clk), .d(n_11402), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__18__u0 ( .ck(ispd_clk), .d(n_11401), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__18__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__18__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__18__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_4__213) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__u0 ( .ck(ispd_clk), .d(n_11399), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__u0 ( .ck(ispd_clk), .d(n_11398), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__u0 ( .ck(ispd_clk), .d(n_11396), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__u0 ( .ck(ispd_clk), .d(n_11394), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__u0 ( .ck(ispd_clk), .d(n_10388), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__u0 ( .ck(ispd_clk), .d(n_11393), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__u0 ( .ck(ispd_clk), .d(n_11391), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__u0 ( .ck(ispd_clk), .d(n_10386), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__u0 ( .ck(ispd_clk), .d(n_11390), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__u0 ( .ck(ispd_clk), .d(n_11388), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__u0 ( .ck(ispd_clk), .d(n_11386), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__u0 ( .ck(ispd_clk), .d(n_11385), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__u0 ( .ck(ispd_clk), .d(n_10385), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__u0 ( .ck(ispd_clk), .d(n_11384), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__u0 ( .ck(ispd_clk), .d(n_11383), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__u0 ( .ck(ispd_clk), .d(n_10803), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__u0 ( .ck(ispd_clk), .d(n_10802), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__34__u0 ( .ck(ispd_clk), .d(n_10298), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__u0 ( .ck(ispd_clk), .d(n_11703), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__u0 ( .ck(ispd_clk), .d(n_8906), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__u0 ( .ck(ispd_clk), .d(n_11382), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__u0 ( .ck(ispd_clk), .d(n_10384), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__u0 ( .ck(ispd_clk), .d(n_10383), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__u0 ( .ck(ispd_clk), .d(n_10381), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__u0 ( .ck(ispd_clk), .d(n_11381), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__u0 ( .ck(ispd_clk), .d(n_11380), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__u0 ( .ck(ispd_clk), .d(n_11379), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__u0 ( .ck(ispd_clk), .d(n_11610), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__u0 ( .ck(ispd_clk), .d(n_11609), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__u0 ( .ck(ispd_clk), .d(n_11607), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__u0 ( .ck(ispd_clk), .d(n_10465), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__u0 ( .ck(ispd_clk), .d(n_11606), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__u0 ( .ck(ispd_clk), .d(n_10464), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__u0 ( .ck(ispd_clk), .d(n_11605), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__u0 ( .ck(ispd_clk), .d(n_11604), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__u0 ( .ck(ispd_clk), .d(n_11603), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__u0 ( .ck(ispd_clk), .d(n_11602), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__u0 ( .ck(ispd_clk), .d(n_11601), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__u0 ( .ck(ispd_clk), .d(n_11600), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__u0 ( .ck(ispd_clk), .d(n_11599), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__u0 ( .ck(ispd_clk), .d(n_11598), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__u0 ( .ck(ispd_clk), .d(n_10463), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__u0 ( .ck(ispd_clk), .d(n_11597), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__u0 ( .ck(ispd_clk), .d(n_11595), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__u0 ( .ck(ispd_clk), .d(n_10462), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__u0 ( .ck(ispd_clk), .d(n_11593), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__u0 ( .ck(ispd_clk), .d(n_11592), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__u0 ( .ck(ispd_clk), .d(n_11590), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__u0 ( .ck(ispd_clk), .d(n_11589), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__u0 ( .ck(ispd_clk), .d(n_10460), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__u0 ( .ck(ispd_clk), .d(n_11588), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__u0 ( .ck(ispd_clk), .d(n_11587), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__u0 ( .ck(ispd_clk), .d(n_10838), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__u0 ( .ck(ispd_clk), .d(n_10836), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__u0 ( .ck(ispd_clk), .d(n_10459), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__u0 ( .ck(ispd_clk), .d(n_11702), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__u0 ( .ck(ispd_clk), .d(n_8904), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__u0 ( .ck(ispd_clk), .d(n_11586), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__u0 ( .ck(ispd_clk), .d(n_10457), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__u0 ( .ck(ispd_clk), .d(n_10455), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__u0 ( .ck(ispd_clk), .d(n_10453), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__u0 ( .ck(ispd_clk), .d(n_11585), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__u0 ( .ck(ispd_clk), .d(n_11584), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__u0 ( .ck(ispd_clk), .d(n_11583), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__u0 ( .ck(ispd_clk), .d(n_11582), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__10__u0 ( .ck(ispd_clk), .d(n_11580), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__u0 ( .ck(ispd_clk), .d(n_11579), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__u0 ( .ck(ispd_clk), .d(n_10451), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__u0 ( .ck(ispd_clk), .d(n_11577), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__u0 ( .ck(ispd_clk), .d(n_10450), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__15__u0 ( .ck(ispd_clk), .d(n_11575), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__u0 ( .ck(ispd_clk), .d(n_11573), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__u0 ( .ck(ispd_clk), .d(n_11572), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__18__u0 ( .ck(ispd_clk), .d(n_11571), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__18__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__18__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__18__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_6__252) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__u0 ( .ck(ispd_clk), .d(n_11570), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__u0 ( .ck(ispd_clk), .d(n_11568), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__u0 ( .ck(ispd_clk), .d(n_11566), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__u0 ( .ck(ispd_clk), .d(n_11565), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__u0 ( .ck(ispd_clk), .d(n_10449), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__u0 ( .ck(ispd_clk), .d(n_11564), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__u0 ( .ck(ispd_clk), .d(n_11562), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__u0 ( .ck(ispd_clk), .d(n_10447), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__u0 ( .ck(ispd_clk), .d(n_11561), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__u0 ( .ck(ispd_clk), .d(n_11560), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__u0 ( .ck(ispd_clk), .d(n_11559), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__u0 ( .ck(ispd_clk), .d(n_11557), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__u0 ( .ck(ispd_clk), .d(n_10446), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__u0 ( .ck(ispd_clk), .d(n_11556), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__31__u0 ( .ck(ispd_clk), .d(n_11555), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__u0 ( .ck(ispd_clk), .d(n_10835), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__u0 ( .ck(ispd_clk), .d(n_10834), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__u0 ( .ck(ispd_clk), .d(n_10445), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__u0 ( .ck(ispd_clk), .d(n_11701), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__u0 ( .ck(ispd_clk), .d(n_8902), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__u0 ( .ck(ispd_clk), .d(n_11553), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__u0 ( .ck(ispd_clk), .d(n_10444), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__u0 ( .ck(ispd_clk), .d(n_10443), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__u0 ( .ck(ispd_clk), .d(n_10440), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__u0 ( .ck(ispd_clk), .d(n_11551), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__8__u0 ( .ck(ispd_clk), .d(n_11549), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__u0 ( .ck(ispd_clk), .d(n_11548), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__u0 ( .ck(ispd_clk), .d(n_11191), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__u0 ( .ck(ispd_clk), .d(n_11190), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__u0 ( .ck(ispd_clk), .d(n_11188), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__u0 ( .ck(ispd_clk), .d(n_10297), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__u0 ( .ck(ispd_clk), .d(n_11187), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__u0 ( .ck(ispd_clk), .d(n_10296), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__15__u0 ( .ck(ispd_clk), .d(n_11186), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__u0 ( .ck(ispd_clk), .d(n_11184), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__u0 ( .ck(ispd_clk), .d(n_11182), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__18__u0 ( .ck(ispd_clk), .d(n_11181), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__18__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__18__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__18__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__291) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__u0 ( .ck(ispd_clk), .d(n_11180), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__u0 ( .ck(ispd_clk), .d(n_11179), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__u0 ( .ck(ispd_clk), .d(n_11178), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__u0 ( .ck(ispd_clk), .d(n_11177), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__u0 ( .ck(ispd_clk), .d(n_10294), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__u0 ( .ck(ispd_clk), .d(n_11175), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__u0 ( .ck(ispd_clk), .d(n_11174), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__u0 ( .ck(ispd_clk), .d(n_10292), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__u0 ( .ck(ispd_clk), .d(n_11173), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__u0 ( .ck(ispd_clk), .d(n_11171), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__u0 ( .ck(ispd_clk), .d(n_11169), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__29__u0 ( .ck(ispd_clk), .d(n_11167), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__u0 ( .ck(ispd_clk), .d(n_10291), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__u0 ( .ck(ispd_clk), .d(n_11165), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__31__u0 ( .ck(ispd_clk), .d(n_11337), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__u0 ( .ck(ispd_clk), .d(n_10800), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__u0 ( .ck(ispd_clk), .d(n_10799), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__u0 ( .ck(ispd_clk), .d(n_10290), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__u0 ( .ck(ispd_clk), .d(n_11164), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__36__u0 ( .ck(ispd_clk), .d(n_9188), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__36__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__36__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__36__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__309) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__u0 ( .ck(ispd_clk), .d(n_11162), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__u0 ( .ck(ispd_clk), .d(n_10289), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__u0 ( .ck(ispd_clk), .d(n_10288), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__u0 ( .ck(ispd_clk), .d(n_10286), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__u0 ( .ck(ispd_clk), .d(n_11161), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__8__u0 ( .ck(ispd_clk), .d(n_11159), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__u0 ( .ck(ispd_clk), .d(n_11158), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__u0 ( .ck(ispd_clk), .d(n_11377), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__u0 ( .ck(ispd_clk), .d(n_11375), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__u0 ( .ck(ispd_clk), .d(n_11373), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__u0 ( .ck(ispd_clk), .d(n_10380), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__u0 ( .ck(ispd_clk), .d(n_11372), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__u0 ( .ck(ispd_clk), .d(n_10378), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__u0 ( .ck(ispd_clk), .d(n_11370), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__u0 ( .ck(ispd_clk), .d(n_11369), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__u0 ( .ck(ispd_clk), .d(n_11367), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__u0 ( .ck(ispd_clk), .d(n_11365), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__u0 ( .ck(ispd_clk), .d(n_11363), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__u0 ( .ck(ispd_clk), .d(n_11362), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__u0 ( .ck(ispd_clk), .d(n_11361), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__u0 ( .ck(ispd_clk), .d(n_11359), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__u0 ( .ck(ispd_clk), .d(n_10377), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__u0 ( .ck(ispd_clk), .d(n_11357), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__u0 ( .ck(ispd_clk), .d(n_11355), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__u0 ( .ck(ispd_clk), .d(n_10376), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__u0 ( .ck(ispd_clk), .d(n_11353), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__u0 ( .ck(ispd_clk), .d(n_11352), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__u0 ( .ck(ispd_clk), .d(n_11350), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__u0 ( .ck(ispd_clk), .d(n_11349), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__u0 ( .ck(ispd_clk), .d(n_10374), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__u0 ( .ck(ispd_clk), .d(n_11347), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__u0 ( .ck(ispd_clk), .d(n_11345), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__u0 ( .ck(ispd_clk), .d(n_10797), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__u0 ( .ck(ispd_clk), .d(n_10795), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__u0 ( .ck(ispd_clk), .d(n_10285), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__u0 ( .ck(ispd_clk), .d(n_11700), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__u0 ( .ck(ispd_clk), .d(n_8957), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__u0 ( .ck(ispd_clk), .d(n_11344), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__u0 ( .ck(ispd_clk), .d(n_10372), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__u0 ( .ck(ispd_clk), .d(n_10370), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__u0 ( .ck(ispd_clk), .d(n_10368), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__u0 ( .ck(ispd_clk), .d(n_11342), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__u0 ( .ck(ispd_clk), .d(n_11340), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__u0 ( .ck(ispd_clk), .d(n_11338), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__u0 ( .ck(ispd_clk), .d(n_11547), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__u0 ( .ck(ispd_clk), .d(n_11546), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__u0 ( .ck(ispd_clk), .d(n_11545), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__u0 ( .ck(ispd_clk), .d(n_10439), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__u0 ( .ck(ispd_clk), .d(n_11544), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__u0 ( .ck(ispd_clk), .d(n_10438), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__u0 ( .ck(ispd_clk), .d(n_11543), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__u0 ( .ck(ispd_clk), .d(n_11542), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__u0 ( .ck(ispd_clk), .d(n_11540), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__u0 ( .ck(ispd_clk), .d(n_11538), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__u0 ( .ck(ispd_clk), .d(n_11536), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__u0 ( .ck(ispd_clk), .d(n_11535), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__u0 ( .ck(ispd_clk), .d(n_11534), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__u0 ( .ck(ispd_clk), .d(n_11533), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__u0 ( .ck(ispd_clk), .d(n_10436), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__u0 ( .ck(ispd_clk), .d(n_11532), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__u0 ( .ck(ispd_clk), .d(n_11531), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__u0 ( .ck(ispd_clk), .d(n_10434), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__u0 ( .ck(ispd_clk), .d(n_11530), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__u0 ( .ck(ispd_clk), .d(n_11528), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__u0 ( .ck(ispd_clk), .d(n_11526), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__u0 ( .ck(ispd_clk), .d(n_11524), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__u0 ( .ck(ispd_clk), .d(n_10433), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__u0 ( .ck(ispd_clk), .d(n_11521), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__u0 ( .ck(ispd_clk), .d(n_11523), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__u0 ( .ck(ispd_clk), .d(n_10833), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__u0 ( .ck(ispd_clk), .d(n_10832), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__u0 ( .ck(ispd_clk), .d(n_10432), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__u0 ( .ck(ispd_clk), .d(n_11699), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__u0 ( .ck(ispd_clk), .d(n_9191), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__u0 ( .ck(ispd_clk), .d(n_11519), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__u0 ( .ck(ispd_clk), .d(n_10430), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__u0 ( .ck(ispd_clk), .d(n_10428), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__u0 ( .ck(ispd_clk), .d(n_10426), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__u0 ( .ck(ispd_clk), .d(n_11517), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__8__u0 ( .ck(ispd_clk), .d(n_11516), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__u0 ( .ck(ispd_clk), .d(n_11515), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_0__u0 ( .ck(ispd_clk), .d(n_8917), .o(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_0__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_0__u1 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_0__Q), .o(wishbone_slave_unit_fifos_wbw_inTransactionCount_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_1__u0 ( .ck(ispd_clk), .d(n_9146), .o(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_1__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_1__u1 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_1__Q), .o(wishbone_slave_unit_fifos_wbw_inTransactionCount_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__u0 ( .ck(ispd_clk), .d(n_8921), .o(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_0__u0 ( .ck(ispd_clk), .d(n_8588), .o(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_0__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_0__u1 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_0__Q), .o(wishbone_slave_unit_fifos_wbw_outTransactionCount_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_1__u0 ( .ck(ispd_clk), .d(n_8669), .o(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_1__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_1__u1 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_1__Q), .o(wishbone_slave_unit_fifos_wbw_outTransactionCount_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__u0 ( .ck(ispd_clk), .d(n_8591), .o(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_bc_out_reg_0__u0 ( .ck(ispd_clk), .d(n_13499), .o(conf_wb_err_bc_in) );
ms00f80 wishbone_slave_unit_pci_initiator_if_bc_out_reg_1__u0 ( .ck(ispd_clk), .d(n_7714), .o(conf_wb_err_bc_in_846) );
ms00f80 wishbone_slave_unit_pci_initiator_if_bc_out_reg_2__u0 ( .ck(ispd_clk), .d(n_13502), .o(conf_wb_err_bc_in_847) );
ms00f80 wishbone_slave_unit_pci_initiator_if_bc_out_reg_3__u0 ( .ck(ispd_clk), .d(n_13500), .o(conf_wb_err_bc_in_848) );
ms00f80 wishbone_slave_unit_pci_initiator_if_be_out_reg_0__u0 ( .ck(ispd_clk), .d(n_13824), .o(n_1111) );
ms00f80 wishbone_slave_unit_pci_initiator_if_be_out_reg_1__u0 ( .ck(ispd_clk), .d(n_7212), .o(wishbone_slave_unit_pcim_sm_be_in_557) );
ms00f80 wishbone_slave_unit_pci_initiator_if_be_out_reg_2__u0 ( .ck(ispd_clk), .d(n_13827), .o(wishbone_slave_unit_pcim_sm_be_in_558) );
ms00f80 wishbone_slave_unit_pci_initiator_if_be_out_reg_3__u0 ( .ck(ispd_clk), .d(n_13826), .o(wishbone_slave_unit_pcim_sm_be_in_559) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_byte_address_reg_0__u0 ( .ck(ispd_clk), .d(n_13497), .o(wishbone_slave_unit_pci_initiator_if_current_byte_address) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_byte_address_reg_1__u0 ( .ck(ispd_clk), .d(n_13496), .o(wishbone_slave_unit_pci_initiator_if_current_byte_address_36) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_0__u0 ( .ck(ispd_clk), .d(n_13556), .o(conf_wb_err_addr_in_943) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_10__u0 ( .ck(ispd_clk), .d(n_13512), .o(conf_wb_err_addr_in_953) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_11__u0 ( .ck(ispd_clk), .d(n_13511), .o(conf_wb_err_addr_in_954) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_12__u0 ( .ck(ispd_clk), .d(n_13648), .o(conf_wb_err_addr_in_955) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_13__u0 ( .ck(ispd_clk), .d(n_13509), .o(conf_wb_err_addr_in_956) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_14__u0 ( .ck(ispd_clk), .d(n_13647), .o(conf_wb_err_addr_in_957) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_15__u0 ( .ck(ispd_clk), .d(n_13508), .o(conf_wb_err_addr_in_958) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_16__u0 ( .ck(ispd_clk), .d(n_13552), .o(conf_wb_err_addr_in_959) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_17__u0 ( .ck(ispd_clk), .d(n_13646), .o(conf_wb_err_addr_in_960) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_18__u0 ( .ck(ispd_clk), .d(n_13645), .o(conf_wb_err_addr_in_961) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_19__u0 ( .ck(ispd_clk), .d(n_13559), .o(conf_wb_err_addr_in_962) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_1__u0 ( .ck(ispd_clk), .d(n_13506), .o(conf_wb_err_addr_in_944) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_20__u0 ( .ck(ispd_clk), .d(n_13643), .o(conf_wb_err_addr_in_963) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_21__u0 ( .ck(ispd_clk), .d(n_13642), .o(conf_wb_err_addr_in_964) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_22__u0 ( .ck(ispd_clk), .d(n_13641), .o(conf_wb_err_addr_in_965) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_23__u0 ( .ck(ispd_clk), .d(n_13558), .o(conf_wb_err_addr_in_966) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_24__u0 ( .ck(ispd_clk), .d(n_13695), .o(conf_wb_err_addr_in_967) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_25__u0 ( .ck(ispd_clk), .d(n_13640), .o(conf_wb_err_addr_in_968) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_26__u0 ( .ck(ispd_clk), .d(n_13638), .o(conf_wb_err_addr_in_969) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_27__u0 ( .ck(ispd_clk), .d(n_13636), .o(conf_wb_err_addr_in_970) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_28__u0 ( .ck(ispd_clk), .d(n_13557), .o(conf_wb_err_addr_in_971) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__u0 ( .ck(ispd_clk), .d(n_13635), .o(wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_2__u0 ( .ck(ispd_clk), .d(n_13634), .o(conf_wb_err_addr_in_945) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_3__u0 ( .ck(ispd_clk), .d(n_13632), .o(conf_wb_err_addr_in_946) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_4__u0 ( .ck(ispd_clk), .d(n_13631), .o(conf_wb_err_addr_in_947) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_5__u0 ( .ck(ispd_clk), .d(n_13629), .o(conf_wb_err_addr_in_948) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_6__u0 ( .ck(ispd_clk), .d(n_13505), .o(conf_wb_err_addr_in_949) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_7__u0 ( .ck(ispd_clk), .d(n_13628), .o(conf_wb_err_addr_in_950) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_8__u0 ( .ck(ispd_clk), .d(n_13504), .o(conf_wb_err_addr_in_951) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_9__u0 ( .ck(ispd_clk), .d(n_13503), .o(conf_wb_err_addr_in_952) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_last_reg_u0 ( .ck(ispd_clk), .d(n_7539), .o(wishbone_slave_unit_pcim_sm_last_in) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_7783), .o(wishbone_slave_unit_pcim_sm_data_in) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_10__u0 ( .ck(ispd_clk), .d(n_7782), .o(wishbone_slave_unit_pcim_sm_data_in_644) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_11__u0 ( .ck(ispd_clk), .d(n_7781), .o(wishbone_slave_unit_pcim_sm_data_in_645) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_12__u0 ( .ck(ispd_clk), .d(n_7780), .o(wishbone_slave_unit_pcim_sm_data_in_646) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_13__u0 ( .ck(ispd_clk), .d(n_7779), .o(wishbone_slave_unit_pcim_sm_data_in_647) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_14__u0 ( .ck(ispd_clk), .d(n_7777), .o(wishbone_slave_unit_pcim_sm_data_in_648) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_15__u0 ( .ck(ispd_clk), .d(n_7776), .o(wishbone_slave_unit_pcim_sm_data_in_649) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_16__u0 ( .ck(ispd_clk), .d(n_7774), .o(wishbone_slave_unit_pcim_sm_data_in_650) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_17__u0 ( .ck(ispd_clk), .d(n_7773), .o(wishbone_slave_unit_pcim_sm_data_in_651) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_18__u0 ( .ck(ispd_clk), .d(n_7771), .o(wishbone_slave_unit_pcim_sm_data_in_652) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_19__u0 ( .ck(ispd_clk), .d(n_7769), .o(wishbone_slave_unit_pcim_sm_data_in_653) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_1__u0 ( .ck(ispd_clk), .d(n_7768), .o(wishbone_slave_unit_pcim_sm_data_in_635) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_20__u0 ( .ck(ispd_clk), .d(n_7767), .o(wishbone_slave_unit_pcim_sm_data_in_654) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_21__u0 ( .ck(ispd_clk), .d(n_7766), .o(wishbone_slave_unit_pcim_sm_data_in_655) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_22__u0 ( .ck(ispd_clk), .d(n_7764), .o(wishbone_slave_unit_pcim_sm_data_in_656) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_23__u0 ( .ck(ispd_clk), .d(n_7762), .o(wishbone_slave_unit_pcim_sm_data_in_657) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_24__u0 ( .ck(ispd_clk), .d(n_7761), .o(wishbone_slave_unit_pcim_sm_data_in_658) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_25__u0 ( .ck(ispd_clk), .d(n_7760), .o(wishbone_slave_unit_pcim_sm_data_in_659) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_26__u0 ( .ck(ispd_clk), .d(n_7759), .o(wishbone_slave_unit_pcim_sm_data_in_660) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_27__u0 ( .ck(ispd_clk), .d(n_7757), .o(wishbone_slave_unit_pcim_sm_data_in_661) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_28__u0 ( .ck(ispd_clk), .d(n_7756), .o(wishbone_slave_unit_pcim_sm_data_in_662) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_29__u0 ( .ck(ispd_clk), .d(n_7755), .o(wishbone_slave_unit_pcim_sm_data_in_663) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_2__u0 ( .ck(ispd_clk), .d(n_7754), .o(wishbone_slave_unit_pcim_sm_data_in_636) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_30__u0 ( .ck(ispd_clk), .d(n_7753), .o(wishbone_slave_unit_pcim_sm_data_in_664) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_31__u0 ( .ck(ispd_clk), .d(n_7752), .o(wishbone_slave_unit_pcim_sm_data_in_665) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_3__u0 ( .ck(ispd_clk), .d(n_7751), .o(wishbone_slave_unit_pcim_sm_data_in_637) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_4__u0 ( .ck(ispd_clk), .d(n_7750), .o(wishbone_slave_unit_pcim_sm_data_in_638) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_5__u0 ( .ck(ispd_clk), .d(n_7749), .o(wishbone_slave_unit_pcim_sm_data_in_639) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_6__u0 ( .ck(ispd_clk), .d(n_7747), .o(wishbone_slave_unit_pcim_sm_data_in_640) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_7__u0 ( .ck(ispd_clk), .d(n_7746), .o(wishbone_slave_unit_pcim_sm_data_in_641) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_8__u0 ( .ck(ispd_clk), .d(n_7745), .o(wishbone_slave_unit_pcim_sm_data_in_642) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_9__u0 ( .ck(ispd_clk), .d(n_7744), .o(wishbone_slave_unit_pcim_sm_data_in_643) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_source_reg_u0 ( .ck(ispd_clk), .d(n_4884), .o(wishbone_slave_unit_pci_initiator_if_data_source) );
ms00f80 wishbone_slave_unit_pci_initiator_if_del_read_req_reg_u0 ( .ck(ispd_clk), .d(n_8535), .o(wishbone_slave_unit_pci_initiator_if_del_read_req) );
ms00f80 wishbone_slave_unit_pci_initiator_if_del_write_req_reg_u0 ( .ck(ispd_clk), .d(n_4693), .o(wishbone_slave_unit_pci_initiator_if_del_write_req) );
ms00f80 wishbone_slave_unit_pci_initiator_if_err_recovery_reg_u0 ( .ck(ispd_clk), .d(n_7300), .o(wishbone_slave_unit_pci_initiator_if_err_recovery) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__u0 ( .ck(ispd_clk), .d(n_13550), .o(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__u0 ( .ck(ispd_clk), .d(n_7621), .o(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__u0 ( .ck(ispd_clk), .d(n_13546), .o(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__u0 ( .ck(ispd_clk), .d(n_13543), .o(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__u0 ( .ck(ispd_clk), .d(n_13540), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__u0 ( .ck(ispd_clk), .d(n_13539), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__u0 ( .ck(ispd_clk), .d(n_13538), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__u0 ( .ck(ispd_clk), .d(n_13537), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__u0 ( .ck(ispd_clk), .d(n_13536), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__u0 ( .ck(ispd_clk), .d(n_13535), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__u0 ( .ck(ispd_clk), .d(n_13534), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__u0 ( .ck(ispd_clk), .d(n_13533), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__u0 ( .ck(ispd_clk), .d(n_13532), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__u0 ( .ck(ispd_clk), .d(n_13531), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__u0 ( .ck(ispd_clk), .d(n_13530), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__u0 ( .ck(ispd_clk), .d(n_13529), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__u0 ( .ck(ispd_clk), .d(n_13528), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__u0 ( .ck(ispd_clk), .d(n_13470), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__u0 ( .ck(ispd_clk), .d(n_13527), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__u0 ( .ck(ispd_clk), .d(n_13526), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__u0 ( .ck(ispd_clk), .d(n_13525), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__u0 ( .ck(ispd_clk), .d(n_13469), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__u0 ( .ck(ispd_clk), .d(n_13627), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__u0 ( .ck(ispd_clk), .d(n_13524), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__u0 ( .ck(ispd_clk), .d(n_13523), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__u0 ( .ck(ispd_clk), .d(n_13522), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__u0 ( .ck(ispd_clk), .d(n_13521), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__u0 ( .ck(ispd_clk), .d(n_13468), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__u0 ( .ck(ispd_clk), .d(n_13520), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__u0 ( .ck(ispd_clk), .d(n_13519), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__u0 ( .ck(ispd_clk), .d(n_13518), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__u0 ( .ck(ispd_clk), .d(n_13517), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__u0 ( .ck(ispd_clk), .d(n_13516), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__u0 ( .ck(ispd_clk), .d(n_13515), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__u0 ( .ck(ispd_clk), .d(n_13514), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__u0 ( .ck(ispd_clk), .d(n_13513), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_last_reg_u0 ( .ck(ispd_clk), .d(n_7625), .o(n_16763) );
ms00f80 wishbone_slave_unit_pci_initiator_if_last_transfered_reg_u0 ( .ck(ispd_clk), .d(n_3081), .o(wishbone_slave_unit_fifos_wbr_control_in) );
ms00f80 wishbone_slave_unit_pci_initiator_if_posted_write_req_reg_u0 ( .ck(ispd_clk), .d(n_7028), .o(wishbone_slave_unit_pci_initiator_if_posted_write_req) );
ms00f80 wishbone_slave_unit_pci_initiator_if_rdy_out_reg_u0 ( .ck(ispd_clk), .d(n_2801), .o(wishbone_slave_unit_pcim_sm_rdy_in) );
ms00f80 wishbone_slave_unit_pci_initiator_if_read_bound_reg_u0 ( .ck(ispd_clk), .d(n_4870), .o(wishbone_slave_unit_pci_initiator_if_read_bound) );
ms00f80 wishbone_slave_unit_pci_initiator_if_read_count_reg_0__u0 ( .ck(ispd_clk), .d(n_4861), .o(wishbone_slave_unit_pci_initiator_if_read_count_0_) );
ms00f80 wishbone_slave_unit_pci_initiator_if_read_count_reg_1__u0 ( .ck(ispd_clk), .d(n_4860), .o(wishbone_slave_unit_pci_initiator_if_read_count_1_) );
ms00f80 wishbone_slave_unit_pci_initiator_if_read_count_reg_2__u0 ( .ck(ispd_clk), .d(n_7333), .o(wishbone_slave_unit_pci_initiator_if_read_count_2_) );
ms00f80 wishbone_slave_unit_pci_initiator_if_read_count_reg_3__u0 ( .ck(ispd_clk), .d(n_7544), .o(wishbone_slave_unit_pci_initiator_if_read_count_reg_3__Q) );
in01s01 wishbone_slave_unit_pci_initiator_if_read_count_reg_3__u1 ( .a(wishbone_slave_unit_pci_initiator_if_read_count_reg_3__Q), .o(wishbone_slave_unit_pci_initiator_if_read_count_3_) );
ms00f80 wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg_u0 ( .ck(ispd_clk), .d(n_3119), .o(wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg_Q) );
in01s01 wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg_u1 ( .a(wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg_Q), .o(conf_target_abort_recv_in) );
ms00f80 wishbone_slave_unit_pci_initiator_if_write_req_int_reg_u0 ( .ck(ispd_clk), .d(n_15859), .o(wishbone_slave_unit_pci_initiator_if_write_req_int) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_cur_state_reg_0__u0 ( .ck(ispd_clk), .d(n_7617), .o(wishbone_slave_unit_pci_initiator_sm_cur_state_0_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_cur_state_reg_1__u0 ( .ck(ispd_clk), .d(n_7616), .o(wishbone_slave_unit_pci_initiator_sm_cur_state_1_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_cur_state_reg_2__u0 ( .ck(ispd_clk), .d(n_7620), .o(wishbone_slave_unit_pci_initiator_sm_cur_state_2_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_cur_state_reg_3__u0 ( .ck(ispd_clk), .d(n_7619), .o(wishbone_slave_unit_pci_initiator_sm_cur_state_3_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_decode_count_reg_0__u0 ( .ck(ispd_clk), .d(n_4537), .o(wishbone_slave_unit_pci_initiator_sm_decode_count_0_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_decode_count_reg_1__u0 ( .ck(ispd_clk), .d(n_4534), .o(wishbone_slave_unit_pci_initiator_sm_decode_count_1_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_decode_count_reg_2__u0 ( .ck(ispd_clk), .d(n_4746), .o(wishbone_slave_unit_pci_initiator_sm_decode_count_2_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_0__u0 ( .ck(ispd_clk), .d(n_6982), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_0_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_1__u0 ( .ck(ispd_clk), .d(n_6984), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_1_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_2__u0 ( .ck(ispd_clk), .d(n_6987), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_2_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_3__u0 ( .ck(ispd_clk), .d(n_5748), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_3_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_4__u0 ( .ck(ispd_clk), .d(n_5644), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_4_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_5__u0 ( .ck(ispd_clk), .d(n_6985), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_5_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_6__u0 ( .ck(ispd_clk), .d(n_5713), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_6_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_7__u0 ( .ck(ispd_clk), .d(n_4892), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_7_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_mabort1_reg_u0 ( .ck(ispd_clk), .d(n_2684), .o(wishbone_slave_unit_pci_initiator_sm_mabort1) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_mabort2_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_pci_initiator_sm_mabort1), .o(wishbone_slave_unit_pci_initiator_sm_mabort2) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg_0__u0 ( .ck(ispd_clk), .d(n_7615), .o(wishbone_slave_unit_pci_initiator_sm_rdata_selector) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg_1__u0 ( .ck(ispd_clk), .d(n_7614), .o(wishbone_slave_unit_pci_initiator_sm_rdata_selector_14) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_timeout_reg_u0 ( .ck(ispd_clk), .d(n_4679), .o(wishbone_slave_unit_pci_initiator_sm_timeout) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_transfer_reg_u0 ( .ck(ispd_clk), .d(n_3812), .o(wishbone_slave_unit_pci_initiator_sm_transfer) );
ms00f80 wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg_u0 ( .ck(ispd_clk), .d(n_14483), .o(wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg_Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_c_state_reg_0__u0 ( .ck(ispd_clk), .d(n_14628), .o(wishbone_slave_unit_wishbone_slave_c_state) );
ms00f80 wishbone_slave_unit_wishbone_slave_c_state_reg_1__u0 ( .ck(ispd_clk), .d(n_7330), .o(wishbone_slave_unit_wishbone_slave_c_state_1) );
ms00f80 wishbone_slave_unit_wishbone_slave_c_state_reg_2__u0 ( .ck(ispd_clk), .d(n_14619), .o(wishbone_slave_unit_wishbone_slave_c_state_2) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_0__u0 ( .ck(ispd_clk), .d(n_8641), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_0__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_10__u0 ( .ck(ispd_clk), .d(n_8640), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_10__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_11__u0 ( .ck(ispd_clk), .d(n_8638), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_11__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_12__u0 ( .ck(ispd_clk), .d(n_8637), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_12__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_13__u0 ( .ck(ispd_clk), .d(n_8636), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_13__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_14__u0 ( .ck(ispd_clk), .d(n_8635), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_14__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_15__u0 ( .ck(ispd_clk), .d(n_8634), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_15__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_16__u0 ( .ck(ispd_clk), .d(n_8633), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_16__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_17__u0 ( .ck(ispd_clk), .d(n_8632), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_17__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_18__u0 ( .ck(ispd_clk), .d(n_8631), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_18__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_19__u0 ( .ck(ispd_clk), .d(n_8630), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_19__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_1__u0 ( .ck(ispd_clk), .d(n_8629), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_1__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_20__u0 ( .ck(ispd_clk), .d(n_8628), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_20__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_21__u0 ( .ck(ispd_clk), .d(n_8627), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_21__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_22__u0 ( .ck(ispd_clk), .d(n_8626), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_22__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_23__u0 ( .ck(ispd_clk), .d(n_8625), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_23__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_24__u0 ( .ck(ispd_clk), .d(n_8624), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_24__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_25__u0 ( .ck(ispd_clk), .d(n_8623), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_25__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_26__u0 ( .ck(ispd_clk), .d(n_8622), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_26__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_27__u0 ( .ck(ispd_clk), .d(n_8621), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_27__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_28__u0 ( .ck(ispd_clk), .d(n_8620), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_28__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_29__u0 ( .ck(ispd_clk), .d(n_8619), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_29__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_2__u0 ( .ck(ispd_clk), .d(n_8618), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_2__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_30__u0 ( .ck(ispd_clk), .d(n_8617), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_30__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_31__u0 ( .ck(ispd_clk), .d(n_8616), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_31__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_32__u0 ( .ck(ispd_clk), .d(n_8615), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_32__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_33__u0 ( .ck(ispd_clk), .d(n_8613), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_33__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_34__u0 ( .ck(ispd_clk), .d(n_8611), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_34__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_35__u0 ( .ck(ispd_clk), .d(n_8609), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_35__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_3__u0 ( .ck(ispd_clk), .d(n_8607), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_3__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_4__u0 ( .ck(ispd_clk), .d(n_8606), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_4__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_5__u0 ( .ck(ispd_clk), .d(n_8605), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_5__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_6__u0 ( .ck(ispd_clk), .d(n_8604), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_6__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_7__u0 ( .ck(ispd_clk), .d(n_8603), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_7__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_8__u0 ( .ck(ispd_clk), .d(n_8602), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_8__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_9__u0 ( .ck(ispd_clk), .d(n_8601), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_9__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_del_addr_hit_reg_u0 ( .ck(ispd_clk), .d(n_7723), .o(wishbone_slave_unit_wishbone_slave_del_addr_hit) );
ms00f80 wishbone_slave_unit_wishbone_slave_del_completion_allow_reg_u0 ( .ck(ispd_clk), .d(n_7701), .o(wishbone_slave_unit_wishbone_slave_del_completion_allow) );
ms00f80 wishbone_slave_unit_wishbone_slave_do_del_request_reg_u0 ( .ck(ispd_clk), .d(n_7722), .o(wishbone_slave_unit_wishbone_slave_do_del_request) );
ms00f80 wishbone_slave_unit_wishbone_slave_img_hit_reg_0__u0 ( .ck(ispd_clk), .d(n_7541), .o(wishbone_slave_unit_wishbone_slave_img_hit_0_) );
ms00f80 wishbone_slave_unit_wishbone_slave_img_hit_reg_1__u0 ( .ck(ispd_clk), .d(n_7540), .o(wishbone_slave_unit_wishbone_slave_img_hit_1_) );
ms00f80 wishbone_slave_unit_wishbone_slave_img_hit_reg_2__u0 ( .ck(ispd_clk), .d(n_5741), .o(wishbone_slave_unit_wishbone_slave_img_hit_2_) );
ms00f80 wishbone_slave_unit_wishbone_slave_img_hit_reg_3__u0 ( .ck(ispd_clk), .d(n_5740), .o(wishbone_slave_unit_wishbone_slave_img_hit_3_) );
ms00f80 wishbone_slave_unit_wishbone_slave_img_hit_reg_4__u0 ( .ck(ispd_clk), .d(n_5733), .o(wishbone_slave_unit_wishbone_slave_img_hit_4_) );
ms00f80 wishbone_slave_unit_wishbone_slave_img_wallow_reg_u0 ( .ck(ispd_clk), .d(n_7721), .o(wishbone_slave_unit_wishbone_slave_img_wallow) );
ms00f80 wishbone_slave_unit_wishbone_slave_map_reg_u0 ( .ck(ispd_clk), .d(n_7542), .o(wishbone_slave_unit_wishbone_slave_map) );
ms00f80 wishbone_slave_unit_wishbone_slave_mrl_en_reg_u0 ( .ck(ispd_clk), .d(n_7719), .o(wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_pref_en_reg_u0 ( .ck(ispd_clk), .d(n_7718), .o(wishbone_slave_unit_wishbone_slave_pref_en_reg_Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_wb_conf_hit_reg_u0 ( .ck(ispd_clk), .d(n_5736), .o(wishbone_slave_unit_wishbone_slave_wb_conf_hit) );
ms00f80 wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg_u0 ( .ck(ispd_clk), .d(n_8525), .o(wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg_Q) );
in01s40 wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg_u1 ( .a(wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg_Q), .o(n_8831) );
in01s06 TIMEBOOST_cell_0 ( .a(TIMEBOOST_net_0), .o(FE_OFN1094_g64577_p) );
in01s02 TIMEBOOST_cell_1 ( .a(TIMEBOOST_net_1), .o(TIMEBOOST_net_0) );
in01f08 TIMEBOOST_cell_2 ( .a(TIMEBOOST_net_2), .o(FE_OFN1061_n_16720) );
in01f04 TIMEBOOST_cell_3 ( .a(TIMEBOOST_net_3), .o(TIMEBOOST_net_2) );
in01f10 TIMEBOOST_cell_4 ( .a(TIMEBOOST_net_4), .o(FE_OCPN1845_n_16427) );
in01f06 TIMEBOOST_cell_5 ( .a(TIMEBOOST_net_5), .o(TIMEBOOST_net_4) );
na02f02 TIMEBOOST_cell_41490 ( .a(TIMEBOOST_net_12983), .b(g57369_sb), .o(n_11381) );

endmodule
