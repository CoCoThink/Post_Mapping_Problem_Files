module s1196 (
G1,
G11,
G8,
G5,
G9,
G3,
G13,
G4,
G12,
G2,
blif_clk_net,
G7,
blif_reset_net,
G10,
G0,
G6,
G549,
G542,
G530,
G552,
G45,
G547,
G548,
G537,
G551,
G532,
G539,
G546,
G535,
G550
);

// Start PIs
input G1;
input G11;
input G8;
input G5;
input G9;
input G3;
input G13;
input G4;
input G12;
input G2;
input blif_clk_net;
input G7;
input blif_reset_net;
input G10;
input G0;
input G6;

// Start POs
output G549;
output G542;
output G530;
output G552;
output G45;
output G547;
output G548;
output G537;
output G551;
output G532;
output G539;
output G546;
output G535;
output G550;

// Start wires
wire G1;
wire G11;
wire G8;
wire G5;
wire G9;
wire G3;
wire G13;
wire G4;
wire G12;
wire G2;
wire blif_clk_net;
wire G7;
wire blif_reset_net;
wire G10;
wire G0;
wire G6;
wire G549;
wire G542;
wire G530;
wire G552;
wire G45;
wire G547;
wire G548;
wire G537;
wire G551;
wire G532;
wire G539;
wire G546;
wire G535;
wire G550;
wire net_568;
wire net_47;
wire net_416;
wire net_215;
wire net_54;
wire net_526;
wire net_429;
wire net_557;
wire net_129;
wire net_373;
wire net_119;
wire net_98;
wire net_151;
wire net_356;
wire net_53;
wire net_452;
wire net_210;
wire TIMEBOOST_net_18;
wire net_284;
wire net_168;
wire net_560;
wire net_477;
wire net_439;
wire net_385;
wire net_259;
wire net_269;
wire net_548;
wire net_469;
wire net_501;
wire net_187;
wire net_111;
wire net_264;
wire net_90;
wire net_225;
wire net_283;
wire net_85;
wire net_263;
wire TIMEBOOST_net_54;
wire net_124;
wire net_404;
wire net_240;
wire net_160;
wire TIMEBOOST_net_55;
wire net_511;
wire net_4;
wire net_420;
wire TIMEBOOST_net_26;
wire net_295;
wire net_410;
wire net_508;
wire net_390;
wire net_307;
wire net_35;
wire net_586;
wire net_344;
wire net_16;
wire net_239;
wire net_193;
wire net_257;
wire net_310;
wire net_233;
wire net_474;
wire net_120;
wire net_292;
wire net_201;
wire net_472;
wire net_109;
wire net_80;
wire net_65;
wire net_96;
wire net_484;
wire net_167;
wire net_207;
wire net_136;
wire net_280;
wire net_126;
wire net_495;
wire net_278;
wire net_34;
wire net_458;
wire net_108;
wire net_598;
wire net_571;
wire net_63;
wire net_593;
wire net_617;
wire net_601;
wire net_274;
wire net_554;
wire net_425;
wire net_321;
wire net_287;
wire net_189;
wire net_490;
wire net_99;
wire net_46;
wire net_480;
wire net_216;
wire net_433;
wire net_584;
wire net_544;
wire net_368;
wire net_224;
wire net_52;
wire net_538;
wire net_165;
wire net_608;
wire net_510;
wire net_370;
wire net_464;
wire net_366;
wire net_13;
wire net_413;
wire net_446;
wire net_114;
wire net_248;
wire net_384;
wire net_36;
wire net_198;
wire net_253;
wire net_311;
wire net_276;
wire net_494;
wire net_209;
wire net_3;
wire net_547;
wire net_294;
wire net_154;
wire net_507;
wire net_616;
wire net_238;
wire net_529;
wire net_28;
wire net_587;
wire net_485;
wire net_97;
wire net_192;
wire net_503;
wire net_256;
wire net_460;
wire net_82;
wire net_64;
wire net_457;
wire net_291;
wire net_121;
wire net_597;
wire net_200;
wire net_308;
wire net_75;
wire net_515;
wire net_600;
wire net_396;
wire net_206;
wire net_195;
wire net_125;
wire net_397;
wire net_107;
wire net_166;
wire net_223;
wire net_235;
wire net_530;
wire net_606;
wire net_623;
wire net_603;
wire net_594;
wire net_320;
wire net_271;
wire net_23;
wire net_117;
wire net_74;
wire net_579;
wire net_401;
wire net_250;
wire net_205;
wire net_242;
wire net_312;
wire net_130;
wire net_572;
wire net_359;
wire TIMEBOOST_net_25;
wire net_286;
wire net_147;
wire net_481;
wire net_369;
wire net_470;
wire net_26;
wire net_403;
wire net_334;
wire net_32;
wire net_430;
wire net_365;
wire net_282;
wire net_426;
wire net_380;
wire net_141;
wire TIMEBOOST_net_28;
wire net_83;
wire net_609;
wire TIMEBOOST_net_24;
wire net_414;
wire net_372;
wire net_437;
wire net_528;
wire net_56;
wire net_566;
wire net_456;
wire net_155;
wire net_335;
wire net_506;
wire TIMEBOOST_net_52;
wire net_336;
wire net_624;
wire net_349;
wire net_39;
wire net_555;
wire net_245;
wire net_2;
wire net_9;
wire net_395;
wire net_331;
wire net_298;
wire net_493;
wire net_475;
wire net_563;
wire net_386;
wire net_605;
wire TIMEBOOST_net_19;
wire net_199;
wire net_502;
wire net_431;
wire net_89;
wire net_290;
wire net_338;
wire net_243;
wire net_400;
wire net_222;
wire net_602;
wire net_313;
wire net_152;
wire net_489;
wire net_175;
wire net_106;
wire net_607;
wire net_258;
wire net_140;
wire net_247;
wire TIMEBOOST_net_56;
wire net_279;
wire net_148;
wire net_419;
wire net_25;
wire net_70;
wire net_251;
wire net_194;
wire net_615;
wire net_478;
wire net_244;
wire net_585;
wire net_441;
wire net_128;
wire net_596;
wire net_138;
wire net_333;
wire net_549;
wire net_374;
wire net_411;
wire net_170;
wire net_531;
wire net_471;
wire net_565;
wire net_499;
wire net_77;
wire net_214;
wire TIMEBOOST_net_14;
wire net_20;
wire net_49;
wire net_518;
wire net_15;
wire net_57;
wire net_71;
wire net_156;
wire net_394;
wire net_92;
wire net_1;
wire net_112;
wire net_139;
wire net_551;
wire net_537;
wire net_332;
wire net_180;
wire net_409;
wire net_367;
wire net_169;
wire net_51;
wire net_171;
wire net_492;
wire net_463;
wire net_432;
wire net_88;
wire net_197;
wire net_513;
wire net_204;
wire net_81;
wire net_604;
wire net_163;
wire net_402;
wire net_67;
wire TIMEBOOST_net_13;
wire net_268;
wire net_110;
wire net_459;
wire net_483;
wire net_48;
wire net_33;
wire net_8;
wire net_203;
wire net_450;
wire TIMEBOOST_net_12;
wire net_505;
wire net_621;
wire TIMEBOOST_net_27;
wire net_176;
wire net_137;
wire net_296;
wire net_132;
wire net_613;
wire net_237;
wire net_105;
wire net_614;
wire net_532;
wire net_12;
wire net_93;
wire net_578;
wire net_302;
wire net_569;
wire net_127;
wire net_327;
wire TIMEBOOST_net_16;
wire net_348;
wire net_76;
wire net_626;
wire net_101;
wire net_388;
wire net_326;
wire TIMEBOOST_net_23;
wire net_589;
wire net_519;
wire net_100;
wire net_412;
wire net_536;
wire net_455;
wire net_221;
wire net_115;
wire net_393;
wire net_442;
wire net_17;
wire net_319;
wire net_542;
wire net_575;
wire net_595;
wire net_581;
wire net_378;
wire net_164;
wire net_408;
wire net_377;
wire net_87;
wire net_0;
wire TIMEBOOST_net_53;
wire TIMEBOOST_net_57;
wire net_328;
wire net_157;
wire net_540;
wire net_512;
wire net_42;
wire net_50;
wire net_234;
wire net_38;
wire net_66;
wire TIMEBOOST_net_29;
wire net_342;
wire net_612;
wire net_19;
wire net_443;
wire net_504;
wire net_522;
wire net_270;
wire net_183;
wire net_618;
wire net_150;
wire net_303;
wire TIMEBOOST_net_21;
wire net_352;
wire net_491;
wire net_30;
wire net_436;
wire net_24;
wire net_392;
wire net_622;
wire net_186;
wire TIMEBOOST_net_11;
wire TIMEBOOST_net_58;
wire net_146;
wire net_550;
wire net_122;
wire net_417;
wire net_7;
wire net_172;
wire net_94;
wire net_246;
wire net_461;
wire net_219;
wire net_18;
wire net_309;
wire net_482;
wire net_131;
wire net_196;
wire net_29;
wire net_358;
wire net_142;
wire net_149;
wire net_516;
wire net_31;
wire net_387;
wire net_330;
wire net_535;
wire net_498;
wire net_158;
wire net_41;
wire net_577;
wire net_360;
wire net_570;
wire net_525;
wire net_444;
wire net_213;
wire net_325;
wire TIMEBOOST_net_20;
wire net_260;
wire net_299;
wire net_438;
wire net_580;
wire net_314;
wire net_182;
wire net_521;
wire net_60;
wire net_590;
wire net_337;
wire net_267;
wire net_273;
wire net_424;
wire net_468;
wire net_58;
wire net_576;
wire net_488;
wire net_73;
wire net_86;
wire net_177;
wire net_523;
wire net_407;
wire net_476;
wire net_564;
wire net_382;
wire net_179;
wire net_159;
wire net_61;
wire net_583;
wire net_449;
wire net_383;
wire net_62;
wire net_6;
wire net_553;
wire net_534;
wire net_217;
wire net_351;
wire net_427;
wire net_486;
wire net_135;
wire net_340;
wire net_265;
wire net_517;
wire net_434;
wire net_406;
wire net_220;
wire net_14;
wire net_293;
wire net_324;
wire net_113;
wire net_497;
wire net_454;
wire net_418;
wire net_462;
wire net_40;
wire net_69;
wire net_543;
wire net_161;
wire net_625;
wire net_300;
wire net_339;
wire net_95;
wire net_173;
wire net_361;
wire net_78;
wire net_27;
wire net_317;
wire net_305;
wire net_514;
wire net_191;
wire net_261;
wire net_22;
wire TIMEBOOST_net_22;
wire net_558;
wire net_354;
wire net_524;
wire net_144;
wire net_102;
wire net_227;
wire net_59;
wire net_363;
wire net_445;
wire net_573;
wire net_162;
wire net_44;
wire net_230;
wire net_520;
wire net_422;
wire net_134;
wire net_546;
wire net_561;
wire net_567;
wire net_45;
wire net_381;
wire net_591;
wire net_185;
wire net_588;
wire net_272;
wire net_178;
wire TIMEBOOST_net_15;
wire net_236;
wire TIMEBOOST_net_10;
wire net_212;
wire net_315;
wire net_552;
wire net_415;
wire net_116;
wire net_556;
wire net_347;
wire net_91;
wire net_297;
wire net_346;
wire net_55;
wire net_559;
wire net_255;
wire net_266;
wire net_345;
wire net_104;
wire net_620;
wire net_448;
wire net_619;
wire net_72;
wire net_350;
wire net_229;
wire net_398;
wire net_306;
wire net_241;
wire net_5;
wire net_405;
wire net_500;
wire net_355;
wire net_184;
wire net_599;
wire net_11;
wire net_610;
wire net_123;
wire net_527;
wire net_262;
wire net_362;
wire net_389;
wire net_68;
wire net_318;
wire net_451;
wire net_323;
wire net_275;
wire net_539;
wire net_399;
wire net_153;
wire net_316;
wire net_218;
wire net_84;
wire net_174;
wire net_611;
wire net_231;
wire net_562;
wire net_103;
wire net_375;
wire TIMEBOOST_net_17;
wire net_364;
wire net_43;
wire net_10;
wire net_228;
wire net_592;
wire net_21;
wire net_79;
wire net_143;
wire net_190;
wire net_391;
wire net_533;
wire net_145;
wire net_285;
wire net_281;
wire net_254;
wire net_37;
wire net_582;
wire net_188;
wire net_496;
wire net_509;
wire net_574;
wire net_479;
wire net_211;
wire net_133;
wire TIMEBOOST_net_0;
wire TIMEBOOST_net_1;
wire TIMEBOOST_net_2;
wire TIMEBOOST_net_3;
wire TIMEBOOST_net_4;
wire TIMEBOOST_net_5;
wire TIMEBOOST_net_6;
wire TIMEBOOST_net_7;
wire TIMEBOOST_net_8;
wire TIMEBOOST_net_9;
wire TIMEBOOST_net_30;
wire TIMEBOOST_net_31;
wire TIMEBOOST_net_32;
wire TIMEBOOST_net_33;
wire TIMEBOOST_net_34;
wire TIMEBOOST_net_35;
wire TIMEBOOST_net_36;
wire TIMEBOOST_net_37;
wire TIMEBOOST_net_38;
wire TIMEBOOST_net_39;
wire TIMEBOOST_net_40;
wire TIMEBOOST_net_41;
wire TIMEBOOST_net_42;
wire TIMEBOOST_net_43;
wire TIMEBOOST_net_44;
wire TIMEBOOST_net_45;
wire TIMEBOOST_net_46;
wire TIMEBOOST_net_47;
wire TIMEBOOST_net_48;
wire TIMEBOOST_net_49;
wire TIMEBOOST_net_50;
wire TIMEBOOST_net_51;

// Start cells
INV_X1 inst_537 ( .A(net_244), .ZN(net_245) );
INV_X1 inst_481 ( .A(net_195), .ZN(net_162) );
DFFR_X1 inst_551 ( .D(net_264), .RN(net_464), .CK(TIMEBOOST_net_8), .Q(net_8) );
NAND2_X1 inst_228 ( .A1(net_22), .A2(net_50), .ZN(net_141) );
NAND4_X1 inst_125 ( .A1(net_479), .A2(net_429), .A3(net_480), .A4(net_438), .ZN(net_568) );
INV_X2 inst_486 ( .A(net_227), .ZN(net_220) );
INV_X1 inst_506 ( .A(net_536), .ZN(net_535) );
INV_X4 inst_495 ( .A(net_374), .ZN(net_381) );
INV_X2 inst_353 ( .A(net_562), .ZN(net_561) );
NAND3_X1 inst_159 ( .A1(net_151), .A2(net_527), .A3(net_522), .ZN(net_481) );
INV_X16 inst_395 ( .A(G7), .ZN(net_478) );
NAND3_X1 inst_134 ( .A1(net_53), .A2(net_133), .A3(net_519), .ZN(net_144) );
NAND2_X1 inst_244 ( .A1(net_99), .A2(net_148), .ZN(net_173) );
NOR2_X1 TIMEBOOST_cell_42 ( .A1(net_335), .A2(net_263), .ZN(TIMEBOOST_net_16) );
INV_X1 inst_452 ( .A(net_76), .ZN(net_77) );
INV_X4 inst_430 ( .A(net_334), .ZN(net_169) );
NAND3_X1 inst_131 ( .A1(net_543), .A2(net_544), .A3(net_469), .ZN(net_551) );
INV_X2 inst_406 ( .A(net_72), .ZN(net_26) );
NAND2_X2 inst_214 ( .A1(net_415), .A2(net_538), .ZN(net_430) );
INV_X4 inst_462 ( .A(net_99), .ZN(net_145) );
AND3_X2 TIMEBOOST_cell_68 ( .A1(net_414), .A2(net_427), .A3(G12), .ZN(TIMEBOOST_net_29) );
NAND2_X1 inst_328 ( .A1(net_531), .A2(net_442), .ZN(net_444) );
NOR2_X2 inst_47 ( .A1(net_520), .A2(G4), .ZN(net_66) );
OR2_X4 inst_19 ( .A1(net_381), .A2(net_2), .ZN(net_537) );
DFFR_X1 inst_548 ( .D(net_236), .RN(net_464), .CK(net_622), .QN(net_527) );
INV_X32 inst_515 ( .A(G6), .ZN(net_507) );
OR2_X1 inst_8 ( .A1(net_158), .A2(net_213), .ZN(net_230) );
INV_X1 inst_370 ( .A(net_501), .ZN(net_502) );
AND2_X1 inst_573 ( .A1(net_206), .A2(net_354), .ZN(net_355) );
NOR2_X1 inst_100 ( .A1(net_335), .A2(net_321), .ZN(net_336) );
INV_X1 inst_459 ( .A(net_180), .ZN(net_262) );
NAND2_X1 inst_279 ( .A1(net_166), .A2(net_225), .ZN(net_291) );
INV_X1 inst_445 ( .A(net_206), .ZN(net_96) );
NOR3_X1 TIMEBOOST_cell_117 ( .A1(TIMEBOOST_net_16), .A2(net_293), .A3(net_105), .ZN(net_348) );
NOR2_X2 inst_81 ( .A1(net_59), .A2(net_160), .ZN(net_235) );
CLKBUF_X1 inst_612 ( .A(net_597), .Z(net_598) );
CLKBUF_X1 inst_606 ( .A(net_591), .Z(net_592) );
INV_X4 inst_367 ( .A(G6), .ZN(net_548) );
INV_X2 inst_525 ( .A(net_42), .ZN(net_33) );
NAND3_X1 inst_139 ( .A1(net_238), .A2(net_169), .A3(net_217), .ZN(net_241) );
DFFR_X1 inst_559 ( .D(net_377), .RN(net_464), .CK(TIMEBOOST_net_53), .QN(net_9) );
CLKBUF_X1 inst_584 ( .A(blif_clk_net), .Z(net_570) );
INV_X1 inst_521 ( .A(net_496), .ZN(net_495) );
INV_X4 inst_434 ( .A(net_49), .ZN(net_80) );
INV_X2 inst_470 ( .A(net_124), .ZN(net_160) );
INV_X1 inst_535 ( .A(net_164), .ZN(net_242) );
INV_X4 inst_450 ( .A(net_68), .ZN(net_270) );
INV_X1 inst_520 ( .A(net_498), .ZN(net_497) );
NAND2_X1 inst_237 ( .A1(net_559), .A2(net_169), .ZN(net_106) );
NAND3_X1 inst_148 ( .A1(net_110), .A2(net_229), .A3(net_275), .ZN(net_300) );
DFFR_X1 inst_554 ( .D(net_330), .RN(net_464), .CK(TIMEBOOST_net_4), .Q(net_5) );
INV_X32 inst_377 ( .A(G8), .ZN(net_14) );
NAND2_X1 TIMEBOOST_cell_72 ( .A1(net_449), .A2(net_347), .ZN(TIMEBOOST_net_31) );
NOR2_X1 inst_51 ( .A1(net_15), .A2(net_562), .ZN(net_213) );
NAND3_X1 inst_142 ( .A1(net_115), .A2(net_212), .A3(net_254), .ZN(net_475) );
NAND2_X1 inst_315 ( .A1(net_386), .A2(net_392), .ZN(net_407) );
NOR2_X1 inst_80 ( .A1(net_107), .A2(net_188), .ZN(net_189) );
NAND2_X2 inst_216 ( .A1(net_432), .A2(net_486), .ZN(net_488) );
NOR2_X1 inst_78 ( .A1(net_136), .A2(net_178), .ZN(net_179) );
NAND2_X1 inst_241 ( .A1(net_115), .A2(net_493), .ZN(net_116) );
NAND2_X1 TIMEBOOST_cell_74 ( .A1(net_260), .A2(net_259), .ZN(TIMEBOOST_net_32) );
NAND3_X1 inst_183 ( .A1(net_395), .A2(net_436), .A3(net_454), .ZN(net_458) );
NAND3_X1 inst_151 ( .A1(net_241), .A2(net_332), .A3(net_291), .ZN(net_333) );
NOR2_X1 inst_64 ( .A1(net_148), .A2(net_128), .ZN(net_129) );
INV_X8 inst_415 ( .A(net_37), .ZN(net_49) );
CLKBUF_X1 inst_615 ( .A(net_596), .Z(net_601) );
INV_X32 inst_393 ( .A(G4), .ZN(net_37) );
NOR2_X1 inst_107 ( .A1(net_186), .A2(net_351), .ZN(net_359) );
NAND2_X2 TIMEBOOST_cell_98 ( .A1(net_50), .A2(net_210), .ZN(TIMEBOOST_net_44) );
MUX2_X2 inst_345 ( .A(net_101), .B(net_120), .S(net_18), .Z(net_102) );
NAND2_X2 inst_223 ( .A1(net_13), .A2(G3), .ZN(net_70) );
INV_X1 inst_402 ( .A(net_28), .ZN(net_25) );
NAND3_X1 TIMEBOOST_cell_50 ( .A1(net_120), .A2(net_566), .A3(net_5), .ZN(TIMEBOOST_net_20) );
INV_X2 inst_494 ( .A(net_363), .ZN(net_378) );
INV_X1 inst_487 ( .A(net_187), .ZN(net_239) );
NAND2_X2 inst_329 ( .A1(net_333), .A2(net_426), .ZN(net_445) );
AND2_X1 inst_574 ( .A1(net_420), .A2(net_383), .ZN(net_393) );
INV_X1 inst_386 ( .A(net_19), .ZN(net_15) );
NAND3_X1 inst_158 ( .A1(net_485), .A2(net_74), .A3(net_72), .ZN(net_544) );
NAND3_X1 inst_141 ( .A1(net_149), .A2(net_334), .A3(net_242), .ZN(net_243) );
NAND2_X2 inst_200 ( .A1(net_54), .A2(net_521), .ZN(net_90) );
INV_X1 inst_507 ( .A(net_535), .ZN(net_533) );
AND2_X2 inst_571 ( .A1(net_493), .A2(G11), .ZN(net_212) );
NOR2_X2 inst_57 ( .A1(net_133), .A2(net_85), .ZN(net_86) );
NAND4_X1 TIMEBOOST_cell_135 ( .A1(net_242), .A2(net_324), .A3(net_449), .A4(net_170), .ZN(net_366) );
DFFR_X1 inst_552 ( .D(net_305), .RN(net_464), .CK(net_612), .Q(net_12) );
CLKBUF_X1 inst_599 ( .A(net_584), .Z(net_585) );
INV_X4 inst_417 ( .A(net_42), .ZN(net_115) );
AND2_X1 inst_579 ( .A1(net_79), .A2(net_141), .ZN(net_142) );
OR2_X2 inst_21 ( .A1(net_378), .A2(net_436), .ZN(net_437) );
INV_X2 inst_469 ( .A(net_178), .ZN(net_215) );
NAND2_X1 inst_281 ( .A1(net_500), .A2(net_237), .ZN(net_299) );
CLKBUF_X1 inst_585 ( .A(net_570), .Z(net_571) );
OR2_X2 inst_18 ( .A1(net_538), .A2(net_332), .ZN(net_375) );
INV_X1 inst_541 ( .A(net_365), .ZN(net_358) );
INV_X4 inst_410 ( .A(net_29), .ZN(net_312) );
NAND2_X1 inst_208 ( .A1(net_474), .A2(net_75), .ZN(net_522) );
NOR2_X1 inst_88 ( .A1(net_416), .A2(net_129), .ZN(net_234) );
NAND2_X1 inst_316 ( .A1(net_366), .A2(net_411), .ZN(net_412) );
NAND2_X4 inst_220 ( .A1(G3), .A2(G1), .ZN(net_520) );
OR2_X2 inst_9 ( .A1(net_527), .A2(net_14), .ZN(net_539) );
NOR2_X1 inst_113 ( .A1(net_383), .A2(net_384), .ZN(net_390) );
INV_X4 inst_505 ( .A(net_555), .ZN(net_554) );
INV_X1 inst_356 ( .A(net_555), .ZN(net_553) );
INV_X8 inst_383 ( .A(net_44), .ZN(net_22) );
INV_X1 inst_360 ( .A(net_529), .ZN(net_528) );
NAND2_X2 inst_198 ( .A1(net_37), .A2(net_494), .ZN(net_117) );
NOR2_X2 inst_50 ( .A1(net_42), .A2(net_34), .ZN(net_526) );
NAND2_X1 inst_245 ( .A1(net_50), .A2(net_123), .ZN(net_195) );
AND2_X4 inst_569 ( .A1(G9), .A2(G11), .ZN(net_35) );
CLKBUF_X1 inst_624 ( .A(net_609), .Z(net_610) );
NAND2_X1 inst_260 ( .A1(net_173), .A2(net_61), .ZN(net_194) );
NAND3_X1 TIMEBOOST_cell_27 ( .A1(net_538), .A2(net_424), .A3(net_337), .ZN(net_479) );
NAND2_X1 inst_313 ( .A1(net_98), .A2(net_4), .ZN(net_486) );
NAND3_X1 TIMEBOOST_cell_123 ( .A1(TIMEBOOST_net_50), .A2(net_430), .A3(net_375), .ZN(net_567) );
CLKBUF_X1 inst_636 ( .A(net_621), .Z(net_622) );
CLKBUF_X1 inst_632 ( .A(net_595), .Z(net_618) );
DFFR_X1 inst_549 ( .D(net_290), .RN(net_464), .CK(net_619), .QN(net_1) );
NAND2_X4 inst_234 ( .A1(net_45), .A2(net_508), .ZN(net_84) );
XNOR2_X1 inst_0 ( .A(net_263), .B(net_262), .ZN(net_264) );
INV_X32 inst_522 ( .A(G2), .ZN(net_13) );
NAND3_X1 TIMEBOOST_cell_120 ( .A1(TIMEBOOST_net_28), .A2(net_407), .A3(TIMEBOOST_net_34), .ZN(G550) );
NAND2_X4 inst_236 ( .A1(net_200), .A2(G6), .ZN(net_168) );
INV_X4 inst_433 ( .A(net_70), .ZN(net_200) );
DFFR_X1 inst_553 ( .D(net_303), .RN(net_464), .CK(net_607), .Q(net_547) );
INV_X1 inst_478 ( .A(net_159), .ZN(net_187) );
NOR2_X1 inst_65 ( .A1(net_525), .A2(net_507), .ZN(net_130) );
INV_X1 inst_536 ( .A(net_218), .ZN(net_219) );
NOR3_X1 TIMEBOOST_cell_13 ( .A1(net_139), .A2(net_163), .A3(net_272), .ZN(net_273) );
INV_X2 inst_516 ( .A(net_507), .ZN(net_506) );
NAND3_X1 TIMEBOOST_cell_118 ( .A1(net_245), .A2(net_314), .A3(net_502), .ZN(TIMEBOOST_net_38) );
NAND2_X1 inst_263 ( .A1(net_178), .A2(net_209), .ZN(net_211) );
NAND4_X2 TIMEBOOST_cell_124 ( .A1(net_462), .A2(net_455), .A3(net_449), .A4(net_445), .ZN(G537) );
CLKBUF_X1 TIMEBOOST_cell_126 ( .A(TIMEBOOST_net_1), .Z(TIMEBOOST_net_53) );
OR2_X1 inst_13 ( .A1(net_169), .A2(net_168), .ZN(net_170) );
NOR2_X1 inst_75 ( .A1(net_96), .A2(net_132), .ZN(net_171) );
OR2_X2 TIMEBOOST_cell_46 ( .A1(net_234), .A2(net_317), .ZN(TIMEBOOST_net_18) );
NAND3_X1 inst_166 ( .A1(net_318), .A2(net_420), .A3(net_396), .ZN(net_402) );
NOR2_X1 inst_116 ( .A1(net_140), .A2(net_495), .ZN(net_175) );
CLKBUF_X1 inst_598 ( .A(net_583), .Z(net_584) );
INV_X1 inst_416 ( .A(net_72), .ZN(net_36) );
NAND2_X1 TIMEBOOST_cell_64 ( .A1(net_77), .A2(net_312), .ZN(TIMEBOOST_net_27) );
INV_X4 inst_471 ( .A(net_134), .ZN(net_192) );
INV_X1 inst_394 ( .A(net_35), .ZN(net_31) );
NOR2_X1 inst_79 ( .A1(net_185), .A2(net_154), .ZN(net_186) );
INV_X4 inst_422 ( .A(net_39), .ZN(net_57) );
NAND2_X4 inst_219 ( .A1(G5), .A2(G3), .ZN(net_24) );
NAND2_X1 inst_201 ( .A1(net_553), .A2(net_19), .ZN(net_88) );
CLKBUF_X1 inst_605 ( .A(net_576), .Z(net_591) );
NOR2_X1 TIMEBOOST_cell_39 ( .A1(TIMEBOOST_net_14), .A2(net_284), .ZN(net_321) );
INV_X1 inst_542 ( .A(net_405), .ZN(net_406) );
NAND2_X1 inst_255 ( .A1(net_203), .A2(net_497), .ZN(net_191) );
INV_X4 inst_453 ( .A(net_79), .ZN(net_335) );
NAND3_X1 inst_128 ( .A1(net_52), .A2(net_92), .A3(net_91), .ZN(net_93) );
NOR2_X1 inst_73 ( .A1(net_334), .A2(net_145), .ZN(net_317) );
INV_X2 inst_493 ( .A(net_340), .ZN(net_350) );
INV_X32 inst_378 ( .A(G1), .ZN(net_19) );
NAND2_X1 TIMEBOOST_cell_56 ( .A1(net_204), .A2(net_384), .ZN(TIMEBOOST_net_23) );
NOR2_X1 TIMEBOOST_cell_49 ( .A1(TIMEBOOST_net_19), .A2(net_336), .ZN(net_372) );
INV_X8 inst_351 ( .A(net_32), .ZN(net_75) );
INV_X1 inst_361 ( .A(net_526), .ZN(net_525) );
INV_X4 inst_408 ( .A(net_210), .ZN(net_148) );
NOR3_X1 TIMEBOOST_cell_134 ( .A1(net_233), .A2(net_313), .A3(TIMEBOOST_net_42), .ZN(net_370) );
INV_X1 inst_461 ( .A(net_335), .ZN(net_95) );
INV_X8 inst_385 ( .A(net_14), .ZN(net_41) );
NAND2_X4 inst_197 ( .A1(net_35), .A2(net_41), .ZN(net_45) );
NAND2_X1 inst_250 ( .A1(G6), .A2(net_89), .ZN(net_157) );
NAND3_X1 TIMEBOOST_cell_114 ( .A1(net_180), .A2(net_114), .A3(net_218), .ZN(TIMEBOOST_net_50) );
NAND2_X1 TIMEBOOST_cell_63 ( .A1(TIMEBOOST_net_26), .A2(net_411), .ZN(net_417) );
NOR2_X2 inst_114 ( .A1(G12), .A2(net_537), .ZN(net_400) );
CLKBUF_X1 inst_617 ( .A(net_602), .Z(net_603) );
NOR2_X1 inst_76 ( .A1(net_200), .A2(net_164), .ZN(net_172) );
INV_X4 inst_397 ( .A(net_21), .ZN(net_48) );
INV_X1 inst_504 ( .A(net_558), .ZN(net_557) );
NAND3_X1 inst_150 ( .A1(net_280), .A2(net_184), .A3(net_276), .ZN(net_331) );
CLKBUF_X1 TIMEBOOST_cell_127 ( .A(TIMEBOOST_net_2), .Z(TIMEBOOST_net_54) );
INV_X1 inst_362 ( .A(net_526), .ZN(net_523) );
NAND3_X1 TIMEBOOST_cell_15 ( .A1(net_511), .A2(net_7), .A3(net_247), .ZN(net_279) );
NOR2_X1 inst_83 ( .A1(net_192), .A2(net_141), .ZN(net_198) );
NAND4_X1 inst_121 ( .A1(net_177), .A2(net_106), .A3(net_168), .A4(net_157), .ZN(net_294) );
INV_X1 inst_534 ( .A(net_135), .ZN(net_136) );
INV_X1 inst_440 ( .A(net_57), .ZN(net_58) );
CLKBUF_X1 TIMEBOOST_cell_130 ( .A(TIMEBOOST_net_7), .Z(TIMEBOOST_net_57) );
OR3_X2 inst_2 ( .A1(net_310), .A2(net_338), .A3(net_337), .ZN(net_339) );
CLKBUF_X1 inst_596 ( .A(net_581), .Z(net_582) );
AND2_X1 inst_578 ( .A1(net_91), .A2(net_137), .ZN(net_138) );
NOR2_X1 inst_52 ( .A1(net_56), .A2(G3), .ZN(net_137) );
NAND3_X1 TIMEBOOST_cell_19 ( .A1(net_126), .A2(net_535), .A3(net_155), .ZN(net_319) );
NAND2_X1 inst_267 ( .A1(net_222), .A2(net_60), .ZN(net_229) );
NAND3_X2 inst_140 ( .A1(net_50), .A2(net_29), .A3(net_199), .ZN(net_267) );
NAND2_X4 inst_221 ( .A1(G5), .A2(net_19), .ZN(net_521) );
DFFR_X1 inst_556 ( .D(net_352), .RN(net_464), .CK(TIMEBOOST_net_5), .QN(net_11) );
CLKBUF_X1 inst_637 ( .A(net_581), .Z(net_623) );
NOR2_X1 TIMEBOOST_cell_30 ( .A1(net_109), .A2(net_137), .ZN(TIMEBOOST_net_10) );
DFFR_X1 inst_547 ( .D(net_248), .RN(net_464), .CK(net_624), .QN(net_6) );
INV_X2 inst_530 ( .A(net_335), .ZN(net_104) );
INV_X4 inst_432 ( .A(net_47), .ZN(net_133) );
INV_X1 inst_420 ( .A(net_50), .ZN(net_542) );
NAND2_X1 inst_282 ( .A1(net_534), .A2(net_554), .ZN(net_332) );
INV_X1 inst_368 ( .A(net_505), .ZN(net_504) );
INV_X1 inst_513 ( .A(net_511), .ZN(net_510) );
NOR2_X2 inst_44 ( .A1(net_551), .A2(net_550), .ZN(net_413) );
NAND3_X1 TIMEBOOST_cell_22 ( .A1(net_298), .A2(net_369), .A3(net_492), .ZN(net_443) );
NAND3_X1 inst_174 ( .A1(net_456), .A2(net_517), .A3(net_406), .ZN(net_422) );
INV_X1 inst_371 ( .A(net_499), .ZN(net_496) );
NAND2_X1 inst_314 ( .A1(net_326), .A2(net_4), .ZN(net_399) );
INV_X4 inst_435 ( .A(net_148), .ZN(net_64) );
NAND2_X1 TIMEBOOST_cell_59 ( .A1(TIMEBOOST_net_24), .A2(net_387), .ZN(net_480) );
CLKBUF_X1 inst_597 ( .A(blif_clk_net), .Z(net_583) );
CLKBUF_X1 inst_621 ( .A(net_606), .Z(net_607) );
NOR2_X1 inst_68 ( .A1(net_58), .A2(net_384), .ZN(net_297) );
NAND2_X4 inst_213 ( .A1(net_517), .A2(net_405), .ZN(net_415) );
CLKBUF_X1 inst_604 ( .A(net_589), .Z(net_590) );
NOR2_X2 inst_53 ( .A1(net_101), .A2(net_507), .ZN(net_247) );
CLKBUF_X1 inst_628 ( .A(net_613), .Z(net_614) );
NAND2_X2 inst_205 ( .A1(net_131), .A2(net_43), .ZN(net_209) );
INV_X2 inst_472 ( .A(net_140), .ZN(net_159) );
INV_X1 inst_447 ( .A(net_117), .ZN(net_65) );
INV_X8 inst_380 ( .A(net_14), .ZN(net_20) );
INV_X1 inst_457 ( .A(net_90), .ZN(net_275) );
NAND2_X1 inst_292 ( .A1(net_194), .A2(net_299), .ZN(net_327) );
INV_X16 inst_379 ( .A(net_13), .ZN(net_50) );
NOR3_X1 TIMEBOOST_cell_80 ( .A1(net_388), .A2(net_416), .A3(net_57), .ZN(TIMEBOOST_net_35) );
NAND3_X2 inst_186 ( .A1(net_404), .A2(net_448), .A3(net_532), .ZN(G542) );
OR2_X2 inst_17 ( .A1(net_44), .A2(net_285), .ZN(net_286) );
INV_X1 inst_413 ( .A(net_31), .ZN(net_46) );
NAND3_X1 inst_146 ( .A1(net_255), .A2(net_275), .A3(net_230), .ZN(net_276) );
NAND2_X1 inst_249 ( .A1(net_152), .A2(net_135), .ZN(net_153) );
NOR2_X1 TIMEBOOST_cell_44 ( .A1(net_112), .A2(net_6), .ZN(TIMEBOOST_net_17) );
NAND3_X1 inst_187 ( .A1(net_532), .A2(net_398), .A3(net_472), .ZN(net_463) );
NAND2_X1 inst_206 ( .A1(net_93), .A2(net_116), .ZN(net_536) );
NAND4_X1 inst_122 ( .A1(net_475), .A2(net_257), .A3(net_214), .A4(net_476), .ZN(net_309) );
NAND2_X1 TIMEBOOST_cell_82 ( .A1(net_311), .A2(net_7), .ZN(TIMEBOOST_net_36) );
INV_X4 inst_354 ( .A(G3), .ZN(net_560) );
INV_X1 inst_405 ( .A(net_25), .ZN(net_40) );
INV_X1 inst_492 ( .A(net_267), .ZN(net_268) );
NAND2_X1 inst_240 ( .A1(net_506), .A2(net_493), .ZN(net_114) );
NAND2_X1 inst_326 ( .A1(net_380), .A2(net_431), .ZN(net_441) );
NOR2_X1 inst_110 ( .A1(net_349), .A2(net_361), .ZN(net_373) );
INV_X1 inst_518 ( .A(net_501), .ZN(net_503) );
NOR2_X1 inst_74 ( .A1(net_87), .A2(net_82), .ZN(net_165) );
NAND2_X1 inst_288 ( .A1(net_558), .A2(net_268), .ZN(net_316) );
INV_X8 inst_396 ( .A(net_56), .ZN(net_210) );
NAND2_X1 inst_229 ( .A1(G6), .A2(net_66), .ZN(net_67) );
NOR2_X1 inst_99 ( .A1(net_295), .A2(net_203), .ZN(net_313) );
NOR2_X1 inst_69 ( .A1(net_43), .A2(net_493), .ZN(net_185) );
INV_X16 inst_373 ( .A(G13), .ZN(net_427) );
NOR2_X1 inst_82 ( .A1(net_514), .A2(net_504), .ZN(net_238) );
NOR2_X1 inst_108 ( .A1(net_344), .A2(net_522), .ZN(net_367) );
CLKBUF_X1 inst_595 ( .A(net_577), .Z(net_581) );
NOR2_X1 TIMEBOOST_cell_31 ( .A1(TIMEBOOST_net_10), .A2(net_78), .ZN(net_156) );
OR2_X2 TIMEBOOST_cell_53 ( .A1(TIMEBOOST_net_21), .A2(net_538), .ZN(net_380) );
NAND2_X1 inst_311 ( .A1(net_243), .A2(net_396), .ZN(net_397) );
INV_X1 inst_460 ( .A(net_94), .ZN(net_272) );
INV_X4 inst_372 ( .A(G6), .ZN(net_494) );
NAND3_X1 inst_169 ( .A1(net_397), .A2(net_389), .A3(net_391), .ZN(net_408) );
NAND2_X2 inst_215 ( .A1(net_492), .A2(net_499), .ZN(net_432) );
NAND2_X1 inst_307 ( .A1(net_200), .A2(net_390), .ZN(net_391) );
CLKBUF_X1 inst_638 ( .A(net_615), .Z(net_624) );
INV_X1 inst_421 ( .A(net_38), .ZN(net_60) );
CLKBUF_X1 TIMEBOOST_cell_129 ( .A(TIMEBOOST_net_6), .Z(TIMEBOOST_net_56) );
DFFR_X1 inst_560 ( .D(net_382), .RN(net_464), .CK(TIMEBOOST_net_57), .Q(net_4) );
CLKBUF_X1 inst_586 ( .A(net_571), .Z(net_572) );
DFFR_X1 inst_555 ( .D(net_348), .RN(net_464), .CK(TIMEBOOST_net_54), .QN(net_0) );
OR2_X2 inst_16 ( .A1(net_176), .A2(net_197), .ZN(net_253) );
NAND2_X1 inst_276 ( .A1(net_281), .A2(net_334), .ZN(net_282) );
INV_X2 inst_431 ( .A(net_46), .ZN(net_231) );
INV_X4 inst_348 ( .A(net_507), .ZN(net_499) );
OR3_X1 inst_3 ( .A1(net_317), .A2(net_174), .A3(net_201), .ZN(net_274) );
NAND2_X1 TIMEBOOST_cell_104 ( .A1(net_195), .A2(net_262), .ZN(TIMEBOOST_net_47) );
AND2_X4 inst_577 ( .A1(net_400), .A2(net_427), .ZN(net_411) );
AND3_X1 inst_566 ( .A1(net_206), .A2(net_495), .A3(net_217), .ZN(net_207) );
NOR2_X1 inst_91 ( .A1(net_259), .A2(net_260), .ZN(net_261) );
NAND3_X2 inst_132 ( .A1(net_120), .A2(net_119), .A3(net_554), .ZN(net_154) );
NOR2_X1 TIMEBOOST_cell_48 ( .A1(net_331), .A2(net_355), .ZN(TIMEBOOST_net_19) );
INV_X1 inst_526 ( .A(net_148), .ZN(net_51) );
NOR3_X1 inst_36 ( .A1(net_2), .A2(G12), .A3(G13), .ZN(net_349) );
INV_X1 inst_463 ( .A(net_335), .ZN(net_100) );
INV_X8 inst_503 ( .A(net_559), .ZN(net_558) );
NOR2_X1 inst_96 ( .A1(net_231), .A2(net_258), .ZN(net_296) );
NOR2_X2 inst_45 ( .A1(net_454), .A2(net_85), .ZN(net_460) );
INV_X2 inst_451 ( .A(net_74), .ZN(net_103) );
NOR2_X2 inst_101 ( .A1(net_1), .A2(net_529), .ZN(net_340) );
NAND2_X2 inst_319 ( .A1(net_554), .A2(net_425), .ZN(net_424) );
NAND2_X1 inst_269 ( .A1(net_239), .A2(net_238), .ZN(net_240) );
INV_X4 inst_458 ( .A(net_203), .ZN(net_140) );
INV_X1 inst_444 ( .A(net_206), .ZN(net_63) );
INV_X4 inst_400 ( .A(net_92), .ZN(net_23) );
CLKBUF_X1 inst_614 ( .A(net_586), .Z(net_600) );
NAND2_X1 inst_261 ( .A1(net_498), .A2(net_195), .ZN(net_196) );
INV_X1 inst_514 ( .A(net_515), .ZN(net_509) );
INV_X2 inst_500 ( .A(net_564), .ZN(net_563) );
INV_X1 inst_510 ( .A(net_520), .ZN(net_518) );
NAND2_X1 inst_268 ( .A1(net_180), .A2(net_193), .ZN(net_237) );
INV_X2 inst_369 ( .A(net_499), .ZN(net_501) );
DFFR_X1 inst_550 ( .D(net_274), .RN(net_464), .CK(net_617), .QN(net_2) );
NOR2_X1 inst_63 ( .A1(net_123), .A2(net_56), .ZN(net_565) );
NAND4_X1 inst_119 ( .A1(net_125), .A2(net_25), .A3(net_217), .A4(net_554), .ZN(net_476) );
CLKBUF_X1 inst_603 ( .A(net_588), .Z(net_589) );
NAND3_X1 TIMEBOOST_cell_36 ( .A1(net_138), .A2(net_247), .A3(net_270), .ZN(TIMEBOOST_net_13) );
NOR2_X1 inst_85 ( .A1(net_223), .A2(net_156), .ZN(net_224) );
NOR3_X1 TIMEBOOST_cell_34 ( .A1(net_497), .A2(net_204), .A3(net_203), .ZN(TIMEBOOST_net_12) );
NAND3_X1 TIMEBOOST_cell_25 ( .A1(net_325), .A2(net_492), .A3(net_403), .ZN(G547) );
INV_X4 inst_473 ( .A(net_145), .ZN(net_255) );
NAND2_X2 inst_217 ( .A1(net_442), .A2(net_530), .ZN(net_454) );
AND2_X2 inst_572 ( .A1(net_507), .A2(net_1), .ZN(net_354) );
NOR2_X1 inst_77 ( .A1(net_173), .A2(net_554), .ZN(net_174) );
NAND2_X1 TIMEBOOST_cell_106 ( .A1(net_292), .A2(net_161), .ZN(TIMEBOOST_net_48) );
DFFR_X1 inst_558 ( .D(net_372), .RN(net_464), .CK(net_590), .Q(net_469) );
INV_X4 inst_427 ( .A(net_50), .ZN(net_76) );
NAND2_X1 inst_257 ( .A1(net_98), .A2(net_101), .ZN(net_306) );
CLKBUF_X1 inst_594 ( .A(net_579), .Z(net_580) );
NAND3_X1 inst_145 ( .A1(net_219), .A2(net_505), .A3(net_493), .ZN(net_266) );
NAND2_X1 inst_290 ( .A1(net_504), .A2(net_282), .ZN(net_324) );
INV_X32 inst_374 ( .A(G9), .ZN(net_17) );
NAND3_X1 TIMEBOOST_cell_29 ( .A1(net_568), .A2(net_456), .A3(net_452), .ZN(G532) );
INV_X32 inst_502 ( .A(G3), .ZN(net_559) );
INV_X2 inst_485 ( .A(net_223), .ZN(net_416) );
AND4_X1 inst_565 ( .A1(net_147), .A2(net_316), .A3(net_144), .A4(net_265), .ZN(net_352) );
NAND2_X1 inst_248 ( .A1(net_152), .A2(net_166), .ZN(net_143) );
CLKBUF_X1 inst_622 ( .A(net_582), .Z(net_608) );
NAND3_X2 inst_138 ( .A1(net_215), .A2(net_47), .A3(net_216), .ZN(net_285) );
INV_X8 inst_389 ( .A(net_17), .ZN(net_477) );
INV_X1 inst_357 ( .A(net_463), .ZN(net_552) );
INV_X4 inst_409 ( .A(net_167), .ZN(net_101) );
NAND3_X1 inst_180 ( .A1(net_412), .A2(net_385), .A3(net_439), .ZN(G552) );
NAND2_X1 TIMEBOOST_cell_57 ( .A1(TIMEBOOST_net_23), .A2(net_387), .ZN(net_386) );
NAND2_X1 inst_312 ( .A1(net_338), .A2(net_4), .ZN(net_398) );
CLKBUF_X1 inst_609 ( .A(net_594), .Z(net_595) );
INV_X2 inst_517 ( .A(net_506), .ZN(net_505) );
NAND2_X1 inst_309 ( .A1(net_393), .A2(net_358), .ZN(net_394) );
NAND2_X4 inst_232 ( .A1(net_75), .A2(net_43), .ZN(net_108) );
MUX2_X2 inst_347 ( .A(net_300), .B(net_335), .S(net_320), .Z(net_347) );
NOR2_X1 TIMEBOOST_cell_38 ( .A1(net_71), .A2(net_320), .ZN(TIMEBOOST_net_14) );
INV_X1 inst_363 ( .A(net_514), .ZN(net_513) );
NAND2_X1 inst_247 ( .A1(net_499), .A2(net_334), .ZN(net_127) );
NAND2_X1 inst_297 ( .A1(net_73), .A2(net_346), .ZN(net_485) );
INV_X32 inst_403 ( .A(G7), .ZN(net_32) );
NAND2_X1 inst_302 ( .A1(net_368), .A2(net_0), .ZN(net_369) );
NAND2_X1 inst_310 ( .A1(net_393), .A2(net_365), .ZN(net_395) );
NOR2_X1 TIMEBOOST_cell_45 ( .A1(TIMEBOOST_net_17), .A2(net_150), .ZN(net_342) );
NOR3_X1 TIMEBOOST_cell_115 ( .A1(net_63), .A2(net_287), .A3(net_159), .ZN(net_310) );
NAND2_X2 inst_211 ( .A1(net_360), .A2(net_374), .ZN(net_383) );
CLKBUF_X1 inst_619 ( .A(net_604), .Z(net_605) );
NAND3_X1 inst_162 ( .A1(net_387), .A2(net_420), .A3(net_327), .ZN(net_385) );
CLKBUF_X1 inst_589 ( .A(net_574), .Z(net_575) );
DFFR_X1 inst_561 ( .D(net_458), .RN(net_464), .CK(TIMEBOOST_net_56), .Q(G45) );
INV_X1 inst_412 ( .A(net_210), .ZN(net_30) );
INV_X2 inst_449 ( .A(net_107), .ZN(net_166) );
CLKBUF_X1 inst_639 ( .A(net_614), .Z(net_625) );
NAND3_X1 inst_155 ( .A1(net_547), .A2(net_562), .A3(net_548), .ZN(net_546) );
INV_X2 inst_464 ( .A(net_123), .ZN(net_134) );
CLKBUF_X1 inst_602 ( .A(net_587), .Z(net_588) );
NOR2_X1 inst_59 ( .A1(net_148), .A2(net_117), .ZN(net_135) );
NAND3_X2 inst_135 ( .A1(net_36), .A2(net_167), .A3(net_166), .ZN(net_482) );
OR2_X2 TIMEBOOST_cell_47 ( .A1(TIMEBOOST_net_18), .A2(net_246), .ZN(net_318) );
NAND2_X4 inst_196 ( .A1(net_34), .A2(G7), .ZN(net_112) );
INV_X1 inst_532 ( .A(net_272), .ZN(net_121) );
NOR2_X2 inst_55 ( .A1(net_72), .A2(net_561), .ZN(net_540) );
NAND2_X1 TIMEBOOST_cell_60 ( .A1(net_388), .A2(net_162), .ZN(TIMEBOOST_net_25) );
INV_X1 inst_498 ( .A(net_418), .ZN(net_419) );
NAND2_X1 inst_264 ( .A1(net_148), .A2(net_222), .ZN(net_281) );
NAND3_X1 TIMEBOOST_cell_17 ( .A1(net_121), .A2(net_187), .A3(net_97), .ZN(net_290) );
AND2_X4 TIMEBOOST_cell_69 ( .A1(net_413), .A2(TIMEBOOST_net_29), .ZN(net_492) );
NAND2_X1 TIMEBOOST_cell_37 ( .A1(TIMEBOOST_net_13), .A2(net_235), .ZN(net_271) );
NOR2_X1 TIMEBOOST_cell_35 ( .A1(TIMEBOOST_net_12), .A2(net_143), .ZN(net_205) );
CLKBUF_X1 inst_611 ( .A(net_596), .Z(net_597) );
NAND2_X4 inst_224 ( .A1(net_41), .A2(net_32), .ZN(net_529) );
NOR2_X1 inst_42 ( .A1(net_103), .A2(net_83), .ZN(net_125) );
NAND2_X1 inst_287 ( .A1(net_312), .A2(net_294), .ZN(net_490) );
NAND2_X1 inst_323 ( .A1(net_9), .A2(net_492), .ZN(net_439) );
CLKBUF_X1 inst_618 ( .A(net_579), .Z(net_604) );
INV_X4 inst_426 ( .A(net_75), .ZN(net_74) );
CLKBUF_X1 inst_588 ( .A(net_573), .Z(net_574) );
INV_X8 inst_350 ( .A(net_20), .ZN(net_42) );
NAND2_X1 inst_231 ( .A1(net_92), .A2(net_91), .ZN(net_73) );
NAND4_X1 TIMEBOOST_cell_119 ( .A1(net_420), .A2(net_408), .A3(net_417), .A4(net_451), .ZN(G551) );
INV_X1 inst_474 ( .A(net_146), .ZN(net_302) );
NAND2_X1 TIMEBOOST_cell_51 ( .A1(TIMEBOOST_net_20), .A2(net_565), .ZN(net_364) );
INV_X1 inst_437 ( .A(net_64), .ZN(net_53) );
INV_X1 inst_490 ( .A(net_220), .ZN(net_221) );
CLKBUF_X1 inst_626 ( .A(net_611), .Z(net_612) );
NOR2_X1 inst_70 ( .A1(net_569), .A2(net_150), .ZN(net_151) );
NAND3_X4 inst_129 ( .A1(net_84), .A2(net_108), .A3(net_350), .ZN(net_374) );
NAND2_X1 TIMEBOOST_cell_102 ( .A1(net_216), .A2(net_270), .ZN(TIMEBOOST_net_46) );
OR2_X1 inst_11 ( .A1(net_100), .A2(net_168), .ZN(net_147) );
CLKBUF_X1 inst_631 ( .A(net_616), .Z(net_617) );
NAND3_X2 inst_188 ( .A1(net_434), .A2(net_461), .A3(net_457), .ZN(G535) );
OR2_X1 inst_14 ( .A1(net_235), .A2(net_165), .ZN(net_236) );
INV_X1 inst_475 ( .A(net_154), .ZN(net_155) );
INV_X1 inst_441 ( .A(net_59), .ZN(net_94) );
NOR3_X1 inst_31 ( .A1(net_179), .A2(net_205), .A3(net_189), .ZN(net_305) );
INV_X1 inst_528 ( .A(net_81), .ZN(net_128) );
NOR3_X1 TIMEBOOST_cell_14 ( .A1(net_302), .A2(net_215), .A3(net_171), .ZN(net_303) );
NOR2_X1 inst_62 ( .A1(net_112), .A2(net_68), .ZN(net_113) );
DFFR_X1 inst_557 ( .D(net_370), .RN(net_464), .CK(TIMEBOOST_net_52), .QN(net_10) );
NAND2_X1 inst_251 ( .A1(net_111), .A2(net_210), .ZN(net_199) );
INV_X32 inst_352 ( .A(G3), .ZN(net_562) );
AND2_X4 inst_575 ( .A1(net_537), .A2(net_427), .ZN(net_517) );
INV_X8 inst_398 ( .A(net_22), .ZN(net_320) );
NAND3_X1 TIMEBOOST_cell_96 ( .A1(net_182), .A2(net_540), .A3(net_546), .ZN(TIMEBOOST_net_43) );
INV_X4 inst_436 ( .A(net_75), .ZN(net_52) );
INV_X2 inst_484 ( .A(net_344), .ZN(net_218) );
CLKBUF_X1 inst_627 ( .A(net_600), .Z(net_613) );
NAND4_X4 TIMEBOOST_cell_136 ( .A1(net_362), .A2(net_286), .A3(net_271), .A4(TIMEBOOST_net_27), .ZN(net_531) );
NOR2_X1 inst_102 ( .A1(net_1), .A2(G6), .ZN(net_474) );
NOR2_X1 TIMEBOOST_cell_55 ( .A1(TIMEBOOST_net_22), .A2(net_307), .ZN(net_377) );
NAND2_X1 inst_344 ( .A1(net_315), .A2(net_430), .ZN(net_431) );
INV_X2 inst_428 ( .A(net_120), .ZN(net_59) );
INV_X2 inst_446 ( .A(net_64), .ZN(net_204) );
INV_X1 inst_364 ( .A(net_514), .ZN(net_512) );
NAND3_X1 inst_144 ( .A1(net_196), .A2(net_519), .A3(net_127), .ZN(net_265) );
CLKBUF_X1 inst_629 ( .A(net_614), .Z(net_615) );
NAND2_X2 inst_195 ( .A1(net_24), .A2(G4), .ZN(net_54) );
INV_X4 inst_407 ( .A(net_320), .ZN(net_39) );
CLKBUF_X1 inst_623 ( .A(net_608), .Z(net_609) );
INV_X2 inst_411 ( .A(net_216), .ZN(net_38) );
NAND3_X1 TIMEBOOST_cell_20 ( .A1(net_533), .A2(net_500), .A3(net_266), .ZN(net_330) );
CLKBUF_X1 inst_616 ( .A(net_601), .Z(net_602) );
NAND4_X1 inst_124 ( .A1(net_522), .A2(net_539), .A3(net_152), .A4(net_167), .ZN(net_543) );
INV_X1 inst_533 ( .A(net_131), .ZN(net_132) );
CLKBUF_X1 inst_620 ( .A(net_605), .Z(net_606) );
NAND3_X2 inst_137 ( .A1(net_507), .A2(net_50), .A3(net_260), .ZN(net_491) );
INV_X4 inst_425 ( .A(net_312), .ZN(net_79) );
INV_X1 inst_545 ( .A(net_432), .ZN(net_433) );
NAND3_X2 inst_130 ( .A1(net_481), .A2(net_356), .A3(net_482), .ZN(net_550) );
NAND2_X4 inst_227 ( .A1(net_83), .A2(net_216), .ZN(net_85) );
INV_X4 inst_399 ( .A(net_92), .ZN(net_167) );
INV_X1 inst_527 ( .A(net_133), .ZN(net_61) );
NAND2_X1 inst_226 ( .A1(net_50), .A2(net_560), .ZN(net_81) );
NAND2_X1 TIMEBOOST_cell_76 ( .A1(net_302), .A2(net_328), .ZN(TIMEBOOST_net_33) );
NOR2_X1 inst_58 ( .A1(net_169), .A2(net_70), .ZN(net_105) );
INV_X4 inst_414 ( .A(net_72), .ZN(net_120) );
NOR2_X1 inst_87 ( .A1(net_227), .A2(net_55), .ZN(net_228) );
NOR2_X1 inst_61 ( .A1(net_526), .A2(net_23), .ZN(net_569) );
DFFR_X1 inst_562 ( .D(net_459), .RN(net_464), .CK(TIMEBOOST_net_55), .QN(net_3) );
INV_X1 inst_531 ( .A(net_108), .ZN(net_489) );
NAND3_X1 TIMEBOOST_cell_11 ( .A1(net_117), .A2(net_69), .A3(net_30), .ZN(net_177) );
NAND2_X4 inst_212 ( .A1(net_484), .A2(net_483), .ZN(net_405) );
INV_X4 inst_499 ( .A(net_562), .ZN(net_564) );
NAND2_X1 inst_335 ( .A1(net_567), .A2(net_456), .ZN(net_455) );
INV_X2 inst_466 ( .A(net_384), .ZN(net_260) );
OR2_X1 inst_10 ( .A1(net_273), .A2(net_296), .ZN(net_326) );
OR3_X2 inst_4 ( .A1(net_224), .A2(net_66), .A3(net_256), .ZN(net_308) );
INV_X1 inst_456 ( .A(net_96), .ZN(net_87) );
AND2_X1 inst_581 ( .A1(net_334), .A2(net_283), .ZN(net_284) );
CLKBUF_X1 inst_600 ( .A(net_585), .Z(net_586) );
NOR3_X1 inst_28 ( .A1(net_227), .A2(net_499), .A3(net_43), .ZN(net_233) );
NAND2_X1 inst_275 ( .A1(net_250), .A2(net_501), .ZN(net_280) );
NOR2_X1 inst_117 ( .A1(net_98), .A2(net_31), .ZN(net_197) );
INV_X2 inst_438 ( .A(net_57), .ZN(net_368) );
INV_X2 inst_501 ( .A(net_562), .ZN(net_566) );
NOR2_X2 inst_49 ( .A1(net_28), .A2(G11), .ZN(net_152) );
NAND2_X1 inst_204 ( .A1(net_88), .A2(net_67), .ZN(net_254) );
CLKBUF_X1 inst_587 ( .A(net_570), .Z(net_573) );
NAND3_X2 inst_154 ( .A1(net_490), .A2(net_267), .A3(net_491), .ZN(net_360) );
CLKBUF_X1 inst_592 ( .A(net_572), .Z(net_578) );
DFFR_X1 inst_546 ( .D(net_113), .RN(net_464), .CK(net_626), .Q(net_7) );
NOR2_X1 TIMEBOOST_cell_41 ( .A1(TIMEBOOST_net_15), .A2(net_221), .ZN(net_307) );
INV_X2 inst_465 ( .A(net_103), .ZN(net_124) );
NAND3_X2 TIMEBOOST_cell_24 ( .A1(net_319), .A2(net_378), .A3(net_542), .ZN(net_483) );
NOR2_X1 inst_54 ( .A1(net_334), .A2(net_70), .ZN(net_71) );
AND2_X2 inst_570 ( .A1(net_35), .A2(net_91), .ZN(net_337) );
INV_X8 inst_390 ( .A(net_83), .ZN(net_29) );
CLKBUF_X1 inst_640 ( .A(net_625), .Z(net_626) );
NOR2_X2 inst_43 ( .A1(net_209), .A2(net_210), .ZN(net_244) );
INV_X2 inst_359 ( .A(net_531), .ZN(net_530) );
NAND2_X1 inst_256 ( .A1(net_192), .A2(net_558), .ZN(net_292) );
NOR2_X1 inst_94 ( .A1(net_228), .A2(net_523), .ZN(net_338) );
INV_X2 inst_454 ( .A(net_80), .ZN(net_123) );
CLKBUF_X1 inst_630 ( .A(net_615), .Z(net_616) );
INV_X8 inst_375 ( .A(G12), .ZN(net_456) );
INV_X4 inst_401 ( .A(net_24), .ZN(net_216) );
NAND3_X1 TIMEBOOST_cell_21 ( .A1(net_503), .A2(net_253), .A3(net_240), .ZN(net_325) );
INV_X1 inst_512 ( .A(net_515), .ZN(net_514) );
INV_X1 inst_355 ( .A(net_557), .ZN(net_556) );
NAND2_X4 inst_243 ( .A1(net_558), .A2(net_270), .ZN(net_122) );
NAND2_X1 TIMEBOOST_cell_33 ( .A1(TIMEBOOST_net_11), .A2(net_212), .ZN(net_214) );
CLKBUF_X1 inst_591 ( .A(net_576), .Z(net_577) );
INV_X1 inst_424 ( .A(net_40), .ZN(net_206) );
INV_X4 inst_497 ( .A(net_415), .ZN(net_425) );
NAND2_X2 inst_218 ( .A1(net_488), .A2(net_489), .ZN(net_532) );
OR2_X1 inst_15 ( .A1(net_247), .A2(net_175), .ZN(net_248) );
NAND2_X1 inst_343 ( .A1(net_564), .A2(net_48), .ZN(net_69) );
OR3_X2 inst_6 ( .A1(net_269), .A2(net_297), .A3(net_261), .ZN(net_328) );
NAND2_X4 inst_194 ( .A1(net_21), .A2(G3), .ZN(net_555) );
INV_X1 inst_543 ( .A(net_436), .ZN(net_426) );
NAND2_X2 inst_337 ( .A1(net_279), .A2(net_460), .ZN(net_462) );
NAND2_X1 TIMEBOOST_cell_61 ( .A1(TIMEBOOST_net_25), .A2(net_387), .ZN(net_389) );
INV_X1 inst_509 ( .A(net_520), .ZN(net_519) );
NAND2_X2 inst_299 ( .A1(net_26), .A2(net_354), .ZN(net_356) );
INV_X2 inst_418 ( .A(net_48), .ZN(net_47) );
INV_X4 inst_476 ( .A(net_98), .ZN(net_344) );
OR2_X2 TIMEBOOST_cell_52 ( .A1(net_185), .A2(net_334), .ZN(TIMEBOOST_net_21) );
NOR2_X1 inst_86 ( .A1(net_227), .A2(net_98), .ZN(net_287) );
NAND3_X1 inst_153 ( .A1(net_527), .A2(net_41), .A3(net_92), .ZN(net_346) );
OR2_X2 inst_20 ( .A1(net_359), .A2(net_436), .ZN(net_434) );
INV_X2 inst_442 ( .A(net_60), .ZN(net_180) );
CLKBUF_X1 inst_613 ( .A(net_598), .Z(net_599) );
NOR2_X4 inst_38 ( .A1(net_20), .A2(net_34), .ZN(net_91) );
INV_X8 inst_381 ( .A(net_17), .ZN(net_92) );
INV_X1 inst_349 ( .A(net_499), .ZN(net_498) );
INV_X2 inst_483 ( .A(net_255), .ZN(net_263) );
AND2_X1 inst_576 ( .A1(net_317), .A2(net_400), .ZN(net_401) );
NAND2_X2 inst_209 ( .A1(net_470), .A2(net_471), .ZN(net_365) );
NAND2_X1 inst_259 ( .A1(net_255), .A2(net_384), .ZN(net_193) );
NOR2_X4 inst_40 ( .A1(net_112), .A2(net_477), .ZN(net_493) );
NAND2_X4 inst_320 ( .A1(net_425), .A2(net_456), .ZN(net_436) );
NAND3_X1 inst_167 ( .A1(net_239), .A2(net_323), .A3(net_4), .ZN(net_403) );
CLKBUF_X1 inst_607 ( .A(net_592), .Z(net_593) );
NAND2_X1 inst_246 ( .A1(net_43), .A2(net_528), .ZN(net_126) );
CLKBUF_X1 inst_635 ( .A(net_620), .Z(net_621) );
NOR2_X1 inst_95 ( .A1(net_287), .A2(net_130), .ZN(net_295) );
XNOR2_X1 inst_1 ( .A(net_251), .B(net_524), .ZN(net_323) );
NOR2_X1 inst_72 ( .A1(net_43), .A2(net_529), .ZN(net_163) );
INV_X1 inst_519 ( .A(net_501), .ZN(net_500) );
INV_X4 inst_439 ( .A(net_55), .ZN(net_203) );
NAND2_X1 inst_331 ( .A1(net_339), .A2(net_433), .ZN(net_448) );
AND2_X1 inst_582 ( .A1(net_281), .A2(net_292), .ZN(net_293) );
NOR4_X1 TIMEBOOST_cell_132 ( .A1(net_512), .A2(net_505), .A3(net_231), .A4(net_272), .ZN(TIMEBOOST_net_42) );
NAND2_X1 inst_235 ( .A1(net_81), .A2(net_54), .ZN(net_89) );
NAND2_X4 inst_210 ( .A1(net_365), .A2(G13), .ZN(net_538) );
NAND2_X1 inst_317 ( .A1(net_414), .A2(net_413), .ZN(net_418) );
NAND3_X1 TIMEBOOST_cell_26 ( .A1(net_10), .A2(net_492), .A3(net_399), .ZN(G548) );
INV_X1 inst_467 ( .A(net_335), .ZN(net_388) );
NAND2_X1 inst_239 ( .A1(G6), .A2(net_80), .ZN(net_111) );
NOR2_X1 inst_105 ( .A1(net_12), .A2(net_558), .ZN(net_351) );
INV_X2 inst_488 ( .A(net_263), .ZN(net_449) );
INV_X4 inst_387 ( .A(net_34), .ZN(net_16) );
CLKBUF_X1 inst_593 ( .A(net_578), .Z(net_579) );
NAND2_X1 TIMEBOOST_cell_112 ( .A1(net_368), .A2(net_308), .ZN(TIMEBOOST_net_51) );
NAND2_X1 inst_254 ( .A1(net_182), .A2(net_212), .ZN(net_183) );
CLKBUF_X1 inst_625 ( .A(net_610), .Z(net_611) );
NAND2_X4 inst_225 ( .A1(net_37), .A2(net_44), .ZN(net_68) );
CLKBUF_X1 inst_601 ( .A(net_586), .Z(net_587) );
NAND3_X1 inst_133 ( .A1(net_40), .A2(net_46), .A3(net_182), .ZN(net_188) );
INV_X1 inst_508 ( .A(net_526), .ZN(net_524) );
AND2_X4 inst_568 ( .A1(G6), .A2(G4), .ZN(net_21) );
NOR2_X1 inst_112 ( .A1(net_95), .A2(net_383), .ZN(net_396) );
INV_X32 inst_523 ( .A(G0), .ZN(net_44) );
INV_X1 inst_365 ( .A(net_512), .ZN(net_511) );
NOR2_X1 inst_67 ( .A1(net_203), .A2(net_509), .ZN(net_139) );
NAND3_X2 inst_181 ( .A1(net_422), .A2(net_394), .A3(net_444), .ZN(G539) );
NOR3_X1 TIMEBOOST_cell_40 ( .A1(net_306), .A2(net_496), .A3(net_94), .ZN(TIMEBOOST_net_15) );
INV_X2 inst_479 ( .A(net_160), .ZN(net_227) );
NAND2_X1 TIMEBOOST_cell_92 ( .A1(net_86), .A2(net_50), .ZN(TIMEBOOST_net_41) );
INV_X4 inst_391 ( .A(net_56), .ZN(net_119) );
CLKBUF_X1 inst_590 ( .A(net_575), .Z(net_576) );
NAND2_X4 inst_202 ( .A1(net_217), .A2(net_515), .ZN(net_178) );
NAND4_X1 inst_126 ( .A1(net_446), .A2(net_468), .A3(net_409), .A4(net_402), .ZN(G549) );
INV_X1 inst_480 ( .A(net_173), .ZN(net_161) );
CLKBUF_X1 inst_634 ( .A(net_616), .Z(net_620) );
INV_X4 inst_419 ( .A(net_101), .ZN(net_55) );
INV_X4 inst_477 ( .A(net_192), .ZN(net_223) );
NAND2_X1 TIMEBOOST_cell_70 ( .A1(net_191), .A2(net_513), .ZN(TIMEBOOST_net_30) );
INV_X1 inst_538 ( .A(net_250), .ZN(net_251) );
INV_X4 inst_423 ( .A(net_115), .ZN(net_62) );
NOR3_X1 inst_35 ( .A1(net_344), .A2(net_505), .A3(net_527), .ZN(net_345) );
INV_X8 inst_382 ( .A(net_19), .ZN(net_83) );
NOR2_X4 inst_48 ( .A1(net_16), .A2(net_17), .ZN(net_43) );
INV_X1 inst_358 ( .A(net_535), .ZN(net_534) );
NOR2_X2 inst_46 ( .A1(net_427), .A2(G12), .ZN(net_420) );
NAND3_X1 inst_136 ( .A1(net_275), .A2(net_368), .A3(net_128), .ZN(net_184) );
NOR3_X1 inst_30 ( .A1(net_142), .A2(net_558), .A3(net_198), .ZN(net_269) );
NAND4_X2 TIMEBOOST_cell_121 ( .A1(net_278), .A2(net_285), .A3(net_364), .A4(net_50), .ZN(net_484) );
CLKBUF_X1 inst_610 ( .A(net_584), .Z(net_596) );
NAND2_X4 inst_233 ( .A1(net_49), .A2(net_83), .ZN(net_384) );
NAND2_X1 TIMEBOOST_cell_66 ( .A1(net_449), .A2(net_420), .ZN(TIMEBOOST_net_28) );
NAND2_X1 inst_271 ( .A1(net_220), .A2(net_524), .ZN(net_258) );
INV_X4 inst_443 ( .A(net_62), .ZN(net_98) );
CLKBUF_X1 inst_633 ( .A(net_618), .Z(net_619) );
NAND2_X1 TIMEBOOST_cell_58 ( .A1(G13), .A2(net_11), .ZN(TIMEBOOST_net_24) );
OR2_X1 inst_12 ( .A1(net_148), .A2(net_168), .ZN(net_149) );
INV_X1 inst_529 ( .A(net_96), .ZN(net_97) );
INV_X32 inst_524 ( .A(G5), .ZN(net_27) );
NOR2_X1 inst_56 ( .A1(net_50), .A2(net_38), .ZN(net_78) );
NOR2_X1 inst_71 ( .A1(net_134), .A2(net_320), .ZN(net_158) );
NAND2_X1 inst_308 ( .A1(net_146), .A2(net_390), .ZN(net_392) );
NOR3_X1 TIMEBOOST_cell_122 ( .A1(net_549), .A2(TIMEBOOST_net_35), .A3(net_401), .ZN(net_459) );
INV_X4 inst_448 ( .A(net_76), .ZN(net_99) );
NOR2_X1 inst_60 ( .A1(net_76), .A2(net_518), .ZN(net_109) );
INV_X1 inst_455 ( .A(net_231), .ZN(net_82) );
NAND3_X1 inst_168 ( .A1(net_306), .A2(net_510), .A3(net_4), .ZN(net_404) );
INV_X16 inst_384 ( .A(net_27), .ZN(net_56) );
NAND2_X1 inst_321 ( .A1(G12), .A2(net_419), .ZN(net_549) );
INV_X1 inst_496 ( .A(net_383), .ZN(net_387) );
CLKBUF_X1 inst_608 ( .A(net_593), .Z(net_594) );
NAND2_X2 inst_336 ( .A1(net_437), .A2(net_450), .ZN(G530) );
DFFR_X1 inst_563 ( .D(net_552), .RN(net_464), .CK(TIMEBOOST_net_58), .QN(G546) );
AND2_X1 inst_583 ( .A1(net_420), .A2(net_360), .ZN(net_361) );
AND2_X1 inst_580 ( .A1(net_200), .A2(net_199), .ZN(net_201) );
AND2_X2 TIMEBOOST_cell_108 ( .A1(net_427), .A2(G12), .ZN(TIMEBOOST_net_49) );
NAND2_X1 inst_258 ( .A1(net_39), .A2(net_558), .ZN(net_259) );
INV_X32 inst_376 ( .A(G10), .ZN(net_34) );
NAND2_X4 inst_199 ( .A1(net_42), .A2(net_478), .ZN(net_107) );
NOR2_X4 inst_41 ( .A1(net_107), .A2(G11), .ZN(net_131) );
INV_X4 inst_511 ( .A(net_516), .ZN(net_515) );
NAND3_X1 inst_143 ( .A1(net_254), .A2(net_337), .A3(net_124), .ZN(net_257) );
NAND2_X1 TIMEBOOST_cell_100 ( .A1(net_427), .A2(net_3), .ZN(TIMEBOOST_net_45) );
NAND2_X1 inst_265 ( .A1(net_153), .A2(net_188), .ZN(net_225) );
INV_X1 inst_482 ( .A(net_192), .ZN(net_222) );
INV_X1 inst_468 ( .A(net_204), .ZN(net_146) );
INV_X1 inst_544 ( .A(blif_reset_net), .ZN(net_464) );
NAND2_X1 inst_238 ( .A1(net_51), .A2(net_519), .ZN(net_110) );
INV_X1 inst_540 ( .A(net_314), .ZN(net_315) );
INV_X1 inst_539 ( .A(net_6), .ZN(net_311) );
INV_X4 inst_429 ( .A(net_45), .ZN(net_217) );
INV_X32 inst_404 ( .A(G11), .ZN(net_72) );
NAND3_X1 TIMEBOOST_cell_78 ( .A1(net_443), .A2(net_468), .A3(net_410), .ZN(TIMEBOOST_net_34) );
NOR2_X1 inst_89 ( .A1(net_64), .A2(net_172), .ZN(net_246) );
NOR2_X1 inst_111 ( .A1(net_381), .A2(net_373), .ZN(net_382) );
NOR2_X2 inst_66 ( .A1(net_558), .A2(net_133), .ZN(net_164) );
INV_X8 inst_388 ( .A(net_34), .ZN(net_28) );
NAND2_X1 TIMEBOOST_cell_62 ( .A1(net_416), .A2(net_8), .ZN(TIMEBOOST_net_26) );
NOR2_X1 TIMEBOOST_cell_90 ( .A1(net_255), .A2(net_558), .ZN(TIMEBOOST_net_40) );
INV_X1 inst_392 ( .A(net_28), .ZN(net_18) );
NOR3_X1 TIMEBOOST_cell_54 ( .A1(net_207), .A2(net_345), .A3(net_367), .ZN(TIMEBOOST_net_22) );
NAND2_X1 inst_273 ( .A1(net_244), .A2(net_554), .ZN(net_278) );
NAND3_X1 TIMEBOOST_cell_32 ( .A1(net_213), .A2(net_65), .A3(net_62), .ZN(TIMEBOOST_net_11) );
NAND2_X4 inst_222 ( .A1(net_28), .A2(G7), .ZN(net_516) );
NAND2_X1 inst_284 ( .A1(net_223), .A2(net_533), .ZN(net_314) );
INV_X2 inst_489 ( .A(net_220), .ZN(net_250) );
NAND2_X1 TIMEBOOST_cell_88 ( .A1(net_503), .A2(net_456), .ZN(TIMEBOOST_net_39) );
NAND2_X1 inst_280 ( .A1(net_556), .A2(net_297), .ZN(net_298) );
INV_X4 inst_366 ( .A(net_516), .ZN(net_508) );
MUX2_X2 inst_346 ( .A(net_102), .B(net_43), .S(net_529), .Z(net_176) );
INV_X1 inst_491 ( .A(net_190), .ZN(net_283) );
NAND3_X1 TIMEBOOST_cell_116 ( .A1(net_117), .A2(net_183), .A3(net_557), .ZN(TIMEBOOST_net_37) );
NAND2_X4 inst_193 ( .A1(net_27), .A2(G4), .ZN(net_334) );
CLKBUF_X1 TIMEBOOST_cell_125 ( .A(TIMEBOOST_net_0), .Z(TIMEBOOST_net_52) );
NOR2_X2 inst_39 ( .A1(net_48), .A2(net_27), .ZN(net_182) );
NAND2_X4 inst_230 ( .A1(net_33), .A2(G11), .ZN(net_150) );
CLKBUF_X1 TIMEBOOST_cell_0 ( .A(net_572), .Z(TIMEBOOST_net_0) );
CLKBUF_X1 TIMEBOOST_cell_1 ( .A(net_586), .Z(TIMEBOOST_net_1) );
CLKBUF_X1 TIMEBOOST_cell_2 ( .A(net_600), .Z(TIMEBOOST_net_2) );
CLKBUF_X1 TIMEBOOST_cell_3 ( .A(net_577), .Z(TIMEBOOST_net_3) );
CLKBUF_X1 TIMEBOOST_cell_4 ( .A(net_603), .Z(TIMEBOOST_net_4) );
CLKBUF_X1 TIMEBOOST_cell_5 ( .A(net_599), .Z(TIMEBOOST_net_5) );
CLKBUF_X1 TIMEBOOST_cell_6 ( .A(net_580), .Z(TIMEBOOST_net_6) );
CLKBUF_X1 TIMEBOOST_cell_7 ( .A(net_582), .Z(TIMEBOOST_net_7) );
CLKBUF_X1 TIMEBOOST_cell_8 ( .A(net_623), .Z(TIMEBOOST_net_8) );
CLKBUF_X1 TIMEBOOST_cell_9 ( .A(net_595), .Z(TIMEBOOST_net_9) );
NAND3_X1 TIMEBOOST_cell_10 ( .A1(net_90), .A2(net_50), .A3(net_563), .ZN(net_190) );
NAND2_X1 TIMEBOOST_cell_71 ( .A1(net_492), .A2(TIMEBOOST_net_30), .ZN(net_472) );
NAND2_X1 TIMEBOOST_cell_73 ( .A1(TIMEBOOST_net_31), .A2(net_492), .ZN(net_450) );
NAND2_X1 TIMEBOOST_cell_75 ( .A1(TIMEBOOST_net_32), .A2(net_492), .ZN(net_446) );
NAND2_X1 TIMEBOOST_cell_77 ( .A1(TIMEBOOST_net_33), .A2(net_492), .ZN(net_451) );
CLKBUF_X1 TIMEBOOST_cell_128 ( .A(TIMEBOOST_net_3), .Z(TIMEBOOST_net_55) );
CLKBUF_X1 TIMEBOOST_cell_131 ( .A(TIMEBOOST_net_9), .Z(TIMEBOOST_net_58) );
NAND2_X2 TIMEBOOST_cell_83 ( .A1(TIMEBOOST_net_36), .A2(net_460), .ZN(net_461) );
NAND2_X1 TIMEBOOST_cell_85 ( .A1(TIMEBOOST_net_37), .A2(net_425), .ZN(net_429) );
NAND2_X1 TIMEBOOST_cell_87 ( .A1(TIMEBOOST_net_38), .A2(net_430), .ZN(net_438) );
NAND2_X1 TIMEBOOST_cell_89 ( .A1(TIMEBOOST_net_39), .A2(net_441), .ZN(net_457) );
NOR2_X1 TIMEBOOST_cell_91 ( .A1(TIMEBOOST_net_40), .A2(net_104), .ZN(net_256) );
NAND2_X1 TIMEBOOST_cell_93 ( .A1(TIMEBOOST_net_41), .A2(net_211), .ZN(net_471) );
NAND2_X1 TIMEBOOST_cell_97 ( .A1(TIMEBOOST_net_43), .A2(net_536), .ZN(net_363) );
NAND2_X1 TIMEBOOST_cell_99 ( .A1(TIMEBOOST_net_44), .A2(net_309), .ZN(net_470) );
NAND2_X1 TIMEBOOST_cell_101 ( .A1(net_556), .A2(TIMEBOOST_net_45), .ZN(net_468) );
NAND2_X1 TIMEBOOST_cell_103 ( .A1(TIMEBOOST_net_46), .A2(net_342), .ZN(net_362) );
NAND2_X1 TIMEBOOST_cell_105 ( .A1(TIMEBOOST_net_47), .A2(net_411), .ZN(net_410) );
NAND2_X1 TIMEBOOST_cell_107 ( .A1(TIMEBOOST_net_48), .A2(net_411), .ZN(net_409) );
AND2_X2 TIMEBOOST_cell_109 ( .A1(TIMEBOOST_net_49), .A2(net_418), .ZN(net_442) );
NAND4_X2 TIMEBOOST_cell_133 ( .A1(net_283), .A2(net_119), .A3(net_122), .A4(net_334), .ZN(net_414) );
NAND2_X1 TIMEBOOST_cell_113 ( .A1(TIMEBOOST_net_51), .A2(net_492), .ZN(net_452) );

endmodule
