module cordic_slow (
beta_0,
beta_1,
beta_10,
beta_11,
beta_12,
beta_13,
beta_14,
beta_15,
beta_16,
beta_17,
beta_18,
beta_19,
beta_2,
beta_20,
beta_21,
beta_22,
beta_23,
beta_24,
beta_25,
beta_26,
beta_27,
beta_28,
beta_29,
beta_3,
beta_30,
beta_31,
beta_4,
beta_5,
beta_6,
beta_7,
beta_8,
beta_9,
ispd_clk,
rst,
cos_out_0,
cos_out_1,
cos_out_10,
cos_out_11,
cos_out_12,
cos_out_13,
cos_out_14,
cos_out_15,
cos_out_16,
cos_out_17,
cos_out_18,
cos_out_19,
cos_out_2,
cos_out_20,
cos_out_21,
cos_out_22,
cos_out_23,
cos_out_24,
cos_out_25,
cos_out_26,
cos_out_27,
cos_out_28,
cos_out_29,
cos_out_3,
cos_out_30,
cos_out_31,
cos_out_4,
cos_out_5,
cos_out_6,
cos_out_7,
cos_out_8,
cos_out_9,
sin_out_0,
sin_out_1,
sin_out_10,
sin_out_11,
sin_out_12,
sin_out_13,
sin_out_14,
sin_out_15,
sin_out_16,
sin_out_17,
sin_out_18,
sin_out_19,
sin_out_2,
sin_out_20,
sin_out_21,
sin_out_22,
sin_out_23,
sin_out_24,
sin_out_25,
sin_out_26,
sin_out_27,
sin_out_28,
sin_out_29,
sin_out_3,
sin_out_30,
sin_out_31,
sin_out_4,
sin_out_5,
sin_out_6,
sin_out_7,
sin_out_8,
sin_out_9
);

// Start PIs
input beta_0;
input beta_1;
input beta_10;
input beta_11;
input beta_12;
input beta_13;
input beta_14;
input beta_15;
input beta_16;
input beta_17;
input beta_18;
input beta_19;
input beta_2;
input beta_20;
input beta_21;
input beta_22;
input beta_23;
input beta_24;
input beta_25;
input beta_26;
input beta_27;
input beta_28;
input beta_29;
input beta_3;
input beta_30;
input beta_31;
input beta_4;
input beta_5;
input beta_6;
input beta_7;
input beta_8;
input beta_9;
input ispd_clk;
input rst;

// Start POs
output cos_out_0;
output cos_out_1;
output cos_out_10;
output cos_out_11;
output cos_out_12;
output cos_out_13;
output cos_out_14;
output cos_out_15;
output cos_out_16;
output cos_out_17;
output cos_out_18;
output cos_out_19;
output cos_out_2;
output cos_out_20;
output cos_out_21;
output cos_out_22;
output cos_out_23;
output cos_out_24;
output cos_out_25;
output cos_out_26;
output cos_out_27;
output cos_out_28;
output cos_out_29;
output cos_out_3;
output cos_out_30;
output cos_out_31;
output cos_out_4;
output cos_out_5;
output cos_out_6;
output cos_out_7;
output cos_out_8;
output cos_out_9;
output sin_out_0;
output sin_out_1;
output sin_out_10;
output sin_out_11;
output sin_out_12;
output sin_out_13;
output sin_out_14;
output sin_out_15;
output sin_out_16;
output sin_out_17;
output sin_out_18;
output sin_out_19;
output sin_out_2;
output sin_out_20;
output sin_out_21;
output sin_out_22;
output sin_out_23;
output sin_out_24;
output sin_out_25;
output sin_out_26;
output sin_out_27;
output sin_out_28;
output sin_out_29;
output sin_out_3;
output sin_out_30;
output sin_out_31;
output sin_out_4;
output sin_out_5;
output sin_out_6;
output sin_out_7;
output sin_out_8;
output sin_out_9;

// Start wires
wire beta_0;
wire beta_1;
wire beta_10;
wire beta_11;
wire beta_12;
wire beta_13;
wire beta_14;
wire beta_15;
wire beta_16;
wire beta_17;
wire beta_18;
wire beta_19;
wire beta_2;
wire beta_20;
wire beta_21;
wire beta_22;
wire beta_23;
wire beta_24;
wire beta_25;
wire beta_26;
wire beta_27;
wire beta_28;
wire beta_29;
wire beta_3;
wire beta_30;
wire beta_31;
wire beta_4;
wire beta_5;
wire beta_6;
wire beta_7;
wire beta_8;
wire beta_9;
wire ispd_clk;
wire rst;
wire cos_out_0;
wire cos_out_1;
wire cos_out_10;
wire cos_out_11;
wire cos_out_12;
wire cos_out_13;
wire cos_out_14;
wire cos_out_15;
wire cos_out_16;
wire cos_out_17;
wire cos_out_18;
wire cos_out_19;
wire cos_out_2;
wire cos_out_20;
wire cos_out_21;
wire cos_out_22;
wire cos_out_23;
wire cos_out_24;
wire cos_out_25;
wire cos_out_26;
wire cos_out_27;
wire cos_out_28;
wire cos_out_29;
wire cos_out_3;
wire cos_out_30;
wire cos_out_31;
wire cos_out_4;
wire cos_out_5;
wire cos_out_6;
wire cos_out_7;
wire cos_out_8;
wire cos_out_9;
wire sin_out_0;
wire sin_out_1;
wire sin_out_10;
wire sin_out_11;
wire sin_out_12;
wire sin_out_13;
wire sin_out_14;
wire sin_out_15;
wire sin_out_16;
wire sin_out_17;
wire sin_out_18;
wire sin_out_19;
wire sin_out_2;
wire sin_out_20;
wire sin_out_21;
wire sin_out_22;
wire sin_out_23;
wire sin_out_24;
wire sin_out_25;
wire sin_out_26;
wire sin_out_27;
wire sin_out_28;
wire sin_out_29;
wire sin_out_3;
wire sin_out_30;
wire sin_out_31;
wire sin_out_4;
wire sin_out_5;
wire sin_out_6;
wire sin_out_7;
wire sin_out_8;
wire sin_out_9;
wire FE_OCPN1043_n_42367;
wire FE_OCPN1044_n_42367;
wire FE_OCPN1047_n_23581;
wire FE_OCPN1048_n_23581;
wire FE_OCPN1049_n_23581;
wire FE_OCPN1050_n_23581;
wire FE_OCPN1051_n_2702;
wire FE_OCPN1052_n_2702;
wire FE_OCPN1055_n_38087;
wire FE_OCPN1056_n_38087;
wire FE_OCPN1061_n_44460;
wire FE_OCPN1063_n_44461;
wire FE_OCPN1064_n_44461;
wire FE_OCPN1065_n_44461;
wire FE_OCPN1066_n_44461;
wire FE_OCPN1067_n_44461;
wire FE_OCPN1068_n_21973;
wire FE_OCPN1070_n_44267;
wire FE_OCPN1071_n_44267;
wire FE_OCPN1072_n_12638;
wire FE_OCPN1073_n_12638;
wire FE_OCPN1077_n_13831;
wire FE_OCPN1078_n_8915;
wire FE_OCPN1079_n_8915;
wire FE_OCPN1080_n_24819;
wire FE_OCPN1081_n_24819;
wire FE_OCPN1082_n_8388;
wire FE_OCPN1083_n_8388;
wire FE_OCPN1084_n_8388;
wire FE_OCPN1085_n_8499;
wire FE_OCPN1086_n_8499;
wire FE_OCPN1087_n_25481;
wire FE_OCPN1088_n_25481;
wire FE_OCPN1089_n_39089;
wire FE_OCPN1090_n_39089;
wire FE_OCPN1091_n_9014;
wire FE_OCPN1092_n_9014;
wire FE_OCPN1093_n_4459;
wire FE_OCPN1094_n_4459;
wire FE_OCPN1095_n_25318;
wire FE_OCPN1096_n_25318;
wire FE_OCPN1201_n_45450;
wire FE_OCPN1202_n_45450;
wire FE_OCPN1203_n_7663;
wire FE_OCPN1204_n_7663;
wire FE_OCPN1205_n_46990;
wire FE_OCPN1206_n_46990;
wire FE_OCPN1207_n_8185;
wire FE_OCPN1208_n_8185;
wire FE_OCPN1209_n_8846;
wire FE_OCPN1210_n_8846;
wire FE_OCPN1212_n_19354;
wire FE_OCPN1213_n_21166;
wire FE_OCPN1214_n_21166;
wire FE_OCPN1215_n_21946;
wire FE_OCPN1216_n_21946;
wire FE_OCPN1217_n_11012;
wire FE_OCPN1218_n_11012;
wire FE_OCPN1219_n_40863;
wire FE_OCPN1220_n_40863;
wire FE_OCPN1221_n_41211;
wire FE_OCPN1222_n_41211;
wire FE_OCPN1223_n_43521;
wire FE_OCPN1224_n_43521;
wire FE_OCPN1226_n_43357;
wire FE_OCPN1227_n_43605;
wire FE_OCPN1228_n_43605;
wire FE_OCPN1229_n_43601;
wire FE_OCPN1230_n_43601;
wire FE_OCPN1233_n_33341;
wire FE_OCPN1234_n_33341;
wire FE_OCPN1235_n_27207;
wire FE_OCPN1236_n_27207;
wire FE_OCPN1237_n_30470;
wire FE_OCPN1238_n_30470;
wire FE_OCPN1239_n_13412;
wire FE_OCPN1240_n_13412;
wire FE_OCPN1241_n_12633;
wire FE_OCPN1242_n_12633;
wire FE_OCPN1243_n_13992;
wire FE_OCPN1244_n_13992;
wire FE_OCPN1245_n_19645;
wire FE_OCPN1246_n_19645;
wire FE_OCPN1247_n_22291;
wire FE_OCPN1248_n_22291;
wire FE_OCPN1249_n_13882;
wire FE_OCPN1250_n_13882;
wire FE_OCPN1251_n_19314;
wire FE_OCPN1252_n_19314;
wire FE_OCPN1253_n_23815;
wire FE_OCPN1256_n_28656;
wire FE_OCPN1257_n_18854;
wire FE_OCPN1258_n_18854;
wire FE_OCPN1263_n_20971;
wire FE_OCPN1267_n_29155;
wire FE_OCPN1268_n_29155;
wire FE_OCPN1269_n_30577;
wire FE_OCPN1270_n_30577;
wire FE_OCPN1271_n_31403;
wire FE_OCPN1272_n_31403;
wire FE_OCPN1274_n_15708;
wire FE_OCPN1275_n_31773;
wire FE_OCPN1276_n_31773;
wire FE_OCPN1277_n_15656;
wire FE_OCPN1278_n_15656;
wire FE_OCPN1279_n_30823;
wire FE_OCPN1280_n_30823;
wire FE_OCPN1281_n_21007;
wire FE_OCPN1287_n_29375;
wire FE_OCPN1288_n_29375;
wire FE_OCPN1289_n_19384;
wire FE_OCPN1290_n_19384;
wire FE_OCPN1291_n_29439;
wire FE_OCPN1293_n_26296;
wire FE_OCPN1294_n_26296;
wire FE_OCPN1295_n_45450;
wire FE_OCPN1296_n_45450;
wire FE_OCPN1297_n_30134;
wire FE_OCPN1298_n_30134;
wire FE_OCPN1299_n_30136;
wire FE_OCPN1300_n_30136;
wire FE_OCPN1302_n_23771;
wire FE_OCPN1303_n_35945;
wire FE_OCPN1304_n_35945;
wire FE_OCPN1306_n_13721;
wire FE_OCPN1307_n_23677;
wire FE_OCPN1309_n_25431;
wire FE_OCPN1310_n_25431;
wire FE_OCPN1311_FE_OCP_RBN1024_n_24125;
wire FE_OCPN1312_FE_OCP_RBN1024_n_24125;
wire FE_OCPN1313_n_25126;
wire FE_OCPN1314_n_25126;
wire FE_OCPN1316_n_20265;
wire FE_OCPN1317_n_24682;
wire FE_OCPN1318_n_24682;
wire FE_OCPN1319_n_31403;
wire FE_OCPN1320_n_31403;
wire FE_OCPN1321_n_33714;
wire FE_OCPN1324_n_14577;
wire FE_OCPN1325_n_45050;
wire FE_OCPN1326_n_45050;
wire FE_OCPN1327_n_16192;
wire FE_OCPN1329_FE_OFN1196_n_27014;
wire FE_OCPN1330_FE_OFN1196_n_27014;
wire FE_OCPN1331_n_30281;
wire FE_OCPN1332_n_30281;
wire FE_OCPN1333_n_23467;
wire FE_OCPN1334_n_23467;
wire FE_OCPN1335_n_25673;
wire FE_OCPN1336_n_25673;
wire FE_OCPN1337_n_25775;
wire FE_OCPN1338_n_25775;
wire FE_OCPN1340_n_27246;
wire FE_OCPN1341_n_11927;
wire FE_OCPN1342_n_11927;
wire FE_OCPN1343_n_12313;
wire FE_OCPN1344_n_12313;
wire FE_OCPN1345_n_24142;
wire FE_OCPN1346_n_24142;
wire FE_OCPN1350_n_35312;
wire FE_OCPN1351_n_26530;
wire FE_OCPN1352_n_26530;
wire FE_OCPN1353_n_22484;
wire FE_OCPN1354_n_22484;
wire FE_OCPN1355_n_23335;
wire FE_OCPN1356_n_23335;
wire FE_OCPN1357_n_17778;
wire FE_OCPN1358_n_17778;
wire FE_OCPN1359_n_12370;
wire FE_OCPN1360_n_12370;
wire FE_OCPN1361_n_23684;
wire FE_OCPN1362_n_23684;
wire FE_OCPN1363_n_29615;
wire FE_OCPN1364_n_29615;
wire FE_OCPN1365_n_29573;
wire FE_OCPN1366_n_29573;
wire FE_OCPN1367_n_23923;
wire FE_OCPN1368_n_23923;
wire FE_OCPN1369_n_34288;
wire FE_OCPN1370_n_34288;
wire FE_OCPN1371_n_13510;
wire FE_OCPN1372_n_13510;
wire FE_OCPN1373_n_34051;
wire FE_OCPN1375_n_30612;
wire FE_OCPN1376_n_30612;
wire FE_OCPN1377_n_17836;
wire FE_OCPN1379_n_33640;
wire FE_OCPN1380_n_33640;
wire FE_OCPN1381_n_45026;
wire FE_OCPN1382_n_45026;
wire FE_OCPN1383_n_21896;
wire FE_OCPN1384_n_21896;
wire FE_OCPN1385_n_21199;
wire FE_OCPN1386_n_21199;
wire FE_OCPN1387_n_20555;
wire FE_OCPN1388_n_20555;
wire FE_OCPN1389_n_26054;
wire FE_OCPN1390_n_26054;
wire FE_OCPN1391_n_15462;
wire FE_OCPN1393_n_22801;
wire FE_OCPN1394_n_22801;
wire FE_OCPN1395_n_27211;
wire FE_OCPN1396_n_27211;
wire FE_OCPN1397_n_14742;
wire FE_OCPN1398_n_14742;
wire FE_OCPN1400_n_28095;
wire FE_OCPN1401_FE_OFN1196_n_27014;
wire FE_OCPN1402_FE_OFN1196_n_27014;
wire FE_OCPN1403_n_30823;
wire FE_OCPN1404_n_30823;
wire FE_OCPN1435_n_21278;
wire FE_OCPN1605_n_45697;
wire FE_OCPN1606_n_45697;
wire FE_OCPN1607_n_18176;
wire FE_OCPN1608_n_18176;
wire FE_OCPN1609_n_23503;
wire FE_OCPN1610_n_23503;
wire FE_OCPN1611_n_44174;
wire FE_OCPN1612_n_44174;
wire FE_OCPN1613_n_7630;
wire FE_OCPN1614_n_7630;
wire FE_OCPN1615_n_12371;
wire FE_OCPN1616_n_12371;
wire FE_OCPN1617_n_8444;
wire FE_OCPN1618_n_8444;
wire FE_OCPN1619_n_3361;
wire FE_OCPN1620_n_3361;
wire FE_OCPN1621_n_36947;
wire FE_OCPN1622_n_36947;
wire FE_OCPN1623_n_37661;
wire FE_OCPN1624_n_37661;
wire FE_OCPN1625_n_38135;
wire FE_OCPN1626_n_38135;
wire FE_OCPN1627_n_34452;
wire FE_OCPN1628_n_34452;
wire FE_OCPN1629_n_33196;
wire FE_OCPN1630_n_33196;
wire FE_OCPN1632_n_1835;
wire FE_OCPN1633_n_33588;
wire FE_OCPN1634_n_33588;
wire FE_OCPN1635_n_18860;
wire FE_OCPN1636_n_18860;
wire FE_OCPN1637_n_45081;
wire FE_OCPN1638_n_45081;
wire FE_OCPN1639_n_35367;
wire FE_OCPN1641_FE_OCP_RBN1596_n_14823;
wire FE_OCPN1642_FE_OCP_RBN1596_n_14823;
wire FE_OCPN1643_n_16866;
wire FE_OCPN1644_n_16866;
wire FE_OCPN1645_n_18860;
wire FE_OCPN1646_n_18860;
wire FE_OCPN1649_n_44734;
wire FE_OCPN1650_n_11918;
wire FE_OCPN1651_n_11918;
wire FE_OCPN1652_n_23078;
wire FE_OCPN1653_n_23078;
wire FE_OCPN1655_n_12488;
wire FE_OCPN1656_n_12368;
wire FE_OCPN1657_n_12368;
wire FE_OCPN1658_n_12488;
wire FE_OCPN1659_n_12488;
wire FE_OCPN1660_n_37661;
wire FE_OCPN1661_n_37661;
wire FE_OCPN1662_n_4556;
wire FE_OCPN1663_n_4556;
wire FE_OCPN1664_FE_OCP_RBN1138_n_19270;
wire FE_OCPN1665_FE_OCP_RBN1138_n_19270;
wire FE_OCPN1666_n_39207;
wire FE_OCPN1667_n_39207;
wire FE_OCPN1668_n_23941;
wire FE_OCPN1669_n_23941;
wire FE_OCPN1670_n_39371;
wire FE_OCPN1671_n_39371;
wire FE_OCPN1672_n_14055;
wire FE_OCPN1674_n_25721;
wire FE_OCPN1675_n_25721;
wire FE_OCPN1676_n_27062;
wire FE_OCPN1677_n_27062;
wire FE_OCPN1679_n_27315;
wire FE_OCPN1680_n_30614;
wire FE_OCPN1681_n_30614;
wire FE_OCPN1682_n_27210;
wire FE_OCPN1683_n_27210;
wire FE_OCPN1684_n_14555;
wire FE_OCPN1685_n_14555;
wire FE_OCPN1686_n_23097;
wire FE_OCPN1687_n_23097;
wire FE_OCPN1688_n_23167;
wire FE_OCPN1689_n_23167;
wire FE_OCPN1690_n_10105;
wire FE_OCPN1692_n_33140;
wire FE_OCPN1693_n_33140;
wire FE_OCPN1694_n_12836;
wire FE_OCPN1695_n_12836;
wire FE_OCPN1696_n_13721;
wire FE_OCPN1698_n_34118;
wire FE_OCPN1699_n_34118;
wire FE_OCPN1700_n_33544;
wire FE_OCPN1701_n_33544;
wire FE_OCPN1702_n_14210;
wire FE_OCPN1703_n_14210;
wire FE_OCPN1704_n_14730;
wire FE_OCPN1705_n_14730;
wire FE_OCPN1706_n_21229;
wire FE_OCPN1707_n_21229;
wire FE_OCPN1708_FE_OFN739_n_17093;
wire FE_OCPN1709_FE_OFN739_n_17093;
wire FE_OCPN1710_n_45073;
wire FE_OCPN1711_n_45073;
wire FE_OCPN1712_n_42306;
wire FE_OCPN1713_n_42306;
wire FE_OCPN1714_n_43449;
wire FE_OCPN1715_n_43449;
wire FE_OCPN1716_n_12311;
wire FE_OCPN1717_n_12311;
wire FE_OCPN1718_n_28065;
wire FE_OCPN1721_n_23818;
wire FE_OCPN1722_n_29060;
wire FE_OCPN1725_n_33136;
wire FE_OCPN1726_n_18099;
wire FE_OCPN1727_n_18099;
wire FE_OCPN1728_n_34096;
wire FE_OCPN1732_n_14524;
wire FE_OCPN1733_n_14524;
wire FE_OCPN1736_n_27009;
wire FE_OCPN1737_n_27009;
wire FE_OCPN1738_n_33968;
wire FE_OCPN1739_n_33968;
wire FE_OCPN1740_n_18591;
wire FE_OCPN1741_n_18591;
wire FE_OCPN1762_n_30708;
wire FE_OCPN1763_n_30708;
wire FE_OCPN1902_n_32712;
wire FE_OCPN1903_n_32554;
wire FE_OCPN1904_n_32554;
wire FE_OCPN1905_n_23322;
wire FE_OCPN1906_n_23322;
wire FE_OCPN1907_n_17921;
wire FE_OCPN1908_n_17921;
wire FE_OCPN1909_n_40921;
wire FE_OCPN1910_n_40921;
wire FE_OCPN1911_n_33907;
wire FE_OCPN1912_n_33907;
wire FE_OCPN1913_n_2669;
wire FE_OCPN1915_n_22111;
wire FE_OCPN1916_n_22111;
wire FE_OCPN1917_n_29571;
wire FE_OCPN1918_n_29571;
wire FE_OCPN1919_n_22393;
wire FE_OCPN1920_n_22393;
wire FE_OCPN1921_n_24962;
wire FE_OCPN1922_n_24962;
wire FE_OCPN1923_n_20430;
wire FE_OCPN1924_n_20430;
wire FE_OCPN1925_n_34516;
wire FE_OCPN1926_n_34516;
wire FE_OCPN1927_n_30385;
wire FE_OCPN1928_n_30385;
wire FE_OCPN1932_n_9114;
wire FE_OCPN1933_n_26801;
wire FE_OCPN1934_n_26801;
wire FE_OCPN1935_n_31676;
wire FE_OCPN1936_n_31676;
wire FE_OCPN1937_n_31719;
wire FE_OCPN1938_n_31719;
wire FE_OCPN1939_delay_sub_ln23_0_unr23_stage8_stallmux_q;
wire FE_OCPN1940_delay_sub_ln23_0_unr23_stage8_stallmux_q;
wire FE_OCPN1941_n_20723;
wire FE_OCPN1942_n_20723;
wire FE_OCPN1946_delay_sub_ln23_0_unr23_stage8_stallmux_q;
wire FE_OCPN1947_delay_sub_ln23_0_unr23_stage8_stallmux_q;
wire FE_OCPN1949_delay_sub_ln23_0_unr23_stage8_stallmux_q;
wire FE_OCPN1950_delay_sub_ln23_0_unr23_stage8_stallmux_q;
wire FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q;
wire FE_OCPN1952_n_36121;
wire FE_OCPN1953_n_36121;
wire FE_OCPN1955_n_36050;
wire FE_OCPN3529_n_28829;
wire FE_OCPN3531_n_26468;
wire FE_OCPN3541_n_32436;
wire FE_OCPN3542_n_32436;
wire FE_OCPN3543_n_1448;
wire FE_OCPN3544_n_1448;
wire FE_OCPN3545_n_1705;
wire FE_OCPN3546_n_1705;
wire FE_OCPN3547_n_28043;
wire FE_OCPN3548_n_28043;
wire FE_OCPN3549_n_28381;
wire FE_OCPN3550_n_28381;
wire FE_OCPN3551_n_33225;
wire FE_OCPN3552_n_33225;
wire FE_OCPN3553_n_12671;
wire FE_OCPN3554_n_12671;
wire FE_OCPN3555_n_40986;
wire FE_OCPN3556_n_40986;
wire FE_OCPN3557_n_7673;
wire FE_OCPN3559_n_2386;
wire FE_OCPN3560_n_2386;
wire FE_OCPN3561_n_3317;
wire FE_OCPN3562_n_3317;
wire FE_OCPN3563_n_38731;
wire FE_OCPN3564_n_38731;
wire FE_OCPN3565_n_10214;
wire FE_OCPN3567_n_8348;
wire FE_OCPN3568_n_8348;
wire FE_OCPN3569_n_19303;
wire FE_OCPN3570_n_19303;
wire FE_OCPN3571_n_4374;
wire FE_OCPN3572_n_4374;
wire FE_OCPN3573_n_30345;
wire FE_OCPN3574_n_30345;
wire FE_OCPN3575_n_3625;
wire FE_OCPN3576_n_3625;
wire FE_OCPN3577_n_23354;
wire FE_OCPN3578_n_23354;
wire FE_OCPN3579_n_25370;
wire FE_OCPN3580_n_25370;
wire FE_OCPN3581_n_39747;
wire FE_OCPN3582_n_39747;
wire FE_OCPN3583_n_4556;
wire FE_OCPN3584_n_4556;
wire FE_OCPN3585_n_31704;
wire FE_OCPN3586_n_31704;
wire FE_OCPN3589_n_21419;
wire FE_OCPN3592_n_45301;
wire FE_OCPN4514_n_21343;
wire FE_OCPN4515_n_21343;
wire FE_OCPN4519_n_32820;
wire FE_OCPN4520_n_32820;
wire FE_OCPN4521_n_13015;
wire FE_OCPN4522_n_13015;
wire FE_OCPN4523_n_7360;
wire FE_OCPN4524_n_7360;
wire FE_OCPN4525_n_8099;
wire FE_OCPN4526_n_8099;
wire FE_OCPN4527_n_18117;
wire FE_OCPN4528_n_18117;
wire FE_OCPN4529_FE_OCP_RBN2748_n_8474;
wire FE_OCPN4532_n_3319;
wire FE_OCPN4533_n_3319;
wire FE_OCPN4534_n_9012;
wire FE_OCPN4535_n_9012;
wire FE_OCPN4536_n_14543;
wire FE_OCPN4538_n_20332;
wire FE_OCPN4539_n_20332;
wire FE_OCPN4542_FE_OCP_RBN2812_n_8835;
wire FE_OCPN4544_FE_OCP_RBN2850_n_3645;
wire FE_OCPN4545_FE_OCP_RBN2850_n_3645;
wire FE_OCPN4546_n_4727;
wire FE_OCPN4547_n_4727;
wire FE_OCPN4548_FE_OCP_RBN3086_n_10015;
wire FE_OCPN4549_FE_OCP_RBN3086_n_10015;
wire FE_OCPN4550_n_10545;
wire FE_OCPN4551_n_10545;
wire FE_OCPN4827_FE_OCP_RBN4275_n_3700;
wire FE_OCPN4828_FE_OCP_RBN4275_n_3700;
wire FE_OCPN4829_n_5603;
wire FE_OCPN4830_n_5603;
wire FE_OCPN4831_n_22294;
wire FE_OCPN4832_n_22294;
wire FE_OCPN4833_n_32863;
wire FE_OCPN4835_n_36034;
wire FE_OCPN4836_n_36034;
wire FE_OCPN4843_FE_OFN4779_n_44490;
wire FE_OCPN4844_FE_OFN4779_n_44490;
wire FE_OCPN4845_FE_OFN4779_n_44490;
wire FE_OCPN4846_FE_OFN4778_n_44490;
wire FE_OCPN4847_FE_OFN4778_n_44490;
wire FE_OCPN4848_n_28460;
wire FE_OCPN4849_n_28460;
wire FE_OCPN4850_n_47235;
wire FE_OCPN4851_n_47235;
wire FE_OCPN4852_n_29502;
wire FE_OCPN4853_n_29502;
wire FE_OCPN4854_n_34369;
wire FE_OCPN4855_n_34369;
wire FE_OCPN4856_n_14317;
wire FE_OCPN4857_n_14317;
wire FE_OCPN4858_n_10369;
wire FE_OCPN4859_n_10369;
wire FE_OCPN4926_n_1452;
wire FE_OCPN4927_n_1452;
wire FE_OCPN4928_n_16143;
wire FE_OCPN4929_n_16143;
wire FE_OCPN4930_n_20275;
wire FE_OCPN4931_n_20275;
wire FE_OCPN4932_n_47023;
wire FE_OCPN4933_n_47023;
wire FE_OCPN4934_n_11993;
wire FE_OCPN4935_n_11993;
wire FE_OCPN4936_n_13570;
wire FE_OCPN4937_n_13570;
wire FE_OCPN5094_n_679;
wire FE_OCPN5095_n_679;
wire FE_OCPN5096_n_694;
wire FE_OCPN5097_n_694;
wire FE_OCPN5098_n_1282;
wire FE_OCPN5099_n_1282;
wire FE_OCPN5100_n_18918;
wire FE_OCPN5101_n_18918;
wire FE_OCPN5102_FE_OCP_RBN5029_n_18678;
wire FE_OCPN5104_n_30371;
wire FE_OCPN5105_n_30371;
wire FE_OCPN5106_n_31804;
wire FE_OCPN5107_n_31804;
wire FE_OCPN5108_n_29715;
wire FE_OCPN5109_n_29715;
wire FE_OCPN5110_n_25973;
wire FE_OCPN5111_n_25973;
wire FE_OCPN5112_n_22249;
wire FE_OCPN5113_n_22249;
wire FE_OCPN5114_n_22249;
wire FE_OCPN5119_n_25595;
wire FE_OCPN5120_n_25595;
wire FE_OCPN5121_n_44438;
wire FE_OCPN5122_n_44438;
wire FE_OCPN5123_n_31197;
wire FE_OCPN5124_n_31197;
wire FE_OCPN5125_n_16111;
wire FE_OCPN5126_n_16111;
wire FE_OCPN5127_n_22280;
wire FE_OCPN5128_n_22280;
wire FE_OCPN5129_FE_OFN1198_n_27014;
wire FE_OCPN5130_FE_OFN1198_n_27014;
wire FE_OCPN5131_n_29081;
wire FE_OCPN5132_n_29081;
wire FE_OCPN5133_n_27667;
wire FE_OCPN5134_n_27667;
wire FE_OCPN5135_n_12795;
wire FE_OCPN5136_n_12795;
wire FE_OCPN5219_n_10300;
wire FE_OCPN5221_FE_OFN753_n_13889;
wire FE_OCPN5222_FE_OFN753_n_13889;
wire FE_OCPN5223_n_10357;
wire FE_OCPN5225_n_25509;
wire FE_OCPN5226_n_25509;
wire FE_OCPN5227_n_33917;
wire FE_OCPN5228_n_33917;
wire FE_OCPN5229_n_30587;
wire FE_OCPN5230_n_30587;
wire FE_OCPN5231_n_35594;
wire FE_OCPN5233_n_27018;
wire FE_OCPN5234_n_27018;
wire FE_OCPN5235_n_44162;
wire FE_OCPN5237_n_22383;
wire FE_OCPN5238_n_22383;
wire FE_OCPN5239_n_26428;
wire FE_OCPN5240_n_26428;
wire FE_OCPN5241_n_30859;
wire FE_OCPN5242_n_30859;
wire FE_OCPN5243_n_21790;
wire FE_OCPN5244_n_21790;
wire FE_OCPN5245_n_18974;
wire FE_OCPN5246_n_18974;
wire FE_OCPN5247_FE_OFN4715_n_18642;
wire FE_OCPN5248_FE_OFN4715_n_18642;
wire FE_OCPN5249_n_20852;
wire FE_OCPN5250_n_20852;
wire FE_OCPN5251_n_30859;
wire FE_OCPN5252_n_30859;
wire FE_OCPN5253_n_31871;
wire FE_OCPN5254_n_31871;
wire FE_OCPN5257_n_13590;
wire FE_OCPN5258_n_13590;
wire FE_OCPN5259_n_30614;
wire FE_OCPN5260_n_30614;
wire FE_OCPN5261_n_27536;
wire FE_OCPN5262_n_27536;
wire FE_OCPN5263_n_14977;
wire FE_OCPN5264_n_14977;
wire FE_OCPN5265_n_20852;
wire FE_OCPN5267_n_34852;
wire FE_OCPN5268_n_34852;
wire FE_OCPN5269_n_18557;
wire FE_OCPN5270_n_18557;
wire FE_OCPN5271_n_21434;
wire FE_OCPN5272_n_21434;
wire FE_OCPN5273_FE_RN_366_0;
wire FE_OCPN5274_FE_RN_366_0;
wire FE_OCPN5275_n_23590;
wire FE_OCPN5276_n_23590;
wire FE_OCPN5277_n_13329;
wire FE_OCPN5279_n_30614;
wire FE_OCPN5280_n_30614;
wire FE_OCPN5281_n_24425;
wire FE_OCPN5283_n_24425;
wire FE_OCPN5284_n_24425;
wire FE_OCPN5285_n_30708;
wire FE_OCPN5286_n_30708;
wire FE_OCPN5287_n_27315;
wire FE_OCPN5288_n_27315;
wire FE_OCPN5289_n_26125;
wire FE_OCPN5290_n_26125;
wire FE_OCPN5291_n_21790;
wire FE_OCPN5292_n_21790;
wire FE_OCPN5293_n_30584;
wire FE_OCPN5294_n_30584;
wire FE_OCPN5295_FE_OCP_RBN1105_n_18746;
wire FE_OCPN5296_FE_OCP_RBN1105_n_18746;
wire FE_OCPN5297_n_29866;
wire FE_OCPN5298_n_29866;
wire FE_OCPN5299_n_27130;
wire FE_OCPN5300_n_27130;
wire FE_OCPN5305_n_22338;
wire FE_OCPN5306_n_22338;
wire FE_OCPN5363_n_24221;
wire FE_OCPN5364_n_24221;
wire FE_OCPN6268_n_30599;
wire FE_OCPN6269_n_30599;
wire FE_OCPN6276_n_45450;
wire FE_OCPN6277_n_45450;
wire FE_OCPN6278_FE_OCP_RBN1594_n_13557;
wire FE_OCPN6279_FE_OCP_RBN1594_n_13557;
wire FE_OCPN6280_n_30612;
wire FE_OCPN6281_n_30612;
wire FE_OCPN6282_FE_OCP_RBN2783_n_8664;
wire FE_OCPN6283_FE_OCP_RBN2783_n_8664;
wire FE_OCPN6284_FE_OCP_RBN1602_n_14638;
wire FE_OCPN6285_FE_OCP_RBN1602_n_14638;
wire FE_OCPN6286_FE_OCP_RBN6082_n_5454;
wire FE_OCPN6287_FE_OCP_RBN6082_n_5454;
wire FE_OCPN6288_FE_OCP_RBN3263_n_5531;
wire FE_OCPN6289_FE_OCP_RBN3263_n_5531;
wire FE_OCPN6900_FE_OCP_RBN4472_n_31819;
wire FE_OCPN6901_FE_OCP_RBN4472_n_31819;
wire FE_OCPN6908_n_32525;
wire FE_OCPN6909_n_32525;
wire FE_OCPN6910_n_1444;
wire FE_OCPN6911_n_1444;
wire FE_OCPN6912_n_1715;
wire FE_OCPN6913_n_1715;
wire FE_OCPN6914_n_23112;
wire FE_OCPN6915_n_23112;
wire FE_OCPN6916_n_28460;
wire FE_OCPN6917_n_28460;
wire FE_OCPN6918_n_7726;
wire FE_OCPN6919_n_7726;
wire FE_OCPN6920_n_3580;
wire FE_OCPN6921_n_3580;
wire FE_OCPN6922_n_39185;
wire FE_OCPN6923_n_39185;
wire FE_OCPN6924_n_45081;
wire FE_OCPN6925_n_45081;
wire FE_OCPN6926_n_26464;
wire FE_OCPN6927_n_26464;
wire FE_OCPN6928_FE_OCP_RBN1152_n_20910;
wire FE_OCPN6929_FE_OCP_RBN1152_n_20910;
wire FE_OCPN6930_n_22156;
wire FE_OCPN6931_n_22156;
wire FE_OCPN6932_FE_OCP_RBN6087_n_10852;
wire FE_OCPN6933_FE_OCP_RBN6087_n_10852;
wire FE_OCPN6934_FE_OCP_RBN6066_n_26081;
wire FE_OCPN6935_FE_OCP_RBN6066_n_26081;
wire FE_OCPN7082_n_28891;
wire FE_OCPN7083_n_28891;
wire FE_OCPN7084_n_45697;
wire FE_OCPN7085_n_45697;
wire FE_OCPN7086_n_6263;
wire FE_OCPN7087_n_6263;
wire FE_OCPN7088_n_20979;
wire FE_OCPN7089_n_20979;
wire FE_OCPN833_n_45450;
wire FE_OCPN835_n_45450;
wire FE_OCPN836_n_45450;
wire FE_OCPN837_n_44672;
wire FE_OCPN838_n_44672;
wire FE_OCPN839_n_44672;
wire FE_OCPN846_n_12799;
wire FE_OCPN847_n_12799;
wire FE_OCPN848_n_7712;
wire FE_OCPN849_n_7712;
wire FE_OCPN850_n_7712;
wire FE_OCPN858_n_7802;
wire FE_OCPN861_n_7743;
wire FE_OCPN865_n_32892;
wire FE_OCPN866_n_45450;
wire FE_OCPN867_n_45450;
wire FE_OCPN868_n_45003;
wire FE_OCPN869_n_45003;
wire FE_OCPN870_n_24098;
wire FE_OCPN871_n_24098;
wire FE_OCPN872_n_42202;
wire FE_OCPN873_n_42202;
wire FE_OCPN877_n_43022;
wire FE_OCPN878_n_43022;
wire FE_OCPN880_n_44593;
wire FE_OCPN881_n_44776;
wire FE_OCPN882_n_44776;
wire FE_OCPN883_n_41540;
wire FE_OCPN884_n_41540;
wire FE_OCPN889_n_44223;
wire FE_OCPN890_n_44223;
wire FE_OCPN893_n_28471;
wire FE_OCPN894_n_28471;
wire FE_OCPN895_n_28506;
wire FE_OCPN896_n_28506;
wire FE_OCPN899_n_16923;
wire FE_OCPN900_n_16923;
wire FE_OCPN901_n_47020;
wire FE_OCPN902_n_47020;
wire FE_OCPN903_n_21955;
wire FE_OCPN904_n_21955;
wire FE_OCPN905_n_21956;
wire FE_OCPN906_n_21956;
wire FE_OCPN907_n_46956;
wire FE_OCPN908_n_46956;
wire FE_OCPN914_n_8091;
wire FE_OCPN916_n_8753;
wire FE_OCPN917_n_8753;
wire FE_OCPN918_n_17042;
wire FE_OCPN919_n_17042;
wire FE_OCPN924_n_13962;
wire FE_OCPN926_n_12914;
wire FE_OCPN928_n_12880;
wire FE_OCPN929_n_12880;
wire FE_OCPN930_n_7817;
wire FE_OCPN931_n_7817;
wire FE_OCPN935_n_7802;
wire FE_OCPN936_n_17684;
wire FE_OCPN937_n_17684;
wire FE_OCPN938_n_23577;
wire FE_OCPN939_n_23577;
wire FE_OCPN940_n_39096;
wire FE_OCPN941_n_39096;
wire FE_OCPN942_n_31466;
wire FE_OCPN943_n_31466;
wire FE_OCPN945_n_27287;
wire FE_OCPN950_n_44180;
wire FE_OCPUNCON1742_n_29375;
wire FE_OCPUNCON1743_n_29375;
wire FE_OCPUNCON1744_n_29420;
wire FE_OCPUNCON1745_n_29420;
wire FE_OCPUNCON1746_n_34137;
wire FE_OCPUNCON1747_n_34137;
wire FE_OCPUNCON1748_n_19807;
wire FE_OCPUNCON1749_n_19807;
wire FE_OCPUNCON1750_n_33904;
wire FE_OCPUNCON1752_n_35382;
wire FE_OCPUNCON1753_n_35382;
wire FE_OCPUNCON1754_n_35420;
wire FE_OCPUNCON1755_n_35420;
wire FE_OCPUNCON1756_n_35482;
wire FE_OCPUNCON1757_n_35482;
wire FE_OCPUNCON1758_n_35644;
wire FE_OCPUNCON1759_n_35644;
wire FE_OCPUNCON3465_n_29391;
wire FE_OCPUNCON3466_n_29391;
wire FE_OCPUNCON3467_n_29644;
wire FE_OCPUNCON3468_n_29644;
wire FE_OCPUNCON3469_n_28654;
wire FE_OCPUNCON3470_n_28654;
wire FE_OCPUNCON3471_n_24962;
wire FE_OCPUNCON3472_n_24962;
wire FE_OCPUNCON3473_n_28656;
wire FE_OCPUNCON3475_n_29812;
wire FE_OCPUNCON3476_n_29812;
wire FE_OCPUNCON3477_n_29844;
wire FE_OCPUNCON3478_n_29844;
wire FE_OCPUNCON3479_n_28872;
wire FE_OCPUNCON3480_n_28872;
wire FE_OCPUNCON3481_n_21058;
wire FE_OCPUNCON3483_n_35500;
wire FE_OCPUNCON3484_n_35500;
wire FE_OCPUNCON3485_n_31012;
wire FE_OCPUNCON3487_n_21458;
wire FE_OCPUNCON3488_n_21458;
wire FE_OCPUNCON3489_n_34327;
wire FE_OCPUNCON3490_n_34327;
wire FE_OCPUNCON3491_n_30322;
wire FE_OCPUNCON4497_n_34182;
wire FE_OCPUNCON4498_n_34182;
wire FE_OCPUNCON5301_n_17836;
wire FE_OCPUNCON5302_n_17836;
wire FE_OCPUNCON6886_n_19961;
wire FE_OCPUNCON6887_n_19961;
wire FE_OCPUNCON7058_n_34058;
wire FE_OCPUNCON7059_n_34058;
wire FE_OCPUNCON7060_n_34222;
wire FE_OCPUNCON7061_n_34222;
wire FE_OCPUNCON7062_n_33904;
wire FE_OCPUNCON7063_n_33904;
wire FE_OCPUNCON7064_n_35500;
wire FE_OCPUNCON7065_n_35500;
wire FE_OCPUNCON7066_n_34151;
wire FE_OCPUNCON7067_n_34151;
wire FE_OCPUNCON7068_n_21493;
wire FE_OCPUNCON7069_n_21493;
wire FE_OCPUNCON7070_n_21788;
wire FE_OCPUNCON7071_n_21788;
wire FE_OCPUNCON7072_n_31583;
wire FE_OCPUNCON7073_n_31583;
wire FE_OCP_DRV_N1405_n_43514;
wire FE_OCP_DRV_N1406_n_43514;
wire FE_OCP_DRV_N1407_n_28550;
wire FE_OCP_DRV_N1409_n_12416;
wire FE_OCP_DRV_N1410_n_12416;
wire FE_OCP_DRV_N1411_n_12570;
wire FE_OCP_DRV_N1412_n_12570;
wire FE_OCP_DRV_N1413_n_33673;
wire FE_OCP_DRV_N1414_n_33673;
wire FE_OCP_DRV_N1416_n_34051;
wire FE_OCP_DRV_N1417_n_32985;
wire FE_OCP_DRV_N1419_n_24747;
wire FE_OCP_DRV_N1420_n_24747;
wire FE_OCP_DRV_N1421_n_35367;
wire FE_OCP_DRV_N1423_n_35292;
wire FE_OCP_DRV_N1424_n_35292;
wire FE_OCP_DRV_N1425_n_24158;
wire FE_OCP_DRV_N1426_n_24158;
wire FE_OCP_DRV_N1427_n_35312;
wire FE_OCP_DRV_N1428_n_35312;
wire FE_OCP_DRV_N1429_n_22126;
wire FE_OCP_DRV_N1430_n_22126;
wire FE_OCP_DRV_N1431_n_26850;
wire FE_OCP_DRV_N1432_n_26850;
wire FE_OCP_DRV_N1433_n_21283;
wire FE_OCP_DRV_N1434_n_21283;
wire FE_OCP_DRV_N1437_n_17643;
wire FE_OCP_DRV_N1438_n_17643;
wire FE_OCP_DRV_N1439_n_19010;
wire FE_OCP_DRV_N1440_n_19010;
wire FE_OCP_DRV_N1441_n_17836;
wire FE_OCP_DRV_N1443_n_19138;
wire FE_OCP_DRV_N1444_n_19138;
wire FE_OCP_DRV_N1445_n_19314;
wire FE_OCP_DRV_N1446_n_19314;
wire FE_OCP_DRV_N1447_n_19354;
wire FE_OCP_DRV_N1448_n_19354;
wire FE_OCP_DRV_N1449_n_19384;
wire FE_OCP_DRV_N1450_n_19384;
wire FE_OCP_DRV_N1451_n_12585;
wire FE_OCP_DRV_N1452_n_12585;
wire FE_OCP_DRV_N1453_n_19590;
wire FE_OCP_DRV_N1454_n_19590;
wire FE_OCP_DRV_N1455_n_19562;
wire FE_OCP_DRV_N1456_n_19562;
wire FE_OCP_DRV_N1457_n_19665;
wire FE_OCP_DRV_N1458_n_19665;
wire FE_OCP_DRV_N1459_n_18111;
wire FE_OCP_DRV_N1460_n_18111;
wire FE_OCP_DRV_N1461_n_29777;
wire FE_OCP_DRV_N1462_n_29777;
wire FE_OCP_DRV_N1463_n_19751;
wire FE_OCP_DRV_N1464_n_19751;
wire FE_OCP_DRV_N1465_n_29860;
wire FE_OCP_DRV_N1466_n_29860;
wire FE_OCP_DRV_N1467_n_28775;
wire FE_OCP_DRV_N1468_n_28775;
wire FE_OCP_DRV_N1469_n_25022;
wire FE_OCP_DRV_N1470_n_25022;
wire FE_OCP_DRV_N1471_n_25044;
wire FE_OCP_DRV_N1472_n_25044;
wire FE_OCP_DRV_N1473_n_23792;
wire FE_OCP_DRV_N1474_n_23792;
wire FE_OCP_DRV_N1475_n_23887;
wire FE_OCP_DRV_N1476_n_23887;
wire FE_OCP_DRV_N1477_n_35106;
wire FE_OCP_DRV_N1478_n_35106;
wire FE_OCP_DRV_N1479_n_30917;
wire FE_OCP_DRV_N1480_n_30917;
wire FE_OCP_DRV_N1481_n_26296;
wire FE_OCP_DRV_N1482_n_26296;
wire FE_OCP_DRV_N1483_n_35427;
wire FE_OCP_DRV_N1484_n_35427;
wire FE_OCP_DRV_N1485_n_21639;
wire FE_OCP_DRV_N1486_n_21639;
wire FE_OCP_DRV_N1487_n_24848;
wire FE_OCP_DRV_N1488_n_24848;
wire FE_OCP_DRV_N1489_n_26656;
wire FE_OCP_DRV_N1490_n_26656;
wire FE_OCP_DRV_N1491_n_31445;
wire FE_OCP_DRV_N1492_n_31445;
wire FE_OCP_DRV_N1493_n_20059;
wire FE_OCP_DRV_N1494_n_20059;
wire FE_OCP_DRV_N1495_n_31473;
wire FE_OCP_DRV_N1496_n_31473;
wire FE_OCP_DRV_N1497_n_34924;
wire FE_OCP_DRV_N1498_n_34924;
wire FE_OCP_DRV_N1499_n_15605;
wire FE_OCP_DRV_N1500_n_15605;
wire FE_OCP_DRV_N1501_n_15979;
wire FE_OCP_DRV_N1502_n_15979;
wire FE_OCP_DRV_N1503_n_16106;
wire FE_OCP_DRV_N1504_n_16106;
wire FE_OCP_DRV_N1505_n_16183;
wire FE_OCP_DRV_N1506_n_16183;
wire FE_OCP_DRV_N1507_n_26491;
wire FE_OCP_DRV_N1508_n_26491;
wire FE_OCP_DRV_N1509_n_36387;
wire FE_OCP_DRV_N1510_n_36387;
wire FE_OCP_DRV_N1511_n_26582;
wire FE_OCP_DRV_N1512_n_26582;
wire FE_OCP_DRV_N1513_n_26786;
wire FE_OCP_DRV_N1514_n_26786;
wire FE_OCP_DRV_N1515_n_21706;
wire FE_OCP_DRV_N1516_n_21706;
wire FE_OCP_DRV_N1517_n_21851;
wire FE_OCP_DRV_N1518_n_21851;
wire FE_OCP_DRV_N1519_n_26761;
wire FE_OCP_DRV_N1520_n_26761;
wire FE_OCP_DRV_N1521_n_26807;
wire FE_OCP_DRV_N1522_n_26807;
wire FE_OCP_DRV_N1523_n_31435;
wire FE_OCP_DRV_N1524_n_31435;
wire FE_OCP_DRV_N1760_n_20145;
wire FE_OCP_DRV_N1761_n_20145;
wire FE_OCP_DRV_N1879_n_28164;
wire FE_OCP_DRV_N1880_n_28164;
wire FE_OCP_DRV_N1881_n_32758;
wire FE_OCP_DRV_N1882_n_32758;
wire FE_OCP_DRV_N1883_n_24361;
wire FE_OCP_DRV_N1884_n_24361;
wire FE_OCP_DRV_N1885_n_34009;
wire FE_OCP_DRV_N1886_n_34009;
wire FE_OCP_DRV_N1887_n_33756;
wire FE_OCP_DRV_N1888_n_33756;
wire FE_OCP_DRV_N1889_n_29317;
wire FE_OCP_DRV_N1891_n_29573;
wire FE_OCP_DRV_N1892_n_29573;
wire FE_OCP_DRV_N1893_n_33221;
wire FE_OCP_DRV_N1894_n_33221;
wire FE_OCP_DRV_N1895_n_19855;
wire FE_OCP_DRV_N1896_n_19855;
wire FE_OCP_DRV_N1897_n_18287;
wire FE_OCP_DRV_N1898_n_18287;
wire FE_OCP_DRV_N1899_n_23668;
wire FE_OCP_DRV_N1900_n_23668;
wire FE_OCP_DRV_N3493_n_40837;
wire FE_OCP_DRV_N3494_n_40837;
wire FE_OCP_DRV_N3495_n_33156;
wire FE_OCP_DRV_N3496_n_33156;
wire FE_OCP_DRV_N3497_n_7233;
wire FE_OCP_DRV_N3498_n_7233;
wire FE_OCP_DRV_N3499_n_7204;
wire FE_OCP_DRV_N3500_n_7204;
wire FE_OCP_DRV_N3501_n_29140;
wire FE_OCP_DRV_N3502_n_29140;
wire FE_OCP_DRV_N3504_FE_OCP_RBN1807_n_13010;
wire FE_OCP_DRV_N3505_n_8189;
wire FE_OCP_DRV_N3506_n_8189;
wire FE_OCP_DRV_N3507_n_13329;
wire FE_OCP_DRV_N3508_n_13329;
wire FE_OCP_DRV_N3509_n_35315;
wire FE_OCP_DRV_N3510_n_35315;
wire FE_OCP_DRV_N3511_n_30318;
wire FE_OCP_DRV_N3512_n_30318;
wire FE_OCP_DRV_N3513_n_14650;
wire FE_OCP_DRV_N3514_n_14650;
wire FE_OCP_DRV_N3515_n_31504;
wire FE_OCP_DRV_N3516_n_31504;
wire FE_OCP_DRV_N3517_n_39785;
wire FE_OCP_DRV_N3518_n_39785;
wire FE_OCP_DRV_N3519_n_43153;
wire FE_OCP_DRV_N3520_n_43153;
wire FE_OCP_DRV_N3521_n_43538;
wire FE_OCP_DRV_N3522_n_43538;
wire FE_OCP_DRV_N3523_FE_OCP_RBN3021_n_15319;
wire FE_OCP_DRV_N3524_FE_OCP_RBN3021_n_15319;
wire FE_OCP_DRV_N3525_n_17031;
wire FE_OCP_DRV_N3526_n_17031;
wire FE_OCP_DRV_N3527_n_17071;
wire FE_OCP_DRV_N3528_n_17071;
wire FE_OCP_DRV_N3533_n_18559;
wire FE_OCP_DRV_N3534_n_18559;
wire FE_OCP_DRV_N3535_n_19053;
wire FE_OCP_DRV_N3536_n_19053;
wire FE_OCP_DRV_N3537_n_21763;
wire FE_OCP_DRV_N3538_n_21763;
wire FE_OCP_DRV_N3539_n_20146;
wire FE_OCP_DRV_N3540_n_20146;
wire FE_OCP_DRV_N4499_n_13785;
wire FE_OCP_DRV_N4500_n_13785;
wire FE_OCP_DRV_N4501_FE_OCP_RBN1807_n_13010;
wire FE_OCP_DRV_N4502_FE_OCP_RBN1807_n_13010;
wire FE_OCP_DRV_N4503_n_28888;
wire FE_OCP_DRV_N4505_n_13476;
wire FE_OCP_DRV_N4507_n_15099;
wire FE_OCP_DRV_N4508_n_15099;
wire FE_OCP_DRV_N4510_n_21343;
wire FE_OCP_DRV_N5140_n_29375;
wire FE_OCP_DRV_N5141_n_29375;
wire FE_OCP_DRV_N5142_n_28426;
wire FE_OCP_DRV_N5143_n_28426;
wire FE_OCP_DRV_N5144_n_28349;
wire FE_OCP_DRV_N5145_n_28349;
wire FE_OCP_DRV_N5146_n_29765;
wire FE_OCP_DRV_N5147_n_29765;
wire FE_OCP_DRV_N5148_n_31125;
wire FE_OCP_DRV_N5149_n_31125;
wire FE_OCP_DRV_N5150_n_31264;
wire FE_OCP_DRV_N5151_n_31264;
wire FE_OCP_DRV_N5152_n_31164;
wire FE_OCP_DRV_N5153_n_31164;
wire FE_OCP_DRV_N5154_n_31206;
wire FE_OCP_DRV_N5155_n_31206;
wire FE_OCP_DRV_N5156_n_25100;
wire FE_OCP_DRV_N5157_n_25100;
wire FE_OCP_DRV_N5158_n_26801;
wire FE_OCP_DRV_N5159_n_26801;
wire FE_OCP_DRV_N5160_n_30322;
wire FE_OCP_DRV_N5161_n_30322;
wire FE_OCP_DRV_N5303_n_29892;
wire FE_OCP_DRV_N5304_n_29892;
wire FE_OCP_DRV_N5353_n_18860;
wire FE_OCP_DRV_N5354_n_18860;
wire FE_OCP_DRV_N5355_n_19010;
wire FE_OCP_DRV_N5356_n_19010;
wire FE_OCP_DRV_N5357_n_12436;
wire FE_OCP_DRV_N5358_n_12436;
wire FE_OCP_DRV_N5359_n_13495;
wire FE_OCP_DRV_N5360_n_13495;
wire FE_OCP_DRV_N5361_n_21732;
wire FE_OCP_DRV_N5362_n_21732;
wire FE_OCP_DRV_N6260_n_37471;
wire FE_OCP_DRV_N6261_n_37471;
wire FE_OCP_DRV_N6262_FE_OCP_RBN5603_n_29056;
wire FE_OCP_DRV_N6263_FE_OCP_RBN5603_n_29056;
wire FE_OCP_DRV_N6264_n_9014;
wire FE_OCP_DRV_N6266_FE_OCP_RBN1823_n_19434;
wire FE_OCP_DRV_N6270_n_13264;
wire FE_OCP_DRV_N6271_n_13264;
wire FE_OCP_DRV_N6272_n_13330;
wire FE_OCP_DRV_N6273_n_13330;
wire FE_OCP_DRV_N6274_n_28582;
wire FE_OCP_DRV_N6275_n_28582;
wire FE_OCP_DRV_N6884_n_28829;
wire FE_OCP_DRV_N6885_n_28829;
wire FE_OCP_DRV_N6888_n_33945;
wire FE_OCP_DRV_N6889_n_33945;
wire FE_OCP_DRV_N6890_n_34296;
wire FE_OCP_DRV_N6891_n_34296;
wire FE_OCP_DRV_N6892_FE_OCPN6281_n_30612;
wire FE_OCP_DRV_N6893_FE_OCPN6281_n_30612;
wire FE_OCP_DRV_N6894_n_15391;
wire FE_OCP_DRV_N6895_n_15391;
wire FE_OCP_DRV_N6896_FE_OCPN1679_n_27315;
wire FE_OCP_DRV_N6897_FE_OCPN1679_n_27315;
wire FE_OCP_DRV_N6898_FE_OCPN5276_n_23590;
wire FE_OCP_DRV_N6899_FE_OCPN5276_n_23590;
wire FE_OCP_DRV_N6902_n_19354;
wire FE_OCP_DRV_N6903_n_19354;
wire FE_OCP_DRV_N6904_n_33945;
wire FE_OCP_DRV_N6906_n_34096;
wire FE_OCP_DRV_N6907_n_34096;
wire FE_OCP_DRV_N7074_n_7116;
wire FE_OCP_DRV_N7076_n_10105;
wire FE_OCP_DRV_N7077_n_10105;
wire FE_OCP_DRV_N7078_n_8992;
wire FE_OCP_DRV_N7079_n_8992;
wire FE_OCP_DRV_N7080_n_27130;
wire FE_OCP_DRV_N7081_n_27130;
wire FE_OCP_RBN1001_n_24079;
wire FE_OCP_RBN1002_n_24079;
wire FE_OCP_RBN1003_n_24079;
wire FE_OCP_RBN1004_n_25545;
wire FE_OCP_RBN1005_n_25545;
wire FE_OCP_RBN1006_n_24094;
wire FE_OCP_RBN1007_n_24175;
wire FE_OCP_RBN1009_n_24175;
wire FE_OCP_RBN1010_n_24175;
wire FE_OCP_RBN1011_n_24246;
wire FE_OCP_RBN1012_n_25826;
wire FE_OCP_RBN1013_n_25826;
wire FE_OCP_RBN1014_n_25826;
wire FE_OCP_RBN1015_n_25826;
wire FE_OCP_RBN1016_n_13601;
wire FE_OCP_RBN1017_n_24165;
wire FE_OCP_RBN1018_n_24165;
wire FE_OCP_RBN1019_n_24165;
wire FE_OCP_RBN1020_n_24181;
wire FE_OCP_RBN1021_n_24181;
wire FE_OCP_RBN1022_n_24181;
wire FE_OCP_RBN1023_n_24125;
wire FE_OCP_RBN1024_n_24125;
wire FE_OCP_RBN1025_n_17417;
wire FE_OCP_RBN1026_n_17417;
wire FE_OCP_RBN1027_n_17417;
wire FE_OCP_RBN1028_n_17417;
wire FE_OCP_RBN1032_n_25844;
wire FE_OCP_RBN1034_n_25844;
wire FE_OCP_RBN1035_FE_RN_557_0;
wire FE_OCP_RBN1036_FE_RN_557_0;
wire FE_OCP_RBN1037_n_45533;
wire FE_OCP_RBN1038_n_45533;
wire FE_OCP_RBN1039_n_45533;
wire FE_OCP_RBN1040_n_26158;
wire FE_OCP_RBN1105_n_18746;
wire FE_OCP_RBN1109_n_44061;
wire FE_OCP_RBN1118_delay_xor_ln22_unr15_stage6_stallmux_q_0_;
wire FE_OCP_RBN1120_delay_xor_ln22_unr12_stage5_stallmux_q_2_;
wire FE_OCP_RBN1121_delay_xor_ln22_unr12_stage5_stallmux_q_2_;
wire FE_OCP_RBN1130_n_18918;
wire FE_OCP_RBN1131_n_19077;
wire FE_OCP_RBN1132_n_19077;
wire FE_OCP_RBN1133_n_19077;
wire FE_OCP_RBN1134_n_19077;
wire FE_OCP_RBN1137_n_19270;
wire FE_OCP_RBN1138_n_19270;
wire FE_OCP_RBN1139_n_19270;
wire FE_OCP_RBN1140_n_19270;
wire FE_OCP_RBN1146_n_19353;
wire FE_OCP_RBN1150_n_18981;
wire FE_OCP_RBN1151_FE_RN_533_0;
wire FE_OCP_RBN1152_n_20910;
wire FE_OCP_RBN1153_n_20910;
wire FE_OCP_RBN1157_n_20336;
wire FE_OCP_RBN1159_n_20763;
wire FE_OCP_RBN1160_n_20763;
wire FE_OCP_RBN1161_n_20763;
wire FE_OCP_RBN1162_n_20763;
wire FE_OCP_RBN1163_n_24471;
wire FE_OCP_RBN1164_n_24471;
wire FE_OCP_RBN1166_n_25889;
wire FE_OCP_RBN1170_n_21318;
wire FE_OCP_RBN1171_n_25817;
wire FE_OCP_RBN1172_n_25817;
wire FE_OCP_RBN1173_n_22476;
wire FE_OCP_RBN1175_n_27593;
wire FE_OCP_RBN1176_n_27593;
wire FE_OCP_RBN1589_n_13460;
wire FE_OCP_RBN1590_n_13557;
wire FE_OCP_RBN1591_n_13557;
wire FE_OCP_RBN1592_n_13557;
wire FE_OCP_RBN1593_n_13557;
wire FE_OCP_RBN1594_n_13557;
wire FE_OCP_RBN1595_n_14823;
wire FE_OCP_RBN1596_n_14823;
wire FE_OCP_RBN1597_n_14763;
wire FE_OCP_RBN1598_n_14763;
wire FE_OCP_RBN1599_n_14763;
wire FE_OCP_RBN1600_n_14763;
wire FE_OCP_RBN1601_n_14638;
wire FE_OCP_RBN1602_n_14638;
wire FE_OCP_RBN1603_n_20995;
wire FE_OCP_RBN1604_n_20995;
wire FE_OCP_RBN1803_n_32647;
wire FE_OCP_RBN1804_n_27825;
wire FE_OCP_RBN1805_n_27934;
wire FE_OCP_RBN1807_n_13010;
wire FE_OCP_RBN1808_n_28968;
wire FE_OCP_RBN1809_n_18754;
wire FE_OCP_RBN1810_n_18754;
wire FE_OCP_RBN1811_n_33750;
wire FE_OCP_RBN1812_n_33750;
wire FE_OCP_RBN1813_n_33846;
wire FE_OCP_RBN1814_n_33846;
wire FE_OCP_RBN1815_n_33873;
wire FE_OCP_RBN1816_n_33873;
wire FE_OCP_RBN1817_n_19178;
wire FE_OCP_RBN1818_n_13858;
wire FE_OCP_RBN1819_n_13858;
wire FE_OCP_RBN1820_n_13858;
wire FE_OCP_RBN1821_n_13858;
wire FE_OCP_RBN1822_n_24473;
wire FE_OCP_RBN1823_n_19434;
wire FE_OCP_RBN1824_n_19434;
wire FE_OCP_RBN1825_n_19513;
wire FE_OCP_RBN1826_n_19513;
wire FE_OCP_RBN1827_n_19538;
wire FE_OCP_RBN1829_n_19528;
wire FE_OCP_RBN1831_n_19663;
wire FE_OCP_RBN1832_n_14197;
wire FE_OCP_RBN1833_n_14197;
wire FE_OCP_RBN1834_n_14664;
wire FE_OCP_RBN1836_n_20209;
wire FE_OCP_RBN1837_n_20215;
wire FE_OCP_RBN1838_n_20273;
wire FE_OCP_RBN1839_n_20273;
wire FE_OCP_RBN1840_n_20439;
wire FE_OCP_RBN1841_FE_RN_442_0;
wire FE_OCP_RBN1842_FE_RN_442_0;
wire FE_OCP_RBN1843_n_20640;
wire FE_OCP_RBN1844_n_20616;
wire FE_OCP_RBN1845_n_30492;
wire FE_OCP_RBN1846_n_30492;
wire FE_OCP_RBN1847_n_30428;
wire FE_OCP_RBN1848_FE_RN_578_0;
wire FE_OCP_RBN1849_FE_RN_578_0;
wire FE_OCP_RBN1850_n_25898;
wire FE_OCP_RBN1851_n_25898;
wire FE_OCP_RBN1855_n_20879;
wire FE_OCP_RBN1856_n_30731;
wire FE_OCP_RBN1857_n_30731;
wire FE_OCP_RBN1859_n_30731;
wire FE_OCP_RBN1862_n_26049;
wire FE_OCP_RBN1864_n_21163;
wire FE_OCP_RBN1865_n_21163;
wire FE_OCP_RBN1866_n_26407;
wire FE_OCP_RBN1867_n_26407;
wire FE_OCP_RBN1868_n_21358;
wire FE_OCP_RBN1869_n_21358;
wire FE_OCP_RBN1871_n_36489;
wire FE_OCP_RBN1872_n_36489;
wire FE_OCP_RBN1875_n_17689;
wire FE_OCP_RBN1876_n_27723;
wire FE_OCP_RBN1877_n_32382;
wire FE_OCP_RBN1878_n_27804;
wire FE_OCP_RBN2028_n_44722;
wire FE_OCP_RBN2029_n_44722;
wire FE_OCP_RBN2030_n_44722;
wire FE_OCP_RBN2034_n_44722;
wire FE_OCP_RBN2037_n_44722;
wire FE_OCP_RBN2038_n_44722;
wire FE_OCP_RBN2039_n_44722;
wire FE_OCP_RBN2040_n_28268;
wire FE_OCP_RBN2041_n_18269;
wire FE_OCP_RBN2042_n_18269;
wire FE_OCP_RBN2043_n_18269;
wire FE_OCP_RBN2044_n_12907;
wire FE_OCP_RBN2045_n_12907;
wire FE_OCP_RBN2046_n_12907;
wire FE_OCP_RBN2049_n_29056;
wire FE_OCP_RBN2050_n_13694;
wire FE_OCP_RBN2055_n_13784;
wire FE_OCP_RBN2056_n_13784;
wire FE_OCP_RBN2057_n_13784;
wire FE_OCP_RBN2058_n_13784;
wire FE_OCP_RBN2059_n_29380;
wire FE_OCP_RBN2060_n_29380;
wire FE_OCP_RBN2061_n_13813;
wire FE_OCP_RBN2062_n_19353;
wire FE_OCP_RBN2063_n_19353;
wire FE_OCP_RBN2064_n_19353;
wire FE_OCP_RBN2065_n_13913;
wire FE_OCP_RBN2066_n_14069;
wire FE_OCP_RBN2067_n_14069;
wire FE_OCP_RBN2068_n_14069;
wire FE_OCP_RBN2069_n_14069;
wire FE_OCP_RBN2070_n_14069;
wire FE_OCP_RBN2071_n_14120;
wire FE_OCP_RBN2073_n_14120;
wire FE_OCP_RBN2074_n_29603;
wire FE_OCP_RBN2075_n_14093;
wire FE_OCP_RBN2076_n_14149;
wire FE_OCP_RBN2077_n_14149;
wire FE_OCP_RBN2078_n_14149;
wire FE_OCP_RBN2079_n_14149;
wire FE_OCP_RBN2080_n_14554;
wire FE_OCP_RBN2081_n_14554;
wire FE_OCP_RBN2082_n_14554;
wire FE_OCP_RBN2083_n_14611;
wire FE_OCP_RBN2084_n_19970;
wire FE_OCP_RBN2085_n_14911;
wire FE_OCP_RBN2086_n_14911;
wire FE_OCP_RBN2087_n_14911;
wire FE_OCP_RBN2089_n_14964;
wire FE_OCP_RBN2090_n_14908;
wire FE_OCP_RBN2091_n_14909;
wire FE_OCP_RBN2092_n_14991;
wire FE_OCP_RBN2093_n_14991;
wire FE_OCP_RBN2094_n_47175;
wire FE_OCP_RBN2095_n_20325;
wire FE_OCP_RBN2096_n_20325;
wire FE_OCP_RBN2097_n_20325;
wire FE_OCP_RBN2098_n_20325;
wire FE_OCP_RBN2101_n_15083;
wire FE_OCP_RBN2102_n_15083;
wire FE_OCP_RBN2103_n_15286;
wire FE_OCP_RBN2104_n_30465;
wire FE_OCP_RBN2105_n_30465;
wire FE_OCP_RBN2106_n_30619;
wire FE_OCP_RBN2107_n_30747;
wire FE_OCP_RBN2108_n_15911;
wire FE_OCP_RBN2109_n_15911;
wire FE_OCP_RBN2110_n_15911;
wire FE_OCP_RBN2111_n_15911;
wire FE_OCP_RBN2112_n_20935;
wire FE_OCP_RBN2113_n_20935;
wire FE_OCP_RBN2114_n_20935;
wire FE_OCP_RBN2115_n_20935;
wire FE_OCP_RBN2118_n_22351;
wire FE_OCP_RBN2250_n_44061;
wire FE_OCP_RBN2258_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN2259_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN2260_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN2261_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN2262_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN2263_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN2264_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN2265_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN2266_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN2267_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN2268_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN2270_delay_xor_ln22_unr15_stage6_stallmux_q_2_;
wire FE_OCP_RBN2271_delay_xor_ln22_unr15_stage6_stallmux_q_5_;
wire FE_OCP_RBN2272_delay_xor_ln22_unr15_stage6_stallmux_q_5_;
wire FE_OCP_RBN2282_delay_sub_ln23_unr21_stage7_stallmux_q_1_;
wire FE_OCP_RBN2311_delay_sub_ln23_unr25_stage8_stallmux_q_1_;
wire FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_;
wire FE_OCP_RBN2337_delay_sub_ln21_0_unr23_stage9_stallmux_q_20_;
wire FE_OCP_RBN2338_delay_sub_ln21_0_unr23_stage9_stallmux_q_20_;
wire FE_OCP_RBN2369_n_44061;
wire FE_OCP_RBN2377_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN2378_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN2382_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN2385_n_22820;
wire FE_OCP_RBN2386_n_22650;
wire FE_OCP_RBN2387_n_23227;
wire FE_OCP_RBN2388_n_23227;
wire FE_OCP_RBN2389_n_23227;
wire FE_OCP_RBN2390_FE_RN_1364_0;
wire FE_OCP_RBN2392_n_16970;
wire FE_OCP_RBN2393_n_45697;
wire FE_OCP_RBN2394_n_45697;
wire FE_OCP_RBN2395_n_45697;
wire FE_OCP_RBN2396_n_45697;
wire FE_OCP_RBN2397_n_45697;
wire FE_OCP_RBN2398_n_45697;
wire FE_OCP_RBN2399_n_45697;
wire FE_OCP_RBN2400_n_45697;
wire FE_OCP_RBN2401_n_45697;
wire FE_OCP_RBN2402_n_45697;
wire FE_OCP_RBN2404_n_45697;
wire FE_OCP_RBN2405_n_45697;
wire FE_OCP_RBN2406_n_45697;
wire FE_OCP_RBN2407_n_6635;
wire FE_OCP_RBN2410_n_40631;
wire FE_OCP_RBN2411_n_44722;
wire FE_OCP_RBN2412_n_44722;
wire FE_OCP_RBN2413_n_44722;
wire FE_OCP_RBN2414_n_44722;
wire FE_OCP_RBN2415_n_44722;
wire FE_OCP_RBN2416_n_44722;
wire FE_OCP_RBN2417_n_44722;
wire FE_OCP_RBN2418_n_44083;
wire FE_OCP_RBN2422_n_23023;
wire FE_OCP_RBN2423_n_32554;
wire FE_OCP_RBN2426_n_11907;
wire FE_OCP_RBN2427_n_11907;
wire FE_OCP_RBN2428_n_37207;
wire FE_OCP_RBN2429_FE_RN_107_0;
wire FE_OCP_RBN2430_FE_RN_107_0;
wire FE_OCP_RBN2431_FE_RN_107_0;
wire FE_OCP_RBN2432_FE_RN_107_0;
wire FE_OCP_RBN2433_FE_RN_107_0;
wire FE_OCP_RBN2434_n_32702;
wire FE_OCP_RBN2435_FE_OCPN833_n_45450;
wire FE_OCP_RBN2436_FE_OCPN833_n_45450;
wire FE_OCP_RBN2437_FE_OCPN833_n_45450;
wire FE_OCP_RBN2438_FE_OCPN833_n_45450;
wire FE_OCP_RBN2439_n_6937;
wire FE_OCP_RBN2440_n_44798;
wire FE_OCP_RBN2441_n_44798;
wire FE_OCP_RBN2442_n_44798;
wire FE_OCP_RBN2443_n_44798;
wire FE_OCP_RBN2444_n_1675;
wire FE_OCP_RBN2445_n_1675;
wire FE_OCP_RBN2446_n_23079;
wire FE_OCP_RBN2447_n_12312;
wire FE_OCP_RBN2448_n_23246;
wire FE_OCP_RBN2449_n_23246;
wire FE_OCP_RBN2450_n_23246;
wire FE_OCP_RBN2451_n_32860;
wire FE_OCP_RBN2452_n_32860;
wire FE_OCP_RBN2453_n_32860;
wire FE_OCP_RBN2454_n_32860;
wire FE_OCP_RBN2460_n_12365;
wire FE_OCP_RBN2461_n_12365;
wire FE_OCP_RBN2462_n_23345;
wire FE_OCP_RBN2463_n_37449;
wire FE_OCP_RBN2464_n_7129;
wire FE_OCP_RBN2467_n_33034;
wire FE_OCP_RBN2468_n_33034;
wire FE_OCP_RBN2469_n_33034;
wire FE_OCP_RBN2476_n_33034;
wire FE_OCP_RBN2477_n_33034;
wire FE_OCP_RBN2478_n_1862;
wire FE_OCP_RBN2479_n_47245;
wire FE_OCP_RBN2480_FE_RN_734_0;
wire FE_OCP_RBN2481_FE_RN_734_0;
wire FE_OCP_RBN2482_n_37509;
wire FE_OCP_RBN2483_FE_RN_657_0;
wire FE_OCP_RBN2484_FE_RN_657_0;
wire FE_OCP_RBN2485_n_41213;
wire FE_OCP_RBN2490_FE_RN_1367_0;
wire FE_OCP_RBN2491_FE_RN_1367_0;
wire FE_OCP_RBN2492_FE_RN_1367_0;
wire FE_OCP_RBN2494_n_7349;
wire FE_OCP_RBN2495_n_18242;
wire FE_OCP_RBN2496_n_18242;
wire FE_OCP_RBN2497_n_18242;
wire FE_OCP_RBN2498_n_37624;
wire FE_OCP_RBN2499_FE_RN_1553_0;
wire FE_OCP_RBN2500_n_28773;
wire FE_OCP_RBN2502_n_33226;
wire FE_OCP_RBN2503_n_33226;
wire FE_OCP_RBN2505_n_33226;
wire FE_OCP_RBN2506_n_33226;
wire FE_OCP_RBN2507_n_37720;
wire FE_OCP_RBN2508_n_37720;
wire FE_OCP_RBN2509_n_41215;
wire FE_OCP_RBN2510_n_12800;
wire FE_OCP_RBN2511_n_12800;
wire FE_OCP_RBN2512_n_12800;
wire FE_OCP_RBN2513_n_28699;
wire FE_OCP_RBN2514_n_28699;
wire FE_OCP_RBN2515_n_45120;
wire FE_OCP_RBN2517_n_45120;
wire FE_OCP_RBN2519_n_12721;
wire FE_OCP_RBN2521_n_12721;
wire FE_OCP_RBN2522_n_12721;
wire FE_OCP_RBN2523_n_29017;
wire FE_OCP_RBN2524_n_28749;
wire FE_OCP_RBN2526_n_2086;
wire FE_OCP_RBN2528_n_2097;
wire FE_OCP_RBN2529_n_12731;
wire FE_OCP_RBN2530_n_13151;
wire FE_OCP_RBN2531_n_33372;
wire FE_OCP_RBN2532_n_33372;
wire FE_OCP_RBN2533_n_33372;
wire FE_OCP_RBN2534_n_33372;
wire FE_OCP_RBN2535_n_33568;
wire FE_OCP_RBN2536_n_12880;
wire FE_OCP_RBN2537_n_12880;
wire FE_OCP_RBN2538_n_12880;
wire FE_OCP_RBN2539_n_12880;
wire FE_OCP_RBN2540_n_12880;
wire FE_OCP_RBN2541_n_12880;
wire FE_OCP_RBN2542_n_12921;
wire FE_OCP_RBN2543_n_33584;
wire FE_OCP_RBN2544_n_33584;
wire FE_OCP_RBN2548_n_44881;
wire FE_OCP_RBN2549_n_44881;
wire FE_OCP_RBN2550_n_33664;
wire FE_OCP_RBN2551_n_33664;
wire FE_OCP_RBN2552_n_33697;
wire FE_OCP_RBN2553_n_33697;
wire FE_OCP_RBN2554_n_13141;
wire FE_OCP_RBN2555_n_13141;
wire FE_OCP_RBN2556_n_13141;
wire FE_OCP_RBN2557_n_13141;
wire FE_OCP_RBN2558_n_7665;
wire FE_OCP_RBN2559_n_13084;
wire FE_OCP_RBN2560_n_13084;
wire FE_OCP_RBN2561_n_13084;
wire FE_OCP_RBN2562_n_13084;
wire FE_OCP_RBN2563_n_13084;
wire FE_OCP_RBN2564_n_29110;
wire FE_OCP_RBN2565_n_29110;
wire FE_OCP_RBN2566_n_29163;
wire FE_OCP_RBN2567_n_29163;
wire FE_OCP_RBN2570_n_33735;
wire FE_OCP_RBN2571_n_2430;
wire FE_OCP_RBN2573_n_2558;
wire FE_OCP_RBN2574_n_2558;
wire FE_OCP_RBN2579_n_13154;
wire FE_OCP_RBN2580_n_13154;
wire FE_OCP_RBN2581_n_37913;
wire FE_OCP_RBN2582_n_29091;
wire FE_OCP_RBN2583_n_29091;
wire FE_OCP_RBN2584_n_29091;
wire FE_OCP_RBN2587_n_7743;
wire FE_OCP_RBN2588_n_7743;
wire FE_OCP_RBN2592_n_7743;
wire FE_OCP_RBN2593_n_7743;
wire FE_OCP_RBN2595_n_7743;
wire FE_OCP_RBN2597_n_7743;
wire FE_OCP_RBN2598_n_7743;
wire FE_OCP_RBN2599_n_7743;
wire FE_OCP_RBN2601_n_13483;
wire FE_OCP_RBN2602_n_13483;
wire FE_OCP_RBN2604_FE_OCPN855_n_7721;
wire FE_OCP_RBN2605_FE_OCPN855_n_7721;
wire FE_OCP_RBN2607_FE_OCPN855_n_7721;
wire FE_OCP_RBN2608_FE_OCPN855_n_7721;
wire FE_OCP_RBN2609_n_47235;
wire FE_OCP_RBN2610_n_29298;
wire FE_OCP_RBN2611_n_29298;
wire FE_OCP_RBN2612_FE_OCPN857_n_7802;
wire FE_OCP_RBN2613_FE_OCPN857_n_7802;
wire FE_OCP_RBN2614_FE_OCPN857_n_7802;
wire FE_OCP_RBN2616_FE_OCPN857_n_7802;
wire FE_OCP_RBN2620_n_24175;
wire FE_OCP_RBN2621_n_24175;
wire FE_OCP_RBN2622_n_24175;
wire FE_OCP_RBN2627_n_2737;
wire FE_OCP_RBN2629_n_2737;
wire FE_OCP_RBN2630_n_2737;
wire FE_OCP_RBN2631_n_9003;
wire FE_OCP_RBN2632_n_9003;
wire FE_OCP_RBN2633_n_9003;
wire FE_OCP_RBN2634_n_9003;
wire FE_OCP_RBN2635_n_29371;
wire FE_OCP_RBN2636_n_29371;
wire FE_OCP_RBN2637_n_33954;
wire FE_OCP_RBN2638_n_33954;
wire FE_OCP_RBN2639_n_13667;
wire FE_OCP_RBN2640_n_13667;
wire FE_OCP_RBN2641_n_13667;
wire FE_OCP_RBN2642_n_13667;
wire FE_OCP_RBN2644_n_13667;
wire FE_OCP_RBN2645_n_2747;
wire FE_OCP_RBN2646_n_2747;
wire FE_OCP_RBN2649_n_8073;
wire FE_OCP_RBN2650_n_29470;
wire FE_OCP_RBN2651_n_29470;
wire FE_OCP_RBN2652_n_29448;
wire FE_OCP_RBN2653_n_29448;
wire FE_OCP_RBN2654_FE_OCPN914_n_8091;
wire FE_OCP_RBN2655_FE_OCPN914_n_8091;
wire FE_OCP_RBN2656_FE_OCPN914_n_8091;
wire FE_OCP_RBN2659_n_2832;
wire FE_OCP_RBN2661_n_9304;
wire FE_OCP_RBN2662_n_19393;
wire FE_OCP_RBN2663_n_19393;
wire FE_OCP_RBN2664_n_24372;
wire FE_OCP_RBN2665_n_24372;
wire FE_OCP_RBN2666_n_24372;
wire FE_OCP_RBN2667_n_24408;
wire FE_OCP_RBN2668_n_29500;
wire FE_OCP_RBN2669_n_29500;
wire FE_OCP_RBN2670_n_46991;
wire FE_OCP_RBN2672_n_38534;
wire FE_OCP_RBN2673_n_38534;
wire FE_OCP_RBN2674_n_8163;
wire FE_OCP_RBN2675_n_8163;
wire FE_OCP_RBN2676_n_8163;
wire FE_OCP_RBN2677_n_8163;
wire FE_OCP_RBN2678_n_8163;
wire FE_OCP_RBN2680_n_38515;
wire FE_OCP_RBN2681_n_38515;
wire FE_OCP_RBN2682_n_38515;
wire FE_OCP_RBN2683_n_13818;
wire FE_OCP_RBN2684_n_13818;
wire FE_OCP_RBN2687_n_44100;
wire FE_OCP_RBN2688_n_44100;
wire FE_OCP_RBN2689_n_44100;
wire FE_OCP_RBN2690_n_8221;
wire FE_OCP_RBN2691_n_8221;
wire FE_OCP_RBN2692_n_8221;
wire FE_OCP_RBN2693_n_24436;
wire FE_OCP_RBN2694_n_24436;
wire FE_OCP_RBN2695_n_24436;
wire FE_OCP_RBN2696_n_13703;
wire FE_OCP_RBN2697_n_13703;
wire FE_OCP_RBN2701_n_8187;
wire FE_OCP_RBN2702_FE_RN_299_0;
wire FE_OCP_RBN2703_FE_RN_984_0;
wire FE_OCP_RBN2704_n_24510;
wire FE_OCP_RBN2705_n_47023;
wire FE_OCP_RBN2706_n_47023;
wire FE_OCP_RBN2708_n_24505;
wire FE_OCP_RBN2709_n_24505;
wire FE_OCP_RBN2711_n_19599;
wire FE_OCP_RBN2712_n_24501;
wire FE_OCP_RBN2713_n_24501;
wire FE_OCP_RBN2714_n_24501;
wire FE_OCP_RBN2715_n_24501;
wire FE_OCP_RBN2716_n_8242;
wire FE_OCP_RBN2717_n_8242;
wire FE_OCP_RBN2719_n_8242;
wire FE_OCP_RBN2720_n_19601;
wire FE_OCP_RBN2721_n_19601;
wire FE_OCP_RBN2722_n_8243;
wire FE_OCP_RBN2723_FE_RN_522_0;
wire FE_OCP_RBN2724_n_14018;
wire FE_OCP_RBN2725_n_14018;
wire FE_OCP_RBN2726_n_14018;
wire FE_OCP_RBN2727_n_14018;
wire FE_OCP_RBN2728_n_14072;
wire FE_OCP_RBN2729_n_14072;
wire FE_OCP_RBN2730_n_14072;
wire FE_OCP_RBN2731_n_14072;
wire FE_OCP_RBN2732_n_29657;
wire FE_OCP_RBN2733_n_29657;
wire FE_OCP_RBN2734_n_8402;
wire FE_OCP_RBN2735_n_8402;
wire FE_OCP_RBN2737_n_8402;
wire FE_OCP_RBN2739_n_8300;
wire FE_OCP_RBN2740_n_8398;
wire FE_OCP_RBN2741_n_14114;
wire FE_OCP_RBN2742_n_14114;
wire FE_OCP_RBN2743_n_14114;
wire FE_OCP_RBN2744_n_14114;
wire FE_OCP_RBN2745_n_19747;
wire FE_OCP_RBN2746_n_19747;
wire FE_OCP_RBN2747_n_8474;
wire FE_OCP_RBN2748_n_8474;
wire FE_OCP_RBN2749_n_14157;
wire FE_OCP_RBN2750_n_14157;
wire FE_OCP_RBN2751_FE_RN_1223_0;
wire FE_OCP_RBN2752_FE_RN_1223_0;
wire FE_OCP_RBN2753_n_3016;
wire FE_OCP_RBN2754_n_3016;
wire FE_OCP_RBN2756_n_13796;
wire FE_OCP_RBN2757_n_13796;
wire FE_OCP_RBN2758_n_13796;
wire FE_OCP_RBN2759_n_13796;
wire FE_OCP_RBN2760_n_13796;
wire FE_OCP_RBN2762_n_13796;
wire FE_OCP_RBN2765_n_38530;
wire FE_OCP_RBN2766_n_38530;
wire FE_OCP_RBN2767_n_3035;
wire FE_OCP_RBN2768_n_3167;
wire FE_OCP_RBN2769_n_3238;
wire FE_OCP_RBN2771_n_4336;
wire FE_OCP_RBN2772_n_45521;
wire FE_OCP_RBN2775_n_8637;
wire FE_OCP_RBN2776_n_8637;
wire FE_OCP_RBN2778_n_8599;
wire FE_OCP_RBN2779_n_8599;
wire FE_OCP_RBN2780_n_8664;
wire FE_OCP_RBN2781_n_8664;
wire FE_OCP_RBN2782_n_8664;
wire FE_OCP_RBN2783_n_8664;
wire FE_OCP_RBN2785_n_8767;
wire FE_OCP_RBN2786_n_8767;
wire FE_OCP_RBN2789_n_8767;
wire FE_OCP_RBN2790_n_8767;
wire FE_OCP_RBN2791_FE_RN_368_0;
wire FE_OCP_RBN2796_n_3250;
wire FE_OCP_RBN2797_n_8530;
wire FE_OCP_RBN2798_n_8817;
wire FE_OCP_RBN2799_n_8817;
wire FE_OCP_RBN2800_n_8817;
wire FE_OCP_RBN2803_n_3220;
wire FE_OCP_RBN2804_n_3261;
wire FE_OCP_RBN2808_n_3338;
wire FE_OCP_RBN2810_n_8542;
wire FE_OCP_RBN2811_n_8542;
wire FE_OCP_RBN2812_n_8835;
wire FE_OCP_RBN2813_n_8835;
wire FE_OCP_RBN2814_n_14441;
wire FE_OCP_RBN2815_n_14441;
wire FE_OCP_RBN2816_n_34509;
wire FE_OCP_RBN2817_n_8939;
wire FE_OCP_RBN2819_n_13962;
wire FE_OCP_RBN2820_n_13962;
wire FE_OCP_RBN2825_n_13962;
wire FE_OCP_RBN2828_n_13962;
wire FE_OCP_RBN2829_n_13962;
wire FE_OCP_RBN2830_n_13962;
wire FE_OCP_RBN2832_n_13962;
wire FE_OCP_RBN2833_n_13962;
wire FE_OCP_RBN2834_n_13962;
wire FE_OCP_RBN2835_n_13962;
wire FE_OCP_RBN2836_n_13962;
wire FE_OCP_RBN2837_n_13962;
wire FE_OCP_RBN2838_n_13962;
wire FE_OCP_RBN2839_n_8974;
wire FE_OCP_RBN2841_n_9044;
wire FE_OCP_RBN2842_n_9044;
wire FE_OCP_RBN2845_n_47018;
wire FE_OCP_RBN2846_n_47018;
wire FE_OCP_RBN2847_n_47018;
wire FE_OCP_RBN2850_n_3645;
wire FE_OCP_RBN2851_n_4905;
wire FE_OCP_RBN2852_n_4905;
wire FE_OCP_RBN2853_n_4905;
wire FE_OCP_RBN2854_n_8692;
wire FE_OCP_RBN2856_n_8755;
wire FE_OCP_RBN2857_n_9082;
wire FE_OCP_RBN2858_n_9082;
wire FE_OCP_RBN2859_n_9082;
wire FE_OCP_RBN2860_n_29800;
wire FE_OCP_RBN2861_n_44921;
wire FE_OCP_RBN2863_n_3468;
wire FE_OCP_RBN2864_n_8714;
wire FE_OCP_RBN2865_n_8850;
wire FE_OCP_RBN2866_n_9347;
wire FE_OCP_RBN2867_n_9347;
wire FE_OCP_RBN2868_n_9188;
wire FE_OCP_RBN2869_n_9188;
wire FE_OCP_RBN2880_n_3539;
wire FE_OCP_RBN2881_n_8872;
wire FE_OCP_RBN2884_n_20127;
wire FE_OCP_RBN2885_n_8806;
wire FE_OCP_RBN2886_n_9017;
wire FE_OCP_RBN2887_n_9492;
wire FE_OCP_RBN2888_n_9492;
wire FE_OCP_RBN2889_n_9492;
wire FE_OCP_RBN2890_n_14460;
wire FE_OCP_RBN2891_n_14460;
wire FE_OCP_RBN2892_n_14460;
wire FE_OCP_RBN2895_n_35003;
wire FE_OCP_RBN2896_n_35003;
wire FE_OCP_RBN2897_n_38750;
wire FE_OCP_RBN2899_n_3807;
wire FE_OCP_RBN2900_n_3807;
wire FE_OCP_RBN2901_n_3643;
wire FE_OCP_RBN2902_n_8902;
wire FE_OCP_RBN2903_n_8902;
wire FE_OCP_RBN2904_n_14590;
wire FE_OCP_RBN2905_n_14590;
wire FE_OCP_RBN2907_n_25238;
wire FE_OCP_RBN2910_n_25178;
wire FE_OCP_RBN2911_n_25178;
wire FE_OCP_RBN2915_n_3878;
wire FE_OCP_RBN2920_n_3878;
wire FE_OCP_RBN2921_n_3878;
wire FE_OCP_RBN2922_n_9030;
wire FE_OCP_RBN2923_n_9070;
wire FE_OCP_RBN2924_n_9198;
wire FE_OCP_RBN2926_n_14684;
wire FE_OCP_RBN2927_n_14684;
wire FE_OCP_RBN2928_n_14923;
wire FE_OCP_RBN2929_n_34971;
wire FE_OCP_RBN2930_n_34971;
wire FE_OCP_RBN2932_n_9075;
wire FE_OCP_RBN2933_n_9075;
wire FE_OCP_RBN2934_n_9075;
wire FE_OCP_RBN2935_n_25401;
wire FE_OCP_RBN2936_n_8981;
wire FE_OCP_RBN2937_n_8981;
wire FE_OCP_RBN2938_n_47013;
wire FE_OCP_RBN2939_n_47013;
wire FE_OCP_RBN2941_n_4101;
wire FE_OCP_RBN2942_n_4101;
wire FE_OCP_RBN2943_n_20242;
wire FE_OCP_RBN2944_n_20242;
wire FE_OCP_RBN2950_n_4158;
wire FE_OCP_RBN2951_n_3867;
wire FE_OCP_RBN2952_n_3867;
wire FE_OCP_RBN2953_n_3841;
wire FE_OCP_RBN2960_n_4046;
wire FE_OCP_RBN2961_n_4046;
wire FE_OCP_RBN2962_n_4046;
wire FE_OCP_RBN2963_n_4046;
wire FE_OCP_RBN2964_n_4046;
wire FE_OCP_RBN2965_n_4046;
wire FE_OCP_RBN2966_n_4046;
wire FE_OCP_RBN2967_n_4046;
wire FE_OCP_RBN2968_n_4046;
wire FE_OCP_RBN2969_n_4046;
wire FE_OCP_RBN2970_n_9676;
wire FE_OCP_RBN2971_n_9676;
wire FE_OCP_RBN2973_n_14768;
wire FE_OCP_RBN2976_n_25295;
wire FE_OCP_RBN2977_n_25509;
wire FE_OCP_RBN2978_n_25562;
wire FE_OCP_RBN2979_n_35213;
wire FE_OCP_RBN2980_n_35213;
wire FE_OCP_RBN2981_n_14814;
wire FE_OCP_RBN2982_n_14814;
wire FE_OCP_RBN2983_n_14814;
wire FE_OCP_RBN2984_n_9247;
wire FE_OCP_RBN2985_n_9247;
wire FE_OCP_RBN2987_n_4238;
wire FE_OCP_RBN2988_n_9182;
wire FE_OCP_RBN2989_n_9182;
wire FE_OCP_RBN2990_n_4041;
wire FE_OCP_RBN2991_n_4041;
wire FE_OCP_RBN2992_n_9413;
wire FE_OCP_RBN2999_n_20374;
wire FE_OCP_RBN3000_n_20374;
wire FE_OCP_RBN3001_n_20400;
wire FE_OCP_RBN3002_n_20400;
wire FE_OCP_RBN3003_n_20432;
wire FE_OCP_RBN3005_n_14905;
wire FE_OCP_RBN3006_n_14905;
wire FE_OCP_RBN3007_n_15206;
wire FE_OCP_RBN3008_n_15206;
wire FE_OCP_RBN3011_n_9565;
wire FE_OCP_RBN3012_n_14985;
wire FE_OCP_RBN3013_n_14985;
wire FE_OCP_RBN3014_n_15055;
wire FE_OCP_RBN3015_n_15300;
wire FE_OCP_RBN3016_n_15300;
wire FE_OCP_RBN3017_n_20404;
wire FE_OCP_RBN3018_n_20404;
wire FE_OCP_RBN3021_n_15319;
wire FE_OCP_RBN3022_n_15319;
wire FE_OCP_RBN3023_n_47011;
wire FE_OCP_RBN3024_n_47011;
wire FE_OCP_RBN3025_n_4065;
wire FE_OCP_RBN3026_n_4699;
wire FE_OCP_RBN3028_n_9584;
wire FE_OCP_RBN3029_n_9584;
wire FE_OCP_RBN3030_n_9624;
wire FE_OCP_RBN3031_n_9624;
wire FE_OCP_RBN3032_n_15150;
wire FE_OCP_RBN3033_n_9629;
wire FE_OCP_RBN3034_n_9629;
wire FE_OCP_RBN3036_n_15079;
wire FE_OCP_RBN3037_n_15079;
wire FE_OCP_RBN3039_n_9494;
wire FE_OCP_RBN3040_n_45139;
wire FE_OCP_RBN3041_n_45139;
wire FE_OCP_RBN3042_n_4296;
wire FE_OCP_RBN3043_n_4296;
wire FE_OCP_RBN3044_n_4449;
wire FE_OCP_RBN3045_n_9621;
wire FE_OCP_RBN3048_n_15200;
wire FE_OCP_RBN3049_n_15200;
wire FE_OCP_RBN3050_n_4376;
wire FE_OCP_RBN3052_n_10100;
wire FE_OCP_RBN3057_n_10100;
wire FE_OCP_RBN3058_n_15595;
wire FE_OCP_RBN3059_n_15595;
wire FE_OCP_RBN3060_n_15595;
wire FE_OCP_RBN3061_n_30575;
wire FE_OCP_RBN3062_n_9859;
wire FE_OCP_RBN3063_n_9859;
wire FE_OCP_RBN3064_n_9892;
wire FE_OCP_RBN3065_n_9892;
wire FE_OCP_RBN3066_n_4294;
wire FE_OCP_RBN3067_n_4294;
wire FE_OCP_RBN3068_n_9910;
wire FE_OCP_RBN3069_n_9910;
wire FE_OCP_RBN3070_n_15275;
wire FE_OCP_RBN3071_n_15433;
wire FE_OCP_RBN3072_n_15433;
wire FE_OCP_RBN3073_n_15706;
wire FE_OCP_RBN3074_n_15706;
wire FE_OCP_RBN3075_n_15706;
wire FE_OCP_RBN3076_n_25816;
wire FE_OCP_RBN3077_n_25816;
wire FE_OCP_RBN3078_n_25816;
wire FE_OCP_RBN3079_n_30643;
wire FE_OCP_RBN3080_n_30643;
wire FE_OCP_RBN3081_n_39514;
wire FE_OCP_RBN3082_n_15314;
wire FE_OCP_RBN3083_n_15314;
wire FE_OCP_RBN3084_n_15314;
wire FE_OCP_RBN3086_n_10015;
wire FE_OCP_RBN3087_n_4458;
wire FE_OCP_RBN3088_n_4458;
wire FE_OCP_RBN3089_n_4872;
wire FE_OCP_RBN3090_n_4872;
wire FE_OCP_RBN3091_n_10023;
wire FE_OCP_RBN3092_n_10023;
wire FE_OCP_RBN3093_n_10023;
wire FE_OCP_RBN3094_n_10023;
wire FE_OCP_RBN3095_n_10023;
wire FE_OCP_RBN3098_n_15561;
wire FE_OCP_RBN3099_n_15561;
wire FE_OCP_RBN3102_n_15768;
wire FE_OCP_RBN3103_n_20710;
wire FE_OCP_RBN3105_n_25819;
wire FE_OCP_RBN3106_n_25849;
wire FE_OCP_RBN3107_n_39531;
wire FE_OCP_RBN3108_n_39531;
wire FE_OCP_RBN3109_n_15817;
wire FE_OCP_RBN3110_n_15817;
wire FE_OCP_RBN3111_n_15817;
wire FE_OCP_RBN3112_n_10025;
wire FE_OCP_RBN3113_n_10195;
wire FE_OCP_RBN3114_n_10198;
wire FE_OCP_RBN3115_n_10198;
wire FE_OCP_RBN3116_n_10198;
wire FE_OCP_RBN3118_n_20812;
wire FE_OCP_RBN3120_n_4751;
wire FE_OCP_RBN3121_n_4751;
wire FE_OCP_RBN3122_n_4784;
wire FE_OCP_RBN3123_n_4784;
wire FE_OCP_RBN3124_n_5121;
wire FE_OCP_RBN3125_n_15856;
wire FE_OCP_RBN3126_n_21051;
wire FE_OCP_RBN3127_n_21051;
wire FE_OCP_RBN3128_n_21051;
wire FE_OCP_RBN3129_n_21051;
wire FE_OCP_RBN3130_n_21051;
wire FE_OCP_RBN3131_n_21051;
wire FE_OCP_RBN3134_n_46982;
wire FE_OCP_RBN3135_n_10274;
wire FE_OCP_RBN3136_n_10274;
wire FE_OCP_RBN3137_n_10326;
wire FE_OCP_RBN3138_n_10326;
wire FE_OCP_RBN3140_n_30849;
wire FE_OCP_RBN3141_n_30849;
wire FE_OCP_RBN3143_n_4858;
wire FE_OCP_RBN3144_n_4858;
wire FE_OCP_RBN3145_n_5085;
wire FE_OCP_RBN3146_n_10369;
wire FE_OCP_RBN3147_n_10369;
wire FE_OCP_RBN3148_n_15584;
wire FE_OCP_RBN3149_n_15553;
wire FE_OCP_RBN3150_n_25925;
wire FE_OCP_RBN3152_n_46962;
wire FE_OCP_RBN3153_n_15804;
wire FE_OCP_RBN3154_n_15804;
wire FE_OCP_RBN3155_n_4925;
wire FE_OCP_RBN3156_n_4925;
wire FE_OCP_RBN3160_n_10399;
wire FE_OCP_RBN3161_n_10399;
wire FE_OCP_RBN3167_n_44211;
wire FE_OCP_RBN3168_n_44211;
wire FE_OCP_RBN3169_n_44211;
wire FE_OCP_RBN3170_n_44211;
wire FE_OCP_RBN3171_n_44211;
wire FE_OCP_RBN3172_n_10134;
wire FE_OCP_RBN3173_n_26178;
wire FE_OCP_RBN3174_n_26158;
wire FE_OCP_RBN3175_n_31001;
wire FE_OCP_RBN3176_n_39640;
wire FE_OCP_RBN3177_n_39640;
wire FE_OCP_RBN3178_n_16088;
wire FE_OCP_RBN3179_n_16088;
wire FE_OCP_RBN3180_n_4959;
wire FE_OCP_RBN3181_n_10477;
wire FE_OCP_RBN3182_n_10477;
wire FE_OCP_RBN3185_n_15599;
wire FE_OCP_RBN3186_n_15599;
wire FE_OCP_RBN3190_n_15599;
wire FE_OCP_RBN3192_n_15599;
wire FE_OCP_RBN3193_n_15599;
wire FE_OCP_RBN3194_n_15599;
wire FE_OCP_RBN3195_n_15599;
wire FE_OCP_RBN3196_n_15599;
wire FE_OCP_RBN3197_n_15599;
wire FE_OCP_RBN3198_n_15599;
wire FE_OCP_RBN3199_n_15599;
wire FE_OCP_RBN3202_n_15900;
wire FE_OCP_RBN3203_n_15900;
wire FE_OCP_RBN3204_n_15900;
wire FE_OCP_RBN3205_n_26042;
wire FE_OCP_RBN3206_n_35517;
wire FE_OCP_RBN3207_n_39662;
wire FE_OCP_RBN3209_n_5221;
wire FE_OCP_RBN3210_n_21203;
wire FE_OCP_RBN3211_n_21203;
wire FE_OCP_RBN3212_n_10568;
wire FE_OCP_RBN3213_n_10568;
wire FE_OCP_RBN3214_n_10568;
wire FE_OCP_RBN3215_n_5003;
wire FE_OCP_RBN3216_n_5003;
wire FE_OCP_RBN3217_n_15758;
wire FE_OCP_RBN3218_n_15992;
wire FE_OCP_RBN3219_n_15992;
wire FE_OCP_RBN3220_n_15992;
wire FE_OCP_RBN3221_n_21242;
wire FE_OCP_RBN3222_n_21242;
wire FE_OCP_RBN3224_n_39575;
wire FE_OCP_RBN3225_n_39575;
wire FE_OCP_RBN3226_n_39575;
wire FE_OCP_RBN3227_n_10644;
wire FE_OCP_RBN3228_n_10644;
wire FE_OCP_RBN3229_n_10644;
wire FE_OCP_RBN3230_n_31107;
wire FE_OCP_RBN3231_n_31107;
wire FE_OCP_RBN3233_n_16041;
wire FE_OCP_RBN3234_n_16041;
wire FE_OCP_RBN3235_n_16041;
wire FE_OCP_RBN3236_n_5130;
wire FE_OCP_RBN3237_n_5130;
wire FE_OCP_RBN3238_n_5307;
wire FE_OCP_RBN3239_n_5307;
wire FE_OCP_RBN3240_n_10612;
wire FE_OCP_RBN3241_n_10612;
wire FE_OCP_RBN3242_n_10676;
wire FE_OCP_RBN3243_n_10676;
wire FE_OCP_RBN3244_n_21269;
wire FE_OCP_RBN3245_n_21351;
wire FE_OCP_RBN3246_n_26169;
wire FE_OCP_RBN3247_n_26169;
wire FE_OCP_RBN3248_n_39697;
wire FE_OCP_RBN3249_n_39697;
wire FE_OCP_RBN3250_n_21312;
wire FE_OCP_RBN3251_n_21312;
wire FE_OCP_RBN3252_n_26276;
wire FE_OCP_RBN3253_n_26276;
wire FE_OCP_RBN3254_n_5478;
wire FE_OCP_RBN3255_n_10454;
wire FE_OCP_RBN3256_n_16113;
wire FE_OCP_RBN3257_n_42998;
wire FE_OCP_RBN3258_n_42998;
wire FE_OCP_RBN3259_n_21360;
wire FE_OCP_RBN3260_n_21360;
wire FE_OCP_RBN3261_n_21360;
wire FE_OCP_RBN3263_n_5531;
wire FE_OCP_RBN3265_n_10852;
wire FE_OCP_RBN3266_n_26160;
wire FE_OCP_RBN3269_n_26160;
wire FE_OCP_RBN3272_n_31239;
wire FE_OCP_RBN3273_n_31239;
wire FE_OCP_RBN3274_n_26464;
wire FE_OCP_RBN3275_n_26464;
wire FE_OCP_RBN3276_n_5284;
wire FE_OCP_RBN3277_n_5284;
wire FE_OCP_RBN3279_FE_RN_1496_0;
wire FE_OCP_RBN3281_n_5614;
wire FE_OCP_RBN3283_n_26316;
wire FE_OCP_RBN3284_n_39674;
wire FE_OCP_RBN3285_n_39674;
wire FE_OCP_RBN3286_n_5656;
wire FE_OCP_RBN3287_n_5656;
wire FE_OCP_RBN3288_n_10915;
wire FE_OCP_RBN3289_n_10915;
wire FE_OCP_RBN3290_n_35539;
wire FE_OCP_RBN3291_n_35539;
wire FE_OCP_RBN3292_n_35539;
wire FE_OCP_RBN3293_n_35539;
wire FE_OCP_RBN3294_n_35539;
wire FE_OCP_RBN3295_n_35539;
wire FE_OCP_RBN3297_n_35539;
wire FE_OCP_RBN3298_n_35539;
wire FE_OCP_RBN3299_n_35539;
wire FE_OCP_RBN3300_n_35539;
wire FE_OCP_RBN3301_n_35539;
wire FE_OCP_RBN3302_n_35539;
wire FE_OCP_RBN3303_n_35539;
wire FE_OCP_RBN3306_n_43022;
wire FE_OCP_RBN3307_n_43022;
wire FE_OCP_RBN3308_n_43022;
wire FE_OCP_RBN3309_n_43022;
wire FE_OCP_RBN3310_n_43022;
wire FE_OCP_RBN3311_n_43022;
wire FE_OCP_RBN3312_n_43022;
wire FE_OCP_RBN3313_n_43022;
wire FE_OCP_RBN3315_n_43022;
wire FE_OCP_RBN3318_n_5555;
wire FE_OCP_RBN3319_n_5555;
wire FE_OCP_RBN3320_n_42959;
wire FE_OCP_RBN3321_n_42959;
wire FE_OCP_RBN3322_n_5586;
wire FE_OCP_RBN3324_n_5813;
wire FE_OCP_RBN3325_n_5813;
wire FE_OCP_RBN3326_n_5813;
wire FE_OCP_RBN3327_n_21616;
wire FE_OCP_RBN3328_n_21616;
wire FE_OCP_RBN3329_n_39685;
wire FE_OCP_RBN3330_n_11087;
wire FE_OCP_RBN3331_n_11087;
wire FE_OCP_RBN3333_n_39942;
wire FE_OCP_RBN3336_n_39942;
wire FE_OCP_RBN3337_n_39942;
wire FE_OCP_RBN3339_n_39942;
wire FE_OCP_RBN3340_n_39942;
wire FE_OCP_RBN3341_n_39942;
wire FE_OCP_RBN3342_n_39942;
wire FE_OCP_RBN3343_n_39942;
wire FE_OCP_RBN3344_n_39942;
wire FE_OCP_RBN3345_n_39942;
wire FE_OCP_RBN3346_n_47269;
wire FE_OCP_RBN3347_n_47269;
wire FE_OCP_RBN3348_n_47269;
wire FE_OCP_RBN3351_n_21812;
wire FE_OCP_RBN3352_FE_OFN760_n_46337;
wire FE_OCP_RBN3355_FE_RN_1058_0;
wire FE_OCP_RBN3356_FE_RN_1058_0;
wire FE_OCP_RBN3357_n_6013;
wire FE_OCP_RBN3358_n_11275;
wire FE_OCP_RBN3359_n_11275;
wire FE_OCP_RBN3360_n_16596;
wire FE_OCP_RBN3361_n_21847;
wire FE_OCP_RBN3362_n_21951;
wire FE_OCP_RBN3365_n_31520;
wire FE_OCP_RBN3368_n_31520;
wire FE_OCP_RBN3369_n_31520;
wire FE_OCP_RBN3370_n_31520;
wire FE_OCP_RBN3371_n_36490;
wire FE_OCP_RBN3372_n_43046;
wire FE_OCP_RBN3373_n_43046;
wire FE_OCP_RBN3374_n_43046;
wire FE_OCP_RBN3375_n_43046;
wire FE_OCP_RBN3377_n_44342;
wire FE_OCP_RBN3380_n_6034;
wire FE_OCP_RBN3381_n_36547;
wire FE_OCP_RBN3382_n_11405;
wire FE_OCP_RBN3383_n_11405;
wire FE_OCP_RBN3384_n_11439;
wire FE_OCP_RBN3386_n_11439;
wire FE_OCP_RBN3387_n_17130;
wire FE_OCP_RBN3388_n_31819;
wire FE_OCP_RBN3390_n_31819;
wire FE_OCP_RBN3391_n_31819;
wire FE_OCP_RBN3394_FE_RN_1094_0;
wire FE_OCP_RBN3395_FE_RN_1094_0;
wire FE_OCP_RBN3396_n_11486;
wire FE_OCP_RBN3398_n_11486;
wire FE_OCP_RBN3401_n_17233;
wire FE_OCP_RBN3402_n_43775;
wire FE_OCP_RBN3403_n_6205;
wire FE_OCP_RBN3404_n_6205;
wire FE_OCP_RBN3405_n_6205;
wire FE_OCP_RBN3406_n_32143;
wire FE_OCP_RBN3407_n_11560;
wire FE_OCP_RBN3408_n_22604;
wire FE_OCP_RBN3409_n_32072;
wire FE_OCP_RBN3410_n_36706;
wire FE_OCP_RBN3411_n_43811;
wire FE_OCP_RBN3412_n_43829;
wire FE_OCP_RBN3413_FE_OCPN891_n_31944;
wire FE_OCP_RBN3414_FE_OCPN891_n_31944;
wire FE_OCP_RBN3416_n_22564;
wire FE_OCP_RBN3417_n_22564;
wire FE_OCP_RBN3418_n_27590;
wire FE_OCP_RBN3419_n_32130;
wire FE_OCP_RBN3420_n_40300;
wire FE_OCP_RBN3421_n_32254;
wire FE_OCP_RBN3424_FE_RN_1622_0;
wire FE_OCP_RBN3425_n_11754;
wire FE_OCP_RBN3426_n_11810;
wire FE_OCP_RBN3427_n_17510;
wire FE_OCP_RBN3428_n_32180;
wire FE_OCP_RBN3429_n_36664;
wire FE_OCP_RBN3430_n_40563;
wire FE_OCP_RBN3431_n_43880;
wire FE_OCP_RBN3432_n_32239;
wire FE_OCP_RBN3434_n_6379;
wire FE_OCP_RBN3435_n_6379;
wire FE_OCP_RBN3436_n_6485;
wire FE_OCP_RBN3437_n_11980;
wire FE_OCP_RBN3438_n_32232;
wire FE_OCP_RBN3441_n_32266;
wire FE_OCP_RBN3442_n_32266;
wire FE_OCP_RBN3443_n_6471;
wire FE_OCP_RBN3444_n_6513;
wire FE_OCP_RBN3445_n_6513;
wire FE_OCP_RBN3446_n_6513;
wire FE_OCP_RBN3449_n_43777;
wire FE_OCP_RBN3450_n_17697;
wire FE_OCP_RBN3451_n_22710;
wire FE_OCP_RBN3453_n_27632;
wire FE_OCP_RBN3454_n_6557;
wire FE_OCP_RBN3455_n_6557;
wire FE_OCP_RBN3456_n_22709;
wire FE_OCP_RBN3458_n_12196;
wire FE_OCP_RBN3463_n_32316;
wire FE_OCP_RBN3464_n_43836;
wire FE_OCP_RBN3702_n_11788;
wire FE_OCP_RBN3703_n_12904;
wire FE_OCP_RBN3706_n_18716;
wire FE_OCP_RBN3707_n_18716;
wire FE_OCP_RBN3709_n_29055;
wire FE_OCP_RBN3710_n_29055;
wire FE_OCP_RBN3711_n_19116;
wire FE_OCP_RBN3713_n_19241;
wire FE_OCP_RBN3714_n_19241;
wire FE_OCP_RBN3715_n_19241;
wire FE_OCP_RBN3716_n_19241;
wire FE_OCP_RBN3717_n_19535;
wire FE_OCP_RBN3718_n_20621;
wire FE_OCP_RBN3719_n_20621;
wire FE_OCP_RBN3720_n_20621;
wire FE_OCP_RBN3721_n_20621;
wire FE_OCP_RBN3722_n_30776;
wire FE_OCP_RBN3723_n_21442;
wire FE_OCP_RBN3762_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN3815_n_45209;
wire FE_OCP_RBN3818_n_45622;
wire FE_OCP_RBN3844_delay_sub_ln23_unr13_stage5_stallmux_q_1_;
wire FE_OCP_RBN3845_delay_sub_ln23_unr13_stage5_stallmux_q_1_;
wire FE_OCP_RBN3871_n_44061;
wire FE_OCP_RBN3879_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN3881_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN3938_n_46254;
wire FE_OCP_RBN3939_n_46254;
wire FE_OCP_RBN3963_delay_sub_ln21_unr24_stage9_stallmux_q_8_;
wire FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_;
wire FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_;
wire FE_OCP_RBN3966_n_44061;
wire FE_OCP_RBN3967_n_44061;
wire FE_OCP_RBN3968_n_44061;
wire FE_OCP_RBN3975_n_45224;
wire FE_OCP_RBN3976_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN3979_n_22972;
wire FE_OCP_RBN3980_n_32436;
wire FE_OCP_RBN3982_n_27911;
wire FE_OCP_RBN3984_n_32791;
wire FE_OCP_RBN3985_FE_RN_158_0;
wire FE_OCP_RBN3986_FE_RN_158_0;
wire FE_OCP_RBN3988_n_32772;
wire FE_OCP_RBN3989_n_32772;
wire FE_OCP_RBN3990_n_32772;
wire FE_OCP_RBN3991_FE_RN_1579_0;
wire FE_OCP_RBN3997_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN3998_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN4002_n_33015;
wire FE_OCP_RBN4003_n_33015;
wire FE_OCP_RBN4004_n_33015;
wire FE_OCP_RBN4005_n_33015;
wire FE_OCP_RBN4006_n_32860;
wire FE_OCP_RBN4007_n_32860;
wire FE_OCP_RBN4008_n_32860;
wire FE_OCP_RBN4009_n_32860;
wire FE_OCP_RBN4011_n_1864;
wire FE_OCP_RBN4012_n_1864;
wire FE_OCP_RBN4013_n_33034;
wire FE_OCP_RBN4014_n_33034;
wire FE_OCP_RBN4015_n_33034;
wire FE_OCP_RBN4016_n_33034;
wire FE_OCP_RBN4017_n_33034;
wire FE_OCP_RBN4018_n_33034;
wire FE_OCP_RBN4019_n_33034;
wire FE_OCP_RBN4020_n_33034;
wire FE_OCP_RBN4021_n_33034;
wire FE_OCP_RBN4022_n_33034;
wire FE_OCP_RBN4023_n_37577;
wire FE_OCP_RBN4024_n_37577;
wire FE_OCP_RBN4025_n_37577;
wire FE_OCP_RBN4026_n_37577;
wire FE_OCP_RBN4027_n_37577;
wire FE_OCP_RBN4028_n_28458;
wire FE_OCP_RBN4030_n_28458;
wire FE_OCP_RBN4031_n_28458;
wire FE_OCP_RBN4032_n_37690;
wire FE_OCP_RBN4033_n_37690;
wire FE_OCP_RBN4034_n_37690;
wire FE_OCP_RBN4035_n_28651;
wire FE_OCP_RBN4036_n_28651;
wire FE_OCP_RBN4037_n_12904;
wire FE_OCP_RBN4038_n_2059;
wire FE_OCP_RBN4040_n_37707;
wire FE_OCP_RBN4041_n_37707;
wire FE_OCP_RBN4042_n_37707;
wire FE_OCP_RBN4043_n_41258;
wire FE_OCP_RBN4044_n_41298;
wire FE_OCP_RBN4045_n_41298;
wire FE_OCP_RBN4046_n_41298;
wire FE_OCP_RBN4047_n_12721;
wire FE_OCP_RBN4048_n_12721;
wire FE_OCP_RBN4049_n_33491;
wire FE_OCP_RBN4052_n_2086;
wire FE_OCP_RBN4053_n_2086;
wire FE_OCP_RBN4054_n_41325;
wire FE_OCP_RBN4055_n_41325;
wire FE_OCP_RBN4058_n_44875;
wire FE_OCP_RBN4059_n_44875;
wire FE_OCP_RBN4060_n_44875;
wire FE_OCP_RBN4061_n_44030;
wire FE_OCP_RBN4062_n_44030;
wire FE_OCP_RBN4063_n_7558;
wire FE_OCP_RBN4064_n_7558;
wire FE_OCP_RBN4065_n_7558;
wire FE_OCP_RBN4066_n_7558;
wire FE_OCP_RBN4067_n_18829;
wire FE_OCP_RBN4068_n_18829;
wire FE_OCP_RBN4070_n_29292;
wire FE_OCP_RBN4071_n_2289;
wire FE_OCP_RBN4072_n_2289;
wire FE_OCP_RBN4073_n_2289;
wire FE_OCP_RBN4074_n_2289;
wire FE_OCP_RBN4075_n_7708;
wire FE_OCP_RBN4080_n_7708;
wire FE_OCP_RBN4081_n_18899;
wire FE_OCP_RBN4082_n_18899;
wire FE_OCP_RBN4083_n_13453;
wire FE_OCP_RBN4084_n_13453;
wire FE_OCP_RBN4087_n_12880;
wire FE_OCP_RBN4088_n_12880;
wire FE_OCP_RBN4089_n_12880;
wire FE_OCP_RBN4090_n_12880;
wire FE_OCP_RBN4091_n_12880;
wire FE_OCP_RBN4092_n_12880;
wire FE_OCP_RBN4093_n_12880;
wire FE_OCP_RBN4094_n_12880;
wire FE_OCP_RBN4095_n_12880;
wire FE_OCP_RBN4096_n_12880;
wire FE_OCP_RBN4097_n_12880;
wire FE_OCP_RBN4098_n_12880;
wire FE_OCP_RBN4099_n_12880;
wire FE_OCP_RBN4100_n_12880;
wire FE_OCP_RBN4101_n_12880;
wire FE_OCP_RBN4102_n_12880;
wire FE_OCP_RBN4103_n_12880;
wire FE_OCP_RBN4104_n_12880;
wire FE_OCP_RBN4105_n_12880;
wire FE_OCP_RBN4106_n_12880;
wire FE_OCP_RBN4107_n_12880;
wire FE_OCP_RBN4108_n_12880;
wire FE_OCP_RBN4109_n_12880;
wire FE_OCP_RBN4110_n_12880;
wire FE_OCP_RBN4111_n_12880;
wire FE_OCP_RBN4112_n_12880;
wire FE_OCP_RBN4113_n_33533;
wire FE_OCP_RBN4114_n_33533;
wire FE_OCP_RBN4115_n_41381;
wire FE_OCP_RBN4118_n_45487;
wire FE_OCP_RBN4120_n_13483;
wire FE_OCP_RBN4130_n_24077;
wire FE_OCP_RBN4131_n_24077;
wire FE_OCP_RBN4132_n_38028;
wire FE_OCP_RBN4133_n_38028;
wire FE_OCP_RBN4135_n_7743;
wire FE_OCP_RBN4136_n_7743;
wire FE_OCP_RBN4137_n_7743;
wire FE_OCP_RBN4138_n_7743;
wire FE_OCP_RBN4139_n_7743;
wire FE_OCP_RBN4140_n_7743;
wire FE_OCP_RBN4141_n_7743;
wire FE_OCP_RBN4142_n_7743;
wire FE_OCP_RBN4143_n_7743;
wire FE_OCP_RBN4144_n_7743;
wire FE_OCP_RBN4145_n_7743;
wire FE_OCP_RBN4146_n_7743;
wire FE_OCP_RBN4147_n_3217;
wire FE_OCP_RBN4148_n_24173;
wire FE_OCP_RBN4149_n_24173;
wire FE_OCP_RBN4150_n_13616;
wire FE_OCP_RBN4151_n_13616;
wire FE_OCP_RBN4152_n_13616;
wire FE_OCP_RBN4153_n_29378;
wire FE_OCP_RBN4154_n_29378;
wire FE_OCP_RBN4156_n_29378;
wire FE_OCP_RBN4157_n_24222;
wire FE_OCP_RBN4158_n_24222;
wire FE_OCP_RBN4159_FE_OCPN857_n_7802;
wire FE_OCP_RBN4160_FE_OCPN857_n_7802;
wire FE_OCP_RBN4161_FE_OCPN857_n_7802;
wire FE_OCP_RBN4162_FE_OCPN857_n_7802;
wire FE_OCP_RBN4163_n_3390;
wire FE_OCP_RBN4164_n_3390;
wire FE_OCP_RBN4165_n_3494;
wire FE_OCP_RBN4166_n_3494;
wire FE_OCP_RBN4167_n_3494;
wire FE_OCP_RBN4168_n_29553;
wire FE_OCP_RBN4169_n_29553;
wire FE_OCP_RBN4170_n_19390;
wire FE_OCP_RBN4171_n_19390;
wire FE_OCP_RBN4172_n_38545;
wire FE_OCP_RBN4173_n_38545;
wire FE_OCP_RBN4174_FE_OCPN1913_n_2669;
wire FE_OCP_RBN4175_n_3626;
wire FE_OCP_RBN4176_n_3626;
wire FE_OCP_RBN4177_n_38586;
wire FE_OCP_RBN4178_n_38586;
wire FE_OCP_RBN4179_n_38592;
wire FE_OCP_RBN4180_n_38592;
wire FE_OCP_RBN4181_n_19599;
wire FE_OCP_RBN4182_n_19599;
wire FE_OCP_RBN4184_n_24467;
wire FE_OCP_RBN4185_n_8288;
wire FE_OCP_RBN4186_n_8288;
wire FE_OCP_RBN4187_n_8621;
wire FE_OCP_RBN4188_n_13765;
wire FE_OCP_RBN4189_n_13765;
wire FE_OCP_RBN4190_n_14279;
wire FE_OCP_RBN4191_n_34285;
wire FE_OCP_RBN4192_n_38537;
wire FE_OCP_RBN4193_n_38537;
wire FE_OCP_RBN4194_n_38683;
wire FE_OCP_RBN4195_n_38683;
wire FE_OCP_RBN4198_n_13796;
wire FE_OCP_RBN4199_n_13796;
wire FE_OCP_RBN4200_n_13796;
wire FE_OCP_RBN4201_n_13796;
wire FE_OCP_RBN4202_n_13796;
wire FE_OCP_RBN4203_n_13796;
wire FE_OCP_RBN4204_n_13796;
wire FE_OCP_RBN4205_n_13796;
wire FE_OCP_RBN4206_n_13796;
wire FE_OCP_RBN4208_n_13796;
wire FE_OCP_RBN4209_n_13796;
wire FE_OCP_RBN4210_n_13796;
wire FE_OCP_RBN4211_n_8767;
wire FE_OCP_RBN4212_n_3343;
wire FE_OCP_RBN4213_n_3386;
wire FE_OCP_RBN4214_FE_OCPN3565_n_10214;
wire FE_OCP_RBN4215_FE_OCPN3565_n_10214;
wire FE_OCP_RBN4216_FE_OCPN3565_n_10214;
wire FE_OCP_RBN4217_n_8597;
wire FE_OCP_RBN4218_n_8597;
wire FE_OCP_RBN4219_n_8594;
wire FE_OCP_RBN4220_n_8594;
wire FE_OCP_RBN4221_n_8732;
wire FE_OCP_RBN4222_n_8732;
wire FE_OCP_RBN4223_n_8784;
wire FE_OCP_RBN4224_n_8799;
wire FE_OCP_RBN4226_n_13962;
wire FE_OCP_RBN4228_n_13962;
wire FE_OCP_RBN4229_n_13962;
wire FE_OCP_RBN4231_n_13962;
wire FE_OCP_RBN4232_n_13962;
wire FE_OCP_RBN4234_n_13962;
wire FE_OCP_RBN4235_n_9089;
wire FE_OCP_RBN4236_n_9089;
wire FE_OCP_RBN4237_n_8781;
wire FE_OCP_RBN4238_n_8781;
wire FE_OCP_RBN4239_n_44594;
wire FE_OCP_RBN4240_n_44594;
wire FE_OCP_RBN4241_n_44594;
wire FE_OCP_RBN4242_n_44594;
wire FE_OCP_RBN4243_n_44594;
wire FE_OCP_RBN4244_n_44594;
wire FE_OCP_RBN4246_n_8904;
wire FE_OCP_RBN4247_n_8904;
wire FE_OCP_RBN4248_n_14573;
wire FE_OCP_RBN4249_n_14697;
wire FE_OCP_RBN4251_n_8687;
wire FE_OCP_RBN4252_n_8687;
wire FE_OCP_RBN4253_n_8687;
wire FE_OCP_RBN4254_n_3705;
wire FE_OCP_RBN4255_n_3705;
wire FE_OCP_RBN4256_n_3705;
wire FE_OCP_RBN4258_n_34921;
wire FE_OCP_RBN4259_n_34921;
wire FE_OCP_RBN4260_n_34921;
wire FE_OCP_RBN4261_n_34878;
wire FE_OCP_RBN4262_n_9009;
wire FE_OCP_RBN4263_n_9009;
wire FE_OCP_RBN4266_FE_RN_998_0;
wire FE_OCP_RBN4269_n_8872;
wire FE_OCP_RBN4270_n_8872;
wire FE_OCP_RBN4274_n_3700;
wire FE_OCP_RBN4280_n_3848;
wire FE_OCP_RBN4281_n_3848;
wire FE_OCP_RBN4282_n_9243;
wire FE_OCP_RBN4283_n_9243;
wire FE_OCP_RBN4288_n_44563;
wire FE_OCP_RBN4289_n_47014;
wire FE_OCP_RBN4290_n_47014;
wire FE_OCP_RBN4291_n_3909;
wire FE_OCP_RBN4292_n_4080;
wire FE_OCP_RBN4293_n_4080;
wire FE_OCP_RBN4294_n_4080;
wire FE_OCP_RBN4295_n_4080;
wire FE_OCP_RBN4296_n_4080;
wire FE_OCP_RBN4298_n_25238;
wire FE_OCP_RBN4302_n_44579;
wire FE_OCP_RBN4303_n_44579;
wire FE_OCP_RBN4304_n_44579;
wire FE_OCP_RBN4305_n_44579;
wire FE_OCP_RBN4307_n_25178;
wire FE_OCP_RBN4309_n_25178;
wire FE_OCP_RBN4311_n_25178;
wire FE_OCP_RBN4314_n_9396;
wire FE_OCP_RBN4315_n_14881;
wire FE_OCP_RBN4316_n_9292;
wire FE_OCP_RBN4317_n_9292;
wire FE_OCP_RBN4319_n_14768;
wire FE_OCP_RBN4322_n_15156;
wire FE_OCP_RBN4323_n_15156;
wire FE_OCP_RBN4324_n_15156;
wire FE_OCP_RBN4325_n_20333;
wire FE_OCP_RBN4326_n_20333;
wire FE_OCP_RBN4327_n_38878;
wire FE_OCP_RBN4328_n_38878;
wire FE_OCP_RBN4329_n_38878;
wire FE_OCP_RBN4330_n_9102;
wire FE_OCP_RBN4334_n_20242;
wire FE_OCP_RBN4335_n_20242;
wire FE_OCP_RBN4337_n_20242;
wire FE_OCP_RBN4338_n_9521;
wire FE_OCP_RBN4339_n_4403;
wire FE_OCP_RBN4340_n_4403;
wire FE_OCP_RBN4341_n_25500;
wire FE_OCP_RBN4342_n_4198;
wire FE_OCP_RBN4343_n_15071;
wire FE_OCP_RBN4344_n_35177;
wire FE_OCP_RBN4345_n_4378;
wire FE_OCP_RBN4347_n_10017;
wire FE_OCP_RBN4348_n_20568;
wire FE_OCP_RBN4349_n_9975;
wire FE_OCP_RBN4350_n_9975;
wire FE_OCP_RBN4351_n_20456;
wire FE_OCP_RBN4352_FE_OCPN1263_n_20971;
wire FE_OCP_RBN4353_FE_OCPN1263_n_20971;
wire FE_OCP_RBN4354_n_4585;
wire FE_OCP_RBN4355_n_10100;
wire FE_OCP_RBN4356_n_10100;
wire FE_OCP_RBN4357_n_10100;
wire FE_OCP_RBN4358_n_10100;
wire FE_OCP_RBN4359_n_10100;
wire FE_OCP_RBN4360_n_20632;
wire FE_OCP_RBN4361_FE_RN_1500_0;
wire FE_OCP_RBN4362_FE_RN_1500_0;
wire FE_OCP_RBN4363_n_39584;
wire FE_OCP_RBN4364_n_20710;
wire FE_OCP_RBN4365_n_4692;
wire FE_OCP_RBN4366_n_4692;
wire FE_OCP_RBN4367_n_25889;
wire FE_OCP_RBN4368_n_25889;
wire FE_OCP_RBN4369_n_46982;
wire FE_OCP_RBN4370_n_46982;
wire FE_OCP_RBN4371_n_5032;
wire FE_OCP_RBN4372_n_5048;
wire FE_OCP_RBN4373_n_5048;
wire FE_OCP_RBN4374_n_5048;
wire FE_OCP_RBN4375_n_15514;
wire FE_OCP_RBN4377_n_15700;
wire FE_OCP_RBN4378_n_4956;
wire FE_OCP_RBN4379_n_4956;
wire FE_OCP_RBN4380_n_5028;
wire FE_OCP_RBN4381_n_5041;
wire FE_OCP_RBN4382_n_39523;
wire FE_OCP_RBN4384_n_5221;
wire FE_OCP_RBN4385_n_10570;
wire FE_OCP_RBN4387_n_5013;
wire FE_OCP_RBN4388_n_26173;
wire FE_OCP_RBN4389_n_26173;
wire FE_OCP_RBN4390_n_26173;
wire FE_OCP_RBN4391_n_16230;
wire FE_OCP_RBN4392_n_26146;
wire FE_OCP_RBN4393_n_10682;
wire FE_OCP_RBN4394_n_16146;
wire FE_OCP_RBN4395_n_16146;
wire FE_OCP_RBN4396_n_16146;
wire FE_OCP_RBN4398_n_39629;
wire FE_OCP_RBN4399_n_5308;
wire FE_OCP_RBN4400_n_5532;
wire FE_OCP_RBN4401_n_16321;
wire FE_OCP_RBN4402_n_43013;
wire FE_OCP_RBN4405_n_26160;
wire FE_OCP_RBN4408_n_26394;
wire FE_OCP_RBN4409_n_16429;
wire FE_OCP_RBN4412_n_26661;
wire FE_OCP_RBN4413_n_31117;
wire FE_OCP_RBN4414_n_31117;
wire FE_OCP_RBN4415_n_31117;
wire FE_OCP_RBN4416_n_31117;
wire FE_OCP_RBN4417_n_31117;
wire FE_OCP_RBN4418_n_31117;
wire FE_OCP_RBN4419_n_31117;
wire FE_OCP_RBN4420_n_31117;
wire FE_OCP_RBN4421_n_31117;
wire FE_OCP_RBN4422_n_31117;
wire FE_OCP_RBN4423_n_31117;
wire FE_OCP_RBN4424_n_31117;
wire FE_OCP_RBN4425_n_31117;
wire FE_OCP_RBN4429_n_39942;
wire FE_OCP_RBN4430_n_39942;
wire FE_OCP_RBN4431_n_39942;
wire FE_OCP_RBN4432_n_26160;
wire FE_OCP_RBN4433_n_26160;
wire FE_OCP_RBN4434_n_26160;
wire FE_OCP_RBN4435_n_26160;
wire FE_OCP_RBN4436_n_26160;
wire FE_OCP_RBN4437_n_26160;
wire FE_OCP_RBN4438_n_26160;
wire FE_OCP_RBN4439_n_26160;
wire FE_OCP_RBN4440_n_5891;
wire FE_OCP_RBN4441_n_5891;
wire FE_OCP_RBN4443_n_46424;
wire FE_OCP_RBN4444_n_5849;
wire FE_OCP_RBN4445_n_43022;
wire FE_OCP_RBN4446_n_43022;
wire FE_OCP_RBN4447_FE_OFN760_n_46337;
wire FE_OCP_RBN4448_FE_OFN760_n_46337;
wire FE_OCP_RBN4451_n_5870;
wire FE_OCP_RBN4454_n_6102;
wire FE_OCP_RBN4455_n_6102;
wire FE_OCP_RBN4456_n_43103;
wire FE_OCP_RBN4457_n_43103;
wire FE_OCP_RBN4458_FE_RN_1190_0;
wire FE_OCP_RBN4459_FE_RN_1190_0;
wire FE_OCP_RBN4462_n_44267;
wire FE_OCP_RBN4464_n_44267;
wire FE_OCP_RBN4466_n_44267;
wire FE_OCP_RBN4467_n_44267;
wire FE_OCP_RBN4468_n_44267;
wire FE_OCP_RBN4471_n_31819;
wire FE_OCP_RBN4472_n_31819;
wire FE_OCP_RBN4476_FE_OCPN913_n_43230;
wire FE_OCP_RBN4477_FE_OCPN913_n_43230;
wire FE_OCP_RBN4478_FE_OCPN913_n_43230;
wire FE_OCP_RBN4479_FE_OCPN913_n_43230;
wire FE_OCP_RBN4480_n_11439;
wire FE_OCP_RBN4481_n_11439;
wire FE_OCP_RBN4482_n_11439;
wire FE_OCP_RBN4483_n_11439;
wire FE_OCP_RBN4484_n_22667;
wire FE_OCP_RBN4485_n_22667;
wire FE_OCP_RBN4486_n_27145;
wire FE_OCP_RBN4487_n_22438;
wire FE_OCP_RBN4488_n_6299;
wire FE_OCP_RBN4489_n_6299;
wire FE_OCP_RBN4490_n_32152;
wire FE_OCP_RBN4492_n_22755;
wire FE_OCP_RBN4494_n_27555;
wire FE_OCP_RBN4495_n_27639;
wire FE_OCP_RBN4496_n_27639;
wire FE_OCP_RBN4590_n_44847;
wire FE_OCP_RBN4593_delay_xor_ln22_unr12_stage5_stallmux_q_1_;
wire FE_OCP_RBN4630_n_44962;
wire FE_OCP_RBN4633_n_44962;
wire FE_OCP_RBN4635_n_33589;
wire FE_OCP_RBN4636_n_18600;
wire FE_OCP_RBN4637_n_18600;
wire FE_OCP_RBN4639_n_18681;
wire FE_OCP_RBN4643_n_35121;
wire FE_OCP_RBN4644_n_20420;
wire FE_OCP_RBN4645_n_20420;
wire FE_OCP_RBN4646_n_22553;
wire FE_OCP_RBN4647_n_22553;
wire FE_OCP_RBN4648_n_22625;
wire FE_OCP_RBN4649_n_22625;
wire FE_OCP_RBN4870_n_35145;
wire FE_OCP_RBN4900_n_29056;
wire FE_OCP_RBN4902_n_44256;
wire FE_OCP_RBN4903_n_44256;
wire FE_OCP_RBN4904_n_44256;
wire FE_OCP_RBN4905_n_44256;
wire FE_OCP_RBN4906_n_44256;
wire FE_OCP_RBN4908_n_44222;
wire FE_OCP_RBN4909_n_44222;
wire FE_OCP_RBN4910_n_44222;
wire FE_OCP_RBN4912_n_33803;
wire FE_OCP_RBN4913_n_33833;
wire FE_OCP_RBN4914_n_33833;
wire FE_OCP_RBN4915_n_33503;
wire FE_OCP_RBN4916_n_33503;
wire FE_OCP_RBN4917_n_33491;
wire FE_OCP_RBN4918_n_33491;
wire FE_OCP_RBN4919_n_32575;
wire FE_OCP_RBN4920_n_33691;
wire FE_OCP_RBN4921_n_33691;
wire FE_OCP_RBN4923_n_34980;
wire FE_OCP_RBN4924_n_34980;
wire FE_OCP_RBN4925_n_34980;
wire FE_OCP_RBN5016_n_12026;
wire FE_OCP_RBN5017_n_12026;
wire FE_OCP_RBN5018_n_16972;
wire FE_OCP_RBN5019_n_13726;
wire FE_OCP_RBN5021_n_13726;
wire FE_OCP_RBN5022_n_29080;
wire FE_OCP_RBN5023_n_29080;
wire FE_OCP_RBN5024_n_29080;
wire FE_OCP_RBN5025_n_29053;
wire FE_OCP_RBN5026_n_29053;
wire FE_OCP_RBN5027_n_18515;
wire FE_OCP_RBN5028_n_18515;
wire FE_OCP_RBN5029_n_18678;
wire FE_OCP_RBN5030_n_18678;
wire FE_OCP_RBN5031_n_18951;
wire FE_OCP_RBN5032_n_18951;
wire FE_OCP_RBN5033_n_18951;
wire FE_OCP_RBN5034_n_19062;
wire FE_OCP_RBN5035_n_19055;
wire FE_OCP_RBN5037_n_13927;
wire FE_OCP_RBN5038_n_13927;
wire FE_OCP_RBN5039_n_13927;
wire FE_OCP_RBN5040_n_27827;
wire FE_OCP_RBN5041_n_14201;
wire FE_OCP_RBN5045_n_14450;
wire FE_OCP_RBN5046_n_14450;
wire FE_OCP_RBN5047_n_29648;
wire FE_OCP_RBN5049_FE_RN_606_0;
wire FE_OCP_RBN5050_FE_RN_606_0;
wire FE_OCP_RBN5051_n_22709;
wire FE_OCP_RBN5053_n_32169;
wire FE_OCP_RBN5055_n_32340;
wire FE_OCP_RBN5058_n_32427;
wire FE_OCP_RBN5175_n_44061;
wire FE_OCP_RBN5179_n_44061;
wire FE_OCP_RBN5180_n_44061;
wire FE_OCP_RBN5181_n_44061;
wire FE_OCP_RBN5196_n_25893;
wire FE_OCP_RBN5197_n_25893;
wire FE_OCP_RBN5198_n_25893;
wire FE_OCP_RBN5199_n_25893;
wire FE_OCP_RBN5200_n_25729;
wire FE_OCP_RBN5201_n_25729;
wire FE_OCP_RBN5202_n_25729;
wire FE_OCP_RBN5203_n_25729;
wire FE_OCP_RBN5204_n_25729;
wire FE_OCP_RBN5205_n_20504;
wire FE_OCP_RBN5206_n_20504;
wire FE_OCP_RBN5207_n_20504;
wire FE_OCP_RBN5208_n_20412;
wire FE_OCP_RBN5209_n_20412;
wire FE_OCP_RBN5210_n_20412;
wire FE_OCP_RBN5211_n_20412;
wire FE_OCP_RBN5212_n_21987;
wire FE_OCP_RBN5213_n_29773;
wire FE_OCP_RBN5214_n_22150;
wire FE_OCP_RBN5215_n_22150;
wire FE_OCP_RBN5216_n_22212;
wire FE_OCP_RBN5217_n_22212;
wire FE_OCP_RBN5218_n_32279;
wire FE_OCP_RBN5322_n_16745;
wire FE_OCP_RBN5323_n_27893;
wire FE_OCP_RBN5324_n_27885;
wire FE_OCP_RBN5325_n_18653;
wire FE_OCP_RBN5326_n_29292;
wire FE_OCP_RBN5327_FE_RN_2034_0;
wire FE_OCP_RBN5328_n_15047;
wire FE_OCP_RBN5329_n_15047;
wire FE_OCP_RBN5330_n_20678;
wire FE_OCP_RBN5331_n_20843;
wire FE_OCP_RBN5333_FE_RN_1490_0;
wire FE_OCP_RBN5334_FE_RN_1490_0;
wire FE_OCP_RBN5335_FE_RN_1144_0;
wire FE_OCP_RBN5336_n_30865;
wire FE_OCP_RBN5337_FE_RN_2064_0;
wire FE_OCP_RBN5338_FE_RN_2064_0;
wire FE_OCP_RBN5340_n_21261;
wire FE_OCP_RBN5341_n_22068;
wire FE_OCP_RBN5342_n_22068;
wire FE_OCP_RBN5343_n_22068;
wire FE_OCP_RBN5344_n_22476;
wire FE_OCP_RBN5345_n_22476;
wire FE_OCP_RBN5346_n_22556;
wire FE_OCP_RBN5347_n_22556;
wire FE_OCP_RBN5348_FE_RN_627_0;
wire FE_OCP_RBN5349_n_32518;
wire FE_OCP_RBN5350_n_22818;
wire FE_OCP_RBN5351_n_22903;
wire FE_OCP_RBN5352_n_32516;
wire FE_OCP_RBN5374_n_28186;
wire FE_OCP_RBN5375_n_28123;
wire FE_OCP_RBN5376_n_28123;
wire FE_OCP_RBN5377_n_19055;
wire FE_OCP_RBN5378_n_19055;
wire FE_OCP_RBN5379_n_19055;
wire FE_OCP_RBN5380_n_19428;
wire FE_OCP_RBN5381_n_20123;
wire FE_OCP_RBN5382_n_20123;
wire FE_OCP_RBN5386_n_20638;
wire FE_OCP_RBN5387_n_22149;
wire FE_OCP_RBN5388_n_22149;
wire FE_OCP_RBN5391_cordic_combinational_sub_ln23_0_unr12_z_0_;
wire FE_OCP_RBN5392_cordic_combinational_sub_ln23_0_unr12_z_0_;
wire FE_OCP_RBN5393_cordic_combinational_sub_ln23_0_unr12_z_0_;
wire FE_OCP_RBN5394_cordic_combinational_sub_ln23_0_unr12_z_0_;
wire FE_OCP_RBN5395_cordic_combinational_sub_ln23_0_unr12_z_0_;
wire FE_OCP_RBN5412_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN5434_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN5435_delay_xor_ln22_unr6_stage3_stallmux_q_0_;
wire FE_OCP_RBN5436_delay_xor_ln22_unr6_stage3_stallmux_q_0_;
wire FE_OCP_RBN5437_delay_xor_ln22_unr6_stage3_stallmux_q_0_;
wire FE_OCP_RBN5438_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_;
wire FE_OCP_RBN5439_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_;
wire FE_OCP_RBN5441_delay_sub_ln23_0_unr8_stage4_stallmux_q_2_;
wire FE_OCP_RBN5442_delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire FE_OCP_RBN5445_delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire FE_OCP_RBN5459_n_44061;
wire FE_OCP_RBN5465_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN5466_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN5467_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire FE_OCP_RBN5498_n_44610;
wire FE_OCP_RBN5503_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN5504_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN5506_n_44061;
wire FE_OCP_RBN5507_n_44061;
wire FE_OCP_RBN5508_FE_RN_1997_0;
wire FE_OCP_RBN5509_FE_RN_1997_0;
wire FE_OCP_RBN5510_FE_RN_1997_0;
wire FE_OCP_RBN5511_n_44365;
wire FE_OCP_RBN5512_n_44365;
wire FE_OCP_RBN5513_n_44365;
wire FE_OCP_RBN5514_n_44365;
wire FE_OCP_RBN5515_n_1472;
wire FE_OCP_RBN5516_n_32436;
wire FE_OCP_RBN5517_n_32436;
wire FE_OCP_RBN5518_n_32436;
wire FE_OCP_RBN5522_n_23078;
wire FE_OCP_RBN5523_n_28058;
wire FE_OCP_RBN5524_n_32752;
wire FE_OCP_RBN5525_n_36921;
wire FE_OCP_RBN5527_n_6760;
wire FE_OCP_RBN5528_n_44061;
wire FE_OCP_RBN5529_n_44061;
wire FE_OCP_RBN5530_n_1541;
wire FE_OCP_RBN5531_n_27941;
wire FE_OCP_RBN5532_n_44083;
wire FE_OCP_RBN5533_n_44083;
wire FE_OCP_RBN5534_n_44083;
wire FE_OCP_RBN5535_n_44083;
wire FE_OCP_RBN5536_n_44083;
wire FE_OCP_RBN5537_n_44083;
wire FE_OCP_RBN5539_n_23307;
wire FE_OCP_RBN5540_n_23307;
wire FE_OCP_RBN5541_n_23044;
wire FE_OCP_RBN5542_n_23044;
wire FE_OCP_RBN5543_n_23044;
wire FE_OCP_RBN5544_n_45145;
wire FE_OCP_RBN5545_n_45145;
wire FE_OCP_RBN5546_n_45145;
wire FE_OCP_RBN5547_n_1733;
wire FE_OCP_RBN5548_FE_OCPN4833_n_32863;
wire FE_OCP_RBN5549_n_28319;
wire FE_OCP_RBN5550_n_17914;
wire FE_OCP_RBN5551_n_17914;
wire FE_OCP_RBN5552_n_23328;
wire FE_OCP_RBN5553_n_1812;
wire FE_OCP_RBN5554_n_1822;
wire FE_OCP_RBN5555_n_1827;
wire FE_OCP_RBN5556_n_37559;
wire FE_OCP_RBN5557_n_37559;
wire FE_OCP_RBN5558_n_37559;
wire FE_OCP_RBN5559_n_1853;
wire FE_OCP_RBN5560_n_1889;
wire FE_OCP_RBN5561_n_33097;
wire FE_OCP_RBN5562_n_33097;
wire FE_OCP_RBN5563_n_37551;
wire FE_OCP_RBN5564_n_37551;
wire FE_OCP_RBN5565_n_2346;
wire FE_OCP_RBN5566_n_2346;
wire FE_OCP_RBN5567_n_2346;
wire FE_OCP_RBN5568_n_2103;
wire FE_OCP_RBN5569_n_2103;
wire FE_OCP_RBN5574_n_12727;
wire FE_OCP_RBN5575_n_12727;
wire FE_OCP_RBN5576_n_12727;
wire FE_OCP_RBN5578_n_12753;
wire FE_OCP_RBN5580_n_12753;
wire FE_OCP_RBN5581_n_12753;
wire FE_OCP_RBN5582_n_12802;
wire FE_OCP_RBN5583_n_12802;
wire FE_OCP_RBN5584_n_12802;
wire FE_OCP_RBN5585_n_33368;
wire FE_OCP_RBN5587_FE_RN_1367_0;
wire FE_OCP_RBN5588_FE_RN_1367_0;
wire FE_OCP_RBN5589_FE_RN_1367_0;
wire FE_OCP_RBN5590_FE_RN_1367_0;
wire FE_OCP_RBN5591_FE_RN_1367_0;
wire FE_OCP_RBN5592_FE_RN_1367_0;
wire FE_OCP_RBN5593_FE_RN_1367_0;
wire FE_OCP_RBN5594_n_45903;
wire FE_OCP_RBN5595_n_45903;
wire FE_OCP_RBN5596_n_45903;
wire FE_OCP_RBN5597_n_45903;
wire FE_OCP_RBN5598_n_2100;
wire FE_OCP_RBN5599_n_2100;
wire FE_OCP_RBN5600_n_44875;
wire FE_OCP_RBN5603_n_29056;
wire FE_OCP_RBN5604_n_29056;
wire FE_OCP_RBN5605_n_2430;
wire FE_OCP_RBN5606_n_7730;
wire FE_OCP_RBN5607_n_7730;
wire FE_OCP_RBN5608_n_7730;
wire FE_OCP_RBN5609_n_7730;
wire FE_OCP_RBN5610_n_7730;
wire FE_OCP_RBN5611_n_7730;
wire FE_OCP_RBN5612_n_7730;
wire FE_OCP_RBN5613_n_7730;
wire FE_OCP_RBN5614_n_7730;
wire FE_OCP_RBN5615_n_24070;
wire FE_OCP_RBN5617_n_18899;
wire FE_OCP_RBN5618_n_18899;
wire FE_OCP_RBN5620_n_18986;
wire FE_OCP_RBN5621_n_18986;
wire FE_OCP_RBN5622_n_18986;
wire FE_OCP_RBN5625_n_2457;
wire FE_OCP_RBN5626_n_2457;
wire FE_OCP_RBN5627_n_33976;
wire FE_OCP_RBN5628_n_33976;
wire FE_OCP_RBN5629_n_33976;
wire FE_OCP_RBN5630_n_33957;
wire FE_OCP_RBN5632_n_7708;
wire FE_OCP_RBN5633_n_7708;
wire FE_OCP_RBN5634_n_7708;
wire FE_OCP_RBN5635_n_7708;
wire FE_OCP_RBN5636_n_7708;
wire FE_OCP_RBN5637_n_41381;
wire FE_OCP_RBN5638_n_41381;
wire FE_OCP_RBN5639_n_41381;
wire FE_OCP_RBN5640_n_19060;
wire FE_OCP_RBN5643_n_33977;
wire FE_OCP_RBN5644_n_2674;
wire FE_OCP_RBN5645_n_29236;
wire FE_OCP_RBN5646_n_33785;
wire FE_OCP_RBN5647_FE_OCPN855_n_7721;
wire FE_OCP_RBN5648_n_2438;
wire FE_OCP_RBN5649_n_2438;
wire FE_OCP_RBN5650_n_2438;
wire FE_OCP_RBN5651_n_2438;
wire FE_OCP_RBN5652_n_2438;
wire FE_OCP_RBN5653_n_2438;
wire FE_OCP_RBN5654_n_2438;
wire FE_OCP_RBN5655_n_2438;
wire FE_OCP_RBN5656_n_2438;
wire FE_OCP_RBN5657_n_2438;
wire FE_OCP_RBN5658_n_2438;
wire FE_OCP_RBN5659_n_2438;
wire FE_OCP_RBN5660_n_2438;
wire FE_OCP_RBN5661_n_2438;
wire FE_OCP_RBN5662_n_2438;
wire FE_OCP_RBN5663_n_2438;
wire FE_OCP_RBN5664_n_13757;
wire FE_OCP_RBN5665_n_19101;
wire FE_OCP_RBN5666_n_19101;
wire FE_OCP_RBN5667_n_19101;
wire FE_OCP_RBN5668_n_19101;
wire FE_OCP_RBN5669_n_19101;
wire FE_OCP_RBN5670_n_24288;
wire FE_OCP_RBN5671_n_24288;
wire FE_OCP_RBN5672_n_29425;
wire FE_OCP_RBN5673_n_41420;
wire FE_OCP_RBN5674_n_41420;
wire FE_OCP_RBN5675_n_41420;
wire FE_OCP_RBN5676_n_41420;
wire FE_OCP_RBN5677_n_19177;
wire FE_OCP_RBN5678_n_19177;
wire FE_OCP_RBN5679_n_19177;
wire FE_OCP_RBN5680_n_19177;
wire FE_OCP_RBN5681_n_19177;
wire FE_OCP_RBN5682_n_19177;
wire FE_OCP_RBN5683_n_38474;
wire FE_OCP_RBN5684_FE_RN_308_0;
wire FE_OCP_RBN5685_FE_RN_308_0;
wire FE_OCP_RBN5686_FE_RN_308_0;
wire FE_OCP_RBN5687_n_24259;
wire FE_OCP_RBN5688_n_24259;
wire FE_OCP_RBN5689_n_38531;
wire FE_OCP_RBN5690_n_38515;
wire FE_OCP_RBN5691_n_2884;
wire FE_OCP_RBN5692_n_2884;
wire FE_OCP_RBN5693_n_8138;
wire FE_OCP_RBN5695_n_8342;
wire FE_OCP_RBN5697_n_8342;
wire FE_OCP_RBN5698_n_38577;
wire FE_OCP_RBN5699_n_42038;
wire FE_OCP_RBN5700_n_45828;
wire FE_OCP_RBN5701_n_13954;
wire FE_OCP_RBN5702_n_29568;
wire FE_OCP_RBN5703_n_19663;
wire FE_OCP_RBN5704_n_19663;
wire FE_OCP_RBN5705_n_19663;
wire FE_OCP_RBN5706_n_24451;
wire FE_OCP_RBN5707_n_24451;
wire FE_OCP_RBN5708_n_3055;
wire FE_OCP_RBN5709_n_3055;
wire FE_OCP_RBN5710_n_13984;
wire FE_OCP_RBN5711_n_13984;
wire FE_OCP_RBN5712_n_44102;
wire FE_OCP_RBN5713_n_44102;
wire FE_OCP_RBN5714_n_44102;
wire FE_OCP_RBN5715_n_44102;
wire FE_OCP_RBN5716_n_8523;
wire FE_OCP_RBN5717_n_24718;
wire FE_OCP_RBN5718_n_24718;
wire FE_OCP_RBN5719_n_29624;
wire FE_OCP_RBN5720_n_29624;
wire FE_OCP_RBN5721_n_24506;
wire FE_OCP_RBN5722_n_24506;
wire FE_OCP_RBN5723_n_47022;
wire FE_OCP_RBN5724_n_47022;
wire FE_OCP_RBN5725_n_14120;
wire FE_OCP_RBN5726_n_14120;
wire FE_OCP_RBN5727_n_14120;
wire FE_OCP_RBN5728_n_14120;
wire FE_OCP_RBN5729_n_4211;
wire FE_OCP_RBN5730_n_4211;
wire FE_OCP_RBN5731_n_4211;
wire FE_OCP_RBN5732_n_19806;
wire FE_OCP_RBN5733_n_19806;
wire FE_OCP_RBN5734_n_8548;
wire FE_OCP_RBN5735_n_38569;
wire FE_OCP_RBN5736_n_38569;
wire FE_OCP_RBN5737_n_8402;
wire FE_OCP_RBN5738_n_8402;
wire FE_OCP_RBN5739_n_8402;
wire FE_OCP_RBN5740_n_4336;
wire FE_OCP_RBN5741_n_4336;
wire FE_OCP_RBN5742_n_8540;
wire FE_OCP_RBN5743_n_34278;
wire FE_OCP_RBN5744_n_42043;
wire FE_OCP_RBN5745_n_24618;
wire FE_OCP_RBN5746_n_8637;
wire FE_OCP_RBN5747_n_8637;
wire FE_OCP_RBN5748_n_8637;
wire FE_OCP_RBN5749_n_8599;
wire FE_OCP_RBN5750_n_8599;
wire FE_OCP_RBN5751_n_4022;
wire FE_OCP_RBN5752_n_4022;
wire FE_OCP_RBN5753_n_4022;
wire FE_OCP_RBN5754_n_4022;
wire FE_OCP_RBN5756_n_34307;
wire FE_OCP_RBN5757_n_14444;
wire FE_OCP_RBN5758_n_14444;
wire FE_OCP_RBN5759_n_14444;
wire FE_OCP_RBN5760_n_14444;
wire FE_OCP_RBN5762_n_19884;
wire FE_OCP_RBN5763_n_19884;
wire FE_OCP_RBN5764_n_19884;
wire FE_OCP_RBN5767_n_3498;
wire FE_OCP_RBN5768_n_3498;
wire FE_OCP_RBN5769_n_3338;
wire FE_OCP_RBN5770_n_3338;
wire FE_OCP_RBN5771_n_3338;
wire FE_OCP_RBN5772_n_34375;
wire FE_OCP_RBN5773_n_34375;
wire FE_OCP_RBN5774_n_13796;
wire FE_OCP_RBN5776_n_13796;
wire FE_OCP_RBN5777_n_13796;
wire FE_OCP_RBN5779_n_44570;
wire FE_OCP_RBN5780_n_44570;
wire FE_OCP_RBN5781_n_44570;
wire FE_OCP_RBN5784_n_8657;
wire FE_OCP_RBN5785_n_30071;
wire FE_OCP_RBN5786_n_3421;
wire FE_OCP_RBN5787_n_3421;
wire FE_OCP_RBN5790_n_13962;
wire FE_OCP_RBN5791_n_13962;
wire FE_OCP_RBN5792_n_13962;
wire FE_OCP_RBN5793_n_13962;
wire FE_OCP_RBN5794_n_13962;
wire FE_OCP_RBN5795_n_13962;
wire FE_OCP_RBN5796_n_13962;
wire FE_OCP_RBN5797_n_13962;
wire FE_OCP_RBN5798_n_13962;
wire FE_OCP_RBN5799_n_13962;
wire FE_OCP_RBN5800_n_13962;
wire FE_OCP_RBN5801_n_13962;
wire FE_OCP_RBN5802_n_13962;
wire FE_OCP_RBN5803_FE_RN_2224_0;
wire FE_OCP_RBN5804_n_47018;
wire FE_OCP_RBN5805_n_47018;
wire FE_OCP_RBN5806_n_47018;
wire FE_OCP_RBN5807_n_47018;
wire FE_OCP_RBN5808_n_47018;
wire FE_OCP_RBN5809_n_3645;
wire FE_OCP_RBN5810_n_3645;
wire FE_OCP_RBN5811_n_3645;
wire FE_OCP_RBN5812_n_9014;
wire FE_OCP_RBN5813_n_9014;
wire FE_OCP_RBN5814_n_20098;
wire FE_OCP_RBN5815_n_24823;
wire FE_OCP_RBN5816_n_38678;
wire FE_OCP_RBN5817_n_8687;
wire FE_OCP_RBN5818_n_8687;
wire FE_OCP_RBN5819_n_8651;
wire FE_OCP_RBN5820_n_3396;
wire FE_OCP_RBN5821_n_3437;
wire FE_OCP_RBN5822_n_8985;
wire FE_OCP_RBN5823_n_14722;
wire FE_OCP_RBN5824_n_14552;
wire FE_OCP_RBN5825_n_8692;
wire FE_OCP_RBN5826_n_8692;
wire FE_OCP_RBN5827_n_44579;
wire FE_OCP_RBN5828_n_44579;
wire FE_OCP_RBN5829_n_44579;
wire FE_OCP_RBN5830_n_44579;
wire FE_OCP_RBN5833_n_44563;
wire FE_OCP_RBN5834_n_44563;
wire FE_OCP_RBN5835_n_44563;
wire FE_OCP_RBN5836_n_44563;
wire FE_OCP_RBN5837_n_44563;
wire FE_OCP_RBN5838_n_44563;
wire FE_OCP_RBN5842_n_44563;
wire FE_OCP_RBN5843_n_9035;
wire FE_OCP_RBN5844_n_42169;
wire FE_OCP_RBN5845_n_42169;
wire FE_OCP_RBN5846_FE_RN_987_0;
wire FE_OCP_RBN5847_FE_RN_987_0;
wire FE_OCP_RBN5848_FE_RN_2187_0;
wire FE_OCP_RBN5849_FE_RN_2187_0;
wire FE_OCP_RBN5850_FE_RN_2187_0;
wire FE_OCP_RBN5851_n_3625;
wire FE_OCP_RBN5852_n_3625;
wire FE_OCP_RBN5853_n_14750;
wire FE_OCP_RBN5854_n_34908;
wire FE_OCP_RBN5855_n_3807;
wire FE_OCP_RBN5856_n_3807;
wire FE_OCP_RBN5857_FE_RN_998_0;
wire FE_OCP_RBN5858_FE_RN_998_0;
wire FE_OCP_RBN5859_FE_RN_998_0;
wire FE_OCP_RBN5860_FE_RN_998_0;
wire FE_OCP_RBN5861_n_3718;
wire FE_OCP_RBN5862_n_3718;
wire FE_OCP_RBN5863_n_3705;
wire FE_OCP_RBN5864_n_3705;
wire FE_OCP_RBN5867_n_3661;
wire FE_OCP_RBN5868_n_3704;
wire FE_OCP_RBN5869_n_3704;
wire FE_OCP_RBN5870_n_3704;
wire FE_OCP_RBN5871_n_3700;
wire FE_OCP_RBN5872_n_3700;
wire FE_OCP_RBN5873_n_3700;
wire FE_OCP_RBN5875_n_3700;
wire FE_OCP_RBN5876_n_3848;
wire FE_OCP_RBN5877_n_3848;
wire FE_OCP_RBN5880_FE_RN_314_0;
wire FE_OCP_RBN5881_FE_RN_314_0;
wire FE_OCP_RBN5882_FE_RN_2220_0;
wire FE_OCP_RBN5883_n_9042;
wire FE_OCP_RBN5884_n_9306;
wire FE_OCP_RBN5885_n_38806;
wire FE_OCP_RBN5890_n_38806;
wire FE_OCP_RBN5892_n_38806;
wire FE_OCP_RBN5893_n_38806;
wire FE_OCP_RBN5894_n_38806;
wire FE_OCP_RBN5895_n_38806;
wire FE_OCP_RBN5896_n_38806;
wire FE_OCP_RBN5897_n_38806;
wire FE_OCP_RBN5898_n_35005;
wire FE_OCP_RBN5899_n_35005;
wire FE_OCP_RBN5900_n_25178;
wire FE_OCP_RBN5901_n_25178;
wire FE_OCP_RBN5902_n_25178;
wire FE_OCP_RBN5903_n_25178;
wire FE_OCP_RBN5904_n_8872;
wire FE_OCP_RBN5905_n_44563;
wire FE_OCP_RBN5906_n_44563;
wire FE_OCP_RBN5907_n_44563;
wire FE_OCP_RBN5908_n_44563;
wire FE_OCP_RBN5909_n_44563;
wire FE_OCP_RBN5910_n_44563;
wire FE_OCP_RBN5911_n_44563;
wire FE_OCP_RBN5912_n_44563;
wire FE_OCP_RBN5913_n_44563;
wire FE_OCP_RBN5914_n_3750;
wire FE_OCP_RBN5915_n_3750;
wire FE_OCP_RBN5916_n_3875;
wire FE_OCP_RBN5917_n_4101;
wire FE_OCP_RBN5918_n_4101;
wire FE_OCP_RBN5919_n_9456;
wire FE_OCP_RBN5920_n_9456;
wire FE_OCP_RBN5921_n_20236;
wire FE_OCP_RBN5922_n_25211;
wire FE_OCP_RBN5923_n_25211;
wire FE_OCP_RBN5924_n_25211;
wire FE_OCP_RBN5925_n_25211;
wire FE_OCP_RBN5926_n_25211;
wire FE_OCP_RBN5927_n_25211;
wire FE_OCP_RBN5929_n_4158;
wire FE_OCP_RBN5930_n_44563;
wire FE_OCP_RBN5931_n_44563;
wire FE_OCP_RBN5932_n_44563;
wire FE_OCP_RBN5933_n_44563;
wire FE_OCP_RBN5934_n_44563;
wire FE_OCP_RBN5935_n_44563;
wire FE_OCP_RBN5936_n_44563;
wire FE_OCP_RBN5937_n_44563;
wire FE_OCP_RBN5938_n_44563;
wire FE_OCP_RBN5939_n_44563;
wire FE_OCP_RBN5940_n_4238;
wire FE_OCP_RBN5941_n_9374;
wire FE_OCP_RBN5942_n_25544;
wire FE_OCP_RBN5943_n_35207;
wire FE_OCP_RBN5944_n_35207;
wire FE_OCP_RBN5945_FE_RN_1231_0;
wire FE_OCP_RBN5946_n_14982;
wire FE_OCP_RBN5947_n_14982;
wire FE_OCP_RBN5948_n_14982;
wire FE_OCP_RBN5949_FE_OFN4772_n_44463;
wire FE_OCP_RBN5950_FE_OFN4772_n_44463;
wire FE_OCP_RBN5951_FE_OFN4772_n_44463;
wire FE_OCP_RBN5952_FE_OFN4772_n_44463;
wire FE_OCP_RBN5953_FE_OFN4772_n_44463;
wire FE_OCP_RBN5954_FE_OFN4772_n_44463;
wire FE_OCP_RBN5955_FE_OFN4772_n_44463;
wire FE_OCP_RBN5956_n_47012;
wire FE_OCP_RBN5957_n_47012;
wire FE_OCP_RBN5958_n_4165;
wire FE_OCP_RBN5959_n_4165;
wire FE_OCP_RBN5960_n_4397;
wire FE_OCP_RBN5961_n_20459;
wire FE_OCP_RBN5962_n_20459;
wire FE_OCP_RBN5963_n_39097;
wire FE_OCP_RBN5964_n_39097;
wire FE_OCP_RBN5965_n_39097;
wire FE_OCP_RBN5966_n_39098;
wire FE_OCP_RBN5967_n_14905;
wire FE_OCP_RBN5968_n_14905;
wire FE_OCP_RBN5969_n_9668;
wire FE_OCP_RBN5970_n_15235;
wire FE_OCP_RBN5971_n_20510;
wire FE_OCP_RBN5972_n_9494;
wire FE_OCP_RBN5973_n_35231;
wire FE_OCP_RBN5974_FE_RN_2033_0;
wire FE_OCP_RBN5975_FE_RN_2033_0;
wire FE_OCP_RBN5976_FE_RN_2033_0;
wire FE_OCP_RBN5977_n_4245;
wire FE_OCP_RBN5978_n_9682;
wire FE_OCP_RBN5979_n_9682;
wire FE_OCP_RBN5980_n_9682;
wire FE_OCP_RBN5981_n_9856;
wire FE_OCP_RBN5982_n_15160;
wire FE_OCP_RBN5983_n_20495;
wire FE_OCP_RBN5984_n_15079;
wire FE_OCP_RBN5985_n_15079;
wire FE_OCP_RBN5987_n_15135;
wire FE_OCP_RBN5988_FE_RN_1865_0;
wire FE_OCP_RBN5989_FE_RN_1865_0;
wire FE_OCP_RBN5990_FE_RN_1865_0;
wire FE_OCP_RBN5991_n_4226;
wire FE_OCP_RBN5992_n_4376;
wire FE_OCP_RBN5993_n_15387;
wire FE_OCP_RBN5994_n_15387;
wire FE_OCP_RBN5995_n_25702;
wire FE_OCP_RBN5996_n_25732;
wire FE_OCP_RBN5997_n_25732;
wire FE_OCP_RBN5998_n_25732;
wire FE_OCP_RBN6000_n_30534;
wire FE_OCP_RBN6001_n_30534;
wire FE_OCP_RBN6002_n_10015;
wire FE_OCP_RBN6003_n_10068;
wire FE_OCP_RBN6004_n_10068;
wire FE_OCP_RBN6005_n_15704;
wire FE_OCP_RBN6006_n_15704;
wire FE_OCP_RBN6008_n_30608;
wire FE_OCP_RBN6009_n_4683;
wire FE_OCP_RBN6010_n_10277;
wire FE_OCP_RBN6011_n_10277;
wire FE_OCP_RBN6012_n_10277;
wire FE_OCP_RBN6013_n_25900;
wire FE_OCP_RBN6015_n_10225;
wire FE_OCP_RBN6016_n_30625;
wire FE_OCP_RBN6017_n_20945;
wire FE_OCP_RBN6018_n_25895;
wire FE_OCP_RBN6019_n_46959;
wire FE_OCP_RBN6020_n_46959;
wire FE_OCP_RBN6021_n_46959;
wire FE_OCP_RBN6022_n_46959;
wire FE_OCP_RBN6023_n_30711;
wire FE_OCP_RBN6024_n_30711;
wire FE_OCP_RBN6025_n_4858;
wire FE_OCP_RBN6026_n_4858;
wire FE_OCP_RBN6027_n_10445;
wire FE_OCP_RBN6028_n_25928;
wire FE_OCP_RBN6029_n_25928;
wire FE_OCP_RBN6031_n_25997;
wire FE_OCP_RBN6032_n_30706;
wire FE_OCP_RBN6033_n_46962;
wire FE_OCP_RBN6034_n_46962;
wire FE_OCP_RBN6035_n_30769;
wire FE_OCP_RBN6036_n_10399;
wire FE_OCP_RBN6037_n_10399;
wire FE_OCP_RBN6038_n_30733;
wire FE_OCP_RBN6039_n_30733;
wire FE_OCP_RBN6040_n_4800;
wire FE_OCP_RBN6041_n_10511;
wire FE_OCP_RBN6044_n_35487;
wire FE_OCP_RBN6045_n_35487;
wire FE_OCP_RBN6046_n_35487;
wire FE_OCP_RBN6047_n_35487;
wire FE_OCP_RBN6048_n_35487;
wire FE_OCP_RBN6049_n_10570;
wire FE_OCP_RBN6050_n_21118;
wire FE_OCP_RBN6051_n_21118;
wire FE_OCP_RBN6053_n_15514;
wire FE_OCP_RBN6055_n_46957;
wire FE_OCP_RBN6056_n_46957;
wire FE_OCP_RBN6057_n_16011;
wire FE_OCP_RBN6058_n_10478;
wire FE_OCP_RBN6059_n_15795;
wire FE_OCP_RBN6060_n_21194;
wire FE_OCP_RBN6061_n_21194;
wire FE_OCP_RBN6062_n_21194;
wire FE_OCP_RBN6063_n_30908;
wire FE_OCP_RBN6064_n_30908;
wire FE_OCP_RBN6065_n_26081;
wire FE_OCP_RBN6066_n_26081;
wire FE_OCP_RBN6067_n_26121;
wire FE_OCP_RBN6068_n_26121;
wire FE_OCP_RBN6069_n_26140;
wire FE_OCP_RBN6070_n_16041;
wire FE_OCP_RBN6071_n_16041;
wire FE_OCP_RBN6072_n_16086;
wire FE_OCP_RBN6073_n_16086;
wire FE_OCP_RBN6074_n_44256;
wire FE_OCP_RBN6075_n_44256;
wire FE_OCP_RBN6076_n_44256;
wire FE_OCP_RBN6077_n_16084;
wire FE_OCP_RBN6078_n_16084;
wire FE_OCP_RBN6079_n_30965;
wire FE_OCP_RBN6080_n_5346;
wire FE_OCP_RBN6081_n_5486;
wire FE_OCP_RBN6082_n_5454;
wire FE_OCP_RBN6083_n_5454;
wire FE_OCP_RBN6084_n_31010;
wire FE_OCP_RBN6085_n_31010;
wire FE_OCP_RBN6086_n_10852;
wire FE_OCP_RBN6087_n_10852;
wire FE_OCP_RBN6088_n_26181;
wire FE_OCP_RBN6089_n_26304;
wire FE_OCP_RBN6090_n_26322;
wire FE_OCP_RBN6091_n_31153;
wire FE_OCP_RBN6092_n_5531;
wire FE_OCP_RBN6093_n_10660;
wire FE_OCP_RBN6094_n_10946;
wire FE_OCP_RBN6095_n_26160;
wire FE_OCP_RBN6096_n_26160;
wire FE_OCP_RBN6097_n_26160;
wire FE_OCP_RBN6098_n_5614;
wire FE_OCP_RBN6101_n_21636;
wire FE_OCP_RBN6102_n_26358;
wire FE_OCP_RBN6104_n_36199;
wire FE_OCP_RBN6105_n_39793;
wire FE_OCP_RBN6106_n_39793;
wire FE_OCP_RBN6108_n_39793;
wire FE_OCP_RBN6109_n_43022;
wire FE_OCP_RBN6110_n_43022;
wire FE_OCP_RBN6111_n_5444;
wire FE_OCP_RBN6112_n_5444;
wire FE_OCP_RBN6113_n_5444;
wire FE_OCP_RBN6114_n_5444;
wire FE_OCP_RBN6115_n_5444;
wire FE_OCP_RBN6116_n_11004;
wire FE_OCP_RBN6117_n_11004;
wire FE_OCP_RBN6118_n_5555;
wire FE_OCP_RBN6119_n_5555;
wire FE_OCP_RBN6120_n_26398;
wire FE_OCP_RBN6121_n_26398;
wire FE_OCP_RBN6122_n_10904;
wire FE_OCP_RBN6123_n_21630;
wire FE_OCP_RBN6124_n_5465;
wire FE_OCP_RBN6127_n_11026;
wire FE_OCP_RBN6128_n_11026;
wire FE_OCP_RBN6129_n_21804;
wire FE_OCP_RBN6130_n_46424;
wire FE_OCP_RBN6131_n_21736;
wire FE_OCP_RBN6132_n_26778;
wire FE_OCP_RBN6133_n_11169;
wire FE_OCP_RBN6134_n_11221;
wire FE_OCP_RBN6135_n_16553;
wire FE_OCP_RBN6136_n_5816;
wire FE_OCP_RBN6137_n_11364;
wire FE_OCP_RBN6138_n_31520;
wire FE_OCP_RBN6139_n_31520;
wire FE_OCP_RBN6144_n_46285;
wire FE_OCP_RBN6149_n_5974;
wire FE_OCP_RBN6150_n_36501;
wire FE_OCP_RBN6151_n_36501;
wire FE_OCP_RBN6152_n_39816;
wire FE_OCP_RBN6153_n_39816;
wire FE_OCP_RBN6154_n_39816;
wire FE_OCP_RBN6155_n_39816;
wire FE_OCP_RBN6156_n_39816;
wire FE_OCP_RBN6157_n_39816;
wire FE_OCP_RBN6158_n_39816;
wire FE_OCP_RBN6159_n_39816;
wire FE_OCP_RBN6160_n_39816;
wire FE_OCP_RBN6161_n_39816;
wire FE_OCP_RBN6162_FE_RN_1136_0;
wire FE_OCP_RBN6163_n_46337;
wire FE_OCP_RBN6164_n_46337;
wire FE_OCP_RBN6165_n_46337;
wire FE_OCP_RBN6166_n_46337;
wire FE_OCP_RBN6167_n_46337;
wire FE_OCP_RBN6168_n_46337;
wire FE_OCP_RBN6169_n_6021;
wire FE_OCP_RBN6170_n_6059;
wire FE_OCP_RBN6171_n_6059;
wire FE_OCP_RBN6172_n_16923;
wire FE_OCP_RBN6173_n_16923;
wire FE_OCP_RBN6174_n_16923;
wire FE_OCP_RBN6175_n_16923;
wire FE_OCP_RBN6176_n_16923;
wire FE_OCP_RBN6177_n_36444;
wire FE_OCP_RBN6178_n_22106;
wire FE_OCP_RBN6179_n_22106;
wire FE_OCP_RBN6182_n_44267;
wire FE_OCP_RBN6183_n_44267;
wire FE_OCP_RBN6184_n_44267;
wire FE_OCP_RBN6185_n_44267;
wire FE_OCP_RBN6186_n_16824;
wire FE_OCP_RBN6187_n_31916;
wire FE_OCP_RBN6188_n_11403;
wire FE_OCP_RBN6189_n_11403;
wire FE_OCP_RBN6190_n_43103;
wire FE_OCP_RBN6191_n_43103;
wire FE_OCP_RBN6192_n_43103;
wire FE_OCP_RBN6193_n_10636;
wire FE_OCP_RBN6194_n_10636;
wire FE_OCP_RBN6195_FE_OFN789_n_46195;
wire FE_OCP_RBN6196_FE_OFN789_n_46195;
wire FE_OCP_RBN6197_FE_OFN789_n_46195;
wire FE_OCP_RBN6198_FE_OFN789_n_46195;
wire FE_OCP_RBN6199_FE_OFN789_n_46195;
wire FE_OCP_RBN6200_FE_OFN789_n_46195;
wire FE_OCP_RBN6201_FE_OFN789_n_46195;
wire FE_OCP_RBN6202_n_31819;
wire FE_OCP_RBN6203_n_31819;
wire FE_OCP_RBN6204_n_31819;
wire FE_OCP_RBN6207_n_11486;
wire FE_OCP_RBN6208_n_11486;
wire FE_OCP_RBN6209_n_11486;
wire FE_OCP_RBN6211_n_22421;
wire FE_OCP_RBN6212_n_16962;
wire FE_OCP_RBN6213_n_27086;
wire FE_OCP_RBN6214_n_27086;
wire FE_OCP_RBN6216_n_27086;
wire FE_OCP_RBN6217_n_27110;
wire FE_OCP_RBN6218_n_27110;
wire FE_OCP_RBN6219_n_27110;
wire FE_OCP_RBN6220_n_27110;
wire FE_OCP_RBN6221_n_27110;
wire FE_OCP_RBN6222_n_27110;
wire FE_OCP_RBN6223_n_27110;
wire FE_OCP_RBN6224_n_32061;
wire FE_OCP_RBN6225_n_11713;
wire FE_OCP_RBN6226_n_32178;
wire FE_OCP_RBN6227_n_32216;
wire FE_OCP_RBN6228_n_40565;
wire FE_OCP_RBN6229_n_36693;
wire FE_OCP_RBN6230_n_43882;
wire FE_OCP_RBN6231_n_22639;
wire FE_OCP_RBN6232_n_22639;
wire FE_OCP_RBN6233_n_27504;
wire FE_OCP_RBN6234_n_36778;
wire FE_OCP_RBN6235_n_36780;
wire FE_OCP_RBN6236_n_40586;
wire FE_OCP_RBN6237_n_11853;
wire FE_OCP_RBN6238_n_22718;
wire FE_OCP_RBN6239_n_6456;
wire FE_OCP_RBN6240_n_6438;
wire FE_OCP_RBN6241_n_22622;
wire FE_OCP_RBN6242_n_27436;
wire FE_OCP_RBN6243_n_32305;
wire FE_OCP_RBN6244_n_6535;
wire FE_OCP_RBN6245_n_17587;
wire FE_OCP_RBN6246_n_17587;
wire FE_OCP_RBN6247_n_6477;
wire FE_OCP_RBN6248_n_6477;
wire FE_OCP_RBN6249_n_6567;
wire FE_OCP_RBN6250_n_6567;
wire FE_OCP_RBN6251_n_12067;
wire FE_OCP_RBN6252_n_12067;
wire FE_OCP_RBN6253_n_12117;
wire FE_OCP_RBN6254_n_17723;
wire FE_OCP_RBN6255_FE_RN_1283_0;
wire FE_OCP_RBN6256_FE_RN_2452_0;
wire FE_OCP_RBN6257_n_43842;
wire FE_OCP_RBN6258_n_27743;
wire FE_OCP_RBN6259_n_27726;
wire FE_OCP_RBN6307_n_45224;
wire FE_OCP_RBN6308_n_45224;
wire FE_OCP_RBN6309_n_45224;
wire FE_OCP_RBN6310_n_45224;
wire FE_OCP_RBN6311_n_45224;
wire FE_OCP_RBN6312_n_45224;
wire FE_OCP_RBN6313_n_45224;
wire FE_OCP_RBN6314_n_45224;
wire FE_OCP_RBN6315_n_45224;
wire FE_OCP_RBN6316_n_45224;
wire FE_OCP_RBN6317_n_45224;
wire FE_OCP_RBN6318_n_45224;
wire FE_OCP_RBN6319_n_45224;
wire FE_OCP_RBN6320_n_45224;
wire FE_OCP_RBN6321_n_45224;
wire FE_OCP_RBN6369_n_27773;
wire FE_OCP_RBN6370_n_17582;
wire FE_OCP_RBN6371_FE_RN_1425_0;
wire FE_OCP_RBN6372_FE_RN_1425_0;
wire FE_OCP_RBN6373_n_19701;
wire FE_OCP_RBN6374_n_19722;
wire FE_OCP_RBN6375_n_14154;
wire FE_OCP_RBN6376_n_14154;
wire FE_OCP_RBN6377_n_14380;
wire FE_OCP_RBN6378_n_14380;
wire FE_OCP_RBN6379_n_14380;
wire FE_OCP_RBN6380_n_20125;
wire FE_OCP_RBN6381_n_30824;
wire FE_OCP_RBN6382_n_21087;
wire FE_OCP_RBN6383_n_21087;
wire FE_OCP_RBN6384_n_21087;
wire FE_OCP_RBN6385_n_21429;
wire FE_OCP_RBN6386_n_21429;
wire FE_OCP_RBN6387_n_32238;
wire FE_OCP_RBN6388_n_32238;
wire FE_OCP_RBN6407_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN6408_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN6409_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN6410_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN6413_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN6435_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN6438_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN6439_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN6440_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN6442_delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire FE_OCP_RBN6444_delay_xor_ln21_unr9_stage4_stallmux_q_1_;
wire FE_OCP_RBN6463_n_44061;
wire FE_OCP_RBN6464_n_44061;
wire FE_OCP_RBN6465_n_44061;
wire FE_OCP_RBN6466_n_44061;
wire FE_OCP_RBN6467_n_44061;
wire FE_OCP_RBN6468_n_44061;
wire FE_OCP_RBN6471_delay_xor_ln21_unr15_stage6_stallmux_q_3_;
wire FE_OCP_RBN6499_n_44610;
wire FE_OCP_RBN6500_n_44610;
wire FE_OCP_RBN6501_n_44610;
wire FE_OCP_RBN6502_n_44610;
wire FE_OCP_RBN6503_n_44610;
wire FE_OCP_RBN6506_delay_add_ln22_unr23_stage9_stallmux_q_24_;
wire FE_OCP_RBN6507_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN6508_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN6509_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN6511_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN6512_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN6513_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN6514_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN6515_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN6516_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN6517_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN6518_n_32706;
wire FE_OCP_RBN6519_n_32706;
wire FE_OCP_RBN6520_n_32706;
wire FE_OCP_RBN6521_n_32706;
wire FE_OCP_RBN6523_n_45224;
wire FE_OCP_RBN6524_n_6649;
wire FE_OCP_RBN6525_n_11829;
wire FE_OCP_RBN6526_n_44962;
wire FE_OCP_RBN6527_n_44962;
wire FE_OCP_RBN6528_n_6745;
wire FE_OCP_RBN6529_n_6745;
wire FE_OCP_RBN6530_n_22822;
wire FE_OCP_RBN6531_n_11780;
wire FE_OCP_RBN6532_n_32791;
wire FE_OCP_RBN6533_n_32436;
wire FE_OCP_RBN6534_n_1577;
wire FE_OCP_RBN6535_n_1602;
wire FE_OCP_RBN6536_n_1602;
wire FE_OCP_RBN6537_n_1614;
wire FE_OCP_RBN6538_n_1614;
wire FE_OCP_RBN6539_n_44083;
wire FE_OCP_RBN6540_n_44083;
wire FE_OCP_RBN6541_n_44083;
wire FE_OCP_RBN6542_n_23186;
wire FE_OCP_RBN6543_n_45145;
wire FE_OCP_RBN6544_n_45145;
wire FE_OCP_RBN6545_n_1672;
wire FE_OCP_RBN6546_n_1672;
wire FE_OCP_RBN6547_n_1725;
wire FE_OCP_RBN6548_n_1725;
wire FE_OCP_RBN6549_n_37377;
wire FE_OCP_RBN6550_n_37377;
wire FE_OCP_RBN6551_n_1905;
wire FE_OCP_RBN6552_n_28458;
wire FE_OCP_RBN6553_n_28458;
wire FE_OCP_RBN6554_n_28458;
wire FE_OCP_RBN6555_n_28458;
wire FE_OCP_RBN6556_n_28458;
wire FE_OCP_RBN6557_n_23572;
wire FE_OCP_RBN6558_n_23572;
wire FE_OCP_RBN6559_n_23572;
wire FE_OCP_RBN6560_n_23572;
wire FE_OCP_RBN6561_n_33208;
wire FE_OCP_RBN6562_n_33208;
wire FE_OCP_RBN6563_n_12753;
wire FE_OCP_RBN6564_n_12753;
wire FE_OCP_RBN6565_n_12753;
wire FE_OCP_RBN6566_n_33368;
wire FE_OCP_RBN6567_n_12714;
wire FE_OCP_RBN6568_n_33803;
wire FE_OCP_RBN6569_n_33803;
wire FE_OCP_RBN6570_n_44875;
wire FE_OCP_RBN6571_n_44875;
wire FE_OCP_RBN6572_n_44875;
wire FE_OCP_RBN6573_n_44875;
wire FE_OCP_RBN6574_n_44875;
wire FE_OCP_RBN6575_n_44875;
wire FE_OCP_RBN6576_n_13011;
wire FE_OCP_RBN6577_n_13011;
wire FE_OCP_RBN6578_n_8676;
wire FE_OCP_RBN6579_n_8676;
wire FE_OCP_RBN6580_n_8676;
wire FE_OCP_RBN6581_n_8021;
wire FE_OCP_RBN6582_n_8021;
wire FE_OCP_RBN6583_n_8021;
wire FE_OCP_RBN6584_n_41491;
wire FE_OCP_RBN6585_n_41491;
wire FE_OCP_RBN6586_n_41491;
wire FE_OCP_RBN6587_n_41491;
wire FE_OCP_RBN6588_n_41491;
wire FE_OCP_RBN6589_n_41491;
wire FE_OCP_RBN6590_n_41491;
wire FE_OCP_RBN6591_n_41491;
wire FE_OCP_RBN6592_n_41491;
wire FE_OCP_RBN6593_n_41491;
wire FE_OCP_RBN6594_n_41491;
wire FE_OCP_RBN6595_n_41491;
wire FE_OCP_RBN6596_n_7708;
wire FE_OCP_RBN6597_n_7708;
wire FE_OCP_RBN6598_n_7708;
wire FE_OCP_RBN6599_n_7708;
wire FE_OCP_RBN6600_n_7708;
wire FE_OCP_RBN6601_n_7708;
wire FE_OCP_RBN6602_n_7881;
wire FE_OCP_RBN6603_n_7881;
wire FE_OCP_RBN6604_n_7881;
wire FE_OCP_RBN6605_n_7881;
wire FE_OCP_RBN6606_n_2289;
wire FE_OCP_RBN6607_n_2289;
wire FE_OCP_RBN6608_n_2289;
wire FE_OCP_RBN6609_n_2289;
wire FE_OCP_RBN6610_n_2289;
wire FE_OCP_RBN6611_n_2289;
wire FE_OCP_RBN6612_n_2289;
wire FE_OCP_RBN6613_n_2289;
wire FE_OCP_RBN6614_n_2289;
wire FE_OCP_RBN6615_n_2289;
wire FE_OCP_RBN6616_n_2289;
wire FE_OCP_RBN6617_n_2289;
wire FE_OCP_RBN6618_n_41381;
wire FE_OCP_RBN6619_n_41381;
wire FE_OCP_RBN6620_n_41381;
wire FE_OCP_RBN6621_n_7821;
wire FE_OCP_RBN6622_n_7943;
wire FE_OCP_RBN6623_n_24175;
wire FE_OCP_RBN6624_n_24175;
wire FE_OCP_RBN6625_n_2537;
wire FE_OCP_RBN6626_n_2537;
wire FE_OCP_RBN6627_n_7832;
wire FE_OCP_RBN6628_n_8269;
wire FE_OCP_RBN6629_n_8269;
wire FE_OCP_RBN6630_n_8269;
wire FE_OCP_RBN6631_n_8111;
wire FE_OCP_RBN6632_n_2633;
wire FE_OCP_RBN6633_n_2633;
wire FE_OCP_RBN6634_n_9304;
wire FE_OCP_RBN6635_n_9304;
wire FE_OCP_RBN6636_n_33983;
wire FE_OCP_RBN6637_n_33983;
wire FE_OCP_RBN6638_n_13726;
wire FE_OCP_RBN6639_n_13726;
wire FE_OCP_RBN6640_n_24268;
wire FE_OCP_RBN6641_n_3502;
wire FE_OCP_RBN6642_n_3502;
wire FE_OCP_RBN6643_n_8342;
wire FE_OCP_RBN6644_n_8342;
wire FE_OCP_RBN6645_n_8342;
wire FE_OCP_RBN6646_n_13818;
wire FE_OCP_RBN6647_n_13818;
wire FE_OCP_RBN6648_n_13818;
wire FE_OCP_RBN6649_n_13818;
wire FE_OCP_RBN6650_n_13818;
wire FE_OCP_RBN6651_n_13818;
wire FE_OCP_RBN6652_n_29494;
wire FE_OCP_RBN6653_n_29494;
wire FE_OCP_RBN6654_n_8187;
wire FE_OCP_RBN6655_n_8187;
wire FE_OCP_RBN6656_n_8187;
wire FE_OCP_RBN6657_n_44352;
wire FE_OCP_RBN6658_n_44352;
wire FE_OCP_RBN6659_n_2829;
wire FE_OCP_RBN6660_n_13884;
wire FE_OCP_RBN6661_n_13702;
wire FE_OCP_RBN6662_n_13702;
wire FE_OCP_RBN6663_n_8355;
wire FE_OCP_RBN6664_n_34297;
wire FE_OCP_RBN6665_n_34297;
wire FE_OCP_RBN6666_n_34297;
wire FE_OCP_RBN6667_n_34297;
wire FE_OCP_RBN6668_n_34297;
wire FE_OCP_RBN6669_n_34297;
wire FE_OCP_RBN6670_n_34297;
wire FE_OCP_RBN6671_n_34297;
wire FE_OCP_RBN6672_n_34297;
wire FE_OCP_RBN6673_n_34297;
wire FE_OCP_RBN6674_n_38519;
wire FE_OCP_RBN6675_n_8288;
wire FE_OCP_RBN6676_n_8288;
wire FE_OCP_RBN6677_n_8288;
wire FE_OCP_RBN6678_n_8288;
wire FE_OCP_RBN6679_n_8288;
wire FE_OCP_RBN6680_n_8448;
wire FE_OCP_RBN6681_n_24648;
wire FE_OCP_RBN6682_FE_OCPN4529_FE_OCP_RBN2748_n_8474;
wire FE_OCP_RBN6683_FE_OCPN4529_FE_OCP_RBN2748_n_8474;
wire FE_OCP_RBN6684_FE_OCPN4529_FE_OCP_RBN2748_n_8474;
wire FE_OCP_RBN6685_FE_OCPN4529_FE_OCP_RBN2748_n_8474;
wire FE_OCP_RBN6686_n_3498;
wire FE_OCP_RBN6687_n_3498;
wire FE_OCP_RBN6688_n_3498;
wire FE_OCP_RBN6689_n_38655;
wire FE_OCP_RBN6690_n_38655;
wire FE_OCP_RBN6691_n_8629;
wire FE_OCP_RBN6692_n_13796;
wire FE_OCP_RBN6693_n_13796;
wire FE_OCP_RBN6694_n_13796;
wire FE_OCP_RBN6695_n_13796;
wire FE_OCP_RBN6696_n_13796;
wire FE_OCP_RBN6697_n_13796;
wire FE_OCP_RBN6698_n_13796;
wire FE_OCP_RBN6699_n_13796;
wire FE_OCP_RBN6700_n_13796;
wire FE_OCP_RBN6701_n_14444;
wire FE_OCP_RBN6702_n_14444;
wire FE_OCP_RBN6703_n_14444;
wire FE_OCP_RBN6704_n_8762;
wire FE_OCP_RBN6705_n_8762;
wire FE_OCP_RBN6706_n_29787;
wire FE_OCP_RBN6707_n_8719;
wire FE_OCP_RBN6708_n_44570;
wire FE_OCP_RBN6709_n_44570;
wire FE_OCP_RBN6710_n_44570;
wire FE_OCP_RBN6711_n_44570;
wire FE_OCP_RBN6712_n_44570;
wire FE_OCP_RBN6713_n_8800;
wire FE_OCP_RBN6714_n_3604;
wire FE_OCP_RBN6715_n_3604;
wire FE_OCP_RBN6716_n_3604;
wire FE_OCP_RBN6717_n_3604;
wire FE_OCP_RBN6718_n_3604;
wire FE_OCP_RBN6719_n_3604;
wire FE_OCP_RBN6720_FE_OCP_DRV_N6264_n_9014;
wire FE_OCP_RBN6721_FE_OCP_DRV_N6264_n_9014;
wire FE_OCP_RBN6722_n_9034;
wire FE_OCP_RBN6723_n_44055;
wire FE_OCP_RBN6724_n_44055;
wire FE_OCP_RBN6725_n_34388;
wire FE_OCP_RBN6726_n_34388;
wire FE_OCP_RBN6727_n_34388;
wire FE_OCP_RBN6728_n_34388;
wire FE_OCP_RBN6729_n_44579;
wire FE_OCP_RBN6730_n_44579;
wire FE_OCP_RBN6731_n_44579;
wire FE_OCP_RBN6732_n_44579;
wire FE_OCP_RBN6733_n_44579;
wire FE_OCP_RBN6734_n_44579;
wire FE_OCP_RBN6735_n_44579;
wire FE_OCP_RBN6736_n_44579;
wire FE_OCP_RBN6737_n_44563;
wire FE_OCP_RBN6738_n_44563;
wire FE_OCP_RBN6739_n_44563;
wire FE_OCP_RBN6740_n_44563;
wire FE_OCP_RBN6741_n_44563;
wire FE_OCP_RBN6742_n_3746;
wire FE_OCP_RBN6743_n_3746;
wire FE_OCP_RBN6744_n_3746;
wire FE_OCP_RBN6745_n_3746;
wire FE_OCP_RBN6746_n_30170;
wire FE_OCP_RBN6747_n_30170;
wire FE_OCP_RBN6748_n_30170;
wire FE_OCP_RBN6749_n_9198;
wire FE_OCP_RBN6750_n_9198;
wire FE_OCP_RBN6751_n_9185;
wire FE_OCP_RBN6752_n_30273;
wire FE_OCP_RBN6753_n_35049;
wire FE_OCP_RBN6754_n_38806;
wire FE_OCP_RBN6755_n_38806;
wire FE_OCP_RBN6756_n_38806;
wire FE_OCP_RBN6757_n_38806;
wire FE_OCP_RBN6758_n_38806;
wire FE_OCP_RBN6759_n_9075;
wire FE_OCP_RBN6760_n_9075;
wire FE_OCP_RBN6761_n_3705;
wire FE_OCP_RBN6762_n_3790;
wire FE_OCP_RBN6763_FE_RN_2259_0;
wire FE_OCP_RBN6764_FE_RN_2259_0;
wire FE_OCP_RBN6765_n_3704;
wire FE_OCP_RBN6766_n_3704;
wire FE_OCP_RBN6767_n_3704;
wire FE_OCP_RBN6768_n_3700;
wire FE_OCP_RBN6769_n_3700;
wire FE_OCP_RBN6770_n_3700;
wire FE_OCP_RBN6771_n_3700;
wire FE_OCP_RBN6772_n_3700;
wire FE_OCP_RBN6773_n_4046;
wire FE_OCP_RBN6774_n_4046;
wire FE_OCP_RBN6775_n_4046;
wire FE_OCP_RBN6776_n_4046;
wire FE_OCP_RBN6777_n_4046;
wire FE_OCP_RBN6778_n_4046;
wire FE_OCP_RBN6779_n_4046;
wire FE_OCP_RBN6780_n_4046;
wire FE_OCP_RBN6781_n_4046;
wire FE_OCP_RBN6782_n_4046;
wire FE_OCP_RBN6783_n_4046;
wire FE_OCP_RBN6784_n_4046;
wire FE_OCP_RBN6785_n_14704;
wire FE_OCP_RBN6786_n_9410;
wire FE_OCP_RBN6787_n_35130;
wire FE_OCP_RBN6788_n_35130;
wire FE_OCP_RBN6789_n_20242;
wire FE_OCP_RBN6790_n_20242;
wire FE_OCP_RBN6791_n_20242;
wire FE_OCP_RBN6792_n_9510;
wire FE_OCP_RBN6793_n_25211;
wire FE_OCP_RBN6794_n_25211;
wire FE_OCP_RBN6795_n_25211;
wire FE_OCP_RBN6796_n_25211;
wire FE_OCP_RBN6797_n_25211;
wire FE_OCP_RBN6798_n_15156;
wire FE_OCP_RBN6799_n_15156;
wire FE_OCP_RBN6800_n_15156;
wire FE_OCP_RBN6801_n_15156;
wire FE_OCP_RBN6802_n_15156;
wire FE_OCP_RBN6803_n_20565;
wire FE_OCP_RBN6804_n_9742;
wire FE_OCP_RBN6805_n_9742;
wire FE_OCP_RBN6806_n_4411;
wire FE_OCP_RBN6807_n_15110;
wire FE_OCP_RBN6808_n_20667;
wire FE_OCP_RBN6809_n_4563;
wire FE_OCP_RBN6810_n_39551;
wire FE_OCP_RBN6811_n_39551;
wire FE_OCP_RBN6812_n_30608;
wire FE_OCP_RBN6813_n_30608;
wire FE_OCP_RBN6814_n_9893;
wire FE_OCP_RBN6815_n_25753;
wire FE_OCP_RBN6816_n_4654;
wire FE_OCP_RBN6817_n_20889;
wire FE_OCP_RBN6818_n_25997;
wire FE_OCP_RBN6819_n_25997;
wire FE_OCP_RBN6820_n_5152;
wire FE_OCP_RBN6821_n_45319;
wire FE_OCP_RBN6822_FE_RN_592_0;
wire FE_OCP_RBN6823_FE_RN_592_0;
wire FE_OCP_RBN6824_n_39542;
wire FE_OCP_RBN6825_n_39542;
wire FE_OCP_RBN6826_n_15514;
wire FE_OCP_RBN6827_n_15514;
wire FE_OCP_RBN6828_n_15514;
wire FE_OCP_RBN6829_n_15514;
wire FE_OCP_RBN6830_n_45484;
wire FE_OCP_RBN6831_n_15676;
wire FE_OCP_RBN6832_n_31073;
wire FE_OCP_RBN6833_n_31073;
wire FE_OCP_RBN6834_n_31073;
wire FE_OCP_RBN6835_n_39577;
wire FE_OCP_RBN6836_n_39577;
wire FE_OCP_RBN6837_FE_RN_586_0;
wire FE_OCP_RBN6838_FE_RN_586_0;
wire FE_OCP_RBN6839_FE_RN_2660_0;
wire FE_OCP_RBN6840_FE_RN_2660_0;
wire FE_OCP_RBN6841_n_31023;
wire FE_OCP_RBN6842_n_5397;
wire FE_OCP_RBN6843_n_31194;
wire FE_OCP_RBN6844_n_15599;
wire FE_OCP_RBN6845_n_15599;
wire FE_OCP_RBN6846_n_15599;
wire FE_OCP_RBN6847_n_15599;
wire FE_OCP_RBN6848_n_15599;
wire FE_OCP_RBN6849_n_26358;
wire FE_OCP_RBN6850_n_26504;
wire FE_OCP_RBN6851_n_39793;
wire FE_OCP_RBN6852_n_39793;
wire FE_OCP_RBN6853_n_39793;
wire FE_OCP_RBN6854_n_5735;
wire FE_OCP_RBN6855_n_5735;
wire FE_OCP_RBN6856_n_26160;
wire FE_OCP_RBN6857_n_26160;
wire FE_OCP_RBN6858_n_26160;
wire FE_OCP_RBN6859_n_26160;
wire FE_OCP_RBN6860_n_26160;
wire FE_OCP_RBN6861_n_46285;
wire FE_OCP_RBN6862_n_46285;
wire FE_OCP_RBN6863_n_46285;
wire FE_OCP_RBN6864_n_46285;
wire FE_OCP_RBN6865_n_46285;
wire FE_OCP_RBN6866_n_5743;
wire FE_OCP_RBN6867_n_16392;
wire FE_OCP_RBN6868_n_16392;
wire FE_OCP_RBN6869_n_5751;
wire FE_OCP_RBN6870_FE_RN_2289_0;
wire FE_OCP_RBN6871_FE_RN_2289_0;
wire FE_OCP_RBN6872_n_31520;
wire FE_OCP_RBN6873_n_31520;
wire FE_OCP_RBN6874_n_31520;
wire FE_OCP_RBN6875_n_31520;
wire FE_OCP_RBN6876_n_16920;
wire FE_OCP_RBN6877_n_16920;
wire FE_OCP_RBN6878_n_44267;
wire FE_OCP_RBN6879_n_31819;
wire FE_OCP_RBN6880_n_31819;
wire FE_OCP_RBN6881_n_31819;
wire FE_OCP_RBN6882_n_11486;
wire FE_OCP_RBN6883_n_11486;
wire FE_OCP_RBN7005_n_44962;
wire FE_OCP_RBN7006_n_44962;
wire FE_OCP_RBN7007_n_44962;
wire FE_OCP_RBN7008_n_44962;
wire FE_OCP_RBN7009_n_44962;
wire FE_OCP_RBN7010_n_44962;
wire FE_OCP_RBN7011_n_44962;
wire FE_OCP_RBN7012_n_44962;
wire FE_OCP_RBN7013_n_44962;
wire FE_OCP_RBN7014_n_44962;
wire FE_OCP_RBN7015_n_44962;
wire FE_OCP_RBN7016_n_32687;
wire FE_OCP_RBN7017_n_32687;
wire FE_OCP_RBN7018_n_32649;
wire FE_OCP_RBN7019_n_28166;
wire FE_OCP_RBN7020_n_17717;
wire FE_OCP_RBN7021_n_33330;
wire FE_OCP_RBN7022_n_18248;
wire FE_OCP_RBN7023_n_18650;
wire FE_OCP_RBN7024_FE_RN_1738_0;
wire FE_OCP_RBN7025_n_18873;
wire FE_OCP_RBN7026_n_18866;
wire FE_OCP_RBN7027_n_18866;
wire FE_OCP_RBN7028_n_18866;
wire FE_OCP_RBN7029_n_44259;
wire FE_OCP_RBN7030_n_44259;
wire FE_OCP_RBN7031_n_18981;
wire FE_OCP_RBN7032_n_18981;
wire FE_OCP_RBN7033_n_18981;
wire FE_OCP_RBN7034_n_18981;
wire FE_OCP_RBN7035_n_18981;
wire FE_OCP_RBN7036_n_18982;
wire FE_OCP_RBN7037_n_18982;
wire FE_OCP_RBN7038_n_34903;
wire FE_OCP_RBN7039_n_34903;
wire FE_OCP_RBN7040_n_20167;
wire FE_OCP_RBN7041_n_20336;
wire FE_OCP_RBN7042_n_20336;
wire FE_OCP_RBN7043_n_20336;
wire FE_OCP_RBN7044_FE_RN_1462_0;
wire FE_OCP_RBN7045_FE_RN_1462_0;
wire FE_OCP_RBN7046_n_20941;
wire FE_OCP_RBN7047_n_20941;
wire FE_OCP_RBN7048_n_20941;
wire FE_OCP_RBN7049_n_20941;
wire FE_OCP_RBN7050_n_20941;
wire FE_OCP_RBN7051_n_20941;
wire FE_OCP_RBN7052_n_20941;
wire FE_OCP_RBN7053_n_30867;
wire FE_OCP_RBN7055_FE_OCPN1068_n_21973;
wire FE_OCP_RBN7056_FE_OCPN1068_n_21973;
wire FE_OCP_RBN7057_n_36677;
wire FE_OCP_RBN7101_n_44365;
wire FE_OCP_RBN7102_n_44365;
wire FE_OCP_RBN7103_n_44365;
wire FE_OCP_RBN7104_n_44365;
wire FE_OCP_RBN7105_n_44365;
wire FE_OCP_RBN7106_n_44365;
wire FE_OCP_RBN7107_n_44365;
wire FE_OCP_RBN7108_n_44365;
wire FE_OCP_RBN7109_n_44365;
wire FE_OCP_RBN7110_n_44365;
wire FE_OCP_RBN7111_n_44365;
wire FE_OCP_RBN7112_n_44365;
wire FE_OCP_RBN7113_n_44365;
wire FE_OCP_RBN7114_n_44365;
wire FE_OCP_RBN7117_delay_xor_ln22_unr12_stage5_stallmux_q_0_;
wire FE_OCP_RBN7118_delay_xor_ln22_unr12_stage5_stallmux_q_0_;
wire FE_OCP_RBN7127_n_44722;
wire FE_OCP_RBN7128_n_44722;
wire FE_OCP_RBN7129_n_44722;
wire FE_OCP_RBN7130_n_29262;
wire FE_OCP_RBN7131_n_29262;
wire FE_OCP_RBN983_n_24262;
wire FE_OCP_RBN984_n_22822;
wire FE_OFN0_n_43918;
wire FE_OFN1178_n_916;
wire FE_OFN1180_n_13195;
wire FE_OFN1181_n_13195;
wire FE_OFN1182_n_24059;
wire FE_OFN1183_n_24059;
wire FE_OFN1185_n_19801;
wire FE_OFN1194_n_27014;
wire FE_OFN1196_n_27014;
wire FE_OFN1198_n_27014;
wire FE_OFN1199_n_27014;
wire FE_OFN1_n_43918;
wire FE_OFN230_n_35655;
wire FE_OFN231_n_35655;
wire FE_OFN2_n_43918;
wire FE_OFN321_n_2929;
wire FE_OFN380_n_9391;
wire FE_OFN381_n_9391;
wire FE_OFN3_n_43918;
wire FE_OFN4650_n_43918;
wire FE_OFN4651_n_43918;
wire FE_OFN4652_n_43918;
wire FE_OFN4653_n_43918;
wire FE_OFN4669_n_16873;
wire FE_OFN4701_n_7702;
wire FE_OFN4714_n_18642;
wire FE_OFN4715_n_18642;
wire FE_OFN4730_n_31403;
wire FE_OFN4731_n_31403;
wire FE_OFN4732_n_29677;
wire FE_OFN4733_n_29677;
wire FE_OFN4755_n_41563;
wire FE_OFN4762_n_3029;
wire FE_OFN4763_n_3029;
wire FE_OFN4764_n_3029;
wire FE_OFN4765_n_3029;
wire FE_OFN4766_n_8309;
wire FE_OFN4767_n_8309;
wire FE_OFN4768_n_8309;
wire FE_OFN4769_n_8309;
wire FE_OFN4770_n_8309;
wire FE_OFN4771_n_8309;
wire FE_OFN4772_n_44463;
wire FE_OFN4774_n_44463;
wire FE_OFN4775_n_44463;
wire FE_OFN4776_n_44463;
wire FE_OFN4777_n_44490;
wire FE_OFN4778_n_44490;
wire FE_OFN4779_n_44490;
wire FE_OFN4780_n_45813;
wire FE_OFN4781_n_45813;
wire FE_OFN4782_n_45813;
wire FE_OFN4783_n_45813;
wire FE_OFN4784_n_45813;
wire FE_OFN4785_n_45813;
wire FE_OFN4786_n_45813;
wire FE_OFN4787_n_46137;
wire FE_OFN4788_n_46137;
wire FE_OFN4789_n_46137;
wire FE_OFN4790_n_13195;
wire FE_OFN4791_n_13195;
wire FE_OFN4792_n_13195;
wire FE_OFN4793_n_13195;
wire FE_OFN4794_n_13195;
wire FE_OFN4795_n_13195;
wire FE_OFN4796_n_13195;
wire FE_OFN4797_n_44498;
wire FE_OFN4798_n_44498;
wire FE_OFN4799_n_44498;
wire FE_OFN4800_n_44498;
wire FE_OFN4801_n_44498;
wire FE_OFN4802_n_44498;
wire FE_OFN4804_n_19384;
wire FE_OFN4805_n_19801;
wire FE_OFN4806_n_7702;
wire FE_OFN4807_n_2432;
wire FE_OFN4808_n_28820;
wire FE_OFN4809_n_41563;
wire FE_OFN4810_n_916;
wire FE_OFN4811_n_902;
wire FE_OFN4812_n_16873;
wire FE_OFN4813_n_19384;
wire FE_OFN4814_n_2432;
wire FE_OFN4815_n_4018;
wire FE_OFN4816_n_47017;
wire FE_OFN4817_n_920;
wire FE_OFN4818_n_920;
wire FE_OFN4_n_43918;
wire FE_OFN5063_n_1545;
wire FE_OFN5064_n_1545;
wire FE_OFN5065_n_8904;
wire FE_OFN5066_n_8904;
wire FE_OFN5069_n_13646;
wire FE_OFN5070_n_13646;
wire FE_OFN5071_n_18287;
wire FE_OFN5072_n_18287;
wire FE_OFN5073_delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire FE_OFN5074_delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire FE_OFN5076_n_31435;
wire FE_OFN5077_n_31435;
wire FE_OFN5078_n_29014;
wire FE_OFN5079_n_29014;
wire FE_OFN5080_n_36439;
wire FE_OFN5081_n_36439;
wire FE_OFN5082_n_36750;
wire FE_OFN5083_n_36750;
wire FE_OFN5084_n_36750;
wire FE_OFN5085_delay_sub_ln23_0_unr22_stage8_stallmux_q;
wire FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q;
wire FE_OFN5087_delay_sub_ln23_0_unr22_stage8_stallmux_q;
wire FE_OFN5088_delay_sub_ln23_0_unr25_stage9_stallmux_q;
wire FE_OFN5089_delay_sub_ln23_0_unr25_stage9_stallmux_q;
wire FE_OFN5090_delay_sub_ln23_0_unr25_stage9_stallmux_q;
wire FE_OFN5091_delay_sub_ln23_0_unr25_stage9_stallmux_q;
wire FE_OFN5092_delay_sub_ln23_0_unr25_stage9_stallmux_q;
wire FE_OFN5093_delay_sub_ln23_0_unr25_stage9_stallmux_q;
wire FE_OFN5_n_43918;
wire FE_OFN620_n_28336;
wire FE_OFN621_n_28336;
wire FE_OFN622_n_28336;
wire FE_OFN735_n_17093;
wire FE_OFN736_n_17093;
wire FE_OFN737_n_17093;
wire FE_OFN738_n_17093;
wire FE_OFN739_n_17093;
wire FE_OFN740_delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire FE_OFN741_delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire FE_OFN742_delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire FE_OFN743_delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire FE_OFN744_n_22641;
wire FE_OFN745_n_22641;
wire FE_OFN747_n_22641;
wire FE_OFN748_n_22641;
wire FE_OFN752_n_13889;
wire FE_OFN753_n_13889;
wire FE_OFN754_n_13889;
wire FE_OFN755_n_44464;
wire FE_OFN756_n_44464;
wire FE_OFN757_n_44464;
wire FE_OFN758_n_45813;
wire FE_OFN759_n_45813;
wire FE_OFN765_n_46337;
wire FE_OFN766_n_46137;
wire FE_OFN767_n_46137;
wire FE_OFN768_n_46137;
wire FE_OFN769_n_46196;
wire FE_OFN770_n_46196;
wire FE_OFN771_n_46196;
wire FE_OFN772_n_25834;
wire FE_OFN773_n_25834;
wire FE_OFN774_n_25834;
wire FE_OFN775_n_25834;
wire FE_OFN776_n_18268;
wire FE_OFN777_n_18268;
wire FE_OFN778_n_23803;
wire FE_OFN779_n_23803;
wire FE_OFN780_n_23803;
wire FE_OFN781_n_47017;
wire FE_OFN787_n_46285;
wire FE_OFN789_n_46195;
wire FE_OFN792_n_1909;
wire FE_OFN793_n_2056;
wire FE_OFN794_n_2929;
wire FE_OFN795_n_19885;
wire FE_OFN796_n_2719;
wire FE_OFN797_n_2285;
wire FE_OFN798_n_2620;
wire FE_OFN799_n_2644;
wire FE_OFN800_n_3771;
wire FE_OFN801_n_3902;
wire FE_OFN802_n_3911;
wire FE_OFN803_n_4142;
wire FE_OFN804_n_4575;
wire FE_OFN805_n_4018;
wire FE_OFN806_n_13742;
wire FE_OFN807_n_4686;
wire FE_OFN808_n_3264;
wire FE_OFN809_n_9939;
wire FE_OFN810_n_9028;
wire FE_OFN812_n_902;
wire FE_OFN813_n_1909;
wire FE_OFN814_n_2056;
wire FE_OFN815_n_19885;
wire FE_OFN816_n_2719;
wire FE_OFN817_n_2644;
wire FE_OFN818_n_2620;
wire FE_OFN819_n_2285;
wire FE_OFN81_n_4117;
wire FE_OFN820_n_3771;
wire FE_OFN821_n_3902;
wire FE_OFN822_n_1045;
wire FE_OFN823_n_1045;
wire FE_OFN824_n_1045;
wire FE_OFN825_n_3911;
wire FE_OFN826_n_4142;
wire FE_OFN827_n_4575;
wire FE_OFN828_n_4686;
wire FE_OFN829_n_13742;
wire FE_OFN82_n_4117;
wire FE_OFN830_n_3264;
wire FE_OFN831_n_9939;
wire FE_OFN832_n_9028;
wire FE_RN_1000_0;
wire FE_RN_1005_0;
wire FE_RN_1007_0;
wire FE_RN_1008_0;
wire FE_RN_1009_0;
wire FE_RN_1010_0;
wire FE_RN_1011_0;
wire FE_RN_1012_0;
wire FE_RN_1013_0;
wire FE_RN_1015_0;
wire FE_RN_1016_0;
wire FE_RN_1017_0;
wire FE_RN_1018_0;
wire FE_RN_1019_0;
wire FE_RN_1021_0;
wire FE_RN_1023_0;
wire FE_RN_1025_0;
wire FE_RN_1026_0;
wire FE_RN_1027_0;
wire FE_RN_1028_0;
wire FE_RN_1029_0;
wire TIMEBOOST_net_880;
wire FE_RN_1032_0;
wire TIMEBOOST_net_8;
wire FE_RN_1034_0;
wire TIMEBOOST_net_2512;
wire FE_RN_1038_0;
wire FE_RN_1040_0;
wire FE_RN_1041_0;
wire FE_RN_1042_0;
wire FE_RN_1043_0;
wire FE_RN_1044_0;
wire FE_RN_1045_0;
wire FE_RN_1046_0;
wire FE_RN_1047_0;
wire FE_RN_1048_0;
wire FE_RN_1051_0;
wire TIMEBOOST_net_1806;
wire TIMEBOOST_net_1578;
wire FE_RN_1054_0;
wire FE_RN_1055_0;
wire FE_RN_1056_0;
wire FE_RN_1058_0;
wire FE_RN_1059_0;
wire FE_RN_105_0;
wire FE_RN_1060_0;
wire FE_RN_1061_0;
wire FE_RN_1062_0;
wire FE_RN_1063_0;
wire FE_RN_1065_0;
wire TIMEBOOST_net_169;
wire FE_RN_1069_0;
wire TIMEBOOST_net_793;
wire FE_RN_1070_0;
wire FE_RN_1071_0;
wire FE_RN_1073_0;
wire FE_RN_1074_0;
wire TIMEBOOST_net_201;
wire FE_RN_1077_0;
wire FE_RN_1078_0;
wire FE_RN_107_0;
wire FE_RN_1082_0;
wire FE_RN_1083_0;
wire FE_RN_1086_0;
wire TIMEBOOST_net_600;
wire FE_RN_1088_0;
wire TIMEBOOST_net_2360;
wire FE_RN_1093_0;
wire FE_RN_1094_0;
wire FE_RN_1095_0;
wire FE_RN_1096_0;
wire FE_RN_1097_0;
wire FE_RN_1098_0;
wire FE_RN_1099_0;
wire FE_RN_109_0;
wire FE_RN_10_0;
wire TIMEBOOST_net_286;
wire FE_RN_1101_0;
wire TIMEBOOST_net_1596;
wire FE_RN_1104_0;
wire TIMEBOOST_net_2044;
wire FE_RN_1106_0;
wire FE_RN_110_0;
wire FE_RN_1112_0;
wire TIMEBOOST_net_1002;
wire FE_RN_1116_0;
wire FE_RN_1117_0;
wire FE_RN_1120_0;
wire FE_RN_1121_0;
wire TIMEBOOST_net_661;
wire FE_RN_1123_0;
wire FE_RN_1124_0;
wire FE_RN_1126_0;
wire TIMEBOOST_net_2066;
wire FE_RN_1128_0;
wire TIMEBOOST_net_1297;
wire FE_RN_1132_0;
wire FE_RN_1133_0;
wire FE_RN_1135_0;
wire FE_RN_1136_0;
wire TIMEBOOST_net_1151;
wire TIMEBOOST_net_2889;
wire FE_RN_1141_0;
wire FE_RN_1144_0;
wire FE_RN_1146_0;
wire TIMEBOOST_net_2251;
wire TIMEBOOST_net_1196;
wire FE_RN_1149_0;
wire FE_RN_114_0;
wire FE_RN_1151_0;
wire FE_RN_1152_0;
wire FE_RN_1154_0;
wire FE_RN_1155_0;
wire FE_RN_1156_0;
wire FE_RN_1158_0;
wire FE_RN_115_0;
wire FE_RN_1161_0;
wire FE_RN_1162_0;
wire FE_RN_1163_0;
wire FE_RN_1164_0;
wire FE_RN_1165_0;
wire FE_RN_116_0;
wire TIMEBOOST_net_1226;
wire FE_RN_1171_0;
wire FE_RN_1172_0;
wire FE_RN_1173_0;
wire TIMEBOOST_net_1368;
wire TIMEBOOST_net_1390;
wire FE_RN_1179_0;
wire FE_RN_117_0;
wire FE_RN_1180_0;
wire TIMEBOOST_net_2084;
wire TIMEBOOST_net_1355;
wire FE_RN_1183_0;
wire FE_RN_1184_0;
wire FE_RN_1185_0;
wire FE_RN_118_0;
wire FE_RN_1190_0;
wire FE_RN_1191_0;
wire FE_RN_1192_0;
wire FE_RN_1193_0;
wire FE_RN_1194_0;
wire FE_RN_1195_0;
wire FE_RN_1197_0;
wire TIMEBOOST_net_618;
wire TIMEBOOST_net_1426;
wire TIMEBOOST_net_62;
wire FE_RN_1203_0;
wire FE_RN_1204_0;
wire FE_RN_1205_0;
wire FE_RN_1206_0;
wire FE_RN_1207_0;
wire FE_RN_1209_0;
wire FE_RN_120_0;
wire FE_RN_1210_0;
wire FE_RN_1213_0;
wire FE_RN_121_0;
wire FE_RN_1220_0;
wire FE_RN_1221_0;
wire FE_RN_1223_0;
wire FE_RN_1224_0;
wire FE_RN_1225_0;
wire FE_RN_1226_0;
wire FE_RN_1227_0;
wire FE_RN_1228_0;
wire FE_RN_1229_0;
wire FE_RN_122_0;
wire FE_RN_1231_0;
wire FE_RN_1232_0;
wire FE_RN_1233_0;
wire FE_RN_1234_0;
wire FE_RN_1236_0;
wire FE_RN_1237_0;
wire FE_RN_123_0;
wire FE_RN_1244_0;
wire FE_RN_1245_0;
wire FE_RN_1246_0;
wire FE_RN_1247_0;
wire FE_RN_1248_0;
wire FE_RN_1249_0;
wire FE_RN_124_0;
wire FE_RN_1250_0;
wire FE_RN_1251_0;
wire FE_RN_1255_0;
wire FE_RN_1256_0;
wire TIMEBOOST_net_39;
wire FE_RN_1258_0;
wire FE_RN_1259_0;
wire FE_RN_125_0;
wire TIMEBOOST_net_2228;
wire FE_RN_1267_0;
wire FE_RN_1268_0;
wire FE_RN_1269_0;
wire TIMEBOOST_net_890;
wire FE_RN_1270_0;
wire FE_RN_1271_0;
wire FE_RN_1273_0;
wire FE_RN_1274_0;
wire FE_RN_1275_0;
wire FE_RN_1276_0;
wire TIMEBOOST_net_2435;
wire FE_RN_1279_0;
wire FE_RN_127_0;
wire TIMEBOOST_net_1217;
wire TIMEBOOST_net_729;
wire FE_RN_1282_0;
wire FE_RN_1283_0;
wire FE_RN_1284_0;
wire FE_RN_1285_0;
wire TIMEBOOST_net_731;
wire FE_RN_1287_0;
wire FE_RN_1288_0;
wire FE_RN_1289_0;
wire FE_RN_128_0;
wire FE_RN_1290_0;
wire FE_RN_1291_0;
wire FE_RN_1292_0;
wire FE_RN_1293_0;
wire FE_RN_1294_0;
wire FE_RN_1295_0;
wire FE_RN_1296_0;
wire FE_RN_1299_0;
wire FE_RN_129_0;
wire FE_RN_12_0;
wire FE_RN_1300_0;
wire FE_RN_1301_0;
wire FE_RN_1302_0;
wire FE_RN_1303_0;
wire FE_RN_1304_0;
wire FE_RN_1305_0;
wire FE_RN_1306_0;
wire FE_RN_1307_0;
wire FE_RN_1308_0;
wire FE_RN_1309_0;
wire FE_RN_130_0;
wire FE_RN_1310_0;
wire FE_RN_1311_0;
wire TIMEBOOST_net_452;
wire FE_RN_1313_0;
wire FE_RN_1314_0;
wire FE_RN_1315_0;
wire FE_RN_1316_0;
wire FE_RN_1317_0;
wire FE_RN_1319_0;
wire TIMEBOOST_net_2212;
wire FE_RN_1322_0;
wire FE_RN_1323_0;
wire FE_RN_1324_0;
wire TIMEBOOST_net_1535;
wire FE_RN_1327_0;
wire FE_RN_1328_0;
wire FE_RN_1329_0;
wire FE_RN_132_0;
wire FE_RN_1330_0;
wire FE_RN_1331_0;
wire FE_RN_1332_0;
wire FE_RN_1333_0;
wire FE_RN_1334_0;
wire FE_RN_133_0;
wire FE_RN_1346_0;
wire FE_RN_1347_0;
wire FE_RN_1348_0;
wire FE_RN_1349_0;
wire TIMEBOOST_net_2810;
wire FE_RN_1350_0;
wire FE_RN_1355_0;
wire FE_RN_1356_0;
wire FE_RN_1357_0;
wire FE_RN_1358_0;
wire FE_RN_1359_0;
wire FE_RN_135_0;
wire FE_RN_1360_0;
wire FE_RN_1364_0;
wire TIMEBOOST_net_2040;
wire FE_RN_136_0;
wire FE_RN_1370_0;
wire FE_RN_1371_0;
wire FE_RN_1372_0;
wire FE_RN_1373_0;
wire FE_RN_1374_0;
wire FE_RN_1375_0;
wire TIMEBOOST_net_848;
wire FE_RN_1377_0;
wire FE_RN_1378_0;
wire FE_RN_137_0;
wire FE_RN_1380_0;
wire TIMEBOOST_net_2079;
wire FE_RN_1384_0;
wire FE_RN_1386_0;
wire FE_RN_1387_0;
wire FE_RN_1388_0;
wire FE_RN_1389_0;
wire FE_RN_138_0;
wire FE_RN_1390_0;
wire FE_RN_1391_0;
wire FE_RN_1396_0;
wire FE_RN_1397_0;
wire TIMEBOOST_net_1464;
wire FE_RN_1399_0;
wire FE_RN_13_0;
wire FE_RN_1400_0;
wire FE_RN_1401_0;
wire FE_RN_1402_0;
wire FE_RN_1404_0;
wire FE_RN_1405_0;
wire FE_RN_1406_0;
wire FE_RN_1409_0;
wire TIMEBOOST_net_2135;
wire FE_RN_1410_0;
wire TIMEBOOST_net_1821;
wire TIMEBOOST_net_2325;
wire FE_RN_1414_0;
wire TIMEBOOST_net_930;
wire FE_RN_1416_0;
wire FE_RN_1417_0;
wire FE_RN_141_0;
wire FE_RN_1420_0;
wire FE_RN_1421_0;
wire FE_RN_1424_0;
wire FE_RN_1425_0;
wire FE_RN_1426_0;
wire FE_RN_1431_0;
wire FE_RN_1434_0;
wire FE_RN_1435_0;
wire FE_RN_1436_0;
wire FE_RN_1438_0;
wire FE_RN_1439_0;
wire TIMEBOOST_net_2742;
wire FE_RN_1440_0;
wire FE_RN_1442_0;
wire FE_RN_1446_0;
wire FE_RN_1447_0;
wire FE_RN_1448_0;
wire FE_RN_1449_0;
wire FE_RN_1450_0;
wire FE_RN_1451_0;
wire FE_RN_1452_0;
wire FE_RN_1453_0;
wire FE_RN_1454_0;
wire FE_RN_1455_0;
wire FE_RN_1456_0;
wire FE_RN_1457_0;
wire FE_RN_1458_0;
wire FE_RN_145_0;
wire FE_RN_1460_0;
wire FE_RN_1461_0;
wire FE_RN_1462_0;
wire FE_RN_1463_0;
wire FE_RN_1466_0;
wire FE_RN_1467_0;
wire FE_RN_1468_0;
wire FE_RN_1469_0;
wire TIMEBOOST_net_2692;
wire FE_RN_1470_0;
wire TIMEBOOST_net_1946;
wire FE_RN_1472_0;
wire FE_RN_1474_0;
wire FE_RN_1475_0;
wire FE_RN_1477_0;
wire FE_RN_1478_0;
wire FE_RN_1479_0;
wire FE_RN_147_0;
wire FE_RN_1480_0;
wire FE_RN_1481_0;
wire TIMEBOOST_net_2865;
wire FE_RN_1486_0;
wire FE_RN_1487_0;
wire FE_RN_1488_0;
wire FE_RN_148_0;
wire FE_RN_1490_0;
wire FE_RN_1491_0;
wire FE_RN_1492_0;
wire FE_RN_1493_0;
wire FE_RN_1494_0;
wire FE_RN_1496_0;
wire FE_RN_1497_0;
wire FE_RN_1498_0;
wire FE_RN_149_0;
wire FE_RN_14_0;
wire FE_RN_1500_0;
wire FE_RN_1505_0;
wire FE_RN_1507_0;
wire FE_RN_1508_0;
wire FE_RN_1509_0;
wire FE_RN_150_0;
wire FE_RN_1511_0;
wire FE_RN_1512_0;
wire FE_RN_1513_0;
wire FE_RN_1514_0;
wire FE_RN_1518_0;
wire FE_RN_1519_0;
wire FE_RN_151_0;
wire FE_RN_1520_0;
wire FE_RN_1523_0;
wire FE_RN_1524_0;
wire FE_RN_1525_0;
wire FE_RN_1528_0;
wire FE_RN_1529_0;
wire FE_RN_152_0;
wire FE_RN_1530_0;
wire FE_RN_1531_0;
wire FE_RN_1532_0;
wire FE_RN_1535_0;
wire FE_RN_153_0;
wire FE_RN_1540_0;
wire FE_RN_1541_0;
wire FE_RN_1542_0;
wire FE_RN_1543_0;
wire FE_RN_1544_0;
wire FE_RN_1545_0;
wire FE_RN_1546_0;
wire TIMEBOOST_net_1774;
wire FE_RN_1548_0;
wire FE_RN_154_0;
wire FE_RN_1550_0;
wire TIMEBOOST_net_2808;
wire FE_RN_1553_0;
wire FE_RN_1554_0;
wire FE_RN_1555_0;
wire TIMEBOOST_net_910;
wire FE_RN_1558_0;
wire TIMEBOOST_net_792;
wire TIMEBOOST_net_2716;
wire TIMEBOOST_net_1460;
wire FE_RN_1561_0;
wire FE_RN_1562_0;
wire FE_RN_1563_0;
wire FE_RN_1564_0;
wire FE_RN_1566_0;
wire FE_RN_1567_0;
wire FE_RN_1568_0;
wire FE_RN_1569_0;
wire TIMEBOOST_net_0;
wire FE_RN_1570_0;
wire FE_RN_1571_0;
wire FE_RN_1572_0;
wire FE_RN_1573_0;
wire FE_RN_1574_0;
wire FE_RN_1577_0;
wire FE_RN_1578_0;
wire FE_RN_1579_0;
wire FE_RN_1580_0;
wire TIMEBOOST_net_1855;
wire TIMEBOOST_net_2802;
wire FE_RN_1584_0;
wire FE_RN_1585_0;
wire FE_RN_1586_0;
wire FE_RN_1587_0;
wire FE_RN_1588_0;
wire FE_RN_1589_0;
wire FE_RN_158_0;
wire FE_RN_1590_0;
wire FE_RN_1591_0;
wire FE_RN_1592_0;
wire TIMEBOOST_net_1450;
wire FE_RN_1594_0;
wire TIMEBOOST_net_2785;
wire FE_RN_1597_0;
wire FE_RN_1598_0;
wire FE_RN_1599_0;
wire FE_RN_1600_0;
wire FE_RN_1601_0;
wire TIMEBOOST_net_1621;
wire FE_RN_1603_0;
wire FE_RN_1604_0;
wire TIMEBOOST_net_2390;
wire FE_RN_1606_0;
wire FE_RN_1607_0;
wire FE_RN_1611_0;
wire FE_RN_1612_0;
wire FE_RN_1613_0;
wire FE_RN_1614_0;
wire FE_RN_1615_0;
wire FE_RN_1616_0;
wire FE_RN_1617_0;
wire FE_RN_1618_0;
wire FE_RN_1620_0;
wire TIMEBOOST_net_1336;
wire FE_RN_1622_0;
wire FE_RN_1623_0;
wire FE_RN_1624_0;
wire TIMEBOOST_net_974;
wire FE_RN_1626_0;
wire FE_RN_1628_0;
wire FE_RN_1629_0;
wire FE_RN_162_0;
wire FE_RN_1630_0;
wire FE_RN_1631_0;
wire TIMEBOOST_net_1496;
wire FE_RN_1639_0;
wire FE_RN_163_0;
wire FE_RN_1640_0;
wire FE_RN_1641_0;
wire FE_RN_1642_0;
wire FE_RN_1644_0;
wire FE_RN_1645_0;
wire FE_RN_1646_0;
wire TIMEBOOST_net_794;
wire FE_RN_1648_0;
wire TIMEBOOST_net_2114;
wire FE_RN_1651_0;
wire TIMEBOOST_net_2741;
wire FE_RN_1654_0;
wire FE_RN_1655_0;
wire FE_RN_1656_0;
wire FE_RN_1657_0;
wire FE_RN_1659_0;
wire FE_RN_1660_0;
wire FE_RN_1661_0;
wire FE_RN_1662_0;
wire FE_RN_1663_0;
wire FE_RN_1664_0;
wire FE_RN_1665_0;
wire FE_RN_1666_0;
wire FE_RN_1667_0;
wire TIMEBOOST_net_126;
wire FE_RN_1669_0;
wire FE_RN_1670_0;
wire FE_RN_1671_0;
wire FE_RN_1672_0;
wire FE_RN_1673_0;
wire TIMEBOOST_net_964;
wire TIMEBOOST_net_135;
wire FE_RN_1680_0;
wire FE_RN_1681_0;
wire TIMEBOOST_net_231;
wire FE_RN_1688_0;
wire FE_RN_1689_0;
wire FE_RN_168_0;
wire FE_RN_1697_0;
wire FE_RN_1699_0;
wire FE_RN_169_0;
wire FE_RN_16_0;
wire FE_RN_1700_0;
wire TIMEBOOST_net_2324;
wire FE_RN_1702_0;
wire FE_RN_170_0;
wire FE_RN_1714_0;
wire FE_RN_1715_0;
wire FE_RN_1716_0;
wire FE_RN_1717_0;
wire FE_RN_1718_0;
wire FE_RN_171_0;
wire TIMEBOOST_net_897;
wire FE_RN_1722_0;
wire FE_RN_172_0;
wire FE_RN_1733_0;
wire FE_RN_1734_0;
wire FE_RN_1735_0;
wire FE_RN_1736_0;
wire FE_RN_1737_0;
wire FE_RN_1738_0;
wire FE_RN_173_0;
wire FE_RN_1741_0;
wire FE_RN_1742_0;
wire FE_RN_1743_0;
wire FE_RN_1744_0;
wire FE_RN_1748_0;
wire FE_RN_1750_0;
wire FE_RN_1751_0;
wire FE_RN_1753_0;
wire FE_RN_1754_0;
wire TIMEBOOST_net_138;
wire FE_RN_1757_0;
wire FE_RN_1758_0;
wire FE_RN_1759_0;
wire FE_RN_1760_0;
wire FE_RN_1761_0;
wire FE_RN_1762_0;
wire FE_RN_1763_0;
wire FE_RN_1764_0;
wire FE_RN_1765_0;
wire FE_RN_1766_0;
wire FE_RN_176_0;
wire FE_RN_1774_0;
wire FE_RN_1775_0;
wire TIMEBOOST_net_345;
wire FE_RN_1778_0;
wire FE_RN_1779_0;
wire FE_RN_177_0;
wire FE_RN_1780_0;
wire FE_RN_1781_0;
wire FE_RN_1784_0;
wire FE_RN_1789_0;
wire FE_RN_1790_0;
wire FE_RN_1791_0;
wire FE_RN_1792_0;
wire FE_RN_1793_0;
wire TIMEBOOST_net_1347;
wire FE_RN_1796_0;
wire FE_RN_1797_0;
wire FE_RN_1798_0;
wire FE_RN_179_0;
wire FE_RN_1805_0;
wire FE_RN_1818_0;
wire FE_RN_1819_0;
wire FE_RN_1820_0;
wire FE_RN_1821_0;
wire FE_RN_1822_0;
wire FE_RN_1823_0;
wire FE_RN_1824_0;
wire FE_RN_1825_0;
wire FE_RN_1826_0;
wire FE_RN_1827_0;
wire FE_RN_1828_0;
wire FE_RN_1829_0;
wire FE_RN_1830_0;
wire TIMEBOOST_net_773;
wire FE_RN_1834_0;
wire FE_RN_1838_0;
wire FE_RN_1839_0;
wire FE_RN_183_0;
wire FE_RN_1840_0;
wire FE_RN_1842_0;
wire FE_RN_1844_0;
wire FE_RN_1845_0;
wire FE_RN_1846_0;
wire FE_RN_1849_0;
wire FE_RN_184_0;
wire FE_RN_1855_0;
wire FE_RN_1856_0;
wire FE_RN_1857_0;
wire FE_RN_1858_0;
wire FE_RN_1859_0;
wire FE_RN_185_0;
wire FE_RN_1860_0;
wire FE_RN_1861_0;
wire FE_RN_1862_0;
wire FE_RN_1863_0;
wire FE_RN_1865_0;
wire FE_RN_1867_0;
wire FE_RN_186_0;
wire FE_RN_1872_0;
wire FE_RN_1873_0;
wire FE_RN_1874_0;
wire FE_RN_1875_0;
wire FE_RN_1876_0;
wire FE_RN_1877_0;
wire FE_RN_1878_0;
wire TIMEBOOST_net_1844;
wire FE_RN_1883_0;
wire FE_RN_1885_0;
wire FE_RN_1886_0;
wire FE_RN_1888_0;
wire FE_RN_1889_0;
wire FE_RN_188_0;
wire FE_RN_1890_0;
wire FE_RN_1894_0;
wire FE_RN_1895_0;
wire FE_RN_1896_0;
wire FE_RN_1897_0;
wire FE_RN_1898_0;
wire FE_RN_1899_0;
wire FE_RN_189_0;
wire FE_RN_18_0;
wire FE_RN_1903_0;
wire FE_RN_1904_0;
wire TIMEBOOST_net_33;
wire TIMEBOOST_net_222;
wire FE_RN_1907_0;
wire FE_RN_1908_0;
wire FE_RN_1909_0;
wire FE_RN_190_0;
wire FE_RN_1910_0;
wire FE_RN_1911_0;
wire FE_RN_1912_0;
wire FE_RN_1913_0;
wire TIMEBOOST_net_2689;
wire FE_RN_1915_0;
wire FE_RN_1916_0;
wire TIMEBOOST_net_2223;
wire FE_RN_1918_0;
wire FE_RN_1919_0;
wire FE_RN_191_0;
wire FE_RN_1920_0;
wire FE_RN_1921_0;
wire FE_RN_1922_0;
wire TIMEBOOST_net_2170;
wire FE_RN_1924_0;
wire FE_RN_1925_0;
wire FE_RN_1926_0;
wire FE_RN_1927_0;
wire FE_RN_1928_0;
wire FE_RN_1929_0;
wire FE_RN_1930_0;
wire FE_RN_1931_0;
wire FE_RN_1932_0;
wire FE_RN_1933_0;
wire FE_RN_1934_0;
wire TIMEBOOST_net_553;
wire FE_RN_1936_0;
wire FE_RN_1937_0;
wire TIMEBOOST_net_2703;
wire FE_RN_1939_0;
wire FE_RN_1940_0;
wire TIMEBOOST_net_552;
wire FE_RN_1942_0;
wire FE_RN_1943_0;
wire FE_RN_1944_0;
wire FE_RN_1954_0;
wire FE_RN_1955_0;
wire FE_RN_1956_0;
wire FE_RN_1957_0;
wire FE_RN_1958_0;
wire FE_RN_1959_0;
wire FE_RN_1960_0;
wire FE_RN_1961_0;
wire TIMEBOOST_net_899;
wire FE_RN_1963_0;
wire FE_RN_1964_0;
wire TIMEBOOST_net_2897;
wire FE_RN_1966_0;
wire FE_RN_1967_0;
wire FE_RN_1968_0;
wire FE_RN_1969_0;
wire FE_RN_1970_0;
wire FE_RN_1971_0;
wire FE_RN_1975_0;
wire FE_RN_1976_0;
wire FE_RN_1977_0;
wire FE_RN_1978_0;
wire FE_RN_1979_0;
wire FE_RN_197_0;
wire TIMEBOOST_net_23;
wire FE_RN_1981_0;
wire FE_RN_1982_0;
wire TIMEBOOST_net_1512;
wire TIMEBOOST_net_2333;
wire FE_RN_198_0;
wire TIMEBOOST_net_1751;
wire FE_RN_1994_0;
wire FE_RN_1995_0;
wire FE_RN_1997_0;
wire FE_RN_199_0;
wire FE_RN_19_0;
wire FE_RN_2000_0;
wire FE_RN_2001_0;
wire FE_RN_2002_0;
wire FE_RN_2003_0;
wire FE_RN_2004_0;
wire FE_RN_2009_0;
wire TIMEBOOST_net_2140;
wire FE_RN_2010_0;
wire FE_RN_2012_0;
wire FE_RN_2013_0;
wire FE_RN_2014_0;
wire FE_RN_2015_0;
wire FE_RN_2016_0;
wire FE_RN_2017_0;
wire FE_RN_2018_0;
wire FE_RN_201_0;
wire TIMEBOOST_net_2110;
wire FE_RN_2021_0;
wire TIMEBOOST_net_1573;
wire FE_RN_2023_0;
wire TIMEBOOST_net_265;
wire FE_RN_2025_0;
wire FE_RN_2027_0;
wire FE_RN_202_0;
wire FE_RN_2031_0;
wire FE_RN_2032_0;
wire FE_RN_2033_0;
wire FE_RN_2034_0;
wire FE_RN_2036_0;
wire FE_RN_2037_0;
wire FE_RN_2038_0;
wire FE_RN_2039_0;
wire TIMEBOOST_net_2308;
wire FE_RN_2040_0;
wire FE_RN_2041_0;
wire TIMEBOOST_net_208;
wire FE_RN_2043_0;
wire FE_RN_2044_0;
wire FE_RN_2045_0;
wire FE_RN_2049_0;
wire FE_RN_204_0;
wire FE_RN_2051_0;
wire FE_RN_2056_0;
wire FE_RN_2059_0;
wire TIMEBOOST_net_50;
wire FE_RN_2060_0;
wire FE_RN_2063_0;
wire FE_RN_2064_0;
wire FE_RN_2067_0;
wire FE_RN_2068_0;
wire FE_RN_2069_0;
wire FE_RN_206_0;
wire FE_RN_2070_0;
wire FE_RN_2074_0;
wire FE_RN_2075_0;
wire FE_RN_2076_0;
wire FE_RN_2077_0;
wire TIMEBOOST_net_2691;
wire FE_RN_2079_0;
wire FE_RN_2080_0;
wire TIMEBOOST_net_829;
wire FE_RN_2082_0;
wire TIMEBOOST_net_110;
wire FE_RN_2084_0;
wire FE_RN_2085_0;
wire FE_RN_2086_0;
wire FE_RN_2087_0;
wire FE_RN_2088_0;
wire FE_RN_2089_0;
wire FE_RN_2090_0;
wire FE_RN_2091_0;
wire FE_RN_2092_0;
wire FE_RN_2093_0;
wire FE_RN_2094_0;
wire FE_RN_2095_0;
wire FE_RN_2097_0;
wire FE_RN_2098_0;
wire TIMEBOOST_net_287;
wire FE_RN_2100_0;
wire FE_RN_2101_0;
wire FE_RN_2103_0;
wire TIMEBOOST_net_782;
wire FE_RN_2105_0;
wire FE_RN_2107_0;
wire FE_RN_2108_0;
wire FE_RN_2109_0;
wire FE_RN_210_0;
wire FE_RN_2110_0;
wire FE_RN_2111_0;
wire FE_RN_2112_0;
wire TIMEBOOST_net_2787;
wire TIMEBOOST_net_1452;
wire FE_RN_2115_0;
wire FE_RN_2116_0;
wire FE_RN_2117_0;
wire FE_RN_211_0;
wire TIMEBOOST_net_1653;
wire FE_RN_2124_0;
wire FE_RN_2125_0;
wire FE_RN_2126_0;
wire FE_RN_2127_0;
wire TIMEBOOST_net_1519;
wire FE_RN_2129_0;
wire FE_RN_212_0;
wire FE_RN_2130_0;
wire TIMEBOOST_net_2932;
wire FE_RN_2132_0;
wire FE_RN_2134_0;
wire FE_RN_2135_0;
wire FE_RN_2136_0;
wire FE_RN_2137_0;
wire FE_RN_2138_0;
wire FE_RN_2139_0;
wire FE_RN_213_0;
wire TIMEBOOST_net_1312;
wire TIMEBOOST_net_2868;
wire FE_RN_2142_0;
wire FE_RN_2143_0;
wire FE_RN_2144_0;
wire FE_RN_2145_0;
wire FE_RN_2149_0;
wire FE_RN_214_0;
wire FE_RN_2150_0;
wire FE_RN_2151_0;
wire FE_RN_2154_0;
wire FE_RN_2156_0;
wire FE_RN_2157_0;
wire FE_RN_2159_0;
wire FE_RN_215_0;
wire TIMEBOOST_net_889;
wire FE_RN_2161_0;
wire FE_RN_2162_0;
wire FE_RN_2164_0;
wire FE_RN_2165_0;
wire FE_RN_2166_0;
wire FE_RN_2167_0;
wire FE_RN_2168_0;
wire FE_RN_2169_0;
wire FE_RN_216_0;
wire FE_RN_2170_0;
wire FE_RN_2171_0;
wire FE_RN_2173_0;
wire FE_RN_2174_0;
wire FE_RN_2175_0;
wire TIMEBOOST_net_1831;
wire FE_RN_2177_0;
wire FE_RN_2178_0;
wire TIMEBOOST_net_2296;
wire FE_RN_2180_0;
wire FE_RN_2181_0;
wire FE_RN_2182_0;
wire FE_RN_2183_0;
wire FE_RN_2184_0;
wire FE_RN_2186_0;
wire FE_RN_2187_0;
wire FE_RN_218_0;
wire FE_RN_2191_0;
wire FE_RN_2192_0;
wire FE_RN_2193_0;
wire FE_RN_2194_0;
wire FE_RN_2195_0;
wire FE_RN_2196_0;
wire FE_RN_2197_0;
wire FE_RN_21_0;
wire FE_RN_2200_0;
wire TIMEBOOST_net_2723;
wire FE_RN_2202_0;
wire FE_RN_2203_0;
wire FE_RN_2204_0;
wire FE_RN_2205_0;
wire FE_RN_2206_0;
wire TIMEBOOST_net_1167;
wire FE_RN_2208_0;
wire FE_RN_220_0;
wire FE_RN_2210_0;
wire FE_RN_2211_0;
wire FE_RN_2212_0;
wire FE_RN_2213_0;
wire FE_RN_2214_0;
wire FE_RN_2215_0;
wire FE_RN_2217_0;
wire FE_RN_2218_0;
wire FE_RN_2219_0;
wire FE_RN_221_0;
wire FE_RN_2220_0;
wire FE_RN_2222_0;
wire FE_RN_2224_0;
wire FE_RN_2225_0;
wire FE_RN_2226_0;
wire FE_RN_2227_0;
wire FE_RN_2228_0;
wire FE_RN_2229_0;
wire FE_RN_222_0;
wire FE_RN_2230_0;
wire FE_RN_2231_0;
wire FE_RN_2232_0;
wire FE_RN_2233_0;
wire FE_RN_2234_0;
wire FE_RN_2235_0;
wire FE_RN_2236_0;
wire FE_RN_2237_0;
wire FE_RN_2238_0;
wire FE_RN_2239_0;
wire FE_RN_223_0;
wire FE_RN_2240_0;
wire FE_RN_2241_0;
wire FE_RN_2242_0;
wire FE_RN_2243_0;
wire FE_RN_2244_0;
wire FE_RN_2245_0;
wire TIMEBOOST_net_280;
wire FE_RN_2247_0;
wire FE_RN_2248_0;
wire FE_RN_2249_0;
wire FE_RN_224_0;
wire FE_RN_2250_0;
wire FE_RN_2251_0;
wire TIMEBOOST_net_1963;
wire FE_RN_2253_0;
wire FE_RN_2254_0;
wire FE_RN_2255_0;
wire FE_RN_2257_0;
wire FE_RN_2258_0;
wire FE_RN_2259_0;
wire FE_RN_2260_0;
wire TIMEBOOST_net_2206;
wire FE_RN_2264_0;
wire TIMEBOOST_net_1089;
wire FE_RN_2266_0;
wire FE_RN_2267_0;
wire FE_RN_2268_0;
wire FE_RN_2269_0;
wire FE_RN_2270_0;
wire FE_RN_2271_0;
wire TIMEBOOST_net_1792;
wire FE_RN_2273_0;
wire FE_RN_2274_0;
wire FE_RN_2275_0;
wire FE_RN_2276_0;
wire FE_RN_2277_0;
wire FE_RN_2278_0;
wire FE_RN_2279_0;
wire FE_RN_2280_0;
wire FE_RN_2281_0;
wire TIMEBOOST_net_1790;
wire FE_RN_2283_0;
wire FE_RN_2284_0;
wire FE_RN_2285_0;
wire FE_RN_2286_0;
wire FE_RN_2287_0;
wire FE_RN_2288_0;
wire FE_RN_2289_0;
wire FE_RN_228_0;
wire FE_RN_2291_0;
wire TIMEBOOST_net_519;
wire TIMEBOOST_net_2015;
wire FE_RN_2294_0;
wire FE_RN_2296_0;
wire FE_RN_2297_0;
wire FE_RN_229_0;
wire FE_RN_22_0;
wire FE_RN_2301_0;
wire TIMEBOOST_net_397;
wire FE_RN_2304_0;
wire FE_RN_2305_0;
wire FE_RN_2306_0;
wire FE_RN_2309_0;
wire FE_RN_230_0;
wire FE_RN_2310_0;
wire FE_RN_2311_0;
wire FE_RN_2312_0;
wire FE_RN_2314_0;
wire FE_RN_2316_0;
wire FE_RN_2317_0;
wire FE_RN_2318_0;
wire FE_RN_2319_0;
wire FE_RN_231_0;
wire FE_RN_2320_0;
wire FE_RN_2321_0;
wire FE_RN_2322_0;
wire FE_RN_2323_0;
wire FE_RN_2324_0;
wire FE_RN_2325_0;
wire FE_RN_2326_0;
wire FE_RN_2327_0;
wire FE_RN_2328_0;
wire FE_RN_2329_0;
wire FE_RN_2330_0;
wire FE_RN_2333_0;
wire FE_RN_2334_0;
wire FE_RN_2335_0;
wire FE_RN_2336_0;
wire TIMEBOOST_net_2945;
wire FE_RN_2344_0;
wire FE_RN_2345_0;
wire TIMEBOOST_net_2152;
wire FE_RN_2347_0;
wire TIMEBOOST_net_1431;
wire FE_RN_234_0;
wire FE_RN_2350_0;
wire FE_RN_2351_0;
wire FE_RN_2352_0;
wire FE_RN_2353_0;
wire FE_RN_2355_0;
wire FE_RN_2356_0;
wire FE_RN_2357_0;
wire TIMEBOOST_net_1839;
wire FE_RN_2359_0;
wire FE_RN_235_0;
wire FE_RN_2360_0;
wire FE_RN_2361_0;
wire TIMEBOOST_net_2492;
wire FE_RN_2366_0;
wire FE_RN_2367_0;
wire FE_RN_2368_0;
wire FE_RN_236_0;
wire TIMEBOOST_net_1867;
wire FE_RN_2375_0;
wire FE_RN_2376_0;
wire TIMEBOOST_net_948;
wire TIMEBOOST_net_2818;
wire TIMEBOOST_net_2853;
wire FE_RN_2380_0;
wire TIMEBOOST_net_988;
wire FE_RN_2382_0;
wire FE_RN_2388_0;
wire FE_RN_2389_0;
wire FE_RN_2390_0;
wire FE_RN_2391_0;
wire FE_RN_2392_0;
wire FE_RN_2393_0;
wire FE_RN_2394_0;
wire FE_RN_2395_0;
wire FE_RN_2396_0;
wire TIMEBOOST_net_870;
wire FE_RN_2398_0;
wire FE_RN_2399_0;
wire FE_RN_239_0;
wire FE_RN_23_0;
wire TIMEBOOST_net_980;
wire FE_RN_2401_0;
wire FE_RN_2402_0;
wire FE_RN_2403_0;
wire FE_RN_2404_0;
wire FE_RN_2407_0;
wire FE_RN_2408_0;
wire FE_RN_240_0;
wire FE_RN_2410_0;
wire FE_RN_2411_0;
wire FE_RN_2412_0;
wire TIMEBOOST_net_226;
wire FE_RN_2414_0;
wire FE_RN_2417_0;
wire FE_RN_2418_0;
wire FE_RN_2419_0;
wire FE_RN_241_0;
wire FE_RN_2420_0;
wire FE_RN_2421_0;
wire FE_RN_2422_0;
wire FE_RN_2423_0;
wire FE_RN_2425_0;
wire FE_RN_2426_0;
wire FE_RN_2428_0;
wire FE_RN_2429_0;
wire FE_RN_242_0;
wire FE_RN_2430_0;
wire FE_RN_2431_0;
wire FE_RN_2432_0;
wire FE_RN_2433_0;
wire FE_RN_2434_0;
wire TIMEBOOST_net_508;
wire TIMEBOOST_net_309;
wire FE_RN_2437_0;
wire FE_RN_2438_0;
wire FE_RN_2439_0;
wire FE_RN_2440_0;
wire FE_RN_2441_0;
wire FE_RN_2442_0;
wire FE_RN_2443_0;
wire FE_RN_2444_0;
wire FE_RN_2445_0;
wire FE_RN_2446_0;
wire FE_RN_2448_0;
wire FE_RN_2449_0;
wire FE_RN_2450_0;
wire FE_RN_2452_0;
wire FE_RN_2453_0;
wire FE_RN_2454_0;
wire FE_RN_2455_0;
wire FE_RN_2456_0;
wire TIMEBOOST_net_2111;
wire FE_RN_2458_0;
wire FE_RN_2459_0;
wire FE_RN_245_0;
wire FE_RN_2460_0;
wire FE_RN_2461_0;
wire FE_RN_2462_0;
wire FE_RN_2463_0;
wire FE_RN_2464_0;
wire TIMEBOOST_net_2855;
wire FE_RN_2466_0;
wire FE_RN_2467_0;
wire FE_RN_2468_0;
wire FE_RN_2469_0;
wire FE_RN_2470_0;
wire FE_RN_2471_0;
wire FE_RN_2472_0;
wire TIMEBOOST_net_516;
wire FE_RN_2477_0;
wire FE_RN_2478_0;
wire FE_RN_2479_0;
wire FE_RN_2480_0;
wire TIMEBOOST_net_2800;
wire FE_RN_2485_0;
wire TIMEBOOST_net_595;
wire FE_RN_2487_0;
wire FE_RN_2488_0;
wire FE_RN_2489_0;
wire FE_RN_248_0;
wire FE_RN_2490_0;
wire FE_RN_2491_0;
wire FE_RN_2492_0;
wire FE_RN_2493_0;
wire FE_RN_2494_0;
wire FE_RN_2495_0;
wire FE_RN_2496_0;
wire FE_RN_2497_0;
wire FE_RN_2498_0;
wire FE_RN_2499_0;
wire FE_RN_249_0;
wire TIMEBOOST_net_2328;
wire FE_RN_2501_0;
wire FE_RN_2502_0;
wire FE_RN_2503_0;
wire FE_RN_2504_0;
wire FE_RN_2505_0;
wire FE_RN_2506_0;
wire FE_RN_2508_0;
wire FE_RN_2509_0;
wire FE_RN_2512_0;
wire TIMEBOOST_net_1459;
wire FE_RN_2514_0;
wire FE_RN_2515_0;
wire FE_RN_2516_0;
wire FE_RN_2517_0;
wire FE_RN_2518_0;
wire FE_RN_2519_0;
wire TIMEBOOST_net_1847;
wire FE_RN_2520_0;
wire FE_RN_2521_0;
wire FE_RN_2522_0;
wire FE_RN_2523_0;
wire FE_RN_2524_0;
wire FE_RN_2526_0;
wire FE_RN_2527_0;
wire FE_RN_2528_0;
wire FE_RN_2529_0;
wire FE_RN_252_0;
wire FE_RN_2530_0;
wire TIMEBOOST_net_838;
wire FE_RN_2532_0;
wire FE_RN_2534_0;
wire FE_RN_2535_0;
wire FE_RN_2536_0;
wire FE_RN_2537_0;
wire TIMEBOOST_net_2205;
wire FE_RN_2539_0;
wire FE_RN_253_0;
wire TIMEBOOST_net_785;
wire FE_RN_2541_0;
wire FE_RN_2542_0;
wire TIMEBOOST_net_873;
wire FE_RN_2544_0;
wire FE_RN_2546_0;
wire FE_RN_2548_0;
wire TIMEBOOST_net_2291;
wire TIMEBOOST_net_1594;
wire FE_RN_2550_0;
wire FE_RN_2551_0;
wire FE_RN_2552_0;
wire FE_RN_2553_0;
wire FE_RN_2554_0;
wire FE_RN_2555_0;
wire FE_RN_2556_0;
wire FE_RN_2557_0;
wire TIMEBOOST_net_787;
wire FE_RN_2559_0;
wire FE_RN_255_0;
wire FE_RN_2560_0;
wire TIMEBOOST_net_1008;
wire FE_RN_2562_0;
wire FE_RN_2563_0;
wire FE_RN_2564_0;
wire TIMEBOOST_net_987;
wire FE_RN_2566_0;
wire FE_RN_2567_0;
wire FE_RN_2568_0;
wire FE_RN_2569_0;
wire FE_RN_256_0;
wire TIMEBOOST_net_1603;
wire FE_RN_2571_0;
wire FE_RN_2574_0;
wire FE_RN_2575_0;
wire FE_RN_2576_0;
wire FE_RN_2577_0;
wire FE_RN_2578_0;
wire FE_RN_2579_0;
wire FE_RN_257_0;
wire FE_RN_2580_0;
wire FE_RN_2581_0;
wire FE_RN_2582_0;
wire FE_RN_2583_0;
wire FE_RN_2584_0;
wire TIMEBOOST_net_1040;
wire FE_RN_2586_0;
wire FE_RN_2587_0;
wire FE_RN_2588_0;
wire FE_RN_2589_0;
wire TIMEBOOST_net_1838;
wire FE_RN_2590_0;
wire FE_RN_2591_0;
wire FE_RN_2592_0;
wire FE_RN_2595_0;
wire FE_RN_2596_0;
wire FE_RN_2597_0;
wire FE_RN_2598_0;
wire FE_RN_2599_0;
wire FE_RN_259_0;
wire FE_RN_2600_0;
wire FE_RN_2601_0;
wire FE_RN_2603_0;
wire FE_RN_2604_0;
wire FE_RN_2605_0;
wire FE_RN_2606_0;
wire FE_RN_2607_0;
wire FE_RN_2608_0;
wire FE_RN_2609_0;
wire FE_RN_260_0;
wire FE_RN_2610_0;
wire FE_RN_2611_0;
wire FE_RN_2612_0;
wire FE_RN_2613_0;
wire FE_RN_2614_0;
wire FE_RN_2615_0;
wire FE_RN_2616_0;
wire FE_RN_2617_0;
wire FE_RN_2618_0;
wire FE_RN_2619_0;
wire FE_RN_2620_0;
wire FE_RN_2621_0;
wire FE_RN_2622_0;
wire FE_RN_2623_0;
wire FE_RN_2624_0;
wire FE_RN_2625_0;
wire FE_RN_2626_0;
wire FE_RN_2627_0;
wire FE_RN_2628_0;
wire FE_RN_2629_0;
wire FE_RN_2630_0;
wire FE_RN_2631_0;
wire FE_RN_2632_0;
wire FE_RN_2633_0;
wire FE_RN_2634_0;
wire FE_RN_2635_0;
wire FE_RN_2636_0;
wire FE_RN_2637_0;
wire FE_RN_2638_0;
wire FE_RN_2639_0;
wire FE_RN_263_0;
wire FE_RN_2640_0;
wire FE_RN_2641_0;
wire FE_RN_2642_0;
wire FE_RN_2643_0;
wire FE_RN_2644_0;
wire FE_RN_2645_0;
wire FE_RN_2646_0;
wire FE_RN_2648_0;
wire FE_RN_2649_0;
wire FE_RN_264_0;
wire TIMEBOOST_net_1308;
wire FE_RN_2652_0;
wire FE_RN_2653_0;
wire FE_RN_2654_0;
wire FE_RN_2655_0;
wire FE_RN_2656_0;
wire FE_RN_2657_0;
wire FE_RN_2658_0;
wire FE_RN_2659_0;
wire FE_RN_265_0;
wire FE_RN_2660_0;
wire FE_RN_2661_0;
wire FE_RN_2662_0;
wire FE_RN_2663_0;
wire FE_RN_2664_0;
wire FE_RN_2665_0;
wire FE_RN_2666_0;
wire TIMEBOOST_net_603;
wire FE_RN_2668_0;
wire FE_RN_2669_0;
wire FE_RN_266_0;
wire FE_RN_2670_0;
wire TIMEBOOST_net_675;
wire FE_RN_2672_0;
wire FE_RN_2673_0;
wire FE_RN_2674_0;
wire FE_RN_2675_0;
wire FE_RN_2676_0;
wire FE_RN_2679_0;
wire FE_RN_267_0;
wire FE_RN_2680_0;
wire FE_RN_2681_0;
wire FE_RN_2682_0;
wire FE_RN_2683_0;
wire TIMEBOOST_net_722;
wire FE_RN_2685_0;
wire FE_RN_2686_0;
wire FE_RN_2687_0;
wire FE_RN_2688_0;
wire FE_RN_2689_0;
wire FE_RN_268_0;
wire FE_RN_2693_0;
wire FE_RN_2694_0;
wire FE_RN_2695_0;
wire TIMEBOOST_net_705;
wire FE_RN_2697_0;
wire FE_RN_2698_0;
wire FE_RN_2699_0;
wire FE_RN_269_0;
wire FE_RN_2700_0;
wire FE_RN_2701_0;
wire FE_RN_2702_0;
wire FE_RN_2703_0;
wire FE_RN_2704_0;
wire TIMEBOOST_net_2598;
wire FE_RN_2706_0;
wire FE_RN_2708_0;
wire FE_RN_2709_0;
wire FE_RN_270_0;
wire FE_RN_2710_0;
wire FE_RN_2711_0;
wire FE_RN_2712_0;
wire FE_RN_2713_0;
wire FE_RN_2714_0;
wire FE_RN_2715_0;
wire FE_RN_2716_0;
wire FE_RN_2717_0;
wire FE_RN_2718_0;
wire FE_RN_2719_0;
wire FE_RN_271_0;
wire TIMEBOOST_net_2188;
wire FE_RN_2721_0;
wire TIMEBOOST_net_104;
wire FE_RN_2725_0;
wire FE_RN_2726_0;
wire FE_RN_2727_0;
wire FE_RN_2728_0;
wire FE_RN_2729_0;
wire TIMEBOOST_net_2525;
wire FE_RN_2730_0;
wire FE_RN_2731_0;
wire FE_RN_2732_0;
wire FE_RN_2733_0;
wire FE_RN_2734_0;
wire TIMEBOOST_net_2184;
wire FE_RN_2736_0;
wire FE_RN_2737_0;
wire FE_RN_2738_0;
wire FE_RN_2739_0;
wire FE_RN_273_0;
wire FE_RN_2740_0;
wire FE_RN_2741_0;
wire FE_RN_2742_0;
wire FE_RN_2743_0;
wire FE_RN_2744_0;
wire FE_RN_2745_0;
wire FE_RN_2746_0;
wire FE_RN_2747_0;
wire FE_RN_2748_0;
wire FE_RN_2749_0;
wire FE_RN_2750_0;
wire FE_RN_2751_0;
wire FE_RN_2752_0;
wire FE_RN_2753_0;
wire FE_RN_2754_0;
wire FE_RN_2758_0;
wire FE_RN_2759_0;
wire TIMEBOOST_net_1852;
wire FE_RN_2760_0;
wire FE_RN_2761_0;
wire FE_RN_2762_0;
wire FE_RN_2763_0;
wire FE_RN_2764_0;
wire FE_RN_2765_0;
wire FE_RN_2766_0;
wire FE_RN_2767_0;
wire FE_RN_2768_0;
wire FE_RN_2769_0;
wire FE_RN_276_0;
wire FE_RN_2770_0;
wire FE_RN_2771_0;
wire FE_RN_2772_0;
wire FE_RN_2773_0;
wire FE_RN_2774_0;
wire FE_RN_2775_0;
wire FE_RN_2776_0;
wire FE_RN_2777_0;
wire FE_RN_2778_0;
wire FE_RN_2779_0;
wire FE_RN_277_0;
wire FE_RN_2780_0;
wire TIMEBOOST_net_1399;
wire FE_RN_2782_0;
wire FE_RN_2783_0;
wire FE_RN_2784_0;
wire FE_RN_2785_0;
wire FE_RN_2786_0;
wire FE_RN_2787_0;
wire FE_RN_2788_0;
wire FE_RN_2789_0;
wire FE_RN_278_0;
wire FE_RN_2790_0;
wire FE_RN_2791_0;
wire FE_RN_2792_0;
wire FE_RN_2793_0;
wire FE_RN_2794_0;
wire FE_RN_2795_0;
wire FE_RN_2796_0;
wire FE_RN_2797_0;
wire FE_RN_2798_0;
wire FE_RN_2799_0;
wire FE_RN_27_0;
wire FE_RN_2800_0;
wire FE_RN_2801_0;
wire FE_RN_2811_0;
wire TIMEBOOST_net_2323;
wire FE_RN_2813_0;
wire TIMEBOOST_net_15;
wire TIMEBOOST_net_1424;
wire FE_RN_2816_0;
wire FE_RN_2817_0;
wire FE_RN_2818_0;
wire FE_RN_2819_0;
wire TIMEBOOST_net_1749;
wire FE_RN_2821_0;
wire FE_RN_2822_0;
wire FE_RN_2823_0;
wire FE_RN_2824_0;
wire FE_RN_2825_0;
wire FE_RN_2826_0;
wire TIMEBOOST_net_2314;
wire FE_RN_2828_0;
wire FE_RN_2829_0;
wire FE_RN_282_0;
wire FE_RN_2830_0;
wire FE_RN_2831_0;
wire FE_RN_2832_0;
wire FE_RN_2833_0;
wire TIMEBOOST_net_1017;
wire FE_RN_2835_0;
wire FE_RN_2836_0;
wire FE_RN_2837_0;
wire FE_RN_2838_0;
wire FE_RN_2839_0;
wire FE_RN_283_0;
wire FE_RN_2840_0;
wire FE_RN_2841_0;
wire FE_RN_2842_0;
wire FE_RN_2843_0;
wire FE_RN_2844_0;
wire FE_RN_2845_0;
wire FE_RN_2846_0;
wire TIMEBOOST_net_1585;
wire FE_RN_2848_0;
wire FE_RN_2849_0;
wire FE_RN_284_0;
wire FE_RN_2850_0;
wire FE_RN_2851_0;
wire FE_RN_2852_0;
wire FE_RN_2853_0;
wire FE_RN_2854_0;
wire FE_RN_2855_0;
wire FE_RN_2856_0;
wire FE_RN_2857_0;
wire FE_RN_2858_0;
wire FE_RN_2859_0;
wire FE_RN_285_0;
wire FE_RN_2861_0;
wire FE_RN_2862_0;
wire FE_RN_2863_0;
wire FE_RN_2864_0;
wire FE_RN_2865_0;
wire FE_RN_2866_0;
wire FE_RN_2867_0;
wire FE_RN_2868_0;
wire FE_RN_2869_0;
wire FE_RN_286_0;
wire FE_RN_2870_0;
wire FE_RN_2871_0;
wire FE_RN_2872_0;
wire FE_RN_2873_0;
wire FE_RN_2874_0;
wire FE_RN_2875_0;
wire FE_RN_2876_0;
wire FE_RN_2877_0;
wire FE_RN_2878_0;
wire FE_RN_2879_0;
wire TIMEBOOST_net_2796;
wire FE_RN_2880_0;
wire TIMEBOOST_net_1438;
wire FE_RN_2882_0;
wire FE_RN_2883_0;
wire FE_RN_2884_0;
wire FE_RN_2885_0;
wire FE_RN_2886_0;
wire FE_RN_2887_0;
wire TIMEBOOST_net_706;
wire FE_RN_288_0;
wire FE_RN_28_0;
wire TIMEBOOST_net_1765;
wire TIMEBOOST_net_175;
wire FE_RN_294_0;
wire FE_RN_295_0;
wire TIMEBOOST_net_2423;
wire TIMEBOOST_net_1056;
wire FE_RN_298_0;
wire FE_RN_299_0;
wire TIMEBOOST_net_1456;
wire FE_RN_303_0;
wire FE_RN_304_0;
wire FE_RN_306_0;
wire FE_RN_307_0;
wire FE_RN_308_0;
wire TIMEBOOST_net_2183;
wire FE_RN_30_0;
wire FE_RN_310_0;
wire FE_RN_311_0;
wire TIMEBOOST_net_2215;
wire FE_RN_314_0;
wire FE_RN_315_0;
wire TIMEBOOST_net_968;
wire FE_RN_317_0;
wire TIMEBOOST_net_1866;
wire FE_RN_319_0;
wire FE_RN_31_0;
wire FE_RN_320_0;
wire TIMEBOOST_net_1647;
wire FE_RN_323_0;
wire FE_RN_324_0;
wire FE_RN_325_0;
wire FE_RN_326_0;
wire FE_RN_327_0;
wire FE_RN_328_0;
wire FE_RN_329_0;
wire FE_RN_32_0;
wire FE_RN_330_0;
wire FE_RN_331_0;
wire TIMEBOOST_net_545;
wire FE_RN_336_0;
wire FE_RN_337_0;
wire FE_RN_338_0;
wire TIMEBOOST_net_1406;
wire TIMEBOOST_net_2894;
wire FE_RN_340_0;
wire FE_RN_341_0;
wire TIMEBOOST_net_2120;
wire FE_RN_344_0;
wire FE_RN_345_0;
wire TIMEBOOST_net_1416;
wire FE_RN_347_0;
wire FE_RN_348_0;
wire FE_RN_349_0;
wire TIMEBOOST_net_2361;
wire FE_RN_354_0;
wire FE_RN_355_0;
wire TIMEBOOST_net_1766;
wire FE_RN_35_0;
wire FE_RN_360_0;
wire FE_RN_361_0;
wire TIMEBOOST_net_840;
wire FE_RN_363_0;
wire FE_RN_364_0;
wire FE_RN_365_0;
wire FE_RN_366_0;
wire FE_RN_367_0;
wire FE_RN_368_0;
wire FE_RN_369_0;
wire TIMEBOOST_net_2125;
wire FE_RN_371_0;
wire FE_RN_372_0;
wire TIMEBOOST_net_2123;
wire FE_RN_374_0;
wire FE_RN_375_0;
wire FE_RN_382_0;
wire FE_RN_383_0;
wire FE_RN_386_0;
wire FE_RN_387_0;
wire FE_RN_388_0;
wire FE_RN_389_0;
wire FE_RN_391_0;
wire FE_RN_392_0;
wire FE_RN_394_0;
wire FE_RN_395_0;
wire TIMEBOOST_net_1820;
wire TIMEBOOST_net_850;
wire FE_RN_398_0;
wire FE_RN_399_0;
wire FE_RN_3_0;
wire FE_RN_400_0;
wire FE_RN_401_0;
wire FE_RN_402_0;
wire FE_RN_403_0;
wire TIMEBOOST_net_1715;
wire FE_RN_405_0;
wire TIMEBOOST_net_1483;
wire FE_RN_424_0;
wire TIMEBOOST_net_2806;
wire FE_RN_426_0;
wire FE_RN_428_0;
wire FE_RN_429_0;
wire FE_RN_42_0;
wire FE_RN_430_0;
wire TIMEBOOST_net_1123;
wire FE_RN_437_0;
wire FE_RN_438_0;
wire FE_RN_439_0;
wire FE_RN_43_0;
wire FE_RN_440_0;
wire FE_RN_442_0;
wire FE_RN_443_0;
wire FE_RN_444_0;
wire FE_RN_445_0;
wire FE_RN_448_0;
wire FE_RN_449_0;
wire TIMEBOOST_net_2900;
wire FE_RN_450_0;
wire FE_RN_453_0;
wire FE_RN_456_0;
wire FE_RN_457_0;
wire FE_RN_459_0;
wire FE_RN_45_0;
wire FE_RN_460_0;
wire FE_RN_462_0;
wire TIMEBOOST_net_863;
wire FE_RN_464_0;
wire FE_RN_466_0;
wire TIMEBOOST_net_114;
wire FE_RN_469_0;
wire FE_RN_46_0;
wire FE_RN_471_0;
wire FE_RN_474_0;
wire FE_RN_476_0;
wire FE_RN_479_0;
wire FE_RN_47_0;
wire FE_RN_480_0;
wire FE_RN_481_0;
wire FE_RN_482_0;
wire FE_RN_485_0;
wire FE_RN_486_0;
wire FE_RN_495_0;
wire FE_RN_496_0;
wire FE_RN_497_0;
wire FE_RN_4_0;
wire FE_RN_510_0;
wire FE_RN_516_0;
wire FE_RN_517_0;
wire FE_RN_519_0;
wire FE_RN_51_0;
wire FE_RN_522_0;
wire FE_RN_525_0;
wire FE_RN_526_0;
wire FE_RN_527_0;
wire FE_RN_528_0;
wire FE_RN_529_0;
wire FE_RN_52_0;
wire FE_RN_530_0;
wire FE_RN_532_0;
wire FE_RN_533_0;
wire FE_RN_535_0;
wire FE_RN_536_0;
wire FE_RN_537_0;
wire FE_RN_538_0;
wire FE_RN_539_0;
wire FE_RN_53_0;
wire FE_RN_541_0;
wire FE_RN_546_0;
wire FE_RN_547_0;
wire FE_RN_552_0;
wire FE_RN_553_0;
wire FE_RN_555_0;
wire FE_RN_557_0;
wire TIMEBOOST_net_1797;
wire FE_RN_559_0;
wire FE_RN_560_0;
wire FE_RN_563_0;
wire FE_RN_564_0;
wire FE_RN_565_0;
wire FE_RN_566_0;
wire FE_RN_567_0;
wire FE_RN_568_0;
wire FE_RN_569_0;
wire FE_RN_570_0;
wire FE_RN_572_0;
wire FE_RN_574_0;
wire TIMEBOOST_net_1255;
wire FE_RN_578_0;
wire FE_RN_579_0;
wire FE_RN_57_0;
wire TIMEBOOST_net_2274;
wire FE_RN_586_0;
wire FE_RN_588_0;
wire FE_RN_58_0;
wire FE_RN_591_0;
wire FE_RN_592_0;
wire FE_RN_595_0;
wire FE_RN_59_0;
wire FE_RN_5_0;
wire TIMEBOOST_net_2717;
wire FE_RN_604_0;
wire FE_RN_606_0;
wire FE_RN_60_0;
wire TIMEBOOST_net_2735;
wire FE_RN_611_0;
wire FE_RN_612_0;
wire FE_RN_614_0;
wire FE_RN_617_0;
wire FE_RN_618_0;
wire FE_RN_61_0;
wire FE_RN_620_0;
wire FE_RN_621_0;
wire FE_RN_622_0;
wire FE_RN_624_0;
wire FE_RN_625_0;
wire FE_RN_627_0;
wire FE_RN_628_0;
wire FE_RN_629_0;
wire FE_RN_62_0;
wire FE_RN_630_0;
wire FE_RN_631_0;
wire FE_RN_632_0;
wire FE_RN_633_0;
wire FE_RN_634_0;
wire FE_RN_635_0;
wire FE_RN_636_0;
wire FE_RN_637_0;
wire TIMEBOOST_net_16;
wire FE_RN_639_0;
wire FE_RN_63_0;
wire FE_RN_640_0;
wire FE_RN_641_0;
wire FE_RN_643_0;
wire FE_RN_644_0;
wire FE_RN_645_0;
wire FE_RN_646_0;
wire TIMEBOOST_net_2913;
wire FE_RN_648_0;
wire TIMEBOOST_net_955;
wire FE_RN_64_0;
wire FE_RN_650_0;
wire TIMEBOOST_net_58;
wire FE_RN_656_0;
wire FE_RN_657_0;
wire FE_RN_658_0;
wire FE_RN_659_0;
wire FE_RN_65_0;
wire FE_RN_660_0;
wire FE_RN_663_0;
wire FE_RN_664_0;
wire FE_RN_665_0;
wire TIMEBOOST_net_1170;
wire TIMEBOOST_net_335;
wire FE_RN_668_0;
wire FE_RN_669_0;
wire TIMEBOOST_net_1473;
wire FE_RN_670_0;
wire TIMEBOOST_net_2077;
wire FE_RN_672_0;
wire FE_RN_673_0;
wire FE_RN_674_0;
wire TIMEBOOST_net_2507;
wire FE_RN_676_0;
wire FE_RN_677_0;
wire FE_RN_678_0;
wire TIMEBOOST_net_359;
wire FE_RN_67_0;
wire FE_RN_681_0;
wire FE_RN_682_0;
wire FE_RN_683_0;
wire FE_RN_686_0;
wire FE_RN_687_0;
wire FE_RN_688_0;
wire FE_RN_689_0;
wire FE_RN_68_0;
wire FE_RN_690_0;
wire TIMEBOOST_net_2837;
wire FE_RN_692_0;
wire FE_RN_693_0;
wire FE_RN_694_0;
wire FE_RN_695_0;
wire FE_RN_696_0;
wire FE_RN_697_0;
wire TIMEBOOST_net_2375;
wire FE_RN_699_0;
wire FE_RN_69_0;
wire FE_RN_6_0;
wire TIMEBOOST_net_241;
wire FE_RN_701_0;
wire FE_RN_702_0;
wire TIMEBOOST_net_356;
wire FE_RN_704_0;
wire TIMEBOOST_net_1094;
wire FE_RN_706_0;
wire FE_RN_707_0;
wire FE_RN_708_0;
wire FE_RN_709_0;
wire TIMEBOOST_net_1854;
wire FE_RN_710_0;
wire FE_RN_71_0;
wire FE_RN_724_0;
wire FE_RN_725_0;
wire TIMEBOOST_net_6;
wire FE_RN_727_0;
wire FE_RN_728_0;
wire TIMEBOOST_net_2780;
wire FE_RN_72_0;
wire TIMEBOOST_net_2784;
wire FE_RN_731_0;
wire FE_RN_732_0;
wire TIMEBOOST_net_806;
wire FE_RN_734_0;
wire FE_RN_735_0;
wire FE_RN_736_0;
wire FE_RN_737_0;
wire FE_RN_738_0;
wire FE_RN_739_0;
wire TIMEBOOST_net_928;
wire FE_RN_741_0;
wire FE_RN_742_0;
wire FE_RN_743_0;
wire TIMEBOOST_net_939;
wire TIMEBOOST_net_852;
wire FE_RN_747_0;
wire FE_RN_748_0;
wire FE_RN_749_0;
wire FE_RN_74_0;
wire FE_RN_751_0;
wire FE_RN_752_0;
wire FE_RN_753_0;
wire FE_RN_754_0;
wire TIMEBOOST_net_158;
wire FE_RN_757_0;
wire TIMEBOOST_net_187;
wire FE_RN_759_0;
wire FE_RN_75_0;
wire FE_RN_760_0;
wire FE_RN_761_0;
wire FE_RN_762_0;
wire TIMEBOOST_net_2404;
wire FE_RN_764_0;
wire FE_RN_765_0;
wire TIMEBOOST_net_776;
wire FE_RN_767_0;
wire FE_RN_768_0;
wire TIMEBOOST_net_41;
wire FE_RN_76_0;
wire FE_RN_770_0;
wire FE_RN_773_0;
wire TIMEBOOST_net_2822;
wire FE_RN_775_0;
wire FE_RN_776_0;
wire TIMEBOOST_net_933;
wire FE_RN_778_0;
wire TIMEBOOST_net_1038;
wire FE_RN_77_0;
wire FE_RN_780_0;
wire FE_RN_781_0;
wire FE_RN_782_0;
wire FE_RN_783_0;
wire TIMEBOOST_net_1829;
wire FE_RN_785_0;
wire FE_RN_786_0;
wire FE_RN_787_0;
wire FE_RN_788_0;
wire FE_RN_789_0;
wire FE_RN_78_0;
wire FE_RN_790_0;
wire FE_RN_791_0;
wire FE_RN_792_0;
wire FE_RN_793_0;
wire FE_RN_794_0;
wire FE_RN_795_0;
wire FE_RN_796_0;
wire FE_RN_797_0;
wire TIMEBOOST_net_2347;
wire TIMEBOOST_net_1843;
wire FE_RN_79_0;
wire FE_RN_7_0;
wire FE_RN_800_0;
wire TIMEBOOST_net_1711;
wire FE_RN_80_0;
wire FE_RN_811_0;
wire FE_RN_812_0;
wire FE_RN_813_0;
wire FE_RN_816_0;
wire FE_RN_818_0;
wire TIMEBOOST_net_1830;
wire FE_RN_821_0;
wire TIMEBOOST_net_2109;
wire FE_RN_824_0;
wire TIMEBOOST_net_1554;
wire FE_RN_826_0;
wire FE_RN_827_0;
wire FE_RN_828_0;
wire FE_RN_829_0;
wire FE_RN_82_0;
wire FE_RN_832_0;
wire FE_RN_833_0;
wire TIMEBOOST_net_1441;
wire FE_RN_835_0;
wire FE_RN_837_0;
wire TIMEBOOST_net_2311;
wire FE_RN_839_0;
wire FE_RN_83_0;
wire TIMEBOOST_net_956;
wire FE_RN_841_0;
wire FE_RN_842_0;
wire FE_RN_843_0;
wire FE_RN_844_0;
wire FE_RN_845_0;
wire FE_RN_846_0;
wire FE_RN_847_0;
wire FE_RN_849_0;
wire TIMEBOOST_net_1900;
wire FE_RN_850_0;
wire FE_RN_851_0;
wire FE_RN_852_0;
wire TIMEBOOST_net_2382;
wire FE_RN_854_0;
wire FE_RN_855_0;
wire FE_RN_856_0;
wire FE_RN_857_0;
wire FE_RN_858_0;
wire FE_RN_859_0;
wire FE_RN_85_0;
wire FE_RN_860_0;
wire TIMEBOOST_net_184;
wire TIMEBOOST_net_2820;
wire TIMEBOOST_net_2379;
wire FE_RN_864_0;
wire FE_RN_865_0;
wire FE_RN_866_0;
wire FE_RN_867_0;
wire FE_RN_86_0;
wire FE_RN_871_0;
wire FE_RN_872_0;
wire FE_RN_873_0;
wire FE_RN_874_0;
wire FE_RN_875_0;
wire FE_RN_876_0;
wire FE_RN_877_0;
wire FE_RN_878_0;
wire FE_RN_879_0;
wire FE_RN_87_0;
wire FE_RN_880_0;
wire FE_RN_881_0;
wire FE_RN_882_0;
wire FE_RN_885_0;
wire FE_RN_886_0;
wire FE_RN_887_0;
wire FE_RN_888_0;
wire FE_RN_889_0;
wire FE_RN_88_0;
wire TIMEBOOST_net_285;
wire FE_RN_891_0;
wire TIMEBOOST_net_1079;
wire FE_RN_893_0;
wire FE_RN_894_0;
wire FE_RN_895_0;
wire FE_RN_896_0;
wire FE_RN_897_0;
wire TIMEBOOST_net_1926;
wire FE_RN_899_0;
wire FE_RN_89_0;
wire TIMEBOOST_net_869;
wire TIMEBOOST_net_1157;
wire FE_RN_901_0;
wire FE_RN_902_0;
wire TIMEBOOST_net_819;
wire FE_RN_904_0;
wire FE_RN_905_0;
wire FE_RN_909_0;
wire FE_RN_90_0;
wire FE_RN_911_0;
wire FE_RN_912_0;
wire FE_RN_916_0;
wire FE_RN_917_0;
wire FE_RN_918_0;
wire FE_RN_919_0;
wire FE_RN_920_0;
wire FE_RN_921_0;
wire FE_RN_922_0;
wire FE_RN_923_0;
wire TIMEBOOST_net_2108;
wire FE_RN_925_0;
wire FE_RN_926_0;
wire FE_RN_927_0;
wire FE_RN_928_0;
wire FE_RN_929_0;
wire TIMEBOOST_net_1087;
wire FE_RN_930_0;
wire FE_RN_931_0;
wire TIMEBOOST_net_2804;
wire FE_RN_933_0;
wire TIMEBOOST_net_1648;
wire TIMEBOOST_net_2773;
wire FE_RN_938_0;
wire FE_RN_939_0;
wire FE_RN_93_0;
wire FE_RN_940_0;
wire FE_RN_941_0;
wire FE_RN_942_0;
wire FE_RN_943_0;
wire TIMEBOOST_net_1570;
wire FE_RN_945_0;
wire FE_RN_946_0;
wire TIMEBOOST_net_2517;
wire FE_RN_948_0;
wire FE_RN_94_0;
wire FE_RN_952_0;
wire TIMEBOOST_net_998;
wire FE_RN_954_0;
wire FE_RN_959_0;
wire TIMEBOOST_net_1703;
wire FE_RN_960_0;
wire FE_RN_961_0;
wire TIMEBOOST_net_2022;
wire FE_RN_964_0;
wire FE_RN_966_0;
wire FE_RN_967_0;
wire FE_RN_968_0;
wire FE_RN_969_0;
wire TIMEBOOST_net_2807;
wire TIMEBOOST_net_844;
wire TIMEBOOST_net_297;
wire FE_RN_974_0;
wire FE_RN_975_0;
wire FE_RN_976_0;
wire FE_RN_977_0;
wire FE_RN_978_0;
wire TIMEBOOST_net_2231;
wire FE_RN_980_0;
wire FE_RN_981_0;
wire FE_RN_982_0;
wire TIMEBOOST_net_1159;
wire FE_RN_984_0;
wire FE_RN_985_0;
wire FE_RN_986_0;
wire FE_RN_987_0;
wire FE_RN_988_0;
wire FE_RN_989_0;
wire TIMEBOOST_net_1377;
wire FE_RN_990_0;
wire FE_RN_991_0;
wire FE_RN_992_0;
wire FE_RN_993_0;
wire FE_RN_994_0;
wire FE_RN_995_0;
wire FE_RN_996_0;
wire FE_RN_997_0;
wire FE_RN_998_0;
wire cordic_combinational_sub_ln23_0_unr12_z_0_;
wire cordic_combinational_sub_ln23_0_unr16_z_0_;
wire cordic_combinational_sub_ln23_0_unr20_z_0_;
wire delay_add_ln22_unr11_stage5_stallmux_q_0_;
wire delay_add_ln22_unr11_stage5_stallmux_q_10_;
wire delay_add_ln22_unr11_stage5_stallmux_q_11_;
wire delay_add_ln22_unr11_stage5_stallmux_q_12_;
wire delay_add_ln22_unr11_stage5_stallmux_q_13_;
wire delay_add_ln22_unr11_stage5_stallmux_q_14_;
wire delay_add_ln22_unr11_stage5_stallmux_q_15_;
wire delay_add_ln22_unr11_stage5_stallmux_q_16_;
wire delay_add_ln22_unr11_stage5_stallmux_q_17_;
wire delay_add_ln22_unr11_stage5_stallmux_q_18_;
wire delay_add_ln22_unr11_stage5_stallmux_q_19_;
wire delay_add_ln22_unr11_stage5_stallmux_q_1_;
wire delay_add_ln22_unr11_stage5_stallmux_q_20_;
wire delay_add_ln22_unr11_stage5_stallmux_q_21_;
wire delay_add_ln22_unr11_stage5_stallmux_q_22_;
wire delay_add_ln22_unr11_stage5_stallmux_q_23_;
wire delay_add_ln22_unr11_stage5_stallmux_q_24_;
wire delay_add_ln22_unr11_stage5_stallmux_q_25_;
wire delay_add_ln22_unr11_stage5_stallmux_q_26_;
wire delay_add_ln22_unr11_stage5_stallmux_q_27_;
wire delay_add_ln22_unr11_stage5_stallmux_q_28_;
wire delay_add_ln22_unr11_stage5_stallmux_q_29_;
wire delay_add_ln22_unr11_stage5_stallmux_q_2_;
wire delay_add_ln22_unr11_stage5_stallmux_q_30_;
wire delay_add_ln22_unr11_stage5_stallmux_q_31_;
wire delay_add_ln22_unr11_stage5_stallmux_q_3_;
wire delay_add_ln22_unr11_stage5_stallmux_q_4_;
wire delay_add_ln22_unr11_stage5_stallmux_q_5_;
wire delay_add_ln22_unr11_stage5_stallmux_q_6_;
wire delay_add_ln22_unr11_stage5_stallmux_q_7_;
wire delay_add_ln22_unr11_stage5_stallmux_q_8_;
wire delay_add_ln22_unr11_stage5_stallmux_q_9_;
wire delay_add_ln22_unr14_stage6_stallmux_q_0_;
wire delay_add_ln22_unr14_stage6_stallmux_q_10_;
wire delay_add_ln22_unr14_stage6_stallmux_q_11_;
wire delay_add_ln22_unr14_stage6_stallmux_q_12_;
wire delay_add_ln22_unr14_stage6_stallmux_q_13_;
wire delay_add_ln22_unr14_stage6_stallmux_q_14_;
wire delay_add_ln22_unr14_stage6_stallmux_q_15_;
wire delay_add_ln22_unr14_stage6_stallmux_q_16_;
wire delay_add_ln22_unr14_stage6_stallmux_q_17_;
wire delay_add_ln22_unr14_stage6_stallmux_q_18_;
wire delay_add_ln22_unr14_stage6_stallmux_q_19_;
wire delay_add_ln22_unr14_stage6_stallmux_q_1_;
wire delay_add_ln22_unr14_stage6_stallmux_q_20_;
wire delay_add_ln22_unr14_stage6_stallmux_q_21_;
wire delay_add_ln22_unr14_stage6_stallmux_q_22_;
wire delay_add_ln22_unr14_stage6_stallmux_q_23_;
wire delay_add_ln22_unr14_stage6_stallmux_q_24_;
wire delay_add_ln22_unr14_stage6_stallmux_q_25_;
wire delay_add_ln22_unr14_stage6_stallmux_q_26_;
wire delay_add_ln22_unr14_stage6_stallmux_q_27_;
wire delay_add_ln22_unr14_stage6_stallmux_q_28_;
wire delay_add_ln22_unr14_stage6_stallmux_q_29_;
wire delay_add_ln22_unr14_stage6_stallmux_q_2_;
wire delay_add_ln22_unr14_stage6_stallmux_q_30_;
wire delay_add_ln22_unr14_stage6_stallmux_q_31_;
wire delay_add_ln22_unr14_stage6_stallmux_q_3_;
wire delay_add_ln22_unr14_stage6_stallmux_q_4_;
wire delay_add_ln22_unr14_stage6_stallmux_q_5_;
wire delay_add_ln22_unr14_stage6_stallmux_q_6_;
wire delay_add_ln22_unr14_stage6_stallmux_q_7_;
wire delay_add_ln22_unr14_stage6_stallmux_q_8_;
wire delay_add_ln22_unr14_stage6_stallmux_q_9_;
wire delay_add_ln22_unr17_stage7_stallmux_q_0_;
wire delay_add_ln22_unr17_stage7_stallmux_q_10_;
wire delay_add_ln22_unr17_stage7_stallmux_q_11_;
wire delay_add_ln22_unr17_stage7_stallmux_q_12_;
wire delay_add_ln22_unr17_stage7_stallmux_q_13_;
wire delay_add_ln22_unr17_stage7_stallmux_q_14_;
wire delay_add_ln22_unr17_stage7_stallmux_q_15_;
wire delay_add_ln22_unr17_stage7_stallmux_q_16_;
wire delay_add_ln22_unr17_stage7_stallmux_q_17_;
wire delay_add_ln22_unr17_stage7_stallmux_q_18_;
wire delay_add_ln22_unr17_stage7_stallmux_q_19_;
wire delay_add_ln22_unr17_stage7_stallmux_q_1_;
wire delay_add_ln22_unr17_stage7_stallmux_q_20_;
wire delay_add_ln22_unr17_stage7_stallmux_q_21_;
wire delay_add_ln22_unr17_stage7_stallmux_q_22_;
wire delay_add_ln22_unr17_stage7_stallmux_q_23_;
wire delay_add_ln22_unr17_stage7_stallmux_q_24_;
wire delay_add_ln22_unr17_stage7_stallmux_q_25_;
wire delay_add_ln22_unr17_stage7_stallmux_q_26_;
wire delay_add_ln22_unr17_stage7_stallmux_q_27_;
wire delay_add_ln22_unr17_stage7_stallmux_q_28_;
wire delay_add_ln22_unr17_stage7_stallmux_q_29_;
wire delay_add_ln22_unr17_stage7_stallmux_q_2_;
wire delay_add_ln22_unr17_stage7_stallmux_q_30_;
wire delay_add_ln22_unr17_stage7_stallmux_q_31_;
wire delay_add_ln22_unr17_stage7_stallmux_q_3_;
wire delay_add_ln22_unr17_stage7_stallmux_q_4_;
wire delay_add_ln22_unr17_stage7_stallmux_q_5_;
wire delay_add_ln22_unr17_stage7_stallmux_q_6_;
wire delay_add_ln22_unr17_stage7_stallmux_q_7_;
wire delay_add_ln22_unr17_stage7_stallmux_q_8_;
wire delay_add_ln22_unr17_stage7_stallmux_q_9_;
wire delay_add_ln22_unr20_stage8_stallmux_q_0_;
wire delay_add_ln22_unr20_stage8_stallmux_q_10_;
wire delay_add_ln22_unr20_stage8_stallmux_q_11_;
wire delay_add_ln22_unr20_stage8_stallmux_q_12_;
wire delay_add_ln22_unr20_stage8_stallmux_q_13_;
wire delay_add_ln22_unr20_stage8_stallmux_q_14_;
wire delay_add_ln22_unr20_stage8_stallmux_q_15_;
wire delay_add_ln22_unr20_stage8_stallmux_q_16_;
wire delay_add_ln22_unr20_stage8_stallmux_q_17_;
wire delay_add_ln22_unr20_stage8_stallmux_q_18_;
wire delay_add_ln22_unr20_stage8_stallmux_q_19_;
wire delay_add_ln22_unr20_stage8_stallmux_q_1_;
wire delay_add_ln22_unr20_stage8_stallmux_q_20_;
wire delay_add_ln22_unr20_stage8_stallmux_q_21_;
wire delay_add_ln22_unr20_stage8_stallmux_q_22_;
wire delay_add_ln22_unr20_stage8_stallmux_q_23_;
wire delay_add_ln22_unr20_stage8_stallmux_q_24_;
wire delay_add_ln22_unr20_stage8_stallmux_q_25_;
wire delay_add_ln22_unr20_stage8_stallmux_q_26_;
wire delay_add_ln22_unr20_stage8_stallmux_q_27_;
wire delay_add_ln22_unr20_stage8_stallmux_q_28_;
wire delay_add_ln22_unr20_stage8_stallmux_q_29_;
wire delay_add_ln22_unr20_stage8_stallmux_q_2_;
wire delay_add_ln22_unr20_stage8_stallmux_q_30_;
wire delay_add_ln22_unr20_stage8_stallmux_q_31_;
wire delay_add_ln22_unr20_stage8_stallmux_q_3_;
wire delay_add_ln22_unr20_stage8_stallmux_q_4_;
wire delay_add_ln22_unr20_stage8_stallmux_q_5_;
wire delay_add_ln22_unr20_stage8_stallmux_q_6_;
wire delay_add_ln22_unr20_stage8_stallmux_q_7_;
wire delay_add_ln22_unr20_stage8_stallmux_q_8_;
wire delay_add_ln22_unr20_stage8_stallmux_q_9_;
wire delay_add_ln22_unr23_stage9_stallmux_q_0_;
wire delay_add_ln22_unr23_stage9_stallmux_q_10_;
wire delay_add_ln22_unr23_stage9_stallmux_q_11_;
wire delay_add_ln22_unr23_stage9_stallmux_q_12_;
wire delay_add_ln22_unr23_stage9_stallmux_q_13_;
wire delay_add_ln22_unr23_stage9_stallmux_q_14_;
wire delay_add_ln22_unr23_stage9_stallmux_q_15_;
wire delay_add_ln22_unr23_stage9_stallmux_q_16_;
wire delay_add_ln22_unr23_stage9_stallmux_q_17_;
wire delay_add_ln22_unr23_stage9_stallmux_q_18_;
wire delay_add_ln22_unr23_stage9_stallmux_q_19_;
wire delay_add_ln22_unr23_stage9_stallmux_q_1_;
wire delay_add_ln22_unr23_stage9_stallmux_q_20_;
wire delay_add_ln22_unr23_stage9_stallmux_q_21_;
wire delay_add_ln22_unr23_stage9_stallmux_q_22_;
wire delay_add_ln22_unr23_stage9_stallmux_q_23_;
wire delay_add_ln22_unr23_stage9_stallmux_q_24_;
wire delay_add_ln22_unr23_stage9_stallmux_q_25_;
wire delay_add_ln22_unr23_stage9_stallmux_q_26_;
wire delay_add_ln22_unr23_stage9_stallmux_q_27_;
wire delay_add_ln22_unr23_stage9_stallmux_q_28_;
wire delay_add_ln22_unr23_stage9_stallmux_q_29_;
wire delay_add_ln22_unr23_stage9_stallmux_q_2_;
wire delay_add_ln22_unr23_stage9_stallmux_q_30_;
wire delay_add_ln22_unr23_stage9_stallmux_q_31_;
wire delay_add_ln22_unr23_stage9_stallmux_q_3_;
wire delay_add_ln22_unr23_stage9_stallmux_q_4_;
wire delay_add_ln22_unr23_stage9_stallmux_q_5_;
wire delay_add_ln22_unr23_stage9_stallmux_q_6_;
wire delay_add_ln22_unr23_stage9_stallmux_q_7_;
wire delay_add_ln22_unr23_stage9_stallmux_q_8_;
wire delay_add_ln22_unr23_stage9_stallmux_q_9_;
wire delay_add_ln22_unr27_stage10_stallmux_q_0_;
wire delay_add_ln22_unr27_stage10_stallmux_q_10_;
wire delay_add_ln22_unr27_stage10_stallmux_q_11_;
wire delay_add_ln22_unr27_stage10_stallmux_q_12_;
wire delay_add_ln22_unr27_stage10_stallmux_q_13_;
wire delay_add_ln22_unr27_stage10_stallmux_q_14_;
wire delay_add_ln22_unr27_stage10_stallmux_q_15_;
wire delay_add_ln22_unr27_stage10_stallmux_q_16_;
wire delay_add_ln22_unr27_stage10_stallmux_q_17_;
wire delay_add_ln22_unr27_stage10_stallmux_q_18_;
wire delay_add_ln22_unr27_stage10_stallmux_q_19_;
wire delay_add_ln22_unr27_stage10_stallmux_q_1_;
wire delay_add_ln22_unr27_stage10_stallmux_q_20_;
wire delay_add_ln22_unr27_stage10_stallmux_q_21_;
wire delay_add_ln22_unr27_stage10_stallmux_q_22_;
wire delay_add_ln22_unr27_stage10_stallmux_q_23_;
wire delay_add_ln22_unr27_stage10_stallmux_q_24_;
wire delay_add_ln22_unr27_stage10_stallmux_q_25_;
wire delay_add_ln22_unr27_stage10_stallmux_q_26_;
wire delay_add_ln22_unr27_stage10_stallmux_q_27_;
wire delay_add_ln22_unr27_stage10_stallmux_q_28_;
wire delay_add_ln22_unr27_stage10_stallmux_q_29_;
wire delay_add_ln22_unr27_stage10_stallmux_q_2_;
wire delay_add_ln22_unr27_stage10_stallmux_q_30_;
wire delay_add_ln22_unr27_stage10_stallmux_q_31_;
wire delay_add_ln22_unr27_stage10_stallmux_q_3_;
wire delay_add_ln22_unr27_stage10_stallmux_q_4_;
wire delay_add_ln22_unr27_stage10_stallmux_q_5_;
wire delay_add_ln22_unr27_stage10_stallmux_q_6_;
wire delay_add_ln22_unr27_stage10_stallmux_q_7_;
wire delay_add_ln22_unr27_stage10_stallmux_q_8_;
wire delay_add_ln22_unr27_stage10_stallmux_q_9_;
wire delay_add_ln22_unr2_stage2_stallmux_q_10_;
wire delay_add_ln22_unr2_stage2_stallmux_q_11_;
wire delay_add_ln22_unr2_stage2_stallmux_q_12_;
wire delay_add_ln22_unr2_stage2_stallmux_q_13_;
wire delay_add_ln22_unr2_stage2_stallmux_q_14_;
wire delay_add_ln22_unr2_stage2_stallmux_q_15_;
wire delay_add_ln22_unr2_stage2_stallmux_q_16_;
wire delay_add_ln22_unr2_stage2_stallmux_q_17_;
wire delay_add_ln22_unr2_stage2_stallmux_q_18_;
wire delay_add_ln22_unr2_stage2_stallmux_q_19_;
wire delay_add_ln22_unr2_stage2_stallmux_q_1_;
wire delay_add_ln22_unr2_stage2_stallmux_q_20_;
wire delay_add_ln22_unr2_stage2_stallmux_q_21_;
wire delay_add_ln22_unr2_stage2_stallmux_q_22_;
wire delay_add_ln22_unr2_stage2_stallmux_q_23_;
wire delay_add_ln22_unr2_stage2_stallmux_q_24_;
wire delay_add_ln22_unr2_stage2_stallmux_q_25_;
wire delay_add_ln22_unr2_stage2_stallmux_q_26_;
wire delay_add_ln22_unr2_stage2_stallmux_q_27_;
wire delay_add_ln22_unr2_stage2_stallmux_q_28_;
wire delay_add_ln22_unr2_stage2_stallmux_q_29_;
wire delay_add_ln22_unr2_stage2_stallmux_q_2_;
wire delay_add_ln22_unr2_stage2_stallmux_q_30_;
wire delay_add_ln22_unr2_stage2_stallmux_q_31_;
wire delay_add_ln22_unr2_stage2_stallmux_q_3_;
wire delay_add_ln22_unr2_stage2_stallmux_q_4_;
wire delay_add_ln22_unr2_stage2_stallmux_q_5_;
wire delay_add_ln22_unr2_stage2_stallmux_q_6_;
wire delay_add_ln22_unr2_stage2_stallmux_q_7_;
wire delay_add_ln22_unr2_stage2_stallmux_q_8_;
wire delay_add_ln22_unr2_stage2_stallmux_q_9_;
wire delay_add_ln22_unr5_stage3_stallmux_q_0_;
wire delay_add_ln22_unr5_stage3_stallmux_q_10_;
wire delay_add_ln22_unr5_stage3_stallmux_q_11_;
wire delay_add_ln22_unr5_stage3_stallmux_q_12_;
wire delay_add_ln22_unr5_stage3_stallmux_q_13_;
wire delay_add_ln22_unr5_stage3_stallmux_q_14_;
wire delay_add_ln22_unr5_stage3_stallmux_q_15_;
wire delay_add_ln22_unr5_stage3_stallmux_q_16_;
wire delay_add_ln22_unr5_stage3_stallmux_q_17_;
wire delay_add_ln22_unr5_stage3_stallmux_q_18_;
wire delay_add_ln22_unr5_stage3_stallmux_q_19_;
wire delay_add_ln22_unr5_stage3_stallmux_q_1_;
wire delay_add_ln22_unr5_stage3_stallmux_q_20_;
wire delay_add_ln22_unr5_stage3_stallmux_q_21_;
wire delay_add_ln22_unr5_stage3_stallmux_q_22_;
wire delay_add_ln22_unr5_stage3_stallmux_q_23_;
wire delay_add_ln22_unr5_stage3_stallmux_q_24_;
wire delay_add_ln22_unr5_stage3_stallmux_q_25_;
wire delay_add_ln22_unr5_stage3_stallmux_q_26_;
wire delay_add_ln22_unr5_stage3_stallmux_q_27_;
wire delay_add_ln22_unr5_stage3_stallmux_q_28_;
wire delay_add_ln22_unr5_stage3_stallmux_q_29_;
wire delay_add_ln22_unr5_stage3_stallmux_q_2_;
wire delay_add_ln22_unr5_stage3_stallmux_q_30_;
wire delay_add_ln22_unr5_stage3_stallmux_q_31_;
wire delay_add_ln22_unr5_stage3_stallmux_q_3_;
wire delay_add_ln22_unr5_stage3_stallmux_q_4_;
wire delay_add_ln22_unr5_stage3_stallmux_q_5_;
wire delay_add_ln22_unr5_stage3_stallmux_q_6_;
wire delay_add_ln22_unr5_stage3_stallmux_q_7_;
wire delay_add_ln22_unr5_stage3_stallmux_q_8_;
wire delay_add_ln22_unr5_stage3_stallmux_q_9_;
wire delay_add_ln22_unr8_stage4_stallmux_q_0_;
wire delay_add_ln22_unr8_stage4_stallmux_q_10_;
wire delay_add_ln22_unr8_stage4_stallmux_q_11_;
wire delay_add_ln22_unr8_stage4_stallmux_q_12_;
wire delay_add_ln22_unr8_stage4_stallmux_q_13_;
wire delay_add_ln22_unr8_stage4_stallmux_q_14_;
wire delay_add_ln22_unr8_stage4_stallmux_q_15_;
wire delay_add_ln22_unr8_stage4_stallmux_q_16_;
wire delay_add_ln22_unr8_stage4_stallmux_q_17_;
wire delay_add_ln22_unr8_stage4_stallmux_q_18_;
wire delay_add_ln22_unr8_stage4_stallmux_q_19_;
wire delay_add_ln22_unr8_stage4_stallmux_q_1_;
wire delay_add_ln22_unr8_stage4_stallmux_q_20_;
wire delay_add_ln22_unr8_stage4_stallmux_q_21_;
wire delay_add_ln22_unr8_stage4_stallmux_q_22_;
wire delay_add_ln22_unr8_stage4_stallmux_q_23_;
wire delay_add_ln22_unr8_stage4_stallmux_q_24_;
wire delay_add_ln22_unr8_stage4_stallmux_q_25_;
wire delay_add_ln22_unr8_stage4_stallmux_q_26_;
wire delay_add_ln22_unr8_stage4_stallmux_q_27_;
wire delay_add_ln22_unr8_stage4_stallmux_q_28_;
wire delay_add_ln22_unr8_stage4_stallmux_q_29_;
wire delay_add_ln22_unr8_stage4_stallmux_q_2_;
wire delay_add_ln22_unr8_stage4_stallmux_q_30_;
wire delay_add_ln22_unr8_stage4_stallmux_q_31_;
wire delay_add_ln22_unr8_stage4_stallmux_q_3_;
wire delay_add_ln22_unr8_stage4_stallmux_q_4_;
wire delay_add_ln22_unr8_stage4_stallmux_q_5_;
wire delay_add_ln22_unr8_stage4_stallmux_q_6_;
wire delay_add_ln22_unr8_stage4_stallmux_q_7_;
wire delay_add_ln22_unr8_stage4_stallmux_q_8_;
wire delay_add_ln22_unr8_stage4_stallmux_q_9_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_0_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_10_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_11_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_12_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_13_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_14_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_15_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_16_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_17_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_18_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_19_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_1_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_20_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_21_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_22_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_23_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_24_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_25_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_26_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_27_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_28_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_29_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_2_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_30_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_31_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_3_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_4_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_5_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_6_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_7_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_8_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_9_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_0_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_10_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_11_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_12_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_13_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_14_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_15_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_16_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_17_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_18_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_19_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_1_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_20_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_21_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_22_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_23_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_24_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_25_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_26_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_27_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_28_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_29_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_2_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_30_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_31_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_3_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_4_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_5_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_6_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_7_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_8_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_9_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_0_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_10_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_11_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_12_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_13_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_14_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_15_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_16_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_17_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_18_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_19_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_1_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_20_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_21_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_22_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_23_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_24_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_25_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_26_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_27_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_28_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_29_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_2_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_30_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_31_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_3_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_4_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_5_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_6_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_7_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_8_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_9_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_0_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_10_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_11_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_12_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_13_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_14_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_15_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_16_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_17_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_18_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_19_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_1_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_20_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_21_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_22_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_23_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_24_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_25_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_26_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_27_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_28_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_29_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_2_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_30_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_31_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_3_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_4_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_5_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_6_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_7_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_8_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_9_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_0_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_10_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_11_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_12_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_13_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_14_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_15_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_16_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_17_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_18_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_19_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_1_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_20_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_21_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_22_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_23_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_24_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_25_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_26_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_27_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_28_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_29_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_2_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_30_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_31_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_3_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_4_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_5_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_6_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_7_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_8_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_9_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_0_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_10_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_11_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_12_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_13_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_14_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_15_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_16_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_17_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_18_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_19_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_1_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_20_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_21_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_22_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_23_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_24_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_25_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_26_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_27_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_28_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_29_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_2_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_30_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_31_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_3_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_4_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_5_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_6_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_7_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_8_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_9_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_0_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_10_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_12_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_13_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_15_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_16_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_17_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_18_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_19_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_1_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_20_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_21_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_22_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_23_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_24_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_25_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_26_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_27_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_28_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_29_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_2_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_3_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_4_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_5_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_6_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_7_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_8_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_9_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_0_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_10_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_11_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_12_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_13_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_14_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_15_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_16_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_17_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_18_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_19_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_1_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_20_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_21_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_22_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_23_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_24_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_25_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_26_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_27_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_28_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_29_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_2_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_30_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_31_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_3_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_4_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_5_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_6_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_7_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_8_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_9_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_0_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_10_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_11_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_12_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_13_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_14_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_15_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_16_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_17_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_18_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_19_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_1_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_20_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_21_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_22_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_23_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_24_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_25_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_26_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_27_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_28_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_29_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_2_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_30_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_31_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_3_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_4_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_5_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_6_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_7_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_8_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_9_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_1_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_2_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_3_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_4_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_5_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_6_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_7_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_8_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_0_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_1_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_2_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_3_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_4_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_5_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_6_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_7_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_10_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_11_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_12_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_13_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_14_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_15_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_16_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_17_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_18_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_19_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_1_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_20_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_21_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_22_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_23_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_24_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_25_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_26_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_27_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_28_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_29_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_2_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_30_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_3_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_4_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_5_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_6_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_7_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_8_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_9_;
wire delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_10_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_11_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_12_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_13_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_14_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_15_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_16_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_17_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_18_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_19_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_1_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_20_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_21_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_22_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_23_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_24_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_25_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_26_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_27_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_28_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_29_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_2_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_30_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_3_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_4_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_5_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_6_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_7_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_8_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_9_;
wire delay_sub_ln23_0_unr1_stage2_stallmux_q_0_;
wire delay_sub_ln23_0_unr1_stage2_stallmux_q_1_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_10_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_11_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_12_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_13_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_14_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_15_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_16_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_17_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_18_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_19_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_1_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_20_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_21_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_22_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_23_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_24_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_25_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_26_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_27_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_28_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_29_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_2_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_30_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_3_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_4_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_5_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_6_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_7_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_8_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_9_;
wire delay_sub_ln23_0_unr21_stage8_stallmux_q;
wire delay_sub_ln23_0_unr22_stage8_stallmux_q;
wire delay_sub_ln23_0_unr23_stage8_stallmux_q;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_0_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_10_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_11_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_12_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_13_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_14_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_15_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_16_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_17_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_18_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_19_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_1_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_20_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_21_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_22_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_23_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_24_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_25_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_26_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_27_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_28_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_29_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_2_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_30_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_3_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_4_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_5_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_6_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_7_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_8_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_9_;
wire delay_sub_ln23_0_unr24_stage9_stallmux_q;
wire delay_sub_ln23_0_unr25_stage9_stallmux_q;
wire delay_sub_ln23_0_unr26_stage9_stallmux_q_0_;
wire delay_sub_ln23_0_unr26_stage9_stallmux_q_1_;
wire delay_sub_ln23_0_unr26_stage9_stallmux_q_2_;
wire delay_sub_ln23_0_unr27_stage10_stallmux_z;
wire delay_sub_ln23_0_unr28_stage10_stallmux_q;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_0_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_10_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_11_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_12_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_13_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_14_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_15_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_16_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_17_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_18_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_19_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_1_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_20_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_21_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_22_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_23_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_24_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_25_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_26_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_27_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_28_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_2_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_3_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_4_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_5_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_6_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_7_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_8_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_9_;
wire delay_sub_ln23_0_unr29_stage10_stallmux_q;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_0_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_10_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_11_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_12_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_13_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_14_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_15_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_16_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_17_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_18_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_19_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_1_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_20_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_21_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_22_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_23_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_24_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_25_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_26_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_27_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_28_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_2_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_3_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_4_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_5_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_6_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_7_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_8_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_9_;
wire delay_sub_ln23_0_unr30_stage10_stallmux_q;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_0_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_10_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_11_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_12_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_13_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_14_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_15_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_16_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_17_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_18_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_19_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_1_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_20_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_21_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_22_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_23_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_24_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_25_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_26_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_27_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_28_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_29_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_2_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_30_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_3_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_4_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_5_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_6_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_7_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_8_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_9_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_0_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_10_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_11_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_12_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_13_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_14_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_15_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_16_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_17_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_18_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_19_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_1_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_20_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_21_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_22_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_23_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_24_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_25_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_26_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_27_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_28_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_29_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_2_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_3_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_4_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_5_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_6_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_7_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_8_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_9_;
wire delay_sub_ln23_unr13_stage5_stallmux_q_1_;
wire delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire delay_sub_ln23_unr21_stage7_stallmux_q_1_;
wire delay_sub_ln23_unr25_stage8_stallmux_q_1_;
wire delay_sub_ln23_unr25_stage8_stallmux_q_3_;
wire delay_sub_ln23_unr29_stage9_stallmux_q_2_;
wire delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_10_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_11_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_12_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_13_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_14_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_15_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_16_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_17_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_18_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_19_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_2_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_3_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_4_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_5_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_6_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_7_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_8_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_9_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_0_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_10_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_11_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_12_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_13_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_14_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_15_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_16_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_1_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_2_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_3_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_4_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_5_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_6_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_7_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_8_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_9_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_10_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_11_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_12_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_13_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_2_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_3_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_5_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_6_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_7_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_8_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_9_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_0_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_10_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_1_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_2_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_3_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_4_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_5_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_6_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_7_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_8_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_9_;
wire delay_xor_ln21_unr28_stage10_stallmux_q_0_;
wire delay_xor_ln21_unr28_stage10_stallmux_q_1_;
wire delay_xor_ln21_unr28_stage10_stallmux_q_2_;
wire delay_xor_ln21_unr28_stage10_stallmux_q_3_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_0_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_10_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_11_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_12_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_13_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_14_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_15_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_16_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_17_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_18_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_19_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_1_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_20_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_21_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_22_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_23_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_24_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_25_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_26_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_27_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_28_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_2_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_3_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_4_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_5_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_6_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_7_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_8_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_9_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_0_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_10_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_11_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_12_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_13_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_14_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_15_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_16_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_17_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_18_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_19_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_1_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_20_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_21_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_22_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_23_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_24_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_25_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_2_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_3_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_4_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_5_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_6_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_7_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_8_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_9_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_0_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_10_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_11_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_12_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_13_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_14_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_15_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_16_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_17_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_18_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_19_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_1_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_20_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_21_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_22_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_2_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_3_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_4_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_5_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_6_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_7_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_8_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_9_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_0_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_10_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_11_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_12_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_13_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_14_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_15_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_16_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_17_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_18_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_19_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_1_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_2_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_3_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_4_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_5_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_6_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_7_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_8_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_9_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_0_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_10_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_11_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_12_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_13_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_14_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_15_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_16_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_2_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_3_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_4_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_5_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_6_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_7_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_8_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_9_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_0_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_10_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_11_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_12_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_13_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_1_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_2_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_3_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_4_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_5_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_6_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_7_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_8_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_9_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_0_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_10_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_1_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_2_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_3_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_4_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_5_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_6_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_7_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_8_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_9_;
wire delay_xor_ln22_unr28_stage10_stallmux_q_0_;
wire delay_xor_ln22_unr28_stage10_stallmux_q_1_;
wire delay_xor_ln22_unr28_stage10_stallmux_q_2_;
wire delay_xor_ln22_unr28_stage10_stallmux_q_3_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_0_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_10_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_11_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_12_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_13_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_14_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_15_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_16_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_17_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_18_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_19_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_1_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_20_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_21_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_22_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_23_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_24_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_25_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_26_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_27_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_28_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_2_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_3_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_4_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_5_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_6_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_7_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_8_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_9_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_0_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_10_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_11_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_12_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_13_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_14_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_15_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_16_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_17_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_18_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_19_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_1_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_20_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_21_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_22_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_23_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_24_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_25_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_2_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_3_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_4_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_5_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_6_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_7_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_8_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_9_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_10_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_11_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_12_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_13_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_14_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_15_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_16_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_17_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_18_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_19_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_20_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_21_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_22_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_2_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_3_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_4_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_5_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_6_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_7_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_8_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_9_;
wire delay_xor_ln23_unr3_stage2_stallmux_q;
wire delay_xor_ln23_unr6_stage3_stallmux_q;
wire mux_while_ln12_psv_q_1_;
wire mux_while_ln12_psv_q_2_;
wire mux_while_ln12_psv_q_3_;
wire mux_while_ln12_psv_q_4_;
wire mux_while_ln12_psv_q_5_;
wire mux_while_ln12_psv_q_6_;
wire mux_while_ln12_psv_q_7_;
wire mux_while_ln12_psv_q_8_;
wire n_1;
wire n_100;
wire n_1000;
wire n_10000;
wire n_10001;
wire n_10002;
wire n_10003;
wire n_10004;
wire n_10005;
wire n_10006;
wire n_10007;
wire n_10008;
wire n_1001;
wire n_10010;
wire n_10013;
wire n_10014;
wire n_10015;
wire n_10016;
wire n_10017;
wire n_10019;
wire n_1002;
wire n_10020;
wire n_10021;
wire n_10022;
wire n_10023;
wire n_10025;
wire n_10027;
wire n_10028;
wire n_10029;
wire n_1003;
wire n_10030;
wire n_10031;
wire n_10032;
wire n_10033;
wire n_10034;
wire n_10035;
wire n_10036;
wire n_10037;
wire n_10038;
wire n_10039;
wire n_1004;
wire n_10040;
wire n_10041;
wire n_10042;
wire n_10043;
wire n_10044;
wire n_10045;
wire n_10047;
wire n_10048;
wire n_10049;
wire n_1005;
wire n_10050;
wire n_10051;
wire TIMEBOOST_net_1329;
wire n_10053;
wire n_10054;
wire n_10057;
wire TIMEBOOST_net_477;
wire n_1006;
wire n_10060;
wire n_10061;
wire n_10062;
wire n_10063;
wire n_10065;
wire n_10067;
wire n_10068;
wire n_1007;
wire n_10070;
wire n_10071;
wire n_10072;
wire n_10073;
wire n_10077;
wire n_10078;
wire n_10079;
wire n_1008;
wire n_10081;
wire n_10082;
wire n_10083;
wire n_10085;
wire n_10086;
wire n_10087;
wire n_10088;
wire n_10089;
wire n_1009;
wire n_10090;
wire TIMEBOOST_net_2733;
wire n_10092;
wire n_10094;
wire n_10095;
wire n_10096;
wire n_10098;
wire n_101;
wire n_1010;
wire n_10100;
wire n_10101;
wire n_10102;
wire n_10104;
wire n_10105;
wire n_10106;
wire n_10107;
wire n_10109;
wire n_1011;
wire n_10111;
wire n_10112;
wire n_10113;
wire n_10116;
wire n_10119;
wire n_1012;
wire n_10120;
wire n_10121;
wire n_10122;
wire n_10123;
wire n_10124;
wire n_10125;
wire n_10127;
wire n_10128;
wire n_10129;
wire n_1013;
wire n_10130;
wire n_10131;
wire n_10132;
wire n_10133;
wire n_10134;
wire n_10136;
wire n_10137;
wire n_10138;
wire n_10139;
wire n_1014;
wire n_10140;
wire n_10141;
wire n_10142;
wire n_10145;
wire n_10146;
wire n_10148;
wire n_10149;
wire n_1015;
wire n_10150;
wire TIMEBOOST_net_638;
wire n_10153;
wire n_10154;
wire n_10156;
wire n_10157;
wire n_10158;
wire n_10159;
wire n_1016;
wire n_10160;
wire n_10161;
wire n_10162;
wire n_10163;
wire n_10164;
wire n_10165;
wire n_10166;
wire n_10167;
wire n_10168;
wire n_10169;
wire n_1017;
wire n_10170;
wire n_10171;
wire n_10174;
wire n_10175;
wire n_10176;
wire n_10177;
wire TIMEBOOST_net_610;
wire n_10179;
wire n_1018;
wire n_10180;
wire n_10181;
wire n_10182;
wire n_10183;
wire n_10185;
wire n_10186;
wire n_10188;
wire n_1019;
wire n_10190;
wire n_10191;
wire n_10192;
wire n_10193;
wire n_10194;
wire n_10195;
wire n_10197;
wire n_10198;
wire n_102;
wire n_1020;
wire n_10200;
wire n_10201;
wire n_10203;
wire n_10204;
wire n_10206;
wire n_10207;
wire n_10208;
wire n_10209;
wire n_1021;
wire n_10210;
wire n_10211;
wire n_10212;
wire n_10213;
wire n_10214;
wire n_10215;
wire n_10216;
wire n_10217;
wire n_10218;
wire n_10219;
wire n_1022;
wire n_10220;
wire n_10222;
wire n_10223;
wire n_10225;
wire n_10228;
wire n_1023;
wire n_10230;
wire n_10236;
wire n_10237;
wire n_10238;
wire n_10239;
wire n_1024;
wire n_10240;
wire n_10241;
wire n_10242;
wire n_10243;
wire n_10245;
wire n_10246;
wire n_10247;
wire n_10248;
wire n_10249;
wire n_1025;
wire n_10250;
wire n_10251;
wire n_10252;
wire n_10254;
wire n_10255;
wire n_10256;
wire n_10257;
wire n_10258;
wire n_10259;
wire n_1026;
wire n_10260;
wire n_10261;
wire n_10262;
wire n_10263;
wire n_10264;
wire n_10265;
wire n_10267;
wire n_1027;
wire n_10270;
wire n_10274;
wire n_10276;
wire n_10277;
wire n_10278;
wire n_10279;
wire n_1028;
wire n_10280;
wire n_10282;
wire n_10283;
wire n_10284;
wire n_10285;
wire n_10286;
wire n_10287;
wire n_10288;
wire n_10289;
wire n_1029;
wire n_10290;
wire n_10293;
wire n_10295;
wire n_10296;
wire n_10297;
wire n_103;
wire n_1030;
wire n_10300;
wire n_10301;
wire n_10302;
wire n_10303;
wire n_10304;
wire n_10305;
wire n_10306;
wire n_10307;
wire n_10309;
wire n_1031;
wire n_10310;
wire n_10311;
wire n_10313;
wire n_10317;
wire n_10318;
wire n_10319;
wire n_1032;
wire n_10320;
wire n_10321;
wire n_10322;
wire n_10323;
wire n_10324;
wire n_10325;
wire n_10326;
wire n_10328;
wire n_10329;
wire n_1033;
wire n_10330;
wire n_10331;
wire n_10332;
wire n_10334;
wire n_10337;
wire n_10338;
wire n_10339;
wire n_10340;
wire n_10341;
wire n_10342;
wire n_10343;
wire n_10344;
wire n_10347;
wire n_10349;
wire n_10350;
wire n_10351;
wire n_10352;
wire n_10353;
wire n_10354;
wire n_10355;
wire n_10356;
wire n_10357;
wire n_10359;
wire n_10360;
wire n_10362;
wire n_10363;
wire n_10364;
wire n_10365;
wire n_10366;
wire TIMEBOOST_net_1244;
wire n_10368;
wire n_10369;
wire n_1037;
wire n_10371;
wire TIMEBOOST_net_644;
wire n_10373;
wire n_10374;
wire n_10375;
wire TIMEBOOST_net_1743;
wire n_10377;
wire n_10379;
wire n_1038;
wire n_10380;
wire n_10381;
wire n_10382;
wire n_10383;
wire n_10384;
wire n_10385;
wire n_10386;
wire n_10387;
wire TIMEBOOST_net_1420;
wire n_10389;
wire n_1039;
wire n_10390;
wire n_10391;
wire n_10392;
wire n_10393;
wire n_10394;
wire n_10396;
wire n_10397;
wire n_10398;
wire n_10399;
wire n_104;
wire n_1040;
wire n_10401;
wire n_10402;
wire n_10403;
wire n_10404;
wire n_10405;
wire n_10406;
wire TIMEBOOST_net_648;
wire TIMEBOOST_net_2753;
wire n_1041;
wire n_10410;
wire n_10411;
wire n_10412;
wire n_10413;
wire TIMEBOOST_net_1304;
wire n_10415;
wire n_10416;
wire n_10417;
wire n_10418;
wire n_10419;
wire n_1042;
wire n_10420;
wire n_10421;
wire n_10422;
wire n_10423;
wire n_10424;
wire n_10425;
wire n_10426;
wire n_10428;
wire n_10429;
wire n_1043;
wire n_10430;
wire n_10431;
wire n_10432;
wire n_10433;
wire n_10434;
wire n_10435;
wire TIMEBOOST_net_2063;
wire n_10437;
wire n_1044;
wire n_10440;
wire n_10441;
wire TIMEBOOST_net_456;
wire TIMEBOOST_net_1717;
wire n_10445;
wire n_1045;
wire n_10451;
wire n_10454;
wire n_10456;
wire n_10457;
wire n_10458;
wire TIMEBOOST_net_369;
wire n_1046;
wire n_10461;
wire n_10462;
wire n_10464;
wire n_10465;
wire n_10467;
wire n_10468;
wire n_10469;
wire n_1047;
wire n_10470;
wire n_10471;
wire n_10472;
wire n_10473;
wire n_10474;
wire n_10475;
wire n_10477;
wire n_10478;
wire n_1048;
wire n_10480;
wire n_10481;
wire n_10483;
wire n_10484;
wire n_10485;
wire TIMEBOOST_net_2236;
wire TIMEBOOST_net_1253;
wire n_10489;
wire n_1049;
wire n_10490;
wire n_10491;
wire n_10492;
wire n_10494;
wire n_10495;
wire n_10496;
wire n_10498;
wire n_10499;
wire n_105;
wire n_1050;
wire n_10500;
wire TIMEBOOST_net_2534;
wire n_10503;
wire n_10505;
wire n_10506;
wire n_10507;
wire n_10508;
wire n_1051;
wire TIMEBOOST_net_1754;
wire n_10511;
wire n_10513;
wire n_10514;
wire n_10517;
wire n_10518;
wire n_1052;
wire TIMEBOOST_net_2764;
wire n_10521;
wire n_10522;
wire n_10523;
wire n_10524;
wire n_10525;
wire n_10526;
wire n_10527;
wire n_10529;
wire n_1053;
wire n_10530;
wire n_10531;
wire n_10535;
wire n_10536;
wire n_10537;
wire n_10538;
wire n_1054;
wire n_10541;
wire n_10543;
wire n_10544;
wire n_10545;
wire n_10547;
wire n_10548;
wire n_10549;
wire n_1055;
wire n_10550;
wire n_10551;
wire TIMEBOOST_net_517;
wire n_10554;
wire n_10555;
wire n_10556;
wire n_10557;
wire n_10559;
wire n_1056;
wire n_10560;
wire n_10561;
wire n_10562;
wire n_10563;
wire n_10564;
wire n_10565;
wire n_10566;
wire n_10567;
wire n_10568;
wire n_10569;
wire n_1057;
wire n_10570;
wire n_10571;
wire n_10572;
wire n_10573;
wire TIMEBOOST_net_615;
wire n_10575;
wire n_10576;
wire n_10577;
wire n_10578;
wire n_10579;
wire n_1058;
wire n_10582;
wire n_10584;
wire n_10585;
wire n_10586;
wire n_10587;
wire n_10588;
wire n_1059;
wire TIMEBOOST_net_591;
wire n_10591;
wire n_10592;
wire n_10594;
wire TIMEBOOST_net_2241;
wire n_10597;
wire n_10598;
wire n_10599;
wire n_106;
wire n_1060;
wire TIMEBOOST_net_652;
wire n_10601;
wire n_10603;
wire n_10604;
wire n_10607;
wire n_10608;
wire n_10609;
wire n_1061;
wire n_10610;
wire n_10611;
wire n_10612;
wire n_10613;
wire n_10614;
wire n_10615;
wire n_10616;
wire n_10618;
wire n_10619;
wire n_1062;
wire n_10620;
wire TIMEBOOST_net_1256;
wire n_10624;
wire n_10626;
wire n_10629;
wire n_1063;
wire n_10630;
wire n_10631;
wire n_10632;
wire n_10633;
wire n_10634;
wire n_10635;
wire n_10636;
wire n_10637;
wire n_10638;
wire n_10639;
wire n_1064;
wire n_10640;
wire n_10641;
wire n_10644;
wire n_10647;
wire TIMEBOOST_net_2813;
wire n_1065;
wire n_10650;
wire n_10652;
wire n_10653;
wire n_10654;
wire n_10656;
wire n_10657;
wire n_10658;
wire n_10659;
wire n_1066;
wire n_10660;
wire n_10664;
wire n_10665;
wire n_10666;
wire n_10667;
wire TIMEBOOST_net_1767;
wire n_10669;
wire n_1067;
wire n_10670;
wire n_10671;
wire n_10672;
wire n_10673;
wire TIMEBOOST_net_2292;
wire n_10676;
wire n_10677;
wire n_10678;
wire n_1068;
wire n_10680;
wire n_10681;
wire n_10682;
wire n_10684;
wire n_10686;
wire n_10687;
wire n_10688;
wire n_10689;
wire n_1069;
wire n_10690;
wire n_10691;
wire n_10692;
wire n_10693;
wire n_10694;
wire n_10696;
wire TIMEBOOST_net_1770;
wire n_10699;
wire n_107;
wire n_1070;
wire n_10700;
wire n_10702;
wire n_10704;
wire n_10705;
wire n_10707;
wire n_10708;
wire n_10709;
wire n_1071;
wire n_10710;
wire n_10711;
wire n_10712;
wire n_10713;
wire n_10714;
wire n_10716;
wire n_10717;
wire TIMEBOOST_net_1996;
wire n_10719;
wire n_1072;
wire n_10720;
wire n_10721;
wire n_10722;
wire n_10723;
wire n_10724;
wire n_10725;
wire n_10726;
wire n_10727;
wire n_10729;
wire n_1073;
wire n_10730;
wire n_10731;
wire n_10732;
wire n_10733;
wire n_10734;
wire n_10735;
wire n_10736;
wire n_10737;
wire n_10739;
wire n_1074;
wire n_10740;
wire TIMEBOOST_net_1107;
wire n_10742;
wire n_10744;
wire n_10745;
wire n_10746;
wire n_10747;
wire n_10748;
wire n_10749;
wire n_1075;
wire n_10751;
wire n_10752;
wire n_10753;
wire n_10754;
wire n_10755;
wire n_10756;
wire n_10757;
wire n_10758;
wire n_10759;
wire n_1076;
wire n_10760;
wire n_10761;
wire n_10762;
wire n_10763;
wire n_10764;
wire n_10765;
wire n_10766;
wire n_10767;
wire n_10768;
wire TIMEBOOST_net_2950;
wire n_1077;
wire n_10770;
wire TIMEBOOST_net_2473;
wire n_10772;
wire n_10773;
wire n_10775;
wire n_10776;
wire n_10777;
wire n_10778;
wire n_10779;
wire n_1078;
wire n_10781;
wire n_10782;
wire n_10783;
wire n_10784;
wire n_10785;
wire TIMEBOOST_net_2477;
wire n_10787;
wire n_10788;
wire n_10789;
wire n_1079;
wire n_10790;
wire n_10791;
wire n_10792;
wire TIMEBOOST_net_2857;
wire n_10795;
wire n_10796;
wire n_10797;
wire n_10798;
wire n_10799;
wire n_108;
wire n_1080;
wire n_10800;
wire n_10801;
wire n_10802;
wire n_10803;
wire n_10804;
wire n_10805;
wire n_10806;
wire TIMEBOOST_net_1342;
wire n_10808;
wire n_10809;
wire n_1081;
wire n_10810;
wire n_10811;
wire n_10812;
wire n_10813;
wire n_10814;
wire n_10815;
wire n_10816;
wire n_10817;
wire n_10818;
wire n_1082;
wire TIMEBOOST_net_2722;
wire n_10821;
wire TIMEBOOST_net_2859;
wire n_10823;
wire n_10825;
wire n_10826;
wire n_10827;
wire n_10828;
wire n_10829;
wire n_1083;
wire n_10831;
wire n_10832;
wire n_10833;
wire n_10834;
wire n_10835;
wire n_10836;
wire n_1084;
wire n_10840;
wire n_10841;
wire n_10842;
wire n_10845;
wire n_10846;
wire n_10847;
wire n_10848;
wire n_10849;
wire n_1085;
wire n_10850;
wire n_10851;
wire n_10852;
wire n_10855;
wire n_10856;
wire n_10857;
wire TIMEBOOST_net_533;
wire n_1086;
wire TIMEBOOST_net_1729;
wire n_10861;
wire n_10862;
wire n_10863;
wire n_10864;
wire n_10865;
wire n_10868;
wire n_10869;
wire n_1087;
wire n_10871;
wire n_10872;
wire n_10874;
wire n_10875;
wire TIMEBOOST_net_1204;
wire n_10877;
wire n_10878;
wire n_10879;
wire n_1088;
wire n_10880;
wire n_10881;
wire TIMEBOOST_net_633;
wire n_10883;
wire n_10884;
wire n_10885;
wire TIMEBOOST_net_2661;
wire TIMEBOOST_net_1345;
wire n_10889;
wire n_1089;
wire n_10890;
wire n_10891;
wire n_10892;
wire n_10893;
wire n_10894;
wire TIMEBOOST_net_2285;
wire n_10896;
wire n_10897;
wire n_10898;
wire n_10899;
wire n_109;
wire n_1090;
wire n_10900;
wire n_10902;
wire n_10903;
wire n_10904;
wire n_10906;
wire n_10907;
wire n_10908;
wire TIMEBOOST_net_2697;
wire n_1091;
wire n_10910;
wire n_10912;
wire n_10913;
wire n_10914;
wire n_10915;
wire n_10917;
wire n_10918;
wire n_10919;
wire n_1092;
wire n_10920;
wire n_10921;
wire n_10922;
wire n_10923;
wire n_10925;
wire n_10926;
wire n_10927;
wire n_10928;
wire TIMEBOOST_net_726;
wire n_1093;
wire n_10930;
wire n_10931;
wire n_10932;
wire n_10933;
wire n_10934;
wire n_10935;
wire n_10936;
wire n_10939;
wire n_1094;
wire n_10940;
wire n_10941;
wire n_10942;
wire n_10943;
wire n_10944;
wire n_10945;
wire n_10946;
wire n_10948;
wire n_1095;
wire n_10950;
wire n_10951;
wire n_10952;
wire n_10953;
wire TIMEBOOST_net_1269;
wire n_10955;
wire n_10956;
wire n_10957;
wire n_10958;
wire n_10959;
wire n_1096;
wire n_10962;
wire n_10965;
wire n_10966;
wire TIMEBOOST_net_2644;
wire TIMEBOOST_net_1344;
wire n_1097;
wire n_10970;
wire n_10971;
wire n_10972;
wire n_10974;
wire TIMEBOOST_net_2953;
wire n_10977;
wire n_10978;
wire n_10979;
wire n_1098;
wire n_10980;
wire n_10981;
wire n_10982;
wire n_10983;
wire n_10984;
wire n_10985;
wire n_10986;
wire n_10987;
wire n_10988;
wire n_10989;
wire n_1099;
wire n_10991;
wire n_10992;
wire n_10993;
wire TIMEBOOST_net_1367;
wire n_10995;
wire n_10998;
wire n_11;
wire n_110;
wire n_1100;
wire n_11000;
wire n_11001;
wire n_11003;
wire n_11004;
wire n_11005;
wire n_11006;
wire n_11007;
wire n_11008;
wire n_1101;
wire TIMEBOOST_net_657;
wire n_11012;
wire n_11013;
wire n_11014;
wire n_11015;
wire n_11016;
wire n_11017;
wire n_11018;
wire n_11019;
wire n_1102;
wire n_11022;
wire n_11024;
wire n_11025;
wire n_11026;
wire n_11027;
wire n_11029;
wire n_1103;
wire n_11031;
wire n_11032;
wire n_11033;
wire n_11035;
wire n_11036;
wire n_11037;
wire n_1104;
wire n_11041;
wire n_11042;
wire n_11043;
wire n_11044;
wire n_11045;
wire n_11047;
wire n_11048;
wire n_11049;
wire n_1105;
wire TIMEBOOST_net_1063;
wire n_11052;
wire n_11053;
wire TIMEBOOST_net_1284;
wire n_11055;
wire n_11056;
wire n_11057;
wire n_11058;
wire n_11059;
wire n_1106;
wire n_11061;
wire TIMEBOOST_net_1287;
wire n_11063;
wire n_11064;
wire TIMEBOOST_net_1286;
wire n_11068;
wire n_11069;
wire n_1107;
wire n_11070;
wire n_11071;
wire n_11072;
wire n_11073;
wire n_11074;
wire n_11075;
wire n_11076;
wire n_11078;
wire n_1108;
wire n_11080;
wire n_11081;
wire n_11082;
wire n_11083;
wire n_11084;
wire n_11086;
wire n_11087;
wire n_11089;
wire n_1109;
wire TIMEBOOST_net_673;
wire TIMEBOOST_net_1637;
wire n_11096;
wire n_11097;
wire n_11098;
wire n_111;
wire n_1110;
wire n_11101;
wire n_11102;
wire n_11103;
wire n_11104;
wire n_11106;
wire n_11107;
wire TIMEBOOST_net_1395;
wire n_1111;
wire n_11110;
wire n_11112;
wire n_11113;
wire n_11114;
wire n_11118;
wire n_1112;
wire TIMEBOOST_net_636;
wire n_11122;
wire n_11123;
wire n_11124;
wire TIMEBOOST_net_660;
wire TIMEBOOST_net_728;
wire n_11128;
wire n_11129;
wire n_1113;
wire n_11130;
wire n_11131;
wire n_11132;
wire TIMEBOOST_net_733;
wire n_11134;
wire n_11136;
wire n_11137;
wire n_11138;
wire n_11139;
wire n_1114;
wire TIMEBOOST_net_1370;
wire n_11144;
wire n_11145;
wire n_11146;
wire n_11148;
wire n_1115;
wire TIMEBOOST_net_1356;
wire n_11151;
wire n_11152;
wire n_11153;
wire n_11154;
wire n_11156;
wire n_11157;
wire n_11158;
wire n_11159;
wire n_1116;
wire n_11161;
wire n_11162;
wire n_11164;
wire n_11165;
wire n_11166;
wire n_11167;
wire n_11168;
wire n_11169;
wire n_1117;
wire TIMEBOOST_net_1325;
wire n_11172;
wire n_11173;
wire TIMEBOOST_net_676;
wire n_11175;
wire TIMEBOOST_net_2878;
wire n_11177;
wire n_11178;
wire n_11179;
wire n_1118;
wire n_11180;
wire n_11181;
wire n_11183;
wire n_11184;
wire n_11187;
wire n_11189;
wire n_1119;
wire n_11190;
wire n_11191;
wire n_11192;
wire n_11193;
wire n_11194;
wire n_11195;
wire n_11196;
wire n_11197;
wire n_11198;
wire n_11199;
wire n_112;
wire n_1120;
wire n_11200;
wire n_11201;
wire n_11202;
wire TIMEBOOST_net_2649;
wire n_11205;
wire n_11208;
wire n_11209;
wire n_1121;
wire n_11210;
wire n_11211;
wire n_11212;
wire n_11213;
wire n_11214;
wire n_11215;
wire TIMEBOOST_net_732;
wire n_11217;
wire n_11218;
wire n_1122;
wire n_11220;
wire n_11221;
wire n_11223;
wire TIMEBOOST_net_2765;
wire n_11225;
wire n_11226;
wire n_11227;
wire n_11228;
wire n_11229;
wire n_1123;
wire n_11230;
wire n_11231;
wire n_11232;
wire n_11233;
wire n_11235;
wire n_11236;
wire n_11237;
wire n_11238;
wire n_11239;
wire n_1124;
wire n_11240;
wire n_11241;
wire n_11242;
wire n_11243;
wire n_11244;
wire n_11245;
wire n_11247;
wire TIMEBOOST_net_1371;
wire n_11249;
wire n_1125;
wire n_11251;
wire n_11252;
wire n_11254;
wire n_11256;
wire n_11257;
wire n_11258;
wire n_11259;
wire n_1126;
wire n_11260;
wire n_11261;
wire n_11262;
wire n_11263;
wire n_11264;
wire n_11265;
wire n_11266;
wire n_11267;
wire n_11268;
wire n_11269;
wire n_1127;
wire TIMEBOOST_net_743;
wire n_11271;
wire n_11272;
wire TIMEBOOST_net_2270;
wire n_11274;
wire n_11275;
wire TIMEBOOST_net_669;
wire n_11278;
wire n_1128;
wire n_11280;
wire n_11281;
wire n_11282;
wire n_11283;
wire n_11284;
wire n_11285;
wire n_11286;
wire n_11287;
wire n_11288;
wire n_11289;
wire n_1129;
wire n_11291;
wire n_11292;
wire n_11293;
wire n_11294;
wire n_11295;
wire n_11296;
wire n_11297;
wire n_11298;
wire n_11299;
wire n_113;
wire n_1130;
wire n_11301;
wire TIMEBOOST_net_1337;
wire n_11303;
wire n_11304;
wire n_11305;
wire n_11306;
wire n_11307;
wire n_11308;
wire n_1131;
wire n_11310;
wire n_11312;
wire n_11313;
wire n_11314;
wire n_11315;
wire n_11316;
wire n_11317;
wire n_11318;
wire n_1132;
wire n_11320;
wire n_11323;
wire n_11324;
wire n_11325;
wire n_11326;
wire n_11327;
wire n_11328;
wire n_1133;
wire n_11331;
wire n_11332;
wire n_11333;
wire n_11334;
wire n_11335;
wire n_11336;
wire n_11337;
wire n_11338;
wire n_1134;
wire n_11340;
wire n_11342;
wire n_11344;
wire n_11345;
wire TIMEBOOST_net_687;
wire n_11349;
wire n_1135;
wire n_11350;
wire n_11351;
wire n_11352;
wire n_11353;
wire TIMEBOOST_net_686;
wire n_11355;
wire n_11356;
wire n_11357;
wire n_11358;
wire n_11359;
wire n_1136;
wire n_11360;
wire n_11361;
wire n_11362;
wire n_11363;
wire n_11364;
wire n_11366;
wire n_11367;
wire n_11369;
wire n_1137;
wire n_11370;
wire n_11371;
wire n_11372;
wire n_11374;
wire n_11375;
wire n_11376;
wire n_11377;
wire n_11378;
wire n_11379;
wire n_1138;
wire n_11380;
wire n_11381;
wire n_11383;
wire n_11384;
wire n_11385;
wire n_11386;
wire TIMEBOOST_net_749;
wire n_11388;
wire n_11389;
wire n_1139;
wire TIMEBOOST_net_1506;
wire n_11392;
wire n_11394;
wire n_11395;
wire n_11396;
wire n_11398;
wire n_11399;
wire n_114;
wire n_1140;
wire n_11400;
wire n_11402;
wire n_11403;
wire n_11405;
wire n_11407;
wire n_11409;
wire n_1141;
wire n_11410;
wire n_11411;
wire n_11412;
wire n_11413;
wire n_11414;
wire n_11415;
wire n_11416;
wire n_11419;
wire n_1142;
wire n_11420;
wire n_11422;
wire n_11425;
wire n_11426;
wire n_11427;
wire n_11429;
wire n_1143;
wire n_11430;
wire n_11433;
wire n_11434;
wire n_11435;
wire TIMEBOOST_net_2510;
wire TIMEBOOST_net_683;
wire n_11439;
wire n_1144;
wire n_1145;
wire n_11451;
wire n_11453;
wire n_11454;
wire n_11456;
wire n_11458;
wire n_11459;
wire n_1146;
wire n_11463;
wire n_11464;
wire n_11465;
wire n_1147;
wire n_11473;
wire n_11474;
wire n_11475;
wire n_11476;
wire n_11477;
wire n_11478;
wire n_11479;
wire n_1148;
wire n_11480;
wire n_11481;
wire n_11482;
wire TIMEBOOST_net_2793;
wire n_11484;
wire n_11485;
wire n_11486;
wire n_1149;
wire n_11490;
wire n_11492;
wire n_11494;
wire n_11495;
wire n_11497;
wire n_11498;
wire TIMEBOOST_net_2290;
wire n_115;
wire n_1150;
wire n_11500;
wire n_11501;
wire n_11503;
wire n_11504;
wire n_11507;
wire n_11509;
wire n_1151;
wire n_11510;
wire n_11511;
wire n_11514;
wire n_11516;
wire n_11517;
wire n_11518;
wire TIMEBOOST_net_2881;
wire n_1152;
wire n_11520;
wire n_11523;
wire n_11524;
wire n_11525;
wire n_11527;
wire n_11528;
wire n_1153;
wire n_11530;
wire n_11532;
wire n_11535;
wire n_11537;
wire n_11538;
wire n_1154;
wire n_11542;
wire n_11543;
wire n_11544;
wire n_11546;
wire n_11547;
wire n_11548;
wire n_11549;
wire n_1155;
wire TIMEBOOST_net_752;
wire n_11552;
wire n_11553;
wire n_11555;
wire n_11557;
wire n_1156;
wire n_11560;
wire n_11568;
wire n_11569;
wire n_1157;
wire n_11570;
wire n_11571;
wire n_11575;
wire n_11578;
wire n_11579;
wire n_1158;
wire n_11580;
wire n_11581;
wire n_11582;
wire TIMEBOOST_net_703;
wire TIMEBOOST_net_2782;
wire n_11586;
wire n_11587;
wire n_11588;
wire n_11589;
wire n_1159;
wire n_11590;
wire n_11593;
wire n_11595;
wire n_11596;
wire n_11597;
wire n_11598;
wire n_11599;
wire n_116;
wire n_1160;
wire n_11600;
wire n_11601;
wire n_11602;
wire n_11603;
wire n_11604;
wire n_11605;
wire n_11606;
wire n_11607;
wire n_11608;
wire n_1161;
wire n_11611;
wire n_11613;
wire n_11617;
wire TIMEBOOST_net_2483;
wire n_1162;
wire n_11620;
wire TIMEBOOST_net_1793;
wire n_11622;
wire n_11623;
wire n_11624;
wire n_11626;
wire TIMEBOOST_net_1446;
wire TIMEBOOST_net_2105;
wire n_1163;
wire n_11630;
wire n_11631;
wire n_11632;
wire n_11633;
wire n_11634;
wire n_11635;
wire n_11636;
wire n_11637;
wire n_11638;
wire n_11639;
wire n_1164;
wire n_11640;
wire TIMEBOOST_net_1458;
wire n_11643;
wire TIMEBOOST_net_701;
wire n_11647;
wire n_11648;
wire n_11649;
wire n_1165;
wire TIMEBOOST_net_1794;
wire n_11652;
wire n_11654;
wire n_11655;
wire n_11656;
wire n_11657;
wire n_11658;
wire n_11659;
wire n_1166;
wire n_11661;
wire n_11662;
wire n_11663;
wire n_11664;
wire n_11665;
wire n_11669;
wire n_1167;
wire n_11671;
wire n_11673;
wire TIMEBOOST_net_702;
wire n_11675;
wire n_11676;
wire n_11677;
wire n_11678;
wire n_1168;
wire n_11680;
wire n_11681;
wire n_11682;
wire n_11685;
wire n_11686;
wire n_11687;
wire n_11689;
wire n_1169;
wire n_11693;
wire n_11694;
wire n_11696;
wire TIMEBOOST_net_2738;
wire n_11698;
wire n_11699;
wire n_117;
wire n_1170;
wire n_11700;
wire n_11701;
wire n_11702;
wire n_11704;
wire n_11707;
wire n_11709;
wire n_1171;
wire n_11710;
wire n_11711;
wire n_11712;
wire n_11713;
wire n_11715;
wire n_11716;
wire n_11718;
wire n_1172;
wire n_11723;
wire n_11725;
wire n_11726;
wire n_11727;
wire n_11728;
wire n_11729;
wire n_1173;
wire n_11730;
wire n_11731;
wire n_11734;
wire n_11735;
wire n_11736;
wire n_11737;
wire n_11738;
wire n_11739;
wire n_1174;
wire n_11740;
wire n_11741;
wire n_11742;
wire n_11743;
wire n_11744;
wire n_11745;
wire n_11746;
wire n_11747;
wire n_11748;
wire n_11749;
wire n_1175;
wire n_11750;
wire n_11751;
wire n_11752;
wire n_11753;
wire n_11754;
wire n_11756;
wire n_11757;
wire n_11758;
wire n_11759;
wire n_1176;
wire n_11760;
wire n_11761;
wire n_11762;
wire n_11763;
wire n_11764;
wire n_11765;
wire n_11766;
wire n_11767;
wire n_11769;
wire n_1177;
wire n_11770;
wire n_11771;
wire n_11772;
wire n_11773;
wire n_11774;
wire n_11775;
wire n_11776;
wire n_11777;
wire n_11778;
wire n_1178;
wire n_11780;
wire n_11784;
wire n_11786;
wire n_11787;
wire n_11788;
wire n_1179;
wire TIMEBOOST_net_751;
wire n_11794;
wire n_11795;
wire n_11796;
wire n_11797;
wire n_11798;
wire n_11799;
wire n_118;
wire n_1180;
wire n_11800;
wire n_11801;
wire n_11802;
wire n_11803;
wire n_11804;
wire n_11805;
wire n_11806;
wire n_11807;
wire n_11808;
wire n_11809;
wire n_1181;
wire n_11810;
wire n_11813;
wire n_11814;
wire n_11815;
wire n_11816;
wire n_11817;
wire n_11818;
wire n_11819;
wire n_1182;
wire n_11821;
wire n_11822;
wire n_11823;
wire n_11825;
wire n_11829;
wire n_1183;
wire n_11833;
wire n_11834;
wire n_11835;
wire n_11836;
wire n_11838;
wire n_1184;
wire n_11840;
wire n_11841;
wire n_11842;
wire n_11843;
wire n_11844;
wire n_11845;
wire n_11846;
wire n_11847;
wire n_11848;
wire n_1185;
wire n_11850;
wire n_11852;
wire n_11853;
wire n_11856;
wire n_1186;
wire n_11860;
wire n_11863;
wire n_11866;
wire n_11867;
wire n_11868;
wire n_1187;
wire n_11870;
wire n_11871;
wire n_11872;
wire n_11873;
wire n_11874;
wire n_11875;
wire n_11876;
wire n_11877;
wire n_11878;
wire n_11879;
wire n_1188;
wire n_11880;
wire n_11881;
wire n_11882;
wire n_11883;
wire n_11884;
wire n_11885;
wire n_11886;
wire n_11888;
wire n_11889;
wire n_1189;
wire n_11890;
wire n_11892;
wire n_11893;
wire n_11894;
wire n_11895;
wire n_11896;
wire n_11897;
wire n_11898;
wire n_11899;
wire n_119;
wire n_1190;
wire n_11900;
wire n_11901;
wire n_11907;
wire n_11908;
wire n_11909;
wire n_1191;
wire n_11910;
wire n_11913;
wire n_11914;
wire n_11915;
wire TIMEBOOST_net_718;
wire n_11917;
wire n_11918;
wire n_11919;
wire n_1192;
wire TIMEBOOST_net_2103;
wire n_11922;
wire n_11923;
wire n_11924;
wire n_11925;
wire n_11927;
wire n_11929;
wire TIMEBOOST_net_778;
wire n_11933;
wire n_11934;
wire n_11935;
wire n_11936;
wire n_11938;
wire n_11939;
wire n_1194;
wire n_11941;
wire n_11943;
wire n_11944;
wire n_11945;
wire n_11946;
wire n_11947;
wire n_1195;
wire TIMEBOOST_net_2886;
wire n_11952;
wire n_11953;
wire n_11954;
wire n_11955;
wire n_11956;
wire n_11957;
wire n_11958;
wire n_11959;
wire n_1196;
wire n_11960;
wire n_11962;
wire n_11964;
wire n_11966;
wire TIMEBOOST_net_822;
wire n_11968;
wire n_1197;
wire n_11970;
wire n_11971;
wire n_11972;
wire n_11973;
wire n_11974;
wire n_11975;
wire n_11976;
wire n_11978;
wire n_1198;
wire n_11980;
wire n_11982;
wire n_11983;
wire n_11984;
wire n_11985;
wire n_11986;
wire n_11987;
wire n_11988;
wire n_11989;
wire n_1199;
wire n_11990;
wire n_11991;
wire TIMEBOOST_net_2799;
wire n_11993;
wire n_11994;
wire n_11996;
wire n_11997;
wire n_11998;
wire n_11999;
wire n_12;
wire n_120;
wire n_1200;
wire n_12003;
wire n_12005;
wire n_12007;
wire n_12008;
wire n_1201;
wire n_12011;
wire n_12013;
wire n_12014;
wire n_12016;
wire n_12017;
wire n_12019;
wire n_12020;
wire n_12021;
wire n_12022;
wire n_12023;
wire n_12024;
wire n_12025;
wire n_12026;
wire n_12027;
wire n_12028;
wire n_12029;
wire n_1203;
wire n_12030;
wire n_12031;
wire n_12033;
wire n_12034;
wire n_12035;
wire n_12036;
wire n_12037;
wire n_12038;
wire n_12039;
wire n_1204;
wire n_12041;
wire n_12042;
wire n_12043;
wire n_12046;
wire n_12047;
wire n_12048;
wire n_12049;
wire n_1205;
wire n_12050;
wire n_12051;
wire n_12053;
wire n_12054;
wire n_12055;
wire n_12056;
wire n_12058;
wire n_12059;
wire n_1206;
wire n_12060;
wire n_12061;
wire n_12062;
wire n_12064;
wire n_12065;
wire n_12067;
wire n_12068;
wire n_12069;
wire n_1207;
wire n_12071;
wire n_12072;
wire n_12076;
wire n_12077;
wire n_12078;
wire n_12079;
wire n_1208;
wire n_12080;
wire n_12081;
wire n_12082;
wire n_12083;
wire n_12084;
wire n_12085;
wire n_12086;
wire n_12087;
wire n_12088;
wire n_12089;
wire n_12091;
wire n_12092;
wire n_12093;
wire n_12094;
wire n_12095;
wire n_12096;
wire n_12097;
wire n_12098;
wire n_12099;
wire n_121;
wire n_1210;
wire n_12100;
wire n_12102;
wire n_12104;
wire n_12105;
wire n_12106;
wire n_12108;
wire n_1211;
wire n_12110;
wire n_12111;
wire n_12112;
wire n_12114;
wire n_12115;
wire n_12116;
wire n_12117;
wire n_12119;
wire n_1212;
wire n_12121;
wire n_12122;
wire n_12123;
wire n_12124;
wire n_12125;
wire n_12126;
wire n_12127;
wire n_12128;
wire n_12129;
wire n_1213;
wire n_12130;
wire n_12131;
wire n_12132;
wire n_12133;
wire n_12134;
wire n_12135;
wire n_12136;
wire n_12137;
wire n_12139;
wire n_1214;
wire n_12140;
wire n_12141;
wire n_12144;
wire n_12145;
wire n_12146;
wire n_12147;
wire n_12148;
wire n_12149;
wire n_1215;
wire n_12150;
wire n_12151;
wire n_12153;
wire n_12154;
wire n_12155;
wire n_12157;
wire n_12158;
wire n_1216;
wire n_12161;
wire n_12162;
wire n_12164;
wire n_12165;
wire n_12166;
wire n_12168;
wire n_1217;
wire n_12170;
wire n_12173;
wire n_12174;
wire n_12175;
wire n_12176;
wire n_12177;
wire n_12178;
wire n_12179;
wire n_1218;
wire n_12180;
wire n_12181;
wire n_12182;
wire n_12183;
wire n_12185;
wire n_12186;
wire n_12187;
wire n_12188;
wire n_12189;
wire n_1219;
wire n_12190;
wire n_12191;
wire n_12192;
wire n_12193;
wire n_12195;
wire n_12196;
wire n_12197;
wire n_12198;
wire n_12199;
wire n_122;
wire n_1220;
wire n_12200;
wire n_12201;
wire n_12202;
wire n_12203;
wire n_12204;
wire n_12205;
wire n_12207;
wire n_12208;
wire n_12209;
wire n_12211;
wire n_12212;
wire n_12213;
wire n_12214;
wire n_12215;
wire n_12217;
wire n_12218;
wire n_12219;
wire n_1222;
wire n_12220;
wire n_12221;
wire n_12222;
wire n_12223;
wire n_12224;
wire n_12225;
wire n_12228;
wire n_12229;
wire TIMEBOOST_net_478;
wire n_12230;
wire n_12231;
wire n_12232;
wire n_12233;
wire n_12234;
wire TIMEBOOST_net_1470;
wire TIMEBOOST_net_2127;
wire n_12238;
wire n_12239;
wire n_1224;
wire n_12240;
wire n_12241;
wire n_12242;
wire n_12243;
wire n_12245;
wire n_12247;
wire n_12248;
wire n_12249;
wire n_1225;
wire n_12250;
wire n_12251;
wire n_12252;
wire n_12253;
wire n_12254;
wire n_12255;
wire n_12256;
wire n_12257;
wire n_1226;
wire n_12260;
wire n_12261;
wire n_12262;
wire n_12263;
wire n_12264;
wire n_12265;
wire n_12266;
wire n_12267;
wire n_12268;
wire n_12269;
wire n_12270;
wire n_12271;
wire n_12273;
wire n_12275;
wire n_12278;
wire n_12279;
wire n_1228;
wire n_12281;
wire n_12283;
wire n_12284;
wire n_12285;
wire n_12286;
wire n_12287;
wire n_12288;
wire n_12289;
wire n_1229;
wire n_12290;
wire n_12291;
wire n_12292;
wire n_12293;
wire n_12294;
wire n_12295;
wire n_12296;
wire n_12297;
wire n_12298;
wire n_12299;
wire n_123;
wire n_1230;
wire n_12300;
wire n_12302;
wire n_12309;
wire n_1231;
wire n_12311;
wire n_12312;
wire n_12313;
wire n_12314;
wire n_12315;
wire n_12316;
wire n_12318;
wire n_12319;
wire n_1232;
wire n_12320;
wire n_12321;
wire n_12322;
wire n_12323;
wire n_12324;
wire n_12325;
wire n_12326;
wire n_12327;
wire n_12328;
wire n_12329;
wire n_1233;
wire n_12331;
wire n_12332;
wire n_12333;
wire n_12334;
wire n_12335;
wire n_12336;
wire n_12338;
wire n_12339;
wire n_1234;
wire n_12341;
wire n_12342;
wire n_12345;
wire n_12346;
wire n_12347;
wire n_12349;
wire n_1235;
wire n_12350;
wire n_12352;
wire n_12353;
wire n_12354;
wire n_12355;
wire n_12356;
wire n_12357;
wire n_12358;
wire n_12360;
wire n_12361;
wire n_12362;
wire n_12363;
wire n_12364;
wire n_12365;
wire n_12366;
wire n_12368;
wire n_1237;
wire n_12370;
wire n_12371;
wire n_12372;
wire n_12373;
wire n_12374;
wire n_12376;
wire n_12377;
wire n_12378;
wire n_12379;
wire n_1238;
wire n_12381;
wire TIMEBOOST_net_1493;
wire n_12384;
wire n_12385;
wire n_12386;
wire n_12387;
wire n_12388;
wire n_12389;
wire n_1239;
wire TIMEBOOST_net_831;
wire n_12391;
wire n_12392;
wire n_12393;
wire n_12394;
wire n_12396;
wire n_12398;
wire n_124;
wire TIMEBOOST_net_2847;
wire n_12400;
wire n_12401;
wire n_12402;
wire n_12404;
wire n_12406;
wire n_12408;
wire n_12409;
wire n_1241;
wire n_12411;
wire n_12412;
wire n_12413;
wire n_12414;
wire n_12415;
wire n_12416;
wire TIMEBOOST_net_1697;
wire n_12418;
wire n_12419;
wire n_1242;
wire n_12420;
wire n_12423;
wire n_12424;
wire n_12427;
wire n_12428;
wire n_12429;
wire n_1243;
wire n_12430;
wire n_12431;
wire n_12432;
wire n_12433;
wire n_12434;
wire n_12435;
wire n_12436;
wire n_12437;
wire n_12438;
wire n_1244;
wire n_12440;
wire n_12441;
wire n_12442;
wire n_12443;
wire n_12444;
wire n_12445;
wire n_12447;
wire n_12448;
wire n_12449;
wire n_1245;
wire n_12450;
wire n_12452;
wire n_12453;
wire n_12454;
wire n_12455;
wire n_12456;
wire n_12457;
wire n_12458;
wire n_12459;
wire n_1246;
wire n_12460;
wire n_12461;
wire n_12462;
wire n_12463;
wire n_12464;
wire n_12465;
wire TIMEBOOST_net_892;
wire n_12467;
wire n_12468;
wire n_12469;
wire n_12470;
wire n_12471;
wire n_12472;
wire n_12474;
wire n_12475;
wire n_12476;
wire n_12477;
wire n_12478;
wire n_12479;
wire n_1248;
wire n_12480;
wire n_12481;
wire n_12482;
wire n_12483;
wire n_12484;
wire n_12485;
wire n_12486;
wire n_12487;
wire n_12488;
wire n_12489;
wire n_1249;
wire n_12490;
wire n_12491;
wire n_12492;
wire n_12493;
wire n_12494;
wire n_12495;
wire n_12496;
wire n_12497;
wire n_12498;
wire n_12499;
wire n_125;
wire n_1250;
wire n_12500;
wire n_12501;
wire n_12502;
wire n_12503;
wire n_12504;
wire n_12505;
wire n_12506;
wire n_12507;
wire n_12508;
wire n_12509;
wire n_1251;
wire n_12510;
wire n_12512;
wire n_12513;
wire n_12514;
wire n_12515;
wire n_12516;
wire n_12517;
wire n_12519;
wire n_12520;
wire n_12521;
wire n_12522;
wire n_12523;
wire n_12524;
wire TIMEBOOST_net_915;
wire n_12526;
wire n_12527;
wire n_12528;
wire n_12529;
wire n_1253;
wire n_12530;
wire n_12531;
wire TIMEBOOST_net_902;
wire n_12533;
wire n_12534;
wire n_12535;
wire n_12537;
wire n_12538;
wire n_12539;
wire n_1254;
wire n_12540;
wire n_12541;
wire n_12542;
wire n_12543;
wire n_12544;
wire n_12545;
wire n_12546;
wire n_12547;
wire n_12549;
wire n_1255;
wire n_12550;
wire n_12551;
wire n_12552;
wire n_12553;
wire n_12554;
wire n_12555;
wire n_12558;
wire n_12559;
wire n_1256;
wire n_12560;
wire n_12561;
wire n_12562;
wire n_12563;
wire n_12564;
wire n_12565;
wire n_12567;
wire n_12568;
wire n_12569;
wire n_1257;
wire n_12570;
wire n_12571;
wire n_12572;
wire n_12573;
wire n_12574;
wire n_12575;
wire n_12576;
wire n_12577;
wire n_12578;
wire n_12579;
wire TIMEBOOST_net_515;
wire n_12580;
wire n_12581;
wire TIMEBOOST_net_918;
wire n_12583;
wire n_12584;
wire n_12585;
wire n_12586;
wire n_12587;
wire n_12588;
wire n_12589;
wire n_1259;
wire n_12590;
wire n_12591;
wire n_12592;
wire n_12593;
wire n_12596;
wire n_12597;
wire n_12598;
wire n_12599;
wire n_126;
wire n_1260;
wire n_12600;
wire n_12602;
wire n_12603;
wire n_12604;
wire n_12605;
wire n_12606;
wire n_12607;
wire n_12608;
wire n_1261;
wire n_12610;
wire n_12611;
wire n_12612;
wire n_12613;
wire n_12614;
wire n_12615;
wire n_12616;
wire n_12617;
wire n_12618;
wire n_12619;
wire n_1262;
wire n_12620;
wire n_12621;
wire n_12622;
wire n_12623;
wire n_12627;
wire n_12628;
wire n_12629;
wire n_1263;
wire n_12630;
wire n_12631;
wire n_12632;
wire n_12633;
wire n_12634;
wire n_12635;
wire n_12638;
wire n_1264;
wire n_12640;
wire n_12641;
wire n_12642;
wire n_12643;
wire n_12644;
wire n_12645;
wire n_12646;
wire n_12647;
wire n_12648;
wire n_12651;
wire n_12652;
wire TIMEBOOST_net_957;
wire n_12654;
wire n_12655;
wire n_12656;
wire n_12657;
wire n_12658;
wire n_12659;
wire n_1266;
wire n_12660;
wire n_12662;
wire n_12663;
wire n_12664;
wire n_12666;
wire n_12667;
wire n_12668;
wire TIMEBOOST_net_81;
wire n_1267;
wire TIMEBOOST_net_1469;
wire n_12671;
wire n_12672;
wire n_12673;
wire n_12674;
wire n_12675;
wire n_12676;
wire n_12678;
wire n_12679;
wire n_1268;
wire n_12680;
wire n_12681;
wire n_12682;
wire n_12683;
wire n_12684;
wire TIMEBOOST_net_2543;
wire n_12686;
wire n_12688;
wire n_12689;
wire n_1269;
wire n_12690;
wire n_12691;
wire n_12692;
wire n_12693;
wire n_12694;
wire n_12695;
wire n_12696;
wire n_12697;
wire n_12698;
wire n_12699;
wire n_127;
wire n_1270;
wire n_12700;
wire n_12701;
wire n_12702;
wire n_12703;
wire n_12704;
wire n_12705;
wire n_12706;
wire n_12707;
wire n_12708;
wire n_1271;
wire n_12710;
wire n_12711;
wire n_12712;
wire n_12713;
wire n_12714;
wire n_12716;
wire n_12717;
wire n_12718;
wire n_12719;
wire n_1272;
wire n_12720;
wire n_12722;
wire n_12723;
wire n_12724;
wire n_12725;
wire n_12727;
wire n_12728;
wire n_12729;
wire n_1273;
wire n_12730;
wire n_12731;
wire n_12733;
wire n_12734;
wire n_12735;
wire n_12736;
wire n_12737;
wire n_12738;
wire n_1274;
wire n_12740;
wire n_12741;
wire n_12742;
wire n_12743;
wire n_12744;
wire n_12745;
wire n_12746;
wire n_12747;
wire n_12748;
wire n_12749;
wire n_1275;
wire n_12750;
wire n_12753;
wire n_12755;
wire n_12756;
wire n_12759;
wire n_12760;
wire n_12761;
wire n_12762;
wire n_12763;
wire n_12764;
wire n_12765;
wire n_12766;
wire n_12767;
wire n_12768;
wire TIMEBOOST_net_2569;
wire n_12770;
wire n_12771;
wire n_12772;
wire n_12773;
wire n_12774;
wire n_12775;
wire n_12776;
wire n_12781;
wire n_12782;
wire n_12783;
wire n_12784;
wire n_12786;
wire n_12787;
wire n_12788;
wire n_12789;
wire n_12790;
wire n_12793;
wire n_12794;
wire n_12795;
wire n_12796;
wire TIMEBOOST_net_1882;
wire n_12798;
wire n_12799;
wire n_128;
wire n_12800;
wire TIMEBOOST_net_122;
wire n_12802;
wire n_12803;
wire n_12804;
wire n_12805;
wire n_12807;
wire n_12808;
wire n_12809;
wire n_12810;
wire n_12811;
wire n_12813;
wire n_12815;
wire n_12816;
wire n_12817;
wire TIMEBOOST_net_88;
wire n_12819;
wire n_1282;
wire n_12820;
wire n_12821;
wire n_12822;
wire n_12823;
wire n_12824;
wire n_12825;
wire n_12826;
wire n_12829;
wire n_12830;
wire n_12831;
wire n_12832;
wire n_12834;
wire n_12836;
wire n_12838;
wire n_12840;
wire n_12841;
wire n_12843;
wire n_12844;
wire n_12845;
wire n_12846;
wire n_12847;
wire n_12848;
wire n_12849;
wire n_1285;
wire n_12850;
wire n_12852;
wire n_12853;
wire n_12854;
wire n_12855;
wire n_12856;
wire n_12857;
wire n_1286;
wire n_12860;
wire n_12861;
wire n_12863;
wire n_12864;
wire n_12865;
wire n_12866;
wire n_12867;
wire n_12868;
wire n_12869;
wire n_1287;
wire n_12870;
wire n_12871;
wire n_12873;
wire n_12875;
wire n_12877;
wire n_12879;
wire n_1288;
wire n_12880;
wire n_12881;
wire n_12882;
wire n_12883;
wire n_12884;
wire n_12885;
wire n_12886;
wire n_12887;
wire n_12888;
wire n_12889;
wire n_1289;
wire n_12890;
wire n_12891;
wire n_12892;
wire n_12898;
wire n_12899;
wire n_129;
wire n_12900;
wire n_12902;
wire TIMEBOOST_net_1555;
wire n_12904;
wire n_12905;
wire n_12907;
wire n_12909;
wire n_1291;
wire n_12910;
wire n_12911;
wire n_12916;
wire n_12917;
wire n_12918;
wire n_12919;
wire n_1292;
wire n_12920;
wire n_12921;
wire n_12923;
wire n_12924;
wire n_12925;
wire n_12926;
wire n_12929;
wire n_12932;
wire n_12935;
wire n_12937;
wire n_12938;
wire n_12939;
wire n_1294;
wire n_12940;
wire n_12941;
wire n_12942;
wire n_12943;
wire n_12947;
wire n_12948;
wire n_12949;
wire n_1295;
wire TIMEBOOST_net_2936;
wire n_12951;
wire n_12954;
wire n_12955;
wire n_12956;
wire n_12958;
wire n_12961;
wire n_12962;
wire n_12963;
wire n_12964;
wire n_12965;
wire n_12967;
wire n_12968;
wire n_12969;
wire n_1297;
wire n_12975;
wire TIMEBOOST_net_2168;
wire n_12977;
wire n_12978;
wire n_1298;
wire n_12980;
wire n_12981;
wire n_12982;
wire n_12983;
wire n_12985;
wire n_12986;
wire n_12987;
wire n_12988;
wire n_1299;
wire n_12990;
wire n_12992;
wire n_12993;
wire n_12994;
wire n_12995;
wire n_12996;
wire n_12997;
wire n_12998;
wire n_12999;
wire n_13;
wire n_130;
wire n_1300;
wire n_13000;
wire n_13002;
wire n_13004;
wire n_13005;
wire n_13006;
wire n_13008;
wire n_13009;
wire n_1301;
wire n_13010;
wire n_13011;
wire n_13013;
wire n_13014;
wire n_13015;
wire n_13016;
wire n_13018;
wire n_13019;
wire n_1302;
wire n_13020;
wire n_13022;
wire n_13023;
wire n_13024;
wire n_13025;
wire n_13028;
wire n_13029;
wire n_1303;
wire n_13031;
wire n_13032;
wire n_13033;
wire n_13034;
wire n_13035;
wire n_13036;
wire n_13037;
wire n_13038;
wire n_13039;
wire n_1304;
wire n_13040;
wire n_13041;
wire n_13043;
wire n_13044;
wire n_13045;
wire n_13046;
wire n_13047;
wire n_13048;
wire n_13050;
wire n_13051;
wire n_13052;
wire n_13053;
wire n_13054;
wire n_13055;
wire n_13056;
wire n_13057;
wire n_13058;
wire n_13059;
wire n_1306;
wire n_13060;
wire n_13062;
wire n_13063;
wire n_13064;
wire n_13065;
wire n_13066;
wire n_1307;
wire n_13073;
wire n_13074;
wire n_13075;
wire n_13076;
wire n_13077;
wire n_13078;
wire n_13079;
wire n_1308;
wire n_13080;
wire n_13082;
wire n_13083;
wire n_13084;
wire n_13086;
wire n_13087;
wire n_13088;
wire n_1309;
wire n_13093;
wire n_13094;
wire n_13095;
wire n_13096;
wire n_13097;
wire n_13098;
wire n_13099;
wire n_131;
wire n_13100;
wire n_13101;
wire n_13103;
wire n_13104;
wire n_13109;
wire n_1311;
wire n_13110;
wire n_13111;
wire n_13112;
wire n_13113;
wire n_13114;
wire n_13115;
wire n_13116;
wire n_13118;
wire n_13119;
wire n_1312;
wire n_13120;
wire n_13121;
wire n_13122;
wire n_13124;
wire n_13126;
wire n_13127;
wire n_13129;
wire n_13130;
wire n_13131;
wire n_13132;
wire n_13133;
wire n_13134;
wire n_13135;
wire n_13136;
wire n_13137;
wire n_13138;
wire n_13139;
wire n_1314;
wire n_13140;
wire n_13141;
wire n_13142;
wire n_13143;
wire n_13144;
wire n_13145;
wire n_13146;
wire n_13148;
wire n_1315;
wire n_13150;
wire n_13151;
wire n_13153;
wire n_13154;
wire n_13156;
wire n_13157;
wire n_13159;
wire n_1316;
wire n_13160;
wire n_13161;
wire n_13162;
wire n_13163;
wire n_13164;
wire n_13165;
wire n_13166;
wire n_13167;
wire n_13168;
wire n_1317;
wire n_13171;
wire n_13172;
wire n_13173;
wire n_13175;
wire n_13176;
wire n_13177;
wire n_13178;
wire n_13179;
wire n_13180;
wire n_13183;
wire n_13190;
wire n_13192;
wire n_13193;
wire n_13195;
wire n_13196;
wire n_13197;
wire n_13198;
wire n_13199;
wire n_132;
wire n_1320;
wire n_13200;
wire n_13201;
wire n_13202;
wire n_13203;
wire n_13204;
wire n_13206;
wire n_13207;
wire n_13208;
wire n_13209;
wire n_13210;
wire n_13211;
wire n_13212;
wire n_13213;
wire n_13215;
wire n_13216;
wire n_13217;
wire n_1322;
wire n_13221;
wire n_13222;
wire n_13223;
wire n_13224;
wire n_13225;
wire n_13226;
wire n_13227;
wire n_13228;
wire n_13229;
wire n_13230;
wire TIMEBOOST_net_2816;
wire n_13232;
wire n_13234;
wire n_13235;
wire n_13236;
wire n_13238;
wire n_13239;
wire n_1324;
wire n_13241;
wire n_13242;
wire n_13243;
wire n_13244;
wire n_13245;
wire n_13248;
wire n_13249;
wire n_1325;
wire n_13251;
wire n_13252;
wire n_13253;
wire n_13255;
wire n_13256;
wire n_13257;
wire n_13259;
wire n_13260;
wire n_13261;
wire n_13262;
wire n_13264;
wire n_13265;
wire n_13266;
wire n_13267;
wire n_13268;
wire n_13269;
wire n_1327;
wire n_13270;
wire n_13271;
wire n_13272;
wire n_13273;
wire n_13274;
wire n_13275;
wire n_13277;
wire n_13278;
wire n_13279;
wire n_1328;
wire n_13280;
wire n_13281;
wire n_13282;
wire n_13284;
wire n_13285;
wire n_13286;
wire n_13287;
wire n_13288;
wire n_13289;
wire n_1329;
wire n_13290;
wire n_13291;
wire n_13292;
wire n_13293;
wire n_13294;
wire n_13295;
wire n_13296;
wire n_13297;
wire n_13298;
wire n_13299;
wire n_133;
wire n_13301;
wire n_13302;
wire n_13303;
wire n_13305;
wire n_13306;
wire n_13307;
wire n_13310;
wire TIMEBOOST_net_962;
wire n_13312;
wire n_13313;
wire n_13314;
wire n_13315;
wire n_13316;
wire n_13319;
wire n_1332;
wire n_13320;
wire n_13321;
wire n_13322;
wire n_13323;
wire n_13324;
wire n_13325;
wire TIMEBOOST_net_105;
wire n_13329;
wire n_1333;
wire n_13330;
wire n_13331;
wire n_13332;
wire TIMEBOOST_net_1876;
wire n_13334;
wire n_13335;
wire n_13336;
wire n_13338;
wire n_1334;
wire n_13343;
wire n_13344;
wire n_13346;
wire n_13347;
wire n_13349;
wire n_1335;
wire n_13350;
wire n_13351;
wire n_13352;
wire n_13353;
wire n_13354;
wire n_13355;
wire n_13356;
wire n_13357;
wire n_13358;
wire n_13359;
wire n_1336;
wire n_13360;
wire n_13361;
wire n_13362;
wire n_13363;
wire n_13364;
wire n_13365;
wire n_13366;
wire n_13367;
wire n_13369;
wire n_1337;
wire n_13370;
wire n_13371;
wire n_13375;
wire n_13376;
wire n_13377;
wire n_13378;
wire n_13379;
wire n_1338;
wire n_13380;
wire n_13381;
wire n_13382;
wire n_13383;
wire n_13384;
wire n_13385;
wire n_13386;
wire n_13388;
wire n_13390;
wire n_13391;
wire n_13392;
wire n_13393;
wire n_13394;
wire n_13395;
wire n_13396;
wire n_13397;
wire n_13398;
wire n_13399;
wire n_134;
wire n_1340;
wire n_13400;
wire n_13401;
wire n_13402;
wire n_13403;
wire n_13405;
wire n_13406;
wire n_13407;
wire n_13408;
wire n_13409;
wire n_13410;
wire n_13411;
wire n_13412;
wire n_13413;
wire TIMEBOOST_net_2954;
wire TIMEBOOST_net_2814;
wire n_13417;
wire n_13418;
wire n_13419;
wire n_13420;
wire n_13421;
wire n_13422;
wire n_13423;
wire n_13424;
wire n_13425;
wire n_13426;
wire n_13427;
wire n_13429;
wire n_1343;
wire n_13430;
wire n_13431;
wire TIMEBOOST_net_979;
wire n_13433;
wire n_13434;
wire n_13435;
wire n_13436;
wire n_13437;
wire TIMEBOOST_net_966;
wire n_13440;
wire n_13441;
wire n_13442;
wire n_13443;
wire n_13444;
wire n_13445;
wire n_13446;
wire n_13447;
wire n_13448;
wire n_13449;
wire n_1345;
wire n_13450;
wire n_13451;
wire n_13452;
wire n_13453;
wire TIMEBOOST_net_174;
wire n_13456;
wire n_13458;
wire n_13459;
wire n_1346;
wire n_13460;
wire n_13462;
wire n_13463;
wire n_13464;
wire n_13468;
wire n_13469;
wire n_13470;
wire n_13471;
wire n_13472;
wire n_13473;
wire n_13474;
wire n_13475;
wire n_13476;
wire n_13478;
wire n_13479;
wire n_1348;
wire n_13480;
wire TIMEBOOST_net_172;
wire n_13482;
wire n_13483;
wire n_13487;
wire n_13488;
wire n_13489;
wire n_13490;
wire n_13491;
wire n_13492;
wire n_13493;
wire n_13494;
wire n_13495;
wire n_13496;
wire n_13497;
wire TIMEBOOST_net_1143;
wire n_135;
wire n_1350;
wire n_13500;
wire n_13501;
wire n_13502;
wire TIMEBOOST_net_213;
wire n_13504;
wire n_13505;
wire n_13506;
wire n_13507;
wire n_13508;
wire n_1351;
wire n_13510;
wire n_13511;
wire n_13512;
wire n_13513;
wire n_13514;
wire n_13515;
wire n_13517;
wire n_13518;
wire n_13520;
wire n_13521;
wire n_13522;
wire n_13525;
wire n_13529;
wire n_13530;
wire TIMEBOOST_net_1146;
wire n_13532;
wire n_13533;
wire n_13535;
wire n_13536;
wire TIMEBOOST_net_178;
wire n_13538;
wire n_1354;
wire n_13540;
wire n_13541;
wire n_13542;
wire n_13544;
wire n_13545;
wire n_13546;
wire n_13547;
wire n_13548;
wire n_13549;
wire n_1355;
wire n_13550;
wire n_13552;
wire n_13557;
wire n_13558;
wire n_13559;
wire n_1356;
wire n_13560;
wire n_13562;
wire n_13563;
wire n_13567;
wire n_13568;
wire n_13569;
wire n_1357;
wire n_13570;
wire TIMEBOOST_net_145;
wire n_13573;
wire n_13574;
wire n_13575;
wire n_13576;
wire n_13578;
wire n_13582;
wire n_13583;
wire n_13584;
wire n_13585;
wire n_13586;
wire n_13587;
wire n_13588;
wire n_13589;
wire n_13590;
wire n_13591;
wire TIMEBOOST_net_1525;
wire n_13594;
wire n_13595;
wire n_13597;
wire n_13598;
wire n_13599;
wire n_136;
wire n_1360;
wire n_13601;
wire n_13602;
wire n_13603;
wire n_13606;
wire n_13608;
wire n_13609;
wire n_13610;
wire n_13611;
wire n_13612;
wire n_13613;
wire n_13614;
wire n_13615;
wire n_13616;
wire n_13618;
wire n_13619;
wire n_1362;
wire n_13620;
wire n_13621;
wire TIMEBOOST_net_219;
wire n_13623;
wire n_13624;
wire n_13625;
wire n_13626;
wire n_13628;
wire n_13629;
wire n_1363;
wire n_13630;
wire n_13633;
wire n_13635;
wire n_13636;
wire n_13637;
wire n_13638;
wire n_13639;
wire n_1364;
wire n_13640;
wire n_13642;
wire n_13643;
wire n_13644;
wire n_13645;
wire n_13646;
wire n_13647;
wire n_13649;
wire n_1365;
wire n_13650;
wire n_13651;
wire n_13652;
wire n_13653;
wire n_13657;
wire n_13658;
wire n_13659;
wire n_1366;
wire n_13661;
wire TIMEBOOST_net_1645;
wire n_13664;
wire n_13665;
wire n_13667;
wire n_13668;
wire n_13669;
wire n_1367;
wire n_13670;
wire n_13671;
wire n_13672;
wire n_13673;
wire n_13674;
wire n_13675;
wire n_13676;
wire TIMEBOOST_net_1035;
wire n_13678;
wire n_13679;
wire n_1368;
wire n_13680;
wire n_13681;
wire n_13682;
wire n_13683;
wire n_13684;
wire n_13685;
wire n_13686;
wire n_13689;
wire n_1369;
wire n_13690;
wire TIMEBOOST_net_1539;
wire n_13693;
wire n_13694;
wire n_13695;
wire n_13696;
wire n_13697;
wire n_13698;
wire n_13699;
wire n_137;
wire n_1370;
wire n_13700;
wire n_13701;
wire n_13702;
wire n_13703;
wire n_13704;
wire n_13705;
wire TIMEBOOST_net_2772;
wire n_13707;
wire n_13709;
wire n_1371;
wire n_13711;
wire n_13712;
wire n_13713;
wire n_13714;
wire n_13715;
wire n_13716;
wire n_13717;
wire n_13718;
wire n_13719;
wire n_1372;
wire n_13721;
wire n_13722;
wire n_13724;
wire n_13725;
wire n_13726;
wire TIMEBOOST_net_2851;
wire n_13728;
wire n_13729;
wire n_1373;
wire TIMEBOOST_net_154;
wire n_13731;
wire n_13732;
wire n_13733;
wire n_13734;
wire n_13735;
wire n_13736;
wire n_13737;
wire n_13738;
wire n_13739;
wire n_1374;
wire n_13740;
wire n_13741;
wire n_13742;
wire n_13743;
wire n_13746;
wire n_13747;
wire n_13748;
wire n_13749;
wire n_13750;
wire n_13751;
wire n_13753;
wire n_13754;
wire n_13756;
wire n_13757;
wire n_13759;
wire n_1376;
wire n_13760;
wire n_13761;
wire n_13762;
wire n_13763;
wire n_13764;
wire n_13765;
wire n_13766;
wire n_13767;
wire n_13768;
wire n_13769;
wire n_1377;
wire n_13770;
wire n_13771;
wire n_13774;
wire TIMEBOOST_net_1541;
wire TIMEBOOST_net_909;
wire n_13777;
wire n_13778;
wire n_13779;
wire TIMEBOOST_net_1553;
wire n_13781;
wire TIMEBOOST_net_1034;
wire n_13783;
wire n_13784;
wire n_13785;
wire n_13787;
wire n_13788;
wire n_13789;
wire n_1379;
wire n_13790;
wire n_13791;
wire n_13792;
wire n_13793;
wire n_13794;
wire n_13795;
wire n_13797;
wire n_13798;
wire n_13799;
wire n_138;
wire TIMEBOOST_net_1437;
wire n_13800;
wire n_13801;
wire n_13803;
wire n_13804;
wire n_13805;
wire n_13806;
wire n_13807;
wire TIMEBOOST_net_2844;
wire n_1381;
wire n_13812;
wire n_13813;
wire n_13814;
wire n_13815;
wire n_13816;
wire n_13817;
wire n_13818;
wire TIMEBOOST_net_2322;
wire n_13821;
wire n_13822;
wire n_13823;
wire n_13824;
wire n_13825;
wire n_13826;
wire n_13827;
wire n_13828;
wire n_13829;
wire n_13836;
wire n_13838;
wire n_13839;
wire n_13840;
wire n_13842;
wire n_13846;
wire n_13847;
wire n_13848;
wire n_13849;
wire n_1385;
wire n_13850;
wire n_13851;
wire n_13853;
wire n_13854;
wire n_13855;
wire TIMEBOOST_net_197;
wire n_13857;
wire n_13858;
wire n_13859;
wire n_13860;
wire n_13862;
wire n_13863;
wire n_13864;
wire n_13865;
wire n_13866;
wire n_13869;
wire n_1387;
wire n_13870;
wire n_13875;
wire n_13876;
wire n_13877;
wire n_13878;
wire n_13879;
wire n_13880;
wire n_13882;
wire n_13883;
wire n_13884;
wire n_13886;
wire n_13887;
wire n_13889;
wire n_13890;
wire n_13891;
wire n_13892;
wire n_13893;
wire TIMEBOOST_net_1502;
wire n_13895;
wire n_13897;
wire n_13898;
wire n_13899;
wire n_139;
wire TIMEBOOST_net_1442;
wire n_13900;
wire n_13901;
wire n_13902;
wire n_13903;
wire n_13904;
wire n_13905;
wire n_13906;
wire n_13907;
wire n_13908;
wire n_13909;
wire TIMEBOOST_net_1826;
wire n_13912;
wire n_13913;
wire TIMEBOOST_net_1543;
wire n_13916;
wire n_13918;
wire n_1392;
wire TIMEBOOST_net_195;
wire n_13922;
wire n_13923;
wire n_13924;
wire TIMEBOOST_net_1542;
wire n_13926;
wire n_13927;
wire n_13928;
wire n_13929;
wire n_1393;
wire n_13930;
wire n_13931;
wire n_13934;
wire n_13936;
wire n_13937;
wire n_13938;
wire n_13939;
wire n_13940;
wire n_13941;
wire n_13942;
wire n_13943;
wire n_13944;
wire n_13945;
wire n_13946;
wire n_13947;
wire n_13948;
wire n_13949;
wire n_13950;
wire n_13952;
wire n_13953;
wire n_13954;
wire n_13955;
wire n_13956;
wire n_13957;
wire n_13958;
wire n_13959;
wire n_1396;
wire n_13960;
wire n_13961;
wire n_13966;
wire n_13967;
wire n_1397;
wire n_13970;
wire n_13971;
wire n_13972;
wire n_13973;
wire n_13974;
wire n_13975;
wire n_13976;
wire n_13977;
wire n_1398;
wire n_13980;
wire n_13981;
wire n_13982;
wire n_13984;
wire n_13988;
wire n_13989;
wire n_1399;
wire n_13994;
wire n_13995;
wire n_13996;
wire n_13997;
wire TIMEBOOST_net_919;
wire n_140;
wire n_1400;
wire n_14000;
wire n_14001;
wire n_14002;
wire n_14004;
wire n_14005;
wire n_14006;
wire n_14007;
wire n_14008;
wire n_14009;
wire n_14010;
wire n_14011;
wire n_14012;
wire n_14013;
wire n_14015;
wire n_14016;
wire n_14018;
wire n_14019;
wire n_1402;
wire n_14020;
wire n_14021;
wire n_14022;
wire n_14023;
wire n_14024;
wire n_14025;
wire n_14026;
wire n_14027;
wire n_14028;
wire n_14029;
wire n_1403;
wire n_14030;
wire n_14032;
wire TIMEBOOST_net_2846;
wire n_14034;
wire n_14035;
wire n_14036;
wire n_14037;
wire n_14038;
wire n_14039;
wire TIMEBOOST_net_1825;
wire n_14040;
wire n_14041;
wire n_14042;
wire n_14043;
wire n_14044;
wire n_14049;
wire TIMEBOOST_net_2902;
wire n_14050;
wire n_14051;
wire n_14052;
wire n_14055;
wire n_14056;
wire n_14057;
wire n_14059;
wire n_1406;
wire TIMEBOOST_net_2537;
wire n_14062;
wire n_14063;
wire n_14064;
wire n_14065;
wire n_14066;
wire n_14067;
wire n_14068;
wire n_14069;
wire n_1407;
wire n_14071;
wire n_14072;
wire n_14075;
wire n_14076;
wire n_14077;
wire n_14078;
wire n_14079;
wire n_1408;
wire n_14080;
wire n_14081;
wire TIMEBOOST_net_2729;
wire n_14083;
wire n_14084;
wire n_14085;
wire TIMEBOOST_net_1162;
wire n_14088;
wire n_14089;
wire n_1409;
wire n_14090;
wire n_14091;
wire n_14092;
wire n_14093;
wire TIMEBOOST_net_1879;
wire n_14096;
wire n_14099;
wire n_141;
wire n_14100;
wire n_14101;
wire n_14102;
wire n_14103;
wire n_14104;
wire n_14105;
wire n_14107;
wire n_14108;
wire n_14109;
wire n_14110;
wire n_14111;
wire n_14112;
wire n_14114;
wire n_14115;
wire n_14116;
wire n_14117;
wire n_14118;
wire n_14120;
wire n_14121;
wire n_14122;
wire n_14123;
wire n_14124;
wire n_14125;
wire n_14126;
wire n_14127;
wire n_14128;
wire n_14129;
wire TIMEBOOST_net_204;
wire n_14132;
wire n_14133;
wire n_14135;
wire n_14136;
wire n_14137;
wire n_14138;
wire n_14139;
wire n_14140;
wire n_14141;
wire n_14144;
wire n_14145;
wire n_14146;
wire n_14147;
wire n_14149;
wire n_1415;
wire n_14153;
wire n_14154;
wire n_14155;
wire n_14156;
wire n_14157;
wire TIMEBOOST_net_1112;
wire n_1416;
wire n_14160;
wire n_14161;
wire n_14162;
wire n_14163;
wire TIMEBOOST_net_185;
wire n_14165;
wire n_14168;
wire n_14170;
wire n_14171;
wire n_14172;
wire n_14176;
wire n_14177;
wire n_14178;
wire n_14181;
wire n_14182;
wire TIMEBOOST_net_1899;
wire n_14184;
wire n_14185;
wire n_14186;
wire n_14187;
wire TIMEBOOST_net_2599;
wire n_14190;
wire n_14192;
wire n_14193;
wire n_14194;
wire n_14197;
wire n_14199;
wire n_142;
wire n_1420;
wire n_14200;
wire n_14201;
wire TIMEBOOST_net_1905;
wire n_14203;
wire n_14204;
wire n_14205;
wire n_14206;
wire n_14207;
wire n_14208;
wire n_14209;
wire n_1421;
wire n_14211;
wire n_14212;
wire n_14213;
wire n_14214;
wire n_14215;
wire n_14216;
wire n_14217;
wire n_14218;
wire n_14219;
wire n_1422;
wire n_14220;
wire n_14221;
wire n_14222;
wire n_14225;
wire n_14228;
wire n_14229;
wire n_1423;
wire n_14230;
wire TIMEBOOST_net_2195;
wire n_14233;
wire n_14235;
wire n_14238;
wire n_14239;
wire n_14240;
wire n_14241;
wire TIMEBOOST_net_189;
wire n_14244;
wire n_14245;
wire n_14246;
wire n_14247;
wire n_14248;
wire n_14249;
wire n_14250;
wire n_14251;
wire n_14252;
wire n_14253;
wire n_14254;
wire n_14256;
wire n_14257;
wire n_14258;
wire n_14259;
wire n_1426;
wire n_14260;
wire n_14261;
wire n_14262;
wire n_14265;
wire n_14266;
wire n_14267;
wire n_14268;
wire n_14269;
wire n_1427;
wire n_14270;
wire n_14271;
wire n_14272;
wire n_14273;
wire n_14274;
wire n_14276;
wire n_14277;
wire n_14278;
wire n_14279;
wire n_14281;
wire n_14283;
wire n_14285;
wire n_14286;
wire n_14287;
wire TIMEBOOST_net_1906;
wire n_14291;
wire n_14292;
wire n_14293;
wire n_14294;
wire n_14295;
wire n_14296;
wire n_14297;
wire n_14298;
wire n_14299;
wire n_143;
wire n_14300;
wire n_14301;
wire n_14303;
wire n_14304;
wire n_14306;
wire n_14307;
wire n_14308;
wire n_14309;
wire n_1431;
wire n_14315;
wire n_14317;
wire n_14318;
wire n_14319;
wire n_14321;
wire n_14323;
wire n_14324;
wire n_14326;
wire n_14327;
wire n_14328;
wire n_14329;
wire n_1433;
wire TIMEBOOST_net_319;
wire n_14332;
wire n_14333;
wire n_14334;
wire n_14335;
wire n_14336;
wire n_14338;
wire n_14339;
wire n_1434;
wire n_14340;
wire n_14341;
wire n_14342;
wire n_14343;
wire n_14344;
wire n_14345;
wire n_14346;
wire n_14347;
wire n_14348;
wire n_14349;
wire n_1435;
wire n_14350;
wire n_14351;
wire n_14352;
wire n_14353;
wire n_14354;
wire n_14355;
wire n_14358;
wire n_14359;
wire n_1436;
wire n_14360;
wire TIMEBOOST_net_353;
wire n_14362;
wire n_14363;
wire n_14364;
wire n_14365;
wire n_14366;
wire n_14367;
wire n_14368;
wire n_14369;
wire n_1437;
wire n_14370;
wire n_14372;
wire TIMEBOOST_net_320;
wire TIMEBOOST_net_202;
wire n_14376;
wire n_14377;
wire TIMEBOOST_net_2193;
wire n_14379;
wire n_1438;
wire n_14380;
wire n_14381;
wire n_14382;
wire n_14385;
wire n_14386;
wire n_14387;
wire n_14388;
wire n_14389;
wire n_14390;
wire n_14391;
wire n_14392;
wire n_14393;
wire n_14396;
wire n_14397;
wire n_14398;
wire n_14399;
wire n_144;
wire n_1440;
wire n_14400;
wire n_14402;
wire n_14403;
wire n_14404;
wire n_14407;
wire n_14408;
wire TIMEBOOST_net_2413;
wire n_1441;
wire TIMEBOOST_net_2208;
wire n_14412;
wire n_14413;
wire n_14414;
wire n_14415;
wire n_14416;
wire n_14419;
wire n_1442;
wire n_14420;
wire n_14421;
wire n_14422;
wire n_14423;
wire n_14424;
wire n_14425;
wire n_14426;
wire n_14427;
wire n_14428;
wire n_14429;
wire n_1443;
wire n_14430;
wire n_14431;
wire n_14432;
wire n_14433;
wire n_14434;
wire n_14435;
wire n_14436;
wire n_14437;
wire TIMEBOOST_net_1551;
wire n_14439;
wire n_1444;
wire n_14441;
wire TIMEBOOST_net_2401;
wire n_14444;
wire n_14447;
wire n_14448;
wire n_1445;
wire n_14450;
wire n_14451;
wire n_14452;
wire n_14454;
wire n_14455;
wire n_14456;
wire n_14457;
wire n_1446;
wire n_14460;
wire n_14461;
wire n_14462;
wire n_14466;
wire n_14467;
wire n_14468;
wire n_14469;
wire n_1447;
wire n_14471;
wire n_14472;
wire n_14473;
wire n_14474;
wire n_14475;
wire n_14476;
wire n_14477;
wire n_14478;
wire n_14479;
wire n_1448;
wire TIMEBOOST_net_325;
wire n_14483;
wire n_14485;
wire n_14486;
wire n_14487;
wire n_14488;
wire n_14489;
wire n_14490;
wire n_14491;
wire n_14492;
wire n_14493;
wire n_14494;
wire n_14495;
wire n_14496;
wire n_14498;
wire n_145;
wire n_1450;
wire n_14503;
wire n_14504;
wire n_14505;
wire n_14506;
wire n_14507;
wire n_14508;
wire n_1451;
wire n_14510;
wire n_14511;
wire TIMEBOOST_net_2307;
wire n_14515;
wire n_14516;
wire TIMEBOOST_net_324;
wire n_14519;
wire n_1452;
wire n_14524;
wire n_14525;
wire n_14526;
wire n_14527;
wire n_14528;
wire n_14529;
wire n_1453;
wire n_14530;
wire n_14531;
wire n_14532;
wire n_14533;
wire n_14534;
wire n_14535;
wire n_14536;
wire n_14539;
wire n_1454;
wire n_14540;
wire n_14543;
wire n_14544;
wire n_14545;
wire n_14546;
wire n_14547;
wire n_14549;
wire n_1455;
wire n_14550;
wire n_14551;
wire n_14552;
wire n_14554;
wire n_14555;
wire n_14556;
wire n_14557;
wire n_1456;
wire n_14560;
wire n_14561;
wire n_14562;
wire n_14563;
wire n_14564;
wire n_14565;
wire n_14566;
wire n_14567;
wire n_14568;
wire n_14569;
wire n_14571;
wire n_14572;
wire n_14573;
wire n_14575;
wire n_14576;
wire n_14579;
wire n_14580;
wire TIMEBOOST_net_2829;
wire n_14582;
wire n_14583;
wire n_14584;
wire n_14585;
wire n_14586;
wire n_14587;
wire n_14588;
wire n_14590;
wire n_14591;
wire n_14592;
wire n_14593;
wire n_14598;
wire n_146;
wire n_1460;
wire n_14600;
wire n_14601;
wire n_14602;
wire TIMEBOOST_net_1122;
wire n_14605;
wire TIMEBOOST_net_1922;
wire n_14607;
wire n_14608;
wire TIMEBOOST_net_1651;
wire n_1461;
wire n_14611;
wire n_14612;
wire n_14613;
wire n_14614;
wire n_14615;
wire n_14616;
wire TIMEBOOST_net_2909;
wire n_14618;
wire n_14619;
wire n_1462;
wire n_14620;
wire n_14621;
wire n_14622;
wire n_14625;
wire n_14626;
wire n_14628;
wire TIMEBOOST_net_332;
wire n_1463;
wire TIMEBOOST_net_331;
wire n_14632;
wire n_14633;
wire n_14634;
wire n_14635;
wire n_14636;
wire n_14638;
wire n_14641;
wire n_14642;
wire n_14643;
wire n_14645;
wire n_14646;
wire n_14647;
wire TIMEBOOST_net_2093;
wire TIMEBOOST_net_2760;
wire n_14650;
wire n_14652;
wire n_14653;
wire TIMEBOOST_net_1670;
wire n_14656;
wire n_14657;
wire n_14658;
wire n_14659;
wire n_14660;
wire n_14661;
wire n_14662;
wire TIMEBOOST_net_1652;
wire n_14664;
wire n_14665;
wire n_14666;
wire n_14667;
wire TIMEBOOST_net_2910;
wire n_14669;
wire n_1467;
wire n_14670;
wire n_14672;
wire n_14673;
wire n_14676;
wire n_14677;
wire n_14678;
wire n_14679;
wire n_14681;
wire n_14682;
wire n_14684;
wire n_14685;
wire n_14686;
wire n_14687;
wire n_14689;
wire n_14693;
wire n_14694;
wire TIMEBOOST_net_1942;
wire n_14696;
wire n_14697;
wire n_14698;
wire n_14699;
wire n_147;
wire n_1470;
wire n_14700;
wire n_14701;
wire n_14702;
wire n_14703;
wire n_14704;
wire n_14706;
wire n_14707;
wire n_14709;
wire n_1471;
wire n_14710;
wire n_14711;
wire n_14714;
wire n_14715;
wire n_14716;
wire n_14717;
wire n_14718;
wire n_14719;
wire n_1472;
wire n_14720;
wire n_14721;
wire n_14722;
wire TIMEBOOST_net_2831;
wire n_14727;
wire n_14730;
wire n_14731;
wire n_14732;
wire n_14733;
wire n_14734;
wire n_14735;
wire n_14736;
wire n_14737;
wire n_14738;
wire n_1474;
wire n_14740;
wire n_14741;
wire n_14742;
wire n_14743;
wire n_14744;
wire n_14745;
wire n_14746;
wire n_14747;
wire n_1475;
wire n_14750;
wire n_14751;
wire TIMEBOOST_net_2199;
wire TIMEBOOST_net_2745;
wire n_14754;
wire n_14755;
wire n_14756;
wire n_14757;
wire n_14759;
wire n_1476;
wire n_14760;
wire n_14761;
wire n_14763;
wire n_14764;
wire n_14768;
wire n_1477;
wire n_14770;
wire n_14771;
wire n_14772;
wire n_14773;
wire n_14774;
wire n_14775;
wire n_14779;
wire n_1478;
wire n_14780;
wire n_14781;
wire n_14782;
wire n_14785;
wire n_14786;
wire n_14788;
wire n_14789;
wire n_1479;
wire n_14790;
wire n_14791;
wire n_14792;
wire n_14793;
wire n_14794;
wire n_14795;
wire n_14796;
wire n_14798;
wire n_14799;
wire n_148;
wire n_1480;
wire TIMEBOOST_net_337;
wire n_14801;
wire n_14802;
wire n_14803;
wire TIMEBOOST_net_301;
wire n_14805;
wire n_14808;
wire n_14809;
wire n_14810;
wire n_14811;
wire n_14812;
wire n_14814;
wire n_14815;
wire n_14816;
wire TIMEBOOST_net_2650;
wire n_14818;
wire n_14819;
wire n_1482;
wire n_14821;
wire n_14823;
wire n_14824;
wire n_14826;
wire n_14827;
wire n_14829;
wire n_1483;
wire n_14830;
wire n_14835;
wire n_14836;
wire n_14837;
wire n_14838;
wire n_14839;
wire n_1484;
wire n_14840;
wire n_14841;
wire n_14842;
wire n_14843;
wire n_14845;
wire n_14846;
wire TIMEBOOST_net_1185;
wire n_1485;
wire n_14851;
wire n_14852;
wire n_14853;
wire n_14854;
wire n_14855;
wire n_14856;
wire n_14857;
wire n_14858;
wire n_14859;
wire n_1486;
wire n_14860;
wire n_14861;
wire n_14862;
wire n_14864;
wire n_14865;
wire n_14868;
wire n_14869;
wire n_1487;
wire n_14870;
wire n_14871;
wire n_14872;
wire n_14873;
wire n_14874;
wire n_14875;
wire n_14877;
wire n_14878;
wire TIMEBOOST_net_1970;
wire n_1488;
wire n_14880;
wire n_14881;
wire TIMEBOOST_net_2863;
wire n_14884;
wire n_14885;
wire n_14886;
wire n_14887;
wire TIMEBOOST_net_1943;
wire n_14889;
wire n_1489;
wire n_14890;
wire n_14891;
wire n_14894;
wire n_14895;
wire n_14896;
wire n_14897;
wire n_14898;
wire n_14899;
wire n_149;
wire n_1490;
wire n_14901;
wire n_14902;
wire n_14903;
wire n_14905;
wire n_14906;
wire n_14907;
wire n_14908;
wire n_14909;
wire n_1491;
wire n_14911;
wire n_14912;
wire n_14913;
wire n_14915;
wire n_14916;
wire n_14917;
wire n_14918;
wire n_14919;
wire n_14920;
wire n_14921;
wire n_14923;
wire n_14924;
wire n_14927;
wire n_14928;
wire n_1493;
wire n_14932;
wire n_14935;
wire n_1494;
wire TIMEBOOST_net_2262;
wire n_14942;
wire n_14943;
wire n_14944;
wire n_14947;
wire n_14948;
wire TIMEBOOST_net_304;
wire n_1495;
wire n_14950;
wire n_14953;
wire n_14954;
wire n_14955;
wire n_14956;
wire TIMEBOOST_net_2899;
wire n_14958;
wire n_14959;
wire n_1496;
wire n_14960;
wire n_14962;
wire TIMEBOOST_net_2727;
wire n_14964;
wire n_14966;
wire n_14967;
wire n_14968;
wire n_14969;
wire n_1497;
wire n_14970;
wire n_14971;
wire n_14972;
wire n_14973;
wire TIMEBOOST_net_2471;
wire n_14975;
wire n_14976;
wire n_14977;
wire n_14978;
wire n_14979;
wire n_1498;
wire n_14982;
wire n_14983;
wire n_14985;
wire n_14986;
wire n_14987;
wire n_14988;
wire n_14989;
wire n_1499;
wire n_14991;
wire n_14992;
wire n_14993;
wire n_14994;
wire n_14995;
wire n_14996;
wire n_14997;
wire n_14998;
wire n_14999;
wire n_150;
wire n_1500;
wire n_15000;
wire n_15001;
wire n_15003;
wire n_15004;
wire n_15005;
wire n_15006;
wire n_15008;
wire n_15009;
wire n_1501;
wire n_15010;
wire n_15012;
wire n_15014;
wire TIMEBOOST_net_1634;
wire n_15017;
wire n_15018;
wire n_15019;
wire n_1502;
wire n_15021;
wire n_15022;
wire n_15023;
wire n_15025;
wire n_15026;
wire n_15029;
wire n_1503;
wire n_15030;
wire n_15031;
wire n_15032;
wire n_15033;
wire n_15035;
wire n_15036;
wire n_15037;
wire n_15038;
wire n_15039;
wire n_1504;
wire n_15040;
wire n_15041;
wire n_15042;
wire n_15043;
wire n_15044;
wire n_15045;
wire n_15047;
wire n_15048;
wire n_15049;
wire n_1505;
wire n_15050;
wire TIMEBOOST_net_1659;
wire n_15053;
wire n_15054;
wire n_15055;
wire n_15058;
wire n_15059;
wire n_1506;
wire n_15060;
wire n_15063;
wire n_15064;
wire n_15065;
wire n_15066;
wire n_15067;
wire n_1507;
wire n_15070;
wire n_15071;
wire n_15075;
wire n_15076;
wire n_15077;
wire n_15079;
wire n_1508;
wire n_15081;
wire n_15082;
wire n_15083;
wire n_15084;
wire n_15085;
wire n_15086;
wire n_15087;
wire n_15088;
wire n_15089;
wire n_1509;
wire n_15090;
wire n_15091;
wire n_15092;
wire n_15093;
wire n_15094;
wire n_15097;
wire n_15098;
wire n_15099;
wire n_151;
wire n_1510;
wire n_15103;
wire n_15108;
wire n_15109;
wire n_15110;
wire n_15112;
wire n_15113;
wire n_15114;
wire n_15118;
wire n_1512;
wire n_15123;
wire n_15124;
wire TIMEBOOST_net_2298;
wire TIMEBOOST_net_1733;
wire n_15127;
wire n_15128;
wire n_1513;
wire n_15132;
wire n_15133;
wire n_15136;
wire n_15137;
wire n_15139;
wire n_1514;
wire n_15140;
wire n_15141;
wire n_15142;
wire n_15143;
wire n_15144;
wire n_15149;
wire n_1515;
wire n_15151;
wire n_15153;
wire n_15154;
wire n_15156;
wire n_15157;
wire n_15159;
wire n_1516;
wire n_15160;
wire TIMEBOOST_net_1643;
wire n_15163;
wire n_15164;
wire n_15168;
wire n_1517;
wire n_15170;
wire n_15171;
wire n_15175;
wire n_15177;
wire n_15178;
wire n_1518;
wire n_15180;
wire n_15181;
wire n_15182;
wire TIMEBOOST_net_1690;
wire n_15187;
wire n_15189;
wire n_1519;
wire TIMEBOOST_net_2024;
wire n_15194;
wire n_15195;
wire n_15196;
wire n_15198;
wire n_152;
wire n_1520;
wire n_15200;
wire n_15204;
wire n_15205;
wire n_15206;
wire n_15207;
wire n_15208;
wire n_15209;
wire n_1521;
wire n_15210;
wire n_15211;
wire n_15212;
wire TIMEBOOST_net_308;
wire TIMEBOOST_net_1188;
wire n_15218;
wire n_15219;
wire n_15221;
wire n_15223;
wire n_15224;
wire n_15225;
wire n_15226;
wire n_15227;
wire n_15228;
wire n_15230;
wire n_15231;
wire n_15233;
wire n_15234;
wire n_15235;
wire n_15237;
wire n_15238;
wire n_15239;
wire n_1524;
wire n_15240;
wire n_15241;
wire n_15242;
wire n_15243;
wire n_15244;
wire n_15245;
wire n_15246;
wire n_15247;
wire n_15248;
wire n_1525;
wire n_15250;
wire n_15252;
wire n_15256;
wire n_15257;
wire n_15258;
wire n_15259;
wire n_15263;
wire n_15264;
wire n_15265;
wire n_15266;
wire n_15267;
wire n_15269;
wire n_1527;
wire n_15270;
wire n_15271;
wire n_15272;
wire n_15273;
wire n_15274;
wire n_15275;
wire n_15276;
wire n_15277;
wire n_15278;
wire n_1528;
wire n_15281;
wire n_15282;
wire TIMEBOOST_net_1980;
wire n_15284;
wire TIMEBOOST_net_2864;
wire n_15286;
wire n_15287;
wire n_15288;
wire n_15289;
wire n_1529;
wire n_15290;
wire n_15293;
wire n_15294;
wire n_15295;
wire n_15296;
wire n_15297;
wire n_15298;
wire n_15299;
wire n_153;
wire n_1530;
wire n_15300;
wire n_15302;
wire n_15303;
wire n_15305;
wire n_15306;
wire n_15308;
wire n_15309;
wire n_15310;
wire n_15311;
wire n_15313;
wire n_15314;
wire n_15319;
wire n_15320;
wire n_15321;
wire n_15323;
wire n_15324;
wire n_15325;
wire TIMEBOOST_net_1187;
wire n_1533;
wire n_15330;
wire n_15331;
wire n_15332;
wire n_15333;
wire n_15335;
wire n_15336;
wire n_15337;
wire n_15338;
wire n_15339;
wire n_1534;
wire n_15340;
wire n_15341;
wire n_15342;
wire n_15343;
wire n_15344;
wire n_15345;
wire n_15349;
wire n_1535;
wire n_15352;
wire n_15353;
wire n_15356;
wire n_15357;
wire TIMEBOOST_net_2257;
wire n_15360;
wire n_15361;
wire n_15362;
wire n_15363;
wire n_15366;
wire n_15369;
wire n_1537;
wire n_15370;
wire n_15371;
wire n_15372;
wire n_15373;
wire n_15374;
wire n_15375;
wire n_15376;
wire n_15377;
wire n_15378;
wire n_15379;
wire n_1538;
wire n_15380;
wire n_15381;
wire n_15382;
wire n_15383;
wire n_15384;
wire n_15385;
wire n_15387;
wire TIMEBOOST_net_2688;
wire n_15389;
wire n_1539;
wire n_15390;
wire n_15391;
wire n_15392;
wire n_15394;
wire n_15395;
wire n_15396;
wire n_15397;
wire n_15398;
wire n_15399;
wire n_154;
wire n_1540;
wire n_15402;
wire n_15403;
wire n_15404;
wire n_15405;
wire n_15406;
wire n_15407;
wire n_15408;
wire n_15409;
wire n_1541;
wire n_15410;
wire n_15412;
wire n_15413;
wire n_15414;
wire n_15415;
wire n_15416;
wire n_15417;
wire n_1542;
wire n_15420;
wire n_15421;
wire n_15422;
wire n_15423;
wire n_15425;
wire n_15426;
wire n_15427;
wire n_15429;
wire n_1543;
wire TIMEBOOST_net_398;
wire n_15433;
wire n_15434;
wire n_15437;
wire n_15438;
wire TIMEBOOST_net_2861;
wire n_1544;
wire n_15440;
wire n_15441;
wire n_15442;
wire n_15443;
wire n_15446;
wire TIMEBOOST_net_2258;
wire n_15448;
wire n_15449;
wire n_1545;
wire n_15450;
wire n_15452;
wire n_15453;
wire n_15454;
wire n_15455;
wire n_15457;
wire n_15458;
wire n_15459;
wire n_1546;
wire n_15460;
wire n_15461;
wire n_15462;
wire n_15463;
wire n_15464;
wire n_15465;
wire TIMEBOOST_net_2271;
wire n_15468;
wire n_15469;
wire n_1547;
wire n_15473;
wire TIMEBOOST_net_1153;
wire n_15475;
wire n_15476;
wire TIMEBOOST_net_2852;
wire n_15479;
wire n_1548;
wire n_15481;
wire n_15482;
wire TIMEBOOST_net_2882;
wire n_15486;
wire n_15487;
wire n_15488;
wire n_15489;
wire n_1549;
wire n_15490;
wire n_15491;
wire n_15492;
wire n_15493;
wire n_15494;
wire n_15495;
wire n_15496;
wire n_15497;
wire n_15498;
wire TIMEBOOST_net_1724;
wire n_155;
wire n_1550;
wire n_15500;
wire n_15501;
wire n_15502;
wire n_15503;
wire n_15504;
wire n_1551;
wire n_15510;
wire n_15512;
wire n_15513;
wire n_15514;
wire n_15515;
wire n_15516;
wire n_15517;
wire n_15518;
wire TIMEBOOST_net_2234;
wire n_15520;
wire n_15521;
wire n_15522;
wire n_15523;
wire n_15524;
wire TIMEBOOST_net_311;
wire n_15526;
wire n_15527;
wire n_15528;
wire n_15529;
wire n_1553;
wire n_15530;
wire n_15531;
wire n_15532;
wire n_15533;
wire n_15534;
wire n_15535;
wire n_15536;
wire n_15537;
wire n_15538;
wire n_1554;
wire n_15541;
wire TIMEBOOST_net_1293;
wire n_15543;
wire n_15545;
wire n_15546;
wire n_15547;
wire n_15548;
wire n_15549;
wire n_1555;
wire n_15551;
wire n_15552;
wire n_15553;
wire TIMEBOOST_net_1633;
wire n_15557;
wire n_15559;
wire n_1556;
wire n_15561;
wire n_15563;
wire n_15564;
wire n_15565;
wire n_15566;
wire n_15567;
wire n_15568;
wire n_15569;
wire n_1557;
wire n_15571;
wire n_15572;
wire n_15573;
wire n_15574;
wire n_15575;
wire n_15576;
wire n_15577;
wire n_15578;
wire TIMEBOOST_net_1119;
wire n_1558;
wire n_15580;
wire n_15581;
wire n_15584;
wire n_15586;
wire n_1559;
wire n_15591;
wire n_15592;
wire n_15595;
wire TIMEBOOST_net_374;
wire n_15598;
wire n_156;
wire n_1560;
wire n_15601;
wire n_15602;
wire n_15603;
wire n_15604;
wire n_15605;
wire n_15606;
wire n_15607;
wire n_15608;
wire n_15609;
wire n_1561;
wire n_15610;
wire n_15611;
wire n_15612;
wire n_15613;
wire n_15614;
wire n_15615;
wire n_15619;
wire n_15620;
wire n_15621;
wire n_15622;
wire n_15623;
wire n_15625;
wire n_15627;
wire n_15628;
wire n_15629;
wire n_1563;
wire n_15631;
wire n_15632;
wire n_15633;
wire n_15634;
wire n_15635;
wire n_15636;
wire n_15637;
wire n_15638;
wire n_15639;
wire n_1564;
wire n_15640;
wire n_15641;
wire n_15642;
wire n_15643;
wire n_15644;
wire n_15648;
wire n_15649;
wire n_1565;
wire n_15651;
wire n_15652;
wire TIMEBOOST_net_465;
wire n_15655;
wire n_15656;
wire n_15657;
wire TIMEBOOST_net_1155;
wire n_15660;
wire n_15661;
wire n_15663;
wire n_15664;
wire n_15665;
wire n_15666;
wire n_15667;
wire n_15668;
wire n_15669;
wire n_1567;
wire n_15671;
wire n_15672;
wire n_15673;
wire n_15674;
wire n_15675;
wire n_15676;
wire n_15677;
wire n_15678;
wire n_15679;
wire n_1568;
wire n_15680;
wire n_15683;
wire n_15684;
wire n_15685;
wire n_15686;
wire n_15687;
wire n_15688;
wire n_1569;
wire n_15692;
wire n_15694;
wire TIMEBOOST_net_1229;
wire n_15696;
wire n_15698;
wire n_157;
wire n_1570;
wire n_15700;
wire n_15701;
wire n_15702;
wire n_15704;
wire n_15706;
wire n_15708;
wire n_15709;
wire n_1571;
wire n_15710;
wire n_15711;
wire n_15712;
wire n_15714;
wire n_15715;
wire n_15716;
wire n_15717;
wire n_15718;
wire n_15719;
wire n_1572;
wire TIMEBOOST_net_2239;
wire n_15721;
wire n_15722;
wire n_15723;
wire n_15724;
wire n_15725;
wire n_15726;
wire n_15727;
wire n_15728;
wire n_15730;
wire n_15731;
wire n_15732;
wire n_15734;
wire TIMEBOOST_net_507;
wire n_15736;
wire n_15737;
wire n_15738;
wire n_15739;
wire n_15741;
wire TIMEBOOST_net_445;
wire n_15743;
wire n_15744;
wire n_15745;
wire n_15747;
wire n_15748;
wire n_15749;
wire n_1575;
wire n_15750;
wire n_15751;
wire n_15752;
wire n_15753;
wire n_15754;
wire n_15755;
wire n_15756;
wire n_15757;
wire n_15758;
wire n_15761;
wire n_15762;
wire TIMEBOOST_net_2928;
wire n_15765;
wire n_15767;
wire n_15768;
wire n_1577;
wire n_15770;
wire n_15771;
wire TIMEBOOST_net_446;
wire TIMEBOOST_net_2884;
wire TIMEBOOST_net_1998;
wire n_15778;
wire n_15779;
wire n_15781;
wire n_15783;
wire n_15784;
wire n_15785;
wire n_15786;
wire n_15787;
wire n_15788;
wire n_15789;
wire n_15790;
wire n_15791;
wire n_15792;
wire n_15793;
wire n_15795;
wire n_15797;
wire n_15799;
wire n_158;
wire n_1580;
wire n_15800;
wire n_15801;
wire n_15802;
wire n_15803;
wire n_15804;
wire n_15805;
wire n_15806;
wire TIMEBOOST_net_518;
wire n_15808;
wire n_15809;
wire n_15810;
wire TIMEBOOST_net_448;
wire TIMEBOOST_net_2310;
wire n_15815;
wire n_15817;
wire n_15818;
wire n_15819;
wire n_15820;
wire n_15821;
wire n_15822;
wire n_15823;
wire n_15826;
wire n_15827;
wire n_15828;
wire n_15829;
wire n_15830;
wire n_15832;
wire n_15833;
wire n_15834;
wire n_15835;
wire n_15836;
wire n_15837;
wire n_15838;
wire n_15839;
wire n_1584;
wire n_15840;
wire n_15841;
wire n_15842;
wire n_15843;
wire n_15844;
wire n_15845;
wire n_15847;
wire n_15849;
wire n_1585;
wire n_15850;
wire n_15852;
wire n_15853;
wire n_15854;
wire TIMEBOOST_net_521;
wire n_15856;
wire n_15857;
wire n_15858;
wire n_1586;
wire n_15860;
wire n_15861;
wire n_15862;
wire n_15865;
wire n_15866;
wire n_15867;
wire n_15868;
wire n_15869;
wire n_1587;
wire n_15870;
wire n_15871;
wire n_15872;
wire n_15873;
wire n_15875;
wire n_15876;
wire n_15877;
wire n_15878;
wire n_15879;
wire n_1588;
wire n_15880;
wire n_15881;
wire n_15882;
wire n_15883;
wire n_15884;
wire n_15886;
wire n_15887;
wire n_15888;
wire n_15889;
wire n_15890;
wire n_15891;
wire n_15892;
wire n_15893;
wire n_15895;
wire n_15896;
wire TIMEBOOST_net_1768;
wire n_15898;
wire n_159;
wire n_1590;
wire n_15900;
wire n_15901;
wire n_15905;
wire n_15906;
wire n_15907;
wire n_15908;
wire n_15909;
wire n_1591;
wire n_15911;
wire n_15912;
wire n_15915;
wire n_15917;
wire n_15918;
wire n_15919;
wire TIMEBOOST_net_2939;
wire n_15920;
wire n_15921;
wire n_15922;
wire n_15923;
wire n_15924;
wire n_15925;
wire n_15926;
wire n_15927;
wire n_15928;
wire n_15929;
wire n_1593;
wire n_15930;
wire n_15931;
wire n_15932;
wire n_15933;
wire n_15934;
wire n_15935;
wire n_15937;
wire n_15938;
wire n_15939;
wire n_1594;
wire n_15942;
wire n_15943;
wire n_15944;
wire n_15945;
wire n_15946;
wire n_15948;
wire n_15949;
wire n_1595;
wire TIMEBOOST_net_2922;
wire n_15951;
wire TIMEBOOST_net_571;
wire n_15953;
wire n_15954;
wire n_15957;
wire n_15958;
wire n_15959;
wire n_1596;
wire n_15960;
wire n_15961;
wire n_15962;
wire n_15963;
wire n_15964;
wire n_15965;
wire n_15967;
wire n_15968;
wire n_15969;
wire n_1597;
wire n_15970;
wire n_15971;
wire n_15972;
wire n_15973;
wire n_15974;
wire n_15975;
wire n_15976;
wire n_15977;
wire n_15978;
wire n_15979;
wire n_15980;
wire n_15981;
wire n_15983;
wire n_15984;
wire n_15985;
wire TIMEBOOST_net_1301;
wire n_15987;
wire n_15988;
wire n_15989;
wire n_1599;
wire n_15990;
wire n_15992;
wire n_15993;
wire n_15995;
wire TIMEBOOST_net_1311;
wire n_15998;
wire n_15999;
wire n_160;
wire n_1600;
wire n_16000;
wire n_16001;
wire n_16003;
wire n_16004;
wire TIMEBOOST_net_1755;
wire n_16007;
wire n_16008;
wire TIMEBOOST_net_1698;
wire n_1601;
wire n_16010;
wire n_16011;
wire n_16016;
wire n_16017;
wire n_16018;
wire n_16019;
wire n_1602;
wire n_16020;
wire n_16021;
wire n_16022;
wire n_16023;
wire n_16024;
wire n_16025;
wire n_16026;
wire n_16027;
wire n_16028;
wire n_16029;
wire n_1603;
wire n_16030;
wire n_16031;
wire n_16032;
wire TIMEBOOST_net_575;
wire n_16036;
wire n_16037;
wire n_16038;
wire n_1604;
wire n_16041;
wire n_16044;
wire n_16046;
wire n_16047;
wire n_16048;
wire n_16049;
wire n_16052;
wire n_16053;
wire n_16056;
wire TIMEBOOST_net_451;
wire n_16059;
wire n_16060;
wire n_16061;
wire n_16062;
wire n_16063;
wire n_16064;
wire n_16065;
wire n_16066;
wire n_16067;
wire n_16070;
wire n_16071;
wire n_16072;
wire n_16074;
wire n_16075;
wire TIMEBOOST_net_559;
wire n_16077;
wire TIMEBOOST_net_1725;
wire n_1608;
wire n_16080;
wire n_16084;
wire n_16086;
wire n_16088;
wire n_16089;
wire n_1609;
wire n_16090;
wire TIMEBOOST_net_2233;
wire n_16094;
wire n_16095;
wire n_16098;
wire n_16099;
wire n_161;
wire n_1610;
wire n_16100;
wire n_16101;
wire n_16102;
wire n_16103;
wire n_16104;
wire n_16105;
wire n_16106;
wire n_16107;
wire n_16108;
wire n_16109;
wire n_16110;
wire n_16111;
wire n_16112;
wire n_16113;
wire n_16118;
wire n_16119;
wire n_16122;
wire n_16123;
wire n_16124;
wire n_16125;
wire TIMEBOOST_net_2642;
wire TIMEBOOST_net_2305;
wire n_1613;
wire n_16131;
wire n_16132;
wire n_16133;
wire n_16134;
wire n_16135;
wire n_16136;
wire n_16137;
wire n_16138;
wire n_16139;
wire n_1614;
wire n_16140;
wire n_16141;
wire n_16142;
wire n_16143;
wire n_16144;
wire n_16146;
wire n_16151;
wire n_16154;
wire n_16155;
wire n_16157;
wire n_16158;
wire n_16159;
wire n_1616;
wire n_16160;
wire n_16161;
wire TIMEBOOST_net_1305;
wire TIMEBOOST_net_1744;
wire n_16166;
wire n_16168;
wire n_16169;
wire n_1617;
wire n_16170;
wire n_16171;
wire n_16172;
wire n_16173;
wire n_16174;
wire n_16175;
wire n_16176;
wire n_16177;
wire n_16178;
wire n_16179;
wire n_16180;
wire n_16181;
wire n_16182;
wire n_16183;
wire n_16188;
wire n_16189;
wire n_1619;
wire n_16190;
wire n_16192;
wire n_16193;
wire n_16194;
wire TIMEBOOST_net_529;
wire n_16197;
wire n_162;
wire n_1620;
wire n_16200;
wire n_16201;
wire n_16202;
wire n_16203;
wire n_16204;
wire n_16205;
wire n_16206;
wire n_16207;
wire n_16210;
wire n_16211;
wire n_16212;
wire n_16216;
wire n_16218;
wire n_16219;
wire n_1622;
wire n_16220;
wire n_16221;
wire n_16223;
wire n_16224;
wire n_16225;
wire n_16226;
wire n_16228;
wire n_1623;
wire n_16230;
wire n_16231;
wire n_16232;
wire n_16233;
wire n_16234;
wire TIMEBOOST_net_562;
wire n_16236;
wire n_16237;
wire n_1624;
wire n_16241;
wire n_16244;
wire n_16245;
wire n_16246;
wire n_16249;
wire n_1625;
wire n_16250;
wire n_16253;
wire n_16254;
wire n_16255;
wire n_16256;
wire n_16257;
wire n_16258;
wire n_16259;
wire n_1626;
wire n_16260;
wire n_16261;
wire n_16262;
wire n_16263;
wire n_16264;
wire n_16265;
wire n_16266;
wire n_16267;
wire n_16268;
wire n_16269;
wire n_1627;
wire n_16270;
wire n_16271;
wire n_16272;
wire n_16273;
wire n_16274;
wire n_16277;
wire n_16278;
wire n_16279;
wire n_1628;
wire n_16283;
wire n_16285;
wire n_16286;
wire n_16287;
wire n_16288;
wire n_16289;
wire n_1629;
wire n_16290;
wire n_16291;
wire n_16293;
wire n_16295;
wire n_16296;
wire TIMEBOOST_net_563;
wire n_163;
wire n_1630;
wire n_16300;
wire n_16301;
wire n_16302;
wire n_16303;
wire n_16304;
wire n_16305;
wire n_16306;
wire n_16307;
wire n_16308;
wire n_16309;
wire n_16310;
wire n_16311;
wire n_16312;
wire n_16313;
wire n_16314;
wire n_16316;
wire n_16317;
wire n_16318;
wire n_16319;
wire n_1632;
wire n_16321;
wire n_16322;
wire n_16324;
wire n_16325;
wire n_16328;
wire TIMEBOOST_net_2912;
wire n_1633;
wire n_16330;
wire n_16332;
wire n_16333;
wire TIMEBOOST_net_1303;
wire n_16336;
wire n_16337;
wire n_16339;
wire TIMEBOOST_net_1840;
wire n_16341;
wire n_16342;
wire n_16343;
wire n_16344;
wire n_16345;
wire n_16346;
wire n_16347;
wire n_16348;
wire n_16349;
wire n_1635;
wire n_16350;
wire n_16351;
wire n_16352;
wire n_16353;
wire n_16354;
wire n_16355;
wire n_16356;
wire n_16357;
wire n_16358;
wire n_16359;
wire n_1636;
wire n_16360;
wire n_16361;
wire n_16362;
wire n_16363;
wire n_16364;
wire n_16365;
wire n_16366;
wire n_16367;
wire n_16368;
wire n_16369;
wire n_16370;
wire n_16371;
wire n_16372;
wire n_16373;
wire n_16374;
wire n_16375;
wire n_16376;
wire n_16377;
wire TIMEBOOST_net_2871;
wire n_16379;
wire n_1638;
wire n_16384;
wire n_16385;
wire n_16386;
wire n_16388;
wire n_16389;
wire n_1639;
wire n_16390;
wire n_16391;
wire n_16392;
wire n_16394;
wire n_16396;
wire n_16397;
wire n_16398;
wire n_16399;
wire n_164;
wire n_16401;
wire n_16402;
wire n_16404;
wire n_16405;
wire n_16406;
wire n_16407;
wire n_16408;
wire n_16409;
wire n_16410;
wire n_16411;
wire n_16412;
wire n_16413;
wire n_16414;
wire n_16415;
wire n_16416;
wire n_16417;
wire n_16418;
wire n_16419;
wire n_16422;
wire n_16423;
wire n_16424;
wire n_16425;
wire n_16426;
wire n_16429;
wire n_1643;
wire n_16431;
wire n_16432;
wire n_16433;
wire n_16434;
wire n_16435;
wire n_16436;
wire n_16437;
wire n_16438;
wire n_16439;
wire n_1644;
wire n_16440;
wire n_16441;
wire n_16442;
wire n_16443;
wire n_16444;
wire n_16445;
wire n_16446;
wire n_16447;
wire n_16448;
wire n_16449;
wire n_1645;
wire n_16450;
wire TIMEBOOST_net_1588;
wire n_16452;
wire n_16453;
wire n_16454;
wire n_16455;
wire n_16456;
wire n_16458;
wire n_1646;
wire n_16460;
wire n_16461;
wire n_16462;
wire n_16463;
wire n_16464;
wire n_16465;
wire n_16466;
wire n_16468;
wire n_16469;
wire n_16471;
wire n_16472;
wire n_16474;
wire n_16475;
wire n_16479;
wire n_1648;
wire n_16480;
wire n_16481;
wire n_16482;
wire n_16484;
wire n_16485;
wire n_16486;
wire TIMEBOOST_net_2094;
wire n_16489;
wire n_1649;
wire n_16490;
wire n_16491;
wire n_16493;
wire n_16494;
wire n_16495;
wire TIMEBOOST_net_566;
wire n_16497;
wire TIMEBOOST_net_570;
wire n_16499;
wire n_165;
wire n_1650;
wire n_16500;
wire n_16503;
wire n_16504;
wire n_16505;
wire n_16506;
wire n_16507;
wire n_16508;
wire n_16509;
wire n_16510;
wire TIMEBOOST_net_2162;
wire TIMEBOOST_net_646;
wire n_16513;
wire n_16514;
wire n_16515;
wire n_16516;
wire TIMEBOOST_net_1309;
wire n_16518;
wire n_1652;
wire n_16523;
wire n_16524;
wire n_16526;
wire n_16527;
wire n_16529;
wire n_1653;
wire n_16530;
wire n_16531;
wire n_16532;
wire n_16533;
wire n_16534;
wire n_16535;
wire n_16536;
wire n_16537;
wire n_1654;
wire TIMEBOOST_net_2190;
wire n_16541;
wire n_16542;
wire n_16543;
wire n_16544;
wire n_16545;
wire n_16546;
wire n_16547;
wire n_16548;
wire n_16549;
wire n_16550;
wire n_16551;
wire n_16552;
wire n_16553;
wire n_16555;
wire n_16556;
wire n_16557;
wire n_16558;
wire n_16559;
wire n_1656;
wire n_16560;
wire n_16561;
wire n_16562;
wire n_16563;
wire n_16564;
wire n_16565;
wire n_16566;
wire n_16567;
wire n_16569;
wire n_1657;
wire n_16570;
wire TIMEBOOST_net_479;
wire n_16572;
wire n_16573;
wire n_16574;
wire n_16575;
wire n_16576;
wire n_16578;
wire n_16579;
wire n_1658;
wire n_16580;
wire n_16582;
wire n_16583;
wire n_16585;
wire n_16588;
wire TIMEBOOST_net_573;
wire n_1659;
wire n_16590;
wire n_16591;
wire n_16592;
wire n_16593;
wire n_16594;
wire n_16595;
wire n_16596;
wire n_16598;
wire n_16599;
wire n_166;
wire n_1660;
wire n_16600;
wire n_16601;
wire n_16602;
wire n_16603;
wire n_16604;
wire TIMEBOOST_net_700;
wire TIMEBOOST_net_2097;
wire n_16607;
wire n_16609;
wire n_16611;
wire n_16612;
wire n_16615;
wire n_16616;
wire n_16617;
wire n_16618;
wire n_16619;
wire n_1662;
wire n_16620;
wire n_16622;
wire n_16624;
wire n_16625;
wire n_16626;
wire n_16628;
wire n_16629;
wire n_1663;
wire n_16630;
wire n_16632;
wire n_16633;
wire n_16634;
wire n_16636;
wire n_16637;
wire n_16638;
wire n_16639;
wire n_1664;
wire n_16640;
wire n_16641;
wire TIMEBOOST_net_2917;
wire n_16643;
wire n_16645;
wire n_16646;
wire n_16648;
wire n_16649;
wire n_1665;
wire n_16650;
wire n_16653;
wire TIMEBOOST_net_2732;
wire n_16656;
wire n_16658;
wire n_1666;
wire n_16661;
wire n_16662;
wire TIMEBOOST_net_2336;
wire n_16665;
wire n_16667;
wire n_16668;
wire n_16669;
wire n_1667;
wire n_16670;
wire n_16671;
wire n_16673;
wire TIMEBOOST_net_485;
wire n_16675;
wire n_16676;
wire n_16677;
wire n_16678;
wire n_1668;
wire n_16681;
wire n_16682;
wire TIMEBOOST_net_1357;
wire n_16684;
wire n_16685;
wire n_16686;
wire n_1669;
wire n_16690;
wire n_16699;
wire n_167;
wire n_16700;
wire n_16702;
wire n_16703;
wire n_16705;
wire n_16706;
wire n_16707;
wire n_16708;
wire TIMEBOOST_net_2526;
wire n_1671;
wire TIMEBOOST_net_2098;
wire n_16712;
wire n_16713;
wire n_16714;
wire n_16715;
wire n_16716;
wire n_16717;
wire n_16719;
wire n_1672;
wire n_16721;
wire n_16722;
wire n_16723;
wire n_16725;
wire n_16726;
wire n_16727;
wire n_16728;
wire n_1673;
wire n_16730;
wire n_16731;
wire n_16732;
wire n_16733;
wire n_16734;
wire n_16735;
wire n_16736;
wire n_16737;
wire n_16739;
wire n_1674;
wire n_16741;
wire n_16742;
wire n_16743;
wire n_16744;
wire n_16745;
wire n_16747;
wire n_16748;
wire n_16749;
wire n_1675;
wire n_16750;
wire n_16751;
wire n_16752;
wire n_16753;
wire n_16755;
wire n_16757;
wire n_16758;
wire n_16759;
wire n_16760;
wire n_16761;
wire n_16762;
wire n_16763;
wire n_16764;
wire n_16767;
wire n_16768;
wire n_16770;
wire n_16772;
wire n_16774;
wire n_16777;
wire n_16778;
wire n_16779;
wire n_1678;
wire n_16781;
wire n_16782;
wire n_16784;
wire n_16785;
wire n_16787;
wire n_16789;
wire n_1679;
wire n_16791;
wire TIMEBOOST_net_761;
wire n_16793;
wire n_16796;
wire n_16798;
wire n_16799;
wire n_168;
wire n_16801;
wire n_16802;
wire n_16804;
wire n_16807;
wire n_16808;
wire n_16809;
wire n_1681;
wire n_16810;
wire n_16811;
wire n_16814;
wire n_16815;
wire n_16816;
wire n_16817;
wire n_16818;
wire n_16819;
wire n_1682;
wire n_16820;
wire n_16821;
wire n_16822;
wire n_16823;
wire n_16824;
wire n_16825;
wire n_16826;
wire n_16827;
wire n_16828;
wire n_16829;
wire n_16830;
wire n_16832;
wire n_16833;
wire n_16834;
wire TIMEBOOST_net_2739;
wire n_16836;
wire n_16837;
wire n_16838;
wire n_16839;
wire n_16840;
wire n_16843;
wire n_16846;
wire n_16847;
wire n_16849;
wire n_1685;
wire n_16850;
wire n_16851;
wire n_16852;
wire n_16853;
wire n_16854;
wire n_16855;
wire n_16857;
wire n_1686;
wire n_16863;
wire n_16864;
wire n_16865;
wire n_16866;
wire n_16867;
wire n_16868;
wire n_16869;
wire n_1687;
wire n_16872;
wire n_16873;
wire n_16874;
wire n_16876;
wire n_16879;
wire n_1688;
wire n_16880;
wire n_16882;
wire n_16883;
wire n_16884;
wire n_16885;
wire n_16886;
wire n_16887;
wire n_16888;
wire n_16889;
wire n_1689;
wire n_16890;
wire TIMEBOOST_net_2792;
wire n_16893;
wire n_16894;
wire n_16895;
wire TIMEBOOST_net_2096;
wire n_16899;
wire n_169;
wire n_1690;
wire n_16900;
wire n_16902;
wire n_16903;
wire n_16904;
wire n_16905;
wire n_16908;
wire n_16909;
wire n_1691;
wire n_16910;
wire n_16911;
wire n_16912;
wire TIMEBOOST_net_587;
wire n_16915;
wire n_16916;
wire n_16917;
wire n_16918;
wire n_16919;
wire n_1692;
wire n_16920;
wire n_16921;
wire n_16923;
wire n_16924;
wire n_16925;
wire n_16926;
wire n_16927;
wire n_16928;
wire n_16929;
wire n_16930;
wire n_16931;
wire TIMEBOOST_net_754;
wire n_16936;
wire n_16938;
wire n_1694;
wire n_16940;
wire n_16941;
wire n_16942;
wire n_16943;
wire n_16944;
wire n_16948;
wire n_1695;
wire n_16950;
wire n_16951;
wire n_16952;
wire n_16953;
wire n_16954;
wire n_16957;
wire TIMEBOOST_net_818;
wire n_16960;
wire n_16961;
wire n_16962;
wire n_16967;
wire n_16968;
wire TIMEBOOST_net_1846;
wire n_16970;
wire n_16972;
wire n_16973;
wire n_16976;
wire n_16977;
wire TIMEBOOST_net_651;
wire n_1698;
wire n_16984;
wire n_16986;
wire n_16987;
wire n_16988;
wire n_1699;
wire n_16990;
wire n_16991;
wire n_16993;
wire TIMEBOOST_net_1359;
wire n_16995;
wire n_16996;
wire n_16998;
wire n_16999;
wire n_170;
wire n_1700;
wire n_17001;
wire n_17002;
wire n_17003;
wire n_17004;
wire n_17005;
wire n_17006;
wire n_17007;
wire TIMEBOOST_net_2827;
wire n_17009;
wire n_1701;
wire n_17014;
wire n_17015;
wire n_17017;
wire n_17018;
wire n_1702;
wire n_17020;
wire n_17022;
wire n_17023;
wire n_17025;
wire n_17026;
wire n_17027;
wire n_17029;
wire n_1703;
wire n_17031;
wire n_17032;
wire n_17033;
wire n_17035;
wire n_17036;
wire n_17037;
wire n_17039;
wire n_1704;
wire n_17040;
wire n_17041;
wire n_17042;
wire n_17043;
wire n_17044;
wire n_17045;
wire TIMEBOOST_net_589;
wire TIMEBOOST_net_655;
wire n_17048;
wire n_17049;
wire n_1705;
wire n_17050;
wire n_17054;
wire n_17055;
wire n_17056;
wire n_17057;
wire n_17058;
wire n_1706;
wire n_17061;
wire n_17069;
wire n_1707;
wire n_17070;
wire n_17071;
wire n_17072;
wire n_17073;
wire TIMEBOOST_net_593;
wire n_1708;
wire n_17081;
wire n_17082;
wire n_17083;
wire n_17084;
wire n_17085;
wire n_17086;
wire TIMEBOOST_net_1358;
wire n_17088;
wire n_1709;
wire n_17090;
wire n_17091;
wire TIMEBOOST_net_762;
wire n_17093;
wire n_17096;
wire n_17097;
wire n_17098;
wire n_17099;
wire n_171;
wire n_17100;
wire n_17101;
wire n_17102;
wire n_17103;
wire n_17104;
wire TIMEBOOST_net_786;
wire n_17106;
wire n_17107;
wire n_17108;
wire n_1711;
wire n_17113;
wire n_17114;
wire n_17115;
wire n_17117;
wire n_17118;
wire n_17119;
wire n_1712;
wire n_17120;
wire n_17121;
wire n_17123;
wire n_17125;
wire n_17126;
wire n_17128;
wire n_17129;
wire n_1713;
wire n_17130;
wire n_17132;
wire n_17133;
wire n_17134;
wire n_17135;
wire n_17136;
wire n_17137;
wire n_17139;
wire n_1714;
wire n_17140;
wire n_17142;
wire n_17144;
wire n_17146;
wire n_17147;
wire n_1715;
wire n_17152;
wire n_17153;
wire n_17154;
wire n_17155;
wire n_17156;
wire n_17157;
wire n_17158;
wire n_17159;
wire TIMEBOOST_net_2559;
wire TIMEBOOST_net_2089;
wire TIMEBOOST_net_2749;
wire n_17167;
wire n_17169;
wire n_1717;
wire n_17170;
wire n_17171;
wire n_17172;
wire n_17174;
wire n_17176;
wire n_17177;
wire n_17178;
wire TIMEBOOST_net_594;
wire n_1718;
wire n_17180;
wire n_17185;
wire n_17186;
wire n_17187;
wire n_17188;
wire n_17189;
wire n_1719;
wire n_17190;
wire n_17191;
wire n_17192;
wire n_17193;
wire n_17194;
wire n_17195;
wire TIMEBOOST_net_1802;
wire n_17197;
wire n_17199;
wire n_172;
wire n_1720;
wire n_17200;
wire n_17201;
wire n_17202;
wire n_17207;
wire n_17208;
wire n_1721;
wire n_17210;
wire n_17211;
wire n_17212;
wire n_17213;
wire n_17214;
wire n_17215;
wire n_17216;
wire n_17217;
wire n_1722;
wire TIMEBOOST_net_2769;
wire n_17221;
wire n_17223;
wire n_17224;
wire n_17226;
wire n_17227;
wire n_17228;
wire n_17229;
wire n_17230;
wire n_17231;
wire n_17232;
wire n_17233;
wire n_17234;
wire n_17235;
wire n_17237;
wire n_17238;
wire n_17239;
wire n_1724;
wire n_17240;
wire TIMEBOOST_net_809;
wire n_17243;
wire n_17244;
wire n_17245;
wire n_17247;
wire TIMEBOOST_net_605;
wire n_17249;
wire n_1725;
wire n_17250;
wire n_17252;
wire n_17255;
wire n_17256;
wire n_17257;
wire n_17258;
wire n_17259;
wire n_17260;
wire n_17261;
wire n_17262;
wire n_17263;
wire n_17265;
wire n_17266;
wire n_17268;
wire n_17269;
wire n_1727;
wire n_17272;
wire n_17273;
wire n_17274;
wire n_17275;
wire TIMEBOOST_net_25;
wire n_17279;
wire n_1728;
wire n_17280;
wire n_17281;
wire n_17282;
wire n_17283;
wire n_17284;
wire n_17287;
wire n_17288;
wire n_17289;
wire n_1729;
wire n_17290;
wire n_17291;
wire n_17292;
wire TIMEBOOST_net_764;
wire n_17294;
wire n_17297;
wire n_17298;
wire n_17299;
wire n_173;
wire n_1730;
wire n_17300;
wire n_17301;
wire n_17302;
wire n_17304;
wire n_17305;
wire n_17306;
wire n_17308;
wire n_17309;
wire n_1731;
wire n_17310;
wire n_17311;
wire n_17312;
wire n_17313;
wire n_17314;
wire n_17315;
wire n_17316;
wire n_17317;
wire n_17318;
wire n_17319;
wire n_1732;
wire n_17320;
wire n_17321;
wire n_17322;
wire n_17323;
wire n_17324;
wire n_17325;
wire n_17326;
wire n_17327;
wire n_17328;
wire n_17329;
wire n_1733;
wire n_17330;
wire n_17331;
wire n_17332;
wire n_17333;
wire n_17334;
wire n_17335;
wire n_17336;
wire n_17337;
wire n_17339;
wire n_17340;
wire n_17341;
wire TIMEBOOST_net_813;
wire n_17343;
wire n_17344;
wire n_17345;
wire n_17346;
wire n_17347;
wire n_17348;
wire n_17349;
wire n_1735;
wire n_17350;
wire n_17353;
wire n_17354;
wire n_17355;
wire n_17356;
wire n_17357;
wire n_17358;
wire n_17359;
wire n_1736;
wire n_17360;
wire n_17362;
wire n_17363;
wire n_17364;
wire n_17365;
wire n_17366;
wire n_17367;
wire n_17368;
wire n_17369;
wire n_1737;
wire n_17370;
wire n_17371;
wire n_17372;
wire n_17373;
wire n_17374;
wire n_17375;
wire n_17376;
wire n_17377;
wire n_17378;
wire n_17379;
wire n_17380;
wire n_17381;
wire n_17382;
wire n_17383;
wire n_17384;
wire n_17385;
wire n_17386;
wire n_17387;
wire n_17388;
wire n_17389;
wire n_1739;
wire n_17390;
wire n_17391;
wire n_17392;
wire n_17393;
wire n_17394;
wire n_17395;
wire n_17396;
wire n_17397;
wire n_17398;
wire n_17399;
wire n_174;
wire n_17400;
wire n_17401;
wire n_17402;
wire n_17403;
wire n_17404;
wire n_17405;
wire n_17406;
wire n_17407;
wire n_17409;
wire n_1741;
wire n_17410;
wire TIMEBOOST_net_1481;
wire n_17414;
wire n_17415;
wire n_17416;
wire n_17417;
wire n_17418;
wire n_1742;
wire n_17421;
wire n_17422;
wire n_17423;
wire n_17424;
wire n_17425;
wire n_17426;
wire n_17427;
wire n_17428;
wire n_17429;
wire n_1743;
wire n_17430;
wire n_17431;
wire n_17432;
wire n_17433;
wire n_17434;
wire n_17435;
wire TIMEBOOST_net_1837;
wire n_17437;
wire n_17438;
wire n_17439;
wire n_1744;
wire n_17440;
wire n_17441;
wire n_17442;
wire TIMEBOOST_net_2122;
wire n_17444;
wire n_17445;
wire n_17446;
wire TIMEBOOST_net_2937;
wire n_17449;
wire n_1745;
wire n_17450;
wire n_17451;
wire n_17452;
wire TIMEBOOST_net_757;
wire n_17454;
wire n_17455;
wire n_17456;
wire n_17457;
wire n_17458;
wire n_17459;
wire n_1746;
wire n_17460;
wire n_17462;
wire n_17463;
wire n_17464;
wire n_17465;
wire n_17466;
wire n_17467;
wire n_17468;
wire n_17469;
wire n_17470;
wire n_17471;
wire n_17472;
wire n_17473;
wire n_17474;
wire n_17475;
wire n_17476;
wire n_17477;
wire n_17478;
wire n_17479;
wire n_1748;
wire n_17480;
wire n_17481;
wire n_17482;
wire n_17483;
wire n_17484;
wire n_17485;
wire n_17486;
wire n_17487;
wire n_17489;
wire n_1749;
wire n_17490;
wire n_17492;
wire n_17493;
wire n_17495;
wire n_17496;
wire n_17497;
wire n_17498;
wire n_17499;
wire n_175;
wire n_17502;
wire n_17503;
wire n_17504;
wire n_17505;
wire n_17507;
wire n_17508;
wire n_1751;
wire n_17510;
wire n_17512;
wire n_17513;
wire n_17514;
wire n_17515;
wire n_17516;
wire n_17517;
wire n_1752;
wire n_17522;
wire n_17523;
wire n_17526;
wire n_17527;
wire n_1753;
wire n_17530;
wire n_17531;
wire n_17532;
wire n_17533;
wire n_17535;
wire n_17536;
wire n_17537;
wire n_17539;
wire n_1754;
wire n_17540;
wire n_17541;
wire n_17542;
wire n_17543;
wire n_17544;
wire n_17545;
wire n_17546;
wire n_17547;
wire n_17548;
wire n_17549;
wire n_1755;
wire n_17550;
wire n_17552;
wire n_17553;
wire n_17554;
wire n_17555;
wire n_17556;
wire n_17557;
wire n_17558;
wire n_17559;
wire n_1756;
wire n_17560;
wire n_17561;
wire n_17562;
wire n_17565;
wire n_17566;
wire n_17567;
wire n_17568;
wire n_17572;
wire n_17573;
wire n_17574;
wire n_17575;
wire n_17576;
wire n_17577;
wire n_17578;
wire n_17579;
wire n_1758;
wire n_17580;
wire n_17581;
wire n_17582;
wire n_17584;
wire n_17585;
wire n_17587;
wire n_17588;
wire n_17589;
wire n_1759;
wire n_17590;
wire n_17591;
wire n_17592;
wire n_17593;
wire n_17594;
wire n_17595;
wire n_17597;
wire n_17598;
wire n_176;
wire n_1760;
wire n_17600;
wire n_17601;
wire n_17602;
wire n_17603;
wire n_17604;
wire n_17605;
wire n_17607;
wire n_17608;
wire n_17609;
wire n_1761;
wire n_17610;
wire n_17611;
wire n_17613;
wire n_17614;
wire n_17615;
wire n_17617;
wire n_17619;
wire n_1762;
wire n_17620;
wire n_17621;
wire n_17622;
wire n_17623;
wire n_17624;
wire n_17625;
wire n_17626;
wire n_17627;
wire n_17628;
wire n_17629;
wire n_1763;
wire n_17630;
wire n_17632;
wire n_17633;
wire n_17634;
wire n_17635;
wire n_17636;
wire n_17637;
wire n_17638;
wire n_17639;
wire n_1764;
wire n_17640;
wire n_17641;
wire n_17642;
wire n_17643;
wire n_17644;
wire n_17647;
wire n_17649;
wire n_1765;
wire n_17654;
wire n_17655;
wire n_17656;
wire n_17657;
wire n_17658;
wire n_17659;
wire n_1766;
wire n_17660;
wire n_17661;
wire n_17663;
wire n_17665;
wire n_17667;
wire n_17669;
wire n_1767;
wire n_17672;
wire n_17674;
wire n_17677;
wire n_17678;
wire n_17679;
wire n_1768;
wire n_17680;
wire n_17682;
wire n_17683;
wire n_17684;
wire n_17685;
wire n_17686;
wire n_17687;
wire n_17688;
wire n_17689;
wire n_1769;
wire n_17692;
wire n_17693;
wire n_17694;
wire n_17695;
wire n_17696;
wire n_17697;
wire n_17698;
wire n_177;
wire n_1770;
wire n_17700;
wire n_17702;
wire n_17703;
wire n_17704;
wire n_17705;
wire n_17706;
wire n_17707;
wire n_17708;
wire n_17709;
wire n_1771;
wire n_17710;
wire n_17711;
wire n_17712;
wire n_17713;
wire TIMEBOOST_net_781;
wire n_17715;
wire n_17717;
wire n_17718;
wire n_17719;
wire n_1772;
wire n_17720;
wire n_17721;
wire n_17722;
wire n_17723;
wire n_17724;
wire n_17725;
wire n_17726;
wire n_17727;
wire n_17728;
wire n_17729;
wire n_1773;
wire n_17731;
wire n_17732;
wire n_17734;
wire n_17736;
wire n_17737;
wire n_17738;
wire n_17739;
wire n_1774;
wire n_17740;
wire n_17741;
wire n_17742;
wire n_17743;
wire n_17744;
wire n_17745;
wire n_17746;
wire n_17747;
wire n_17748;
wire n_17749;
wire n_17750;
wire n_17752;
wire n_17753;
wire n_17754;
wire n_17755;
wire n_17756;
wire n_17758;
wire n_17759;
wire n_1776;
wire n_17762;
wire n_17763;
wire n_17765;
wire n_17766;
wire n_17769;
wire n_17770;
wire n_17771;
wire n_17772;
wire n_17773;
wire n_17776;
wire n_17777;
wire n_17778;
wire n_17779;
wire n_1778;
wire n_17780;
wire n_17781;
wire n_17782;
wire n_17783;
wire n_17785;
wire n_17786;
wire n_17787;
wire n_17788;
wire n_17789;
wire n_1779;
wire n_17790;
wire n_17791;
wire n_17792;
wire n_17793;
wire n_17794;
wire n_17795;
wire n_17796;
wire n_17797;
wire n_17798;
wire n_17799;
wire n_178;
wire n_1780;
wire n_17800;
wire n_17801;
wire n_17802;
wire n_17803;
wire TIMEBOOST_net_2809;
wire n_17805;
wire n_17806;
wire n_17808;
wire n_17809;
wire n_1781;
wire n_17811;
wire n_17812;
wire n_17813;
wire n_17815;
wire n_17816;
wire n_17817;
wire n_17818;
wire n_17819;
wire n_1782;
wire n_17820;
wire n_17822;
wire n_17823;
wire n_17824;
wire n_17825;
wire n_17826;
wire n_17827;
wire n_17828;
wire n_17829;
wire n_1783;
wire n_17832;
wire n_17834;
wire n_17835;
wire n_17836;
wire n_17838;
wire n_17839;
wire n_1784;
wire n_17840;
wire n_17841;
wire n_17842;
wire n_17843;
wire n_17845;
wire n_17846;
wire n_17847;
wire n_17848;
wire n_17849;
wire n_1785;
wire n_17850;
wire n_17851;
wire n_17852;
wire n_17855;
wire n_17856;
wire n_17859;
wire n_17860;
wire n_17862;
wire n_17863;
wire n_17864;
wire n_17865;
wire n_17866;
wire n_17867;
wire n_17868;
wire n_17869;
wire n_1787;
wire n_17870;
wire TIMEBOOST_net_2171;
wire n_17872;
wire n_17873;
wire n_17875;
wire n_17878;
wire n_17879;
wire n_17880;
wire n_17881;
wire n_17882;
wire n_17883;
wire n_17884;
wire n_17885;
wire n_17886;
wire n_17887;
wire n_17888;
wire n_17889;
wire n_1789;
wire n_17890;
wire n_17891;
wire n_17892;
wire n_17893;
wire n_17894;
wire n_17895;
wire n_17896;
wire n_17897;
wire n_179;
wire n_1790;
wire n_17900;
wire n_17902;
wire n_17903;
wire n_17904;
wire n_17905;
wire n_17906;
wire n_17907;
wire n_17908;
wire n_17909;
wire n_1791;
wire n_17910;
wire n_17911;
wire n_17912;
wire n_17913;
wire n_17914;
wire n_17915;
wire n_17916;
wire n_17917;
wire n_17918;
wire n_17919;
wire n_1792;
wire n_17920;
wire n_17921;
wire n_17922;
wire n_17923;
wire n_17924;
wire n_17925;
wire n_17926;
wire n_17927;
wire n_17928;
wire n_17929;
wire n_17930;
wire n_17931;
wire n_17932;
wire n_17937;
wire TIMEBOOST_net_2938;
wire n_17939;
wire n_1794;
wire n_17940;
wire n_17941;
wire n_17942;
wire n_17943;
wire n_17944;
wire n_17945;
wire n_17946;
wire n_17947;
wire n_17948;
wire n_17949;
wire n_1795;
wire n_17950;
wire n_17951;
wire n_17952;
wire n_17953;
wire n_17954;
wire n_17958;
wire n_17959;
wire n_17960;
wire n_17961;
wire n_17962;
wire n_17963;
wire n_17964;
wire n_17965;
wire n_17966;
wire n_17967;
wire n_1797;
wire n_17970;
wire n_17971;
wire n_17972;
wire n_17973;
wire n_17975;
wire n_17977;
wire n_1798;
wire n_17980;
wire n_17981;
wire n_17982;
wire n_17983;
wire n_17984;
wire n_17985;
wire n_17986;
wire n_17987;
wire n_17988;
wire n_17989;
wire n_1799;
wire n_17990;
wire n_17991;
wire n_17992;
wire n_17993;
wire n_17994;
wire n_17995;
wire n_17996;
wire n_17997;
wire n_17999;
wire n_18;
wire n_180;
wire n_1800;
wire n_18000;
wire n_18001;
wire n_18002;
wire n_18003;
wire n_18004;
wire n_18005;
wire n_18006;
wire n_18008;
wire n_18009;
wire n_1801;
wire n_18010;
wire n_18013;
wire n_18015;
wire n_18016;
wire n_18017;
wire n_18018;
wire n_18019;
wire n_1802;
wire n_18020;
wire n_18021;
wire n_18022;
wire n_18023;
wire n_18024;
wire n_18025;
wire n_18026;
wire n_1803;
wire n_18032;
wire n_18033;
wire n_18034;
wire n_18035;
wire n_18036;
wire n_18037;
wire n_18038;
wire n_18039;
wire n_1804;
wire n_18040;
wire n_18041;
wire n_18042;
wire n_18043;
wire n_18045;
wire n_18046;
wire TIMEBOOST_net_1687;
wire n_18048;
wire n_18049;
wire n_1805;
wire n_18050;
wire n_18051;
wire n_18052;
wire n_18054;
wire n_18055;
wire n_18056;
wire n_18057;
wire n_18058;
wire n_18059;
wire n_1806;
wire n_18060;
wire n_18061;
wire n_18064;
wire n_18065;
wire n_18066;
wire n_18067;
wire n_18068;
wire n_18069;
wire n_18070;
wire n_18071;
wire n_18072;
wire TIMEBOOST_net_1760;
wire n_18074;
wire n_18075;
wire n_18076;
wire n_18077;
wire n_18078;
wire n_18079;
wire n_1808;
wire n_18080;
wire n_18083;
wire n_18084;
wire n_18085;
wire TIMEBOOST_net_871;
wire n_18087;
wire n_18088;
wire n_18089;
wire n_1809;
wire n_18090;
wire n_18091;
wire n_18092;
wire n_18093;
wire TIMEBOOST_net_1759;
wire n_18095;
wire n_18096;
wire TIMEBOOST_net_51;
wire n_18099;
wire n_181;
wire n_1810;
wire n_18102;
wire n_18103;
wire n_18104;
wire n_18105;
wire n_18106;
wire n_18107;
wire n_18108;
wire n_18109;
wire n_1811;
wire n_18110;
wire n_18111;
wire n_18112;
wire n_18113;
wire n_18114;
wire n_18115;
wire TIMEBOOST_net_2132;
wire n_18117;
wire n_18119;
wire n_1812;
wire n_18123;
wire n_18124;
wire n_18125;
wire n_18126;
wire n_18127;
wire n_18128;
wire n_18129;
wire n_1813;
wire n_18130;
wire n_18133;
wire n_18134;
wire n_18135;
wire n_18136;
wire n_18137;
wire n_18138;
wire n_1814;
wire n_18140;
wire n_18141;
wire n_18142;
wire n_18146;
wire n_18148;
wire n_18149;
wire n_1815;
wire n_18150;
wire n_18152;
wire n_18153;
wire n_18156;
wire n_18157;
wire n_18158;
wire n_18159;
wire n_18160;
wire n_18161;
wire n_18162;
wire n_18163;
wire n_18164;
wire n_18165;
wire TIMEBOOST_net_2312;
wire n_18167;
wire n_18168;
wire n_18169;
wire n_1817;
wire TIMEBOOST_net_894;
wire n_18171;
wire n_18173;
wire n_18174;
wire n_18175;
wire n_18176;
wire n_18177;
wire n_18178;
wire n_18179;
wire n_1818;
wire n_18180;
wire n_18183;
wire n_18184;
wire n_18185;
wire n_18186;
wire n_18187;
wire n_18188;
wire n_18189;
wire n_1819;
wire n_18190;
wire TIMEBOOST_net_1756;
wire n_18193;
wire n_18194;
wire n_18195;
wire n_18196;
wire n_18197;
wire n_18198;
wire n_18199;
wire n_182;
wire n_1820;
wire n_18200;
wire n_18201;
wire n_18202;
wire n_18204;
wire n_18205;
wire n_18206;
wire n_18208;
wire n_1821;
wire n_18210;
wire n_18211;
wire n_18212;
wire n_18213;
wire n_18214;
wire n_18215;
wire n_18216;
wire n_18217;
wire n_18218;
wire n_18219;
wire n_1822;
wire n_18220;
wire n_18221;
wire n_18222;
wire n_18223;
wire n_18224;
wire n_18225;
wire n_18226;
wire TIMEBOOST_net_2009;
wire n_18230;
wire n_18231;
wire n_18232;
wire n_18234;
wire n_18235;
wire n_18236;
wire n_18237;
wire n_18238;
wire n_18239;
wire n_1824;
wire n_18240;
wire n_18241;
wire n_18242;
wire n_18243;
wire n_18244;
wire n_18245;
wire n_18246;
wire n_18247;
wire n_18248;
wire n_1825;
wire n_18251;
wire n_18252;
wire n_18253;
wire n_18254;
wire n_18255;
wire n_18256;
wire n_18257;
wire n_18259;
wire n_18260;
wire n_18261;
wire n_18262;
wire n_18263;
wire n_18264;
wire n_18265;
wire n_18266;
wire n_18267;
wire n_18268;
wire n_18269;
wire n_1827;
wire n_18271;
wire n_18276;
wire n_18277;
wire n_18278;
wire n_18279;
wire n_18280;
wire n_18282;
wire n_18283;
wire n_18284;
wire n_18285;
wire TIMEBOOST_net_2759;
wire n_18287;
wire n_1829;
wire n_18291;
wire n_18293;
wire n_18294;
wire n_18295;
wire n_18298;
wire n_183;
wire n_1830;
wire n_18300;
wire n_18301;
wire n_18302;
wire n_18309;
wire n_18310;
wire n_18311;
wire n_18313;
wire n_18316;
wire n_18317;
wire n_18318;
wire n_18319;
wire n_1832;
wire n_18320;
wire n_18321;
wire n_18322;
wire n_18323;
wire n_18324;
wire n_18326;
wire n_18327;
wire n_18328;
wire n_18329;
wire n_1833;
wire n_18331;
wire n_18332;
wire n_18333;
wire n_18334;
wire n_18335;
wire n_18336;
wire n_18337;
wire n_18339;
wire n_1834;
wire n_18343;
wire n_18345;
wire n_18346;
wire n_18347;
wire n_18348;
wire n_1835;
wire n_18350;
wire n_18351;
wire n_18352;
wire n_18354;
wire n_18355;
wire n_18356;
wire n_18357;
wire n_1836;
wire n_18360;
wire n_18366;
wire n_18367;
wire n_18368;
wire n_1837;
wire n_18370;
wire n_18371;
wire n_18372;
wire n_18373;
wire TIMEBOOST_net_2149;
wire n_18375;
wire n_18376;
wire n_18377;
wire TIMEBOOST_net_87;
wire n_18379;
wire n_1838;
wire n_18380;
wire n_18382;
wire n_18383;
wire n_18384;
wire n_18385;
wire n_18386;
wire n_18387;
wire TIMEBOOST_net_2176;
wire n_18390;
wire n_18391;
wire n_18392;
wire n_18393;
wire n_18394;
wire n_18395;
wire n_18396;
wire n_18397;
wire n_18398;
wire n_1840;
wire TIMEBOOST_net_2798;
wire n_18401;
wire n_18404;
wire n_18405;
wire n_18406;
wire n_18407;
wire n_18408;
wire n_18409;
wire n_18411;
wire n_18412;
wire n_18414;
wire n_18415;
wire n_18416;
wire n_18417;
wire n_18418;
wire n_18419;
wire n_1842;
wire n_18420;
wire n_18421;
wire n_18422;
wire n_18424;
wire n_18425;
wire n_18426;
wire n_18427;
wire n_18428;
wire n_1843;
wire n_18431;
wire n_18432;
wire n_18433;
wire n_18434;
wire n_18435;
wire n_18436;
wire n_18437;
wire n_18438;
wire n_18439;
wire n_1844;
wire n_18440;
wire n_18441;
wire n_18443;
wire n_18444;
wire n_18445;
wire n_18446;
wire n_18448;
wire n_18449;
wire n_1845;
wire n_18450;
wire n_18451;
wire n_18452;
wire n_18453;
wire n_18455;
wire n_18456;
wire n_18457;
wire n_18458;
wire n_18459;
wire n_1846;
wire n_18460;
wire n_18461;
wire n_18462;
wire n_18467;
wire n_18468;
wire n_1847;
wire n_18470;
wire n_18472;
wire n_18473;
wire n_18475;
wire n_18476;
wire n_18477;
wire n_18478;
wire n_18479;
wire n_1848;
wire n_18480;
wire n_18481;
wire n_18482;
wire n_18483;
wire n_18484;
wire n_18487;
wire n_18488;
wire n_18490;
wire n_18492;
wire n_18494;
wire n_18495;
wire n_18496;
wire n_18497;
wire n_18498;
wire n_18499;
wire n_1850;
wire n_18500;
wire n_18501;
wire n_18505;
wire n_18506;
wire n_18507;
wire n_18508;
wire n_18509;
wire n_1851;
wire n_18510;
wire n_18511;
wire n_18512;
wire n_18513;
wire n_18514;
wire n_18515;
wire n_18516;
wire n_18517;
wire n_18518;
wire n_18519;
wire n_1852;
wire n_18520;
wire n_18521;
wire n_18522;
wire n_18523;
wire n_18524;
wire n_18526;
wire n_18528;
wire n_18529;
wire n_1853;
wire n_18531;
wire n_18532;
wire n_18533;
wire n_18534;
wire n_18535;
wire n_18536;
wire n_18537;
wire n_18538;
wire n_18539;
wire n_1854;
wire n_18540;
wire n_18541;
wire n_18544;
wire n_18545;
wire n_18546;
wire n_18547;
wire n_18548;
wire n_18549;
wire n_1855;
wire n_18550;
wire n_18553;
wire n_18554;
wire n_18555;
wire n_18557;
wire n_18559;
wire n_1856;
wire n_18560;
wire n_18561;
wire n_18562;
wire n_18563;
wire n_18564;
wire n_18565;
wire TIMEBOOST_net_100;
wire n_18568;
wire n_18569;
wire n_1857;
wire n_18571;
wire n_18572;
wire n_18574;
wire n_18575;
wire n_18576;
wire n_18577;
wire n_18578;
wire n_18579;
wire n_1858;
wire n_18580;
wire n_18581;
wire n_18582;
wire n_18583;
wire n_18584;
wire n_18585;
wire n_18586;
wire n_18587;
wire n_18589;
wire n_1859;
wire n_18590;
wire n_18591;
wire n_18592;
wire n_18593;
wire n_18594;
wire n_18595;
wire n_18599;
wire n_186;
wire n_1860;
wire n_18600;
wire TIMEBOOST_net_2790;
wire n_18602;
wire n_18607;
wire n_18608;
wire n_18609;
wire n_1861;
wire n_18610;
wire n_18611;
wire n_18612;
wire n_18613;
wire n_18614;
wire n_18615;
wire n_18616;
wire n_18617;
wire n_18618;
wire n_18619;
wire n_1862;
wire n_18620;
wire n_18622;
wire n_18623;
wire n_18624;
wire n_18625;
wire n_18626;
wire n_18627;
wire n_18629;
wire n_1863;
wire n_18630;
wire n_18631;
wire n_18633;
wire n_18634;
wire n_18637;
wire n_18638;
wire n_18639;
wire n_1864;
wire n_18640;
wire n_18641;
wire n_18642;
wire n_18645;
wire n_18646;
wire n_18647;
wire n_18649;
wire n_1865;
wire n_18650;
wire n_18652;
wire n_18653;
wire n_18655;
wire n_18657;
wire n_18658;
wire n_18659;
wire n_1866;
wire n_18660;
wire n_18661;
wire n_18663;
wire n_18664;
wire n_18665;
wire n_18666;
wire n_18667;
wire n_18668;
wire n_18669;
wire n_18670;
wire n_18672;
wire n_18674;
wire n_18675;
wire n_18678;
wire n_18681;
wire n_18682;
wire n_18683;
wire n_18684;
wire n_18688;
wire n_18689;
wire n_1869;
wire n_18692;
wire n_18693;
wire n_18694;
wire n_18695;
wire n_18696;
wire n_18697;
wire n_18698;
wire n_18700;
wire n_18701;
wire n_18702;
wire n_18703;
wire n_18704;
wire n_18705;
wire n_18706;
wire n_18707;
wire n_18708;
wire n_18709;
wire n_1871;
wire n_18710;
wire n_18713;
wire n_18716;
wire n_18717;
wire n_18718;
wire TIMEBOOST_net_140;
wire n_18721;
wire n_18722;
wire n_18723;
wire n_18724;
wire n_18725;
wire n_18726;
wire n_18727;
wire n_18728;
wire n_18729;
wire n_1873;
wire n_18730;
wire n_18731;
wire n_18734;
wire n_18735;
wire n_18736;
wire n_18737;
wire n_18738;
wire n_18739;
wire n_1874;
wire n_18741;
wire n_18742;
wire n_18743;
wire n_18744;
wire n_18745;
wire n_18746;
wire n_18748;
wire n_18749;
wire n_1875;
wire n_18750;
wire n_18754;
wire n_18756;
wire n_18757;
wire n_18758;
wire n_1876;
wire n_18760;
wire n_18761;
wire n_18765;
wire n_18766;
wire n_18767;
wire n_18769;
wire n_1877;
wire n_18771;
wire n_18772;
wire n_18773;
wire n_18774;
wire n_18775;
wire n_18776;
wire n_18777;
wire n_18778;
wire n_18779;
wire n_1878;
wire n_18780;
wire n_18781;
wire n_18784;
wire n_18785;
wire n_18786;
wire n_18787;
wire n_18789;
wire n_1879;
wire n_18791;
wire n_18794;
wire n_18795;
wire n_18797;
wire n_18798;
wire n_18799;
wire n_188;
wire n_1880;
wire n_18801;
wire n_18807;
wire n_18808;
wire n_18809;
wire n_1881;
wire n_18810;
wire n_18811;
wire n_18812;
wire n_18813;
wire n_18814;
wire n_18815;
wire n_18816;
wire n_18817;
wire n_18818;
wire n_1882;
wire n_18820;
wire n_18821;
wire n_18822;
wire n_18824;
wire n_18825;
wire n_18826;
wire n_18828;
wire n_18829;
wire n_1883;
wire n_18831;
wire n_18832;
wire n_18834;
wire n_18835;
wire n_18836;
wire n_18837;
wire n_18838;
wire n_18839;
wire n_1884;
wire n_18840;
wire n_18841;
wire n_18843;
wire n_18845;
wire n_18846;
wire n_18847;
wire n_18848;
wire n_18849;
wire n_1885;
wire n_18850;
wire n_18851;
wire n_18852;
wire n_18853;
wire n_18854;
wire n_18855;
wire TIMEBOOST_net_117;
wire n_18858;
wire n_18859;
wire n_1886;
wire n_18860;
wire n_18861;
wire n_18862;
wire n_18863;
wire n_18864;
wire n_18866;
wire n_18869;
wire n_1887;
wire n_18870;
wire n_18871;
wire TIMEBOOST_net_181;
wire n_18873;
wire n_18875;
wire n_18876;
wire n_1888;
wire n_18882;
wire n_18883;
wire n_18884;
wire n_18885;
wire n_18886;
wire n_18887;
wire n_18888;
wire TIMEBOOST_net_960;
wire n_1889;
wire n_18890;
wire n_18892;
wire n_18893;
wire n_18894;
wire n_18895;
wire n_18896;
wire n_18899;
wire n_189;
wire n_1890;
wire TIMEBOOST_net_190;
wire n_18901;
wire n_1891;
wire n_18910;
wire n_18911;
wire n_18912;
wire n_18913;
wire n_18914;
wire n_18915;
wire n_18916;
wire n_18918;
wire n_18919;
wire n_1892;
wire n_18920;
wire TIMEBOOST_net_1803;
wire TIMEBOOST_net_965;
wire TIMEBOOST_net_193;
wire n_18925;
wire n_18930;
wire n_18931;
wire n_18932;
wire n_18934;
wire n_18935;
wire n_18936;
wire n_18937;
wire n_18938;
wire n_18939;
wire n_1894;
wire n_18940;
wire n_18942;
wire n_18945;
wire n_18947;
wire n_18948;
wire n_18949;
wire n_1895;
wire n_18950;
wire n_18951;
wire n_18952;
wire n_18953;
wire n_18954;
wire n_18955;
wire n_18956;
wire n_18963;
wire n_18964;
wire n_18966;
wire n_18968;
wire n_18969;
wire n_18970;
wire n_18971;
wire n_18974;
wire n_18978;
wire n_1898;
wire n_18980;
wire n_18981;
wire n_18982;
wire n_18984;
wire n_18985;
wire n_18986;
wire n_18987;
wire TIMEBOOST_net_148;
wire n_18989;
wire n_1899;
wire n_18990;
wire n_18992;
wire n_18993;
wire n_18994;
wire n_18995;
wire n_18996;
wire n_18997;
wire n_18998;
wire n_18999;
wire n_190;
wire n_1900;
wire n_19000;
wire n_19002;
wire n_19003;
wire TIMEBOOST_net_1524;
wire n_19005;
wire n_19006;
wire n_19008;
wire TIMEBOOST_net_2888;
wire n_1901;
wire n_19010;
wire n_19011;
wire TIMEBOOST_net_1769;
wire n_19014;
wire TIMEBOOST_net_864;
wire n_19019;
wire n_1902;
wire n_19020;
wire n_19021;
wire n_19022;
wire n_19023;
wire n_19024;
wire n_19025;
wire n_19026;
wire n_19027;
wire n_19028;
wire n_19029;
wire n_1903;
wire n_19030;
wire n_19032;
wire n_19033;
wire n_19035;
wire TIMEBOOST_net_1025;
wire n_19037;
wire n_19038;
wire TIMEBOOST_net_1024;
wire n_1904;
wire n_19041;
wire n_19044;
wire TIMEBOOST_net_1856;
wire n_19046;
wire n_19049;
wire n_1905;
wire n_19050;
wire n_19051;
wire n_19053;
wire n_19054;
wire n_19055;
wire n_19056;
wire n_19058;
wire n_19059;
wire n_19060;
wire n_19062;
wire n_19064;
wire n_19070;
wire n_19071;
wire n_19072;
wire n_19073;
wire TIMEBOOST_net_882;
wire n_19075;
wire n_19076;
wire n_19077;
wire n_19078;
wire n_1908;
wire n_19080;
wire n_19081;
wire n_19082;
wire n_19083;
wire n_19084;
wire n_19087;
wire n_19088;
wire n_19089;
wire n_1909;
wire n_19096;
wire n_19097;
wire n_19098;
wire n_19099;
wire n_1910;
wire n_19101;
wire n_19104;
wire n_19105;
wire n_19106;
wire n_19107;
wire n_19108;
wire n_1911;
wire n_19110;
wire n_19112;
wire TIMEBOOST_net_1058;
wire n_19114;
wire n_19115;
wire n_19116;
wire n_19119;
wire n_19125;
wire n_19126;
wire n_19127;
wire n_19128;
wire n_19129;
wire n_1913;
wire n_19130;
wire n_19133;
wire n_19134;
wire n_19135;
wire n_19138;
wire n_19139;
wire n_19140;
wire n_19141;
wire n_19142;
wire n_19143;
wire n_19144;
wire n_19146;
wire n_19147;
wire n_19148;
wire n_1915;
wire n_19150;
wire TIMEBOOST_net_205;
wire n_19152;
wire n_19153;
wire n_19154;
wire n_19158;
wire n_19159;
wire n_1916;
wire n_19160;
wire n_19161;
wire n_19164;
wire n_19166;
wire n_19167;
wire n_19168;
wire n_19169;
wire n_1917;
wire n_19170;
wire n_19171;
wire n_19172;
wire n_19173;
wire n_19174;
wire n_19175;
wire n_19177;
wire n_19178;
wire n_1918;
wire n_19180;
wire n_19181;
wire n_19182;
wire TIMEBOOST_net_983;
wire n_19184;
wire TIMEBOOST_net_1812;
wire n_19186;
wire n_19187;
wire n_19188;
wire n_1919;
wire n_19191;
wire n_19193;
wire n_19194;
wire n_19195;
wire n_19196;
wire n_19197;
wire n_19198;
wire n_1920;
wire n_19200;
wire n_19201;
wire n_19202;
wire n_19203;
wire n_19206;
wire n_19207;
wire TIMEBOOST_net_2409;
wire n_1921;
wire n_19210;
wire n_19212;
wire n_19213;
wire TIMEBOOST_net_225;
wire n_19215;
wire TIMEBOOST_net_1862;
wire TIMEBOOST_net_1091;
wire n_19218;
wire n_19219;
wire TIMEBOOST_net_1777;
wire n_19222;
wire n_19223;
wire n_19225;
wire n_19228;
wire n_19229;
wire n_1923;
wire n_19230;
wire n_19231;
wire n_19232;
wire n_19233;
wire n_19236;
wire n_19237;
wire n_19238;
wire n_1924;
wire n_19241;
wire n_19243;
wire n_19245;
wire n_19246;
wire n_19247;
wire n_19248;
wire n_19249;
wire n_1925;
wire n_19250;
wire TIMEBOOST_net_1547;
wire TIMEBOOST_net_1930;
wire n_19255;
wire n_19256;
wire n_19262;
wire n_19264;
wire n_19268;
wire n_1927;
wire n_19270;
wire n_19271;
wire n_19272;
wire n_19273;
wire n_19274;
wire TIMEBOOST_net_207;
wire TIMEBOOST_net_209;
wire n_19277;
wire n_19278;
wire n_19279;
wire n_1928;
wire n_19280;
wire n_19281;
wire TIMEBOOST_net_991;
wire TIMEBOOST_net_147;
wire n_19284;
wire n_19285;
wire n_19286;
wire n_19287;
wire n_1929;
wire n_19291;
wire n_19292;
wire n_19293;
wire n_19294;
wire n_19295;
wire n_19296;
wire n_19297;
wire n_193;
wire n_1930;
wire n_19300;
wire n_19301;
wire n_19308;
wire n_19309;
wire n_1931;
wire n_19310;
wire n_19313;
wire n_19314;
wire n_19315;
wire n_19317;
wire n_19318;
wire n_19319;
wire n_1932;
wire TIMEBOOST_net_1099;
wire n_19322;
wire n_19323;
wire n_19324;
wire n_19325;
wire n_19327;
wire n_19328;
wire n_19329;
wire n_1933;
wire n_19330;
wire n_19331;
wire n_19332;
wire n_19333;
wire n_19334;
wire n_19335;
wire n_19337;
wire n_19339;
wire n_1934;
wire n_19342;
wire n_19344;
wire n_19345;
wire n_19346;
wire n_19347;
wire n_19348;
wire n_19349;
wire n_1935;
wire n_19350;
wire TIMEBOOST_net_1610;
wire n_19353;
wire n_19354;
wire n_19355;
wire n_19357;
wire n_19358;
wire n_1936;
wire n_19360;
wire n_19362;
wire n_19363;
wire n_19364;
wire n_19365;
wire TIMEBOOST_net_2794;
wire n_19367;
wire n_19368;
wire n_19369;
wire n_19370;
wire n_19372;
wire n_19374;
wire n_19375;
wire n_19377;
wire n_19378;
wire n_1938;
wire n_19380;
wire n_19381;
wire n_19382;
wire n_19383;
wire n_19384;
wire n_19385;
wire n_19386;
wire n_19387;
wire n_19388;
wire n_1939;
wire n_19390;
wire n_19391;
wire n_19393;
wire n_19398;
wire n_19399;
wire n_194;
wire n_1940;
wire n_19400;
wire n_19401;
wire n_19402;
wire n_19404;
wire n_19405;
wire n_19406;
wire n_19407;
wire n_19408;
wire n_1941;
wire n_19414;
wire n_19416;
wire n_19417;
wire n_19418;
wire n_19419;
wire n_1942;
wire n_19420;
wire n_19421;
wire n_19422;
wire n_19423;
wire TIMEBOOST_net_212;
wire n_19425;
wire n_19427;
wire n_19428;
wire n_1943;
wire n_19430;
wire TIMEBOOST_net_170;
wire n_19434;
wire n_19435;
wire n_19436;
wire n_19437;
wire n_19438;
wire TIMEBOOST_net_1720;
wire TIMEBOOST_net_2326;
wire n_19441;
wire n_19442;
wire n_19445;
wire n_19446;
wire n_19449;
wire n_1945;
wire n_19450;
wire n_19451;
wire n_19453;
wire n_19454;
wire n_19455;
wire n_19456;
wire n_19457;
wire n_19458;
wire TIMEBOOST_net_1030;
wire n_1946;
wire TIMEBOOST_net_1613;
wire n_19461;
wire n_19462;
wire n_19463;
wire n_19465;
wire n_19466;
wire n_19467;
wire n_19468;
wire n_19469;
wire n_1947;
wire n_19470;
wire n_19472;
wire TIMEBOOST_net_2191;
wire n_19474;
wire n_19475;
wire n_19476;
wire n_19477;
wire n_19478;
wire TIMEBOOST_net_879;
wire TIMEBOOST_net_922;
wire n_19485;
wire n_19486;
wire n_19487;
wire n_19488;
wire n_19489;
wire n_1949;
wire n_19490;
wire n_19491;
wire n_19492;
wire n_19493;
wire n_19494;
wire n_19496;
wire n_19497;
wire n_19498;
wire n_19499;
wire n_1950;
wire n_19500;
wire n_19501;
wire n_19502;
wire n_19505;
wire n_19506;
wire n_19507;
wire n_19508;
wire n_19509;
wire n_1951;
wire n_19510;
wire n_19511;
wire n_19512;
wire n_19513;
wire n_19514;
wire n_19516;
wire n_19517;
wire n_19518;
wire n_19519;
wire n_1952;
wire n_19520;
wire n_19521;
wire n_19522;
wire n_19523;
wire n_19524;
wire n_19525;
wire n_19526;
wire n_19528;
wire n_1953;
wire n_19530;
wire n_19531;
wire n_19532;
wire n_19533;
wire n_19534;
wire n_19535;
wire n_19537;
wire n_19538;
wire n_19539;
wire n_19540;
wire n_19541;
wire n_19542;
wire n_19543;
wire n_19544;
wire n_19545;
wire n_19546;
wire n_19547;
wire n_19548;
wire n_19549;
wire n_1955;
wire n_19552;
wire n_19553;
wire n_19555;
wire n_19556;
wire n_1956;
wire n_19561;
wire n_19562;
wire n_19563;
wire n_19564;
wire n_19565;
wire n_19566;
wire TIMEBOOST_net_408;
wire n_19568;
wire n_19569;
wire n_1957;
wire n_19570;
wire n_19571;
wire n_19572;
wire n_19573;
wire n_19574;
wire n_19575;
wire n_19576;
wire n_19577;
wire n_19578;
wire n_19579;
wire n_1958;
wire n_19580;
wire n_19581;
wire n_19583;
wire n_19585;
wire n_19587;
wire n_19588;
wire n_19589;
wire n_1959;
wire n_19590;
wire n_19591;
wire n_19592;
wire n_19593;
wire n_19594;
wire n_19595;
wire TIMEBOOST_net_173;
wire n_19597;
wire n_19599;
wire n_1960;
wire n_19601;
wire n_19602;
wire n_19603;
wire TIMEBOOST_net_1888;
wire n_19605;
wire TIMEBOOST_net_1173;
wire n_19607;
wire n_19608;
wire n_19609;
wire n_1961;
wire n_19610;
wire n_19611;
wire n_19612;
wire n_19613;
wire n_19615;
wire n_19616;
wire n_19617;
wire n_19618;
wire n_1962;
wire n_19621;
wire n_19623;
wire n_19624;
wire n_19625;
wire n_19626;
wire n_19627;
wire TIMEBOOST_net_2839;
wire TIMEBOOST_net_2956;
wire n_19633;
wire n_19634;
wire n_19635;
wire n_19636;
wire n_19637;
wire TIMEBOOST_net_179;
wire n_19639;
wire n_1964;
wire TIMEBOOST_net_2408;
wire n_19641;
wire n_19642;
wire TIMEBOOST_net_1001;
wire n_19645;
wire n_19646;
wire n_19647;
wire n_19648;
wire n_19649;
wire n_1965;
wire n_19650;
wire n_19651;
wire n_19652;
wire n_19653;
wire n_19654;
wire n_19656;
wire n_19658;
wire TIMEBOOST_net_2815;
wire n_19661;
wire n_19663;
wire n_19664;
wire n_19665;
wire n_19666;
wire TIMEBOOST_net_163;
wire n_19669;
wire n_1967;
wire TIMEBOOST_net_162;
wire n_19672;
wire n_19673;
wire n_19676;
wire n_19677;
wire n_19678;
wire n_19679;
wire n_1968;
wire n_19680;
wire n_19681;
wire n_19682;
wire n_19685;
wire n_19686;
wire n_19687;
wire n_19688;
wire n_19689;
wire n_1969;
wire n_19690;
wire n_19691;
wire n_19692;
wire n_19693;
wire n_19694;
wire n_19695;
wire n_19696;
wire n_19698;
wire n_19700;
wire n_19701;
wire n_19703;
wire n_19704;
wire TIMEBOOST_net_2414;
wire TIMEBOOST_net_2653;
wire n_19707;
wire n_19708;
wire n_19709;
wire n_1971;
wire n_19710;
wire n_19711;
wire n_19712;
wire n_19713;
wire n_19714;
wire n_19715;
wire n_19716;
wire n_19718;
wire n_19719;
wire n_1972;
wire n_19720;
wire n_19721;
wire n_19722;
wire n_19724;
wire n_19725;
wire n_19726;
wire n_19728;
wire TIMEBOOST_net_900;
wire n_1973;
wire n_19730;
wire n_19731;
wire n_19732;
wire n_19733;
wire n_19735;
wire n_19736;
wire n_19737;
wire n_19738;
wire n_19739;
wire n_1974;
wire n_19740;
wire n_19741;
wire n_19742;
wire n_19743;
wire n_19744;
wire n_19745;
wire n_19746;
wire n_19747;
wire n_19748;
wire n_19749;
wire n_1975;
wire n_19750;
wire n_19751;
wire n_19752;
wire n_19753;
wire n_19754;
wire n_19755;
wire n_19758;
wire n_1976;
wire n_19760;
wire n_19761;
wire n_19762;
wire n_19763;
wire n_19764;
wire n_19765;
wire n_19766;
wire n_19767;
wire n_19768;
wire n_19769;
wire n_1977;
wire n_19770;
wire n_19771;
wire n_19772;
wire n_19773;
wire n_19774;
wire n_19775;
wire n_19776;
wire n_19778;
wire n_19779;
wire n_1978;
wire n_19783;
wire n_19784;
wire n_19785;
wire n_19786;
wire n_19787;
wire n_19789;
wire n_1979;
wire n_19790;
wire n_19792;
wire n_19793;
wire n_19794;
wire n_19796;
wire n_19797;
wire n_19798;
wire n_19799;
wire n_198;
wire TIMEBOOST_net_2640;
wire n_19801;
wire n_19802;
wire n_19803;
wire n_19804;
wire n_19806;
wire n_19807;
wire n_19808;
wire n_19809;
wire n_1981;
wire n_19810;
wire n_19811;
wire n_19812;
wire n_19813;
wire n_19816;
wire n_19817;
wire n_19818;
wire n_19819;
wire n_1982;
wire n_19820;
wire n_19821;
wire n_19822;
wire n_19823;
wire n_19824;
wire n_19825;
wire n_19826;
wire n_19827;
wire n_19828;
wire n_19829;
wire n_1983;
wire n_19830;
wire n_19832;
wire n_19833;
wire n_19834;
wire n_19835;
wire n_19836;
wire n_19837;
wire n_19838;
wire n_19839;
wire n_1984;
wire n_19842;
wire TIMEBOOST_net_2385;
wire n_19844;
wire n_19845;
wire n_19846;
wire n_19847;
wire n_19848;
wire n_19849;
wire n_19850;
wire n_19851;
wire n_19852;
wire n_19853;
wire n_19854;
wire n_19855;
wire n_19856;
wire n_19859;
wire n_19860;
wire n_19861;
wire n_19862;
wire n_19863;
wire TIMEBOOST_net_253;
wire n_19866;
wire TIMEBOOST_net_2175;
wire n_19868;
wire n_1987;
wire n_19871;
wire n_19872;
wire n_19873;
wire n_19875;
wire n_19876;
wire n_19877;
wire n_19878;
wire n_19879;
wire n_1988;
wire n_19880;
wire n_19881;
wire n_19882;
wire n_19884;
wire n_19885;
wire n_19886;
wire n_19887;
wire n_19888;
wire n_19889;
wire n_19890;
wire n_19891;
wire n_19892;
wire n_19894;
wire n_19895;
wire n_19896;
wire n_19897;
wire n_19899;
wire n_199;
wire n_1990;
wire n_19900;
wire n_19901;
wire n_19902;
wire n_19903;
wire n_19904;
wire n_19905;
wire n_19906;
wire n_19907;
wire n_19909;
wire n_19910;
wire n_19911;
wire n_19912;
wire n_19913;
wire n_19914;
wire n_19915;
wire n_19919;
wire n_1992;
wire n_19920;
wire n_19921;
wire n_19922;
wire n_19924;
wire n_19926;
wire n_19927;
wire n_19928;
wire n_1993;
wire n_19930;
wire n_19931;
wire n_19932;
wire n_19933;
wire n_19934;
wire n_19935;
wire n_19936;
wire n_19938;
wire n_19939;
wire n_1994;
wire n_19940;
wire n_19941;
wire n_19942;
wire n_19943;
wire n_19944;
wire n_19945;
wire n_19946;
wire n_19948;
wire n_19949;
wire n_19950;
wire n_19952;
wire n_19953;
wire n_19954;
wire n_19956;
wire n_19957;
wire n_19958;
wire n_19959;
wire n_1996;
wire n_19960;
wire n_19961;
wire n_19962;
wire n_19963;
wire n_19964;
wire n_19965;
wire n_19967;
wire n_19968;
wire n_19969;
wire n_1997;
wire n_19970;
wire n_19972;
wire n_19973;
wire TIMEBOOST_net_2470;
wire n_19975;
wire n_19976;
wire n_19977;
wire n_19978;
wire n_19979;
wire n_1998;
wire n_19980;
wire n_19981;
wire n_19982;
wire n_19983;
wire n_19984;
wire n_19985;
wire n_19986;
wire n_19988;
wire n_19989;
wire n_1999;
wire n_19990;
wire n_19991;
wire n_19992;
wire n_19993;
wire n_19994;
wire n_19997;
wire n_19998;
wire n_19999;
wire n_200;
wire n_20000;
wire n_20001;
wire n_20002;
wire n_20003;
wire n_20004;
wire n_20005;
wire n_20006;
wire n_20007;
wire n_20009;
wire n_2001;
wire n_20010;
wire n_20011;
wire n_20012;
wire n_20013;
wire n_20014;
wire n_20015;
wire n_20016;
wire n_20017;
wire n_20018;
wire n_2002;
wire n_20020;
wire n_20021;
wire n_20022;
wire TIMEBOOST_net_2226;
wire n_20024;
wire n_20026;
wire TIMEBOOST_net_2242;
wire n_20028;
wire n_20029;
wire n_2003;
wire n_20030;
wire n_20031;
wire n_20032;
wire n_20033;
wire n_20034;
wire n_20036;
wire n_20037;
wire TIMEBOOST_net_999;
wire n_20039;
wire n_2004;
wire n_20040;
wire n_20041;
wire n_20042;
wire TIMEBOOST_net_1191;
wire n_20044;
wire n_20046;
wire n_20047;
wire n_20049;
wire n_2005;
wire n_20050;
wire n_20051;
wire n_20052;
wire n_20053;
wire n_20054;
wire n_20055;
wire TIMEBOOST_net_417;
wire n_20057;
wire n_20058;
wire n_20059;
wire n_2006;
wire n_20062;
wire TIMEBOOST_net_1065;
wire n_20064;
wire n_20065;
wire n_20068;
wire n_20069;
wire n_2007;
wire n_20070;
wire n_20072;
wire n_20073;
wire n_20074;
wire n_20075;
wire n_20076;
wire n_20078;
wire n_20079;
wire n_2008;
wire TIMEBOOST_net_2895;
wire n_20081;
wire n_20082;
wire n_20083;
wire n_20084;
wire n_20085;
wire n_20086;
wire n_20087;
wire n_20088;
wire n_20089;
wire n_2009;
wire n_20090;
wire n_20091;
wire n_20092;
wire n_20093;
wire n_20094;
wire n_20095;
wire n_20096;
wire n_20098;
wire n_2010;
wire TIMEBOOST_net_1597;
wire n_20103;
wire n_20104;
wire n_20105;
wire n_20106;
wire n_20107;
wire n_2011;
wire n_20112;
wire n_20113;
wire n_20114;
wire n_20115;
wire n_20116;
wire n_20117;
wire n_20118;
wire n_20119;
wire n_2012;
wire n_20120;
wire n_20121;
wire n_20122;
wire n_20123;
wire n_20124;
wire n_20125;
wire TIMEBOOST_net_438;
wire n_20127;
wire n_20129;
wire n_2013;
wire n_20133;
wire n_20134;
wire n_20135;
wire n_20136;
wire n_20137;
wire TIMEBOOST_net_2754;
wire n_2014;
wire n_20144;
wire n_20145;
wire n_20146;
wire n_20147;
wire n_20148;
wire n_20149;
wire n_2015;
wire n_20150;
wire n_20151;
wire n_20153;
wire TIMEBOOST_net_1239;
wire n_20155;
wire n_20156;
wire n_20157;
wire n_20160;
wire n_20161;
wire n_20162;
wire n_20163;
wire n_20164;
wire n_20165;
wire n_20167;
wire n_20168;
wire n_20169;
wire n_2017;
wire n_20170;
wire n_20171;
wire n_20172;
wire n_20174;
wire n_20176;
wire n_20177;
wire n_20178;
wire n_20179;
wire n_2018;
wire n_20180;
wire n_20181;
wire n_20182;
wire n_20183;
wire n_20184;
wire n_20186;
wire n_20187;
wire n_20188;
wire n_20189;
wire n_2019;
wire n_20190;
wire n_20191;
wire n_20192;
wire TIMEBOOST_net_474;
wire n_20194;
wire n_20195;
wire n_20196;
wire n_20197;
wire n_20198;
wire n_20199;
wire n_202;
wire n_2020;
wire n_20200;
wire n_20201;
wire n_20202;
wire n_20203;
wire n_20204;
wire n_20205;
wire n_20206;
wire n_20207;
wire n_20208;
wire n_20209;
wire n_2021;
wire n_20211;
wire n_20212;
wire n_20213;
wire n_20214;
wire n_20215;
wire n_20218;
wire n_20219;
wire n_20220;
wire n_20222;
wire n_20224;
wire TIMEBOOST_net_442;
wire n_20226;
wire n_20227;
wire n_20228;
wire n_20229;
wire n_2023;
wire n_20231;
wire n_20234;
wire n_20236;
wire n_20238;
wire n_20239;
wire n_2024;
wire n_20240;
wire n_20241;
wire n_20242;
wire n_20243;
wire n_20244;
wire n_20245;
wire n_20249;
wire n_2025;
wire n_20250;
wire n_20251;
wire n_20252;
wire n_20254;
wire n_20255;
wire n_20256;
wire n_20257;
wire n_2026;
wire n_20261;
wire n_20262;
wire n_20264;
wire n_20265;
wire n_20266;
wire n_20267;
wire n_20269;
wire n_2027;
wire n_20270;
wire n_20271;
wire n_20272;
wire n_20273;
wire n_20275;
wire n_20277;
wire n_20279;
wire n_2028;
wire n_20280;
wire n_20281;
wire n_20282;
wire n_20285;
wire n_20286;
wire n_20288;
wire n_20289;
wire n_2029;
wire n_20290;
wire n_20291;
wire TIMEBOOST_net_2645;
wire n_20293;
wire n_20294;
wire n_20297;
wire TIMEBOOST_net_486;
wire n_20299;
wire n_203;
wire n_2030;
wire n_20301;
wire n_20302;
wire n_20303;
wire n_20304;
wire n_20305;
wire n_20307;
wire n_20309;
wire n_2031;
wire n_20310;
wire n_20311;
wire n_20312;
wire n_20313;
wire n_20314;
wire TIMEBOOST_net_443;
wire n_20317;
wire TIMEBOOST_net_2561;
wire n_2032;
wire n_20320;
wire n_20321;
wire n_20325;
wire n_20327;
wire n_20328;
wire n_20329;
wire n_2033;
wire n_20330;
wire n_20332;
wire n_20333;
wire n_20334;
wire n_20336;
wire n_20337;
wire n_20338;
wire n_2034;
wire n_20340;
wire n_20341;
wire n_20342;
wire n_20343;
wire n_20344;
wire n_20345;
wire n_20348;
wire n_20349;
wire n_2035;
wire n_20353;
wire n_20354;
wire n_20355;
wire n_20356;
wire n_20357;
wire n_20363;
wire n_20366;
wire n_20369;
wire n_20370;
wire n_20371;
wire n_20372;
wire TIMEBOOST_net_453;
wire n_20374;
wire n_20375;
wire n_20376;
wire n_20378;
wire n_20379;
wire n_2038;
wire TIMEBOOST_net_449;
wire n_20383;
wire n_20384;
wire n_20385;
wire n_20386;
wire n_20391;
wire n_20395;
wire n_20396;
wire n_20399;
wire n_204;
wire n_2040;
wire n_20400;
wire n_20404;
wire TIMEBOOST_net_455;
wire n_20406;
wire n_20409;
wire n_2041;
wire n_20412;
wire n_20413;
wire n_20414;
wire n_20415;
wire TIMEBOOST_net_1681;
wire n_20417;
wire n_20418;
wire n_2042;
wire n_20420;
wire TIMEBOOST_net_487;
wire n_20422;
wire n_20423;
wire n_20424;
wire n_20425;
wire n_20426;
wire n_20429;
wire n_2043;
wire n_20430;
wire n_20432;
wire n_20433;
wire n_20434;
wire n_20435;
wire TIMEBOOST_net_2873;
wire n_20439;
wire n_2044;
wire n_20441;
wire n_20442;
wire n_20445;
wire n_20446;
wire n_20447;
wire n_20450;
wire n_20451;
wire n_20456;
wire n_20459;
wire n_2046;
wire n_20460;
wire n_20461;
wire n_20462;
wire n_20463;
wire n_20464;
wire n_20465;
wire n_20466;
wire n_20468;
wire n_20469;
wire n_2047;
wire n_20470;
wire n_20472;
wire n_20473;
wire n_20474;
wire n_20476;
wire n_20477;
wire n_20481;
wire n_20482;
wire n_20485;
wire n_20489;
wire n_2049;
wire n_20491;
wire n_20492;
wire n_20495;
wire n_20499;
wire n_205;
wire n_2050;
wire n_20500;
wire n_20501;
wire n_20502;
wire n_20504;
wire n_20505;
wire n_20506;
wire n_20508;
wire n_2051;
wire n_20510;
wire TIMEBOOST_net_506;
wire n_20512;
wire n_20513;
wire n_20514;
wire n_20515;
wire n_20516;
wire n_20517;
wire n_20518;
wire n_20519;
wire n_2052;
wire n_20523;
wire n_20526;
wire n_20528;
wire n_20529;
wire n_2053;
wire n_20531;
wire n_20532;
wire n_20533;
wire n_20534;
wire n_20535;
wire n_20536;
wire n_20539;
wire n_2054;
wire n_20540;
wire n_20542;
wire n_20545;
wire n_20548;
wire n_20549;
wire n_2055;
wire n_20552;
wire n_20553;
wire n_20555;
wire n_20558;
wire n_20559;
wire n_2056;
wire n_20560;
wire n_20565;
wire n_20567;
wire n_20568;
wire n_2057;
wire n_20570;
wire n_20573;
wire n_20575;
wire TIMEBOOST_net_1592;
wire n_20578;
wire n_20579;
wire TIMEBOOST_net_2189;
wire n_20582;
wire n_20583;
wire n_20587;
wire n_2059;
wire n_20591;
wire n_20594;
wire n_20595;
wire n_20596;
wire n_20597;
wire n_20598;
wire n_20599;
wire n_206;
wire n_20600;
wire n_20603;
wire TIMEBOOST_net_2870;
wire n_20605;
wire n_20606;
wire n_20607;
wire n_20608;
wire n_2061;
wire n_20611;
wire n_20612;
wire n_20614;
wire n_20615;
wire n_20616;
wire TIMEBOOST_net_484;
wire n_20618;
wire n_20619;
wire n_2062;
wire n_20620;
wire n_20621;
wire n_20624;
wire n_20626;
wire n_20628;
wire n_2063;
wire n_20630;
wire TIMEBOOST_net_1135;
wire n_20632;
wire n_20634;
wire n_20635;
wire n_20636;
wire n_20637;
wire n_20638;
wire n_2064;
wire n_20640;
wire n_20641;
wire n_20642;
wire TIMEBOOST_net_2927;
wire n_20647;
wire n_20648;
wire n_2065;
wire n_20650;
wire n_20651;
wire n_20652;
wire n_20653;
wire n_20654;
wire n_20655;
wire n_20657;
wire n_20658;
wire n_20659;
wire n_2066;
wire n_20660;
wire n_20661;
wire TIMEBOOST_net_1224;
wire n_20664;
wire n_20665;
wire n_20666;
wire n_20667;
wire n_20669;
wire n_2067;
wire n_20670;
wire n_20671;
wire n_20672;
wire n_20673;
wire n_20674;
wire n_20675;
wire n_20676;
wire n_20677;
wire n_20678;
wire n_2068;
wire n_20682;
wire n_20683;
wire n_20684;
wire TIMEBOOST_net_1910;
wire n_20687;
wire n_2069;
wire n_20690;
wire n_20691;
wire n_20693;
wire n_20694;
wire TIMEBOOST_net_2771;
wire n_20696;
wire n_20699;
wire n_207;
wire n_2070;
wire n_20700;
wire n_20701;
wire n_20702;
wire n_20703;
wire n_20704;
wire n_20705;
wire n_20708;
wire n_20709;
wire n_2071;
wire n_20710;
wire n_20712;
wire n_20713;
wire n_20714;
wire n_20715;
wire n_20716;
wire n_20717;
wire n_20719;
wire n_20721;
wire n_20722;
wire n_20723;
wire n_20724;
wire TIMEBOOST_net_1208;
wire n_20727;
wire TIMEBOOST_net_2933;
wire n_2073;
wire n_20730;
wire n_20731;
wire n_20732;
wire n_20733;
wire n_20734;
wire n_20735;
wire n_20736;
wire n_20739;
wire n_2074;
wire n_20740;
wire n_20741;
wire n_20742;
wire n_20743;
wire n_20744;
wire n_20745;
wire TIMEBOOST_net_1223;
wire n_20749;
wire n_2075;
wire n_20750;
wire n_20751;
wire n_20752;
wire n_20753;
wire n_20754;
wire n_20755;
wire n_20756;
wire n_20757;
wire n_20759;
wire n_2076;
wire n_20760;
wire n_20761;
wire n_20763;
wire n_20764;
wire n_20767;
wire TIMEBOOST_net_490;
wire n_2077;
wire n_20771;
wire n_20774;
wire n_20775;
wire TIMEBOOST_net_524;
wire n_20777;
wire n_20778;
wire n_20781;
wire n_20782;
wire n_20783;
wire n_20784;
wire n_20785;
wire n_20786;
wire n_20787;
wire TIMEBOOST_net_1727;
wire n_20790;
wire n_20791;
wire n_20793;
wire TIMEBOOST_net_2463;
wire n_20795;
wire TIMEBOOST_net_2915;
wire n_20797;
wire n_20798;
wire n_20799;
wire n_208;
wire TIMEBOOST_net_2935;
wire n_20802;
wire n_20803;
wire n_20804;
wire n_20805;
wire TIMEBOOST_net_1247;
wire n_20809;
wire n_2081;
wire n_20810;
wire n_20811;
wire n_20812;
wire n_20815;
wire TIMEBOOST_net_491;
wire TIMEBOOST_net_2724;
wire n_20819;
wire n_2082;
wire n_20820;
wire n_20821;
wire n_20822;
wire n_20823;
wire n_20825;
wire n_20828;
wire n_20829;
wire n_2083;
wire n_20830;
wire n_20831;
wire n_20834;
wire n_20835;
wire n_20836;
wire n_20837;
wire n_20838;
wire n_2084;
wire n_20841;
wire n_20842;
wire n_20843;
wire n_20846;
wire n_20847;
wire n_20848;
wire n_20849;
wire n_2085;
wire n_20850;
wire TIMEBOOST_net_1901;
wire n_20852;
wire n_20853;
wire n_20854;
wire n_20855;
wire n_20856;
wire n_20857;
wire n_20859;
wire n_2086;
wire n_20861;
wire n_20862;
wire n_20865;
wire n_20866;
wire n_20867;
wire n_20868;
wire n_2087;
wire n_20871;
wire n_20872;
wire n_20873;
wire n_20874;
wire n_20875;
wire n_20876;
wire n_20877;
wire n_20878;
wire n_20879;
wire n_2088;
wire n_20881;
wire n_20882;
wire n_20883;
wire n_20884;
wire n_20885;
wire n_20886;
wire n_20889;
wire n_2089;
wire n_20891;
wire n_20894;
wire n_20895;
wire n_20896;
wire n_20897;
wire n_20898;
wire n_20899;
wire n_209;
wire n_2090;
wire n_20900;
wire n_20901;
wire n_20902;
wire n_20903;
wire n_20904;
wire n_20905;
wire TIMEBOOST_net_1694;
wire n_20907;
wire n_20908;
wire n_2091;
wire n_20910;
wire n_20912;
wire n_20913;
wire n_20914;
wire n_20915;
wire n_20916;
wire n_20917;
wire n_20918;
wire n_20919;
wire n_2092;
wire n_20920;
wire n_20922;
wire n_20924;
wire n_20925;
wire n_20926;
wire n_20927;
wire n_20928;
wire n_20929;
wire n_2093;
wire n_20930;
wire n_20931;
wire n_20932;
wire n_20933;
wire n_20935;
wire n_20936;
wire n_20939;
wire n_2094;
wire n_20941;
wire n_20942;
wire n_20943;
wire n_20944;
wire n_20945;
wire n_20947;
wire n_20948;
wire n_20949;
wire n_2095;
wire n_20950;
wire n_20951;
wire n_20953;
wire n_20954;
wire n_20956;
wire n_20957;
wire n_20958;
wire n_2096;
wire n_20960;
wire n_20961;
wire n_20962;
wire n_20963;
wire n_20966;
wire n_20967;
wire n_20968;
wire n_2097;
wire n_20970;
wire TIMEBOOST_net_504;
wire n_20973;
wire TIMEBOOST_net_1977;
wire n_20976;
wire n_20977;
wire n_20978;
wire n_20979;
wire n_20980;
wire n_20981;
wire n_20982;
wire n_20983;
wire n_20984;
wire n_20985;
wire n_20987;
wire n_20988;
wire n_20989;
wire n_20991;
wire n_20993;
wire n_20995;
wire n_20997;
wire n_20999;
wire n_210;
wire n_2100;
wire n_21000;
wire n_21001;
wire n_21002;
wire n_21003;
wire n_21004;
wire n_21006;
wire n_21007;
wire n_2101;
wire n_21011;
wire n_21012;
wire n_21013;
wire n_21014;
wire n_21015;
wire n_21016;
wire n_21018;
wire n_21019;
wire n_2102;
wire n_21020;
wire n_21021;
wire n_21022;
wire n_21023;
wire n_21024;
wire n_21027;
wire n_21028;
wire n_21029;
wire n_2103;
wire n_21034;
wire n_21035;
wire n_21036;
wire n_21037;
wire n_21039;
wire n_2104;
wire n_21040;
wire n_21041;
wire n_21042;
wire n_21043;
wire n_21044;
wire n_21045;
wire n_21046;
wire TIMEBOOST_net_1275;
wire n_2105;
wire n_21050;
wire n_21051;
wire n_21052;
wire n_21053;
wire n_21054;
wire n_21055;
wire n_21056;
wire n_21058;
wire n_21059;
wire n_2106;
wire n_21061;
wire n_21062;
wire n_21063;
wire n_21064;
wire n_21065;
wire n_21066;
wire n_21067;
wire n_21068;
wire n_21069;
wire TIMEBOOST_net_954;
wire TIMEBOOST_net_510;
wire n_21071;
wire n_21072;
wire n_21074;
wire n_21075;
wire n_21076;
wire n_21077;
wire n_21078;
wire n_2108;
wire n_21080;
wire TIMEBOOST_net_2021;
wire n_21084;
wire n_21087;
wire n_21088;
wire n_21089;
wire n_2109;
wire n_21090;
wire n_21091;
wire n_21092;
wire n_21093;
wire n_21094;
wire n_21095;
wire n_21096;
wire n_21098;
wire n_21099;
wire n_211;
wire n_2110;
wire n_21100;
wire n_21101;
wire n_21102;
wire n_21103;
wire n_21104;
wire n_21105;
wire n_21106;
wire n_21107;
wire n_21108;
wire n_21109;
wire n_2111;
wire n_21110;
wire n_21111;
wire n_21114;
wire n_21115;
wire n_21116;
wire n_21118;
wire n_21119;
wire n_2112;
wire n_21120;
wire n_21121;
wire n_21124;
wire n_21125;
wire n_21127;
wire n_2113;
wire n_21130;
wire n_21131;
wire n_21132;
wire n_21133;
wire n_21134;
wire n_21136;
wire n_21137;
wire n_21138;
wire n_21139;
wire n_2114;
wire n_21140;
wire n_21141;
wire n_21142;
wire n_21143;
wire n_21144;
wire n_21147;
wire n_21148;
wire n_21149;
wire n_2115;
wire n_21150;
wire n_21153;
wire n_21154;
wire TIMEBOOST_net_1320;
wire n_21157;
wire n_21159;
wire n_2116;
wire n_21160;
wire n_21163;
wire n_21164;
wire n_21165;
wire n_21166;
wire n_21169;
wire n_2117;
wire n_21171;
wire n_21172;
wire n_21173;
wire n_21174;
wire n_21175;
wire TIMEBOOST_net_2059;
wire n_21177;
wire n_21178;
wire n_2118;
wire TIMEBOOST_net_542;
wire n_21183;
wire n_21184;
wire n_21185;
wire n_21186;
wire n_21187;
wire n_21188;
wire n_2119;
wire n_21192;
wire n_21194;
wire n_21195;
wire n_21196;
wire n_21197;
wire n_21198;
wire n_21199;
wire n_212;
wire n_2120;
wire n_21200;
wire n_21202;
wire n_21203;
wire n_21205;
wire n_21206;
wire n_21207;
wire n_21208;
wire n_2121;
wire n_21212;
wire n_21214;
wire n_21218;
wire n_21219;
wire n_21220;
wire n_21224;
wire n_21227;
wire n_21229;
wire n_2123;
wire n_21230;
wire n_21232;
wire n_21233;
wire n_21236;
wire n_21237;
wire n_21238;
wire n_2124;
wire n_21240;
wire n_21242;
wire n_21244;
wire n_21246;
wire n_21247;
wire n_21248;
wire n_21249;
wire n_2125;
wire n_21251;
wire n_21252;
wire n_21253;
wire n_21254;
wire n_21255;
wire n_21256;
wire n_21257;
wire n_21258;
wire n_21259;
wire n_2126;
wire n_21260;
wire n_21261;
wire n_21263;
wire n_21264;
wire n_21265;
wire n_21266;
wire n_21268;
wire n_21269;
wire n_2127;
wire n_21271;
wire n_21272;
wire n_21273;
wire n_21276;
wire n_21277;
wire n_21278;
wire n_21279;
wire n_2128;
wire n_21280;
wire n_21281;
wire n_21282;
wire n_21283;
wire n_21285;
wire n_21286;
wire n_21287;
wire n_21288;
wire n_21289;
wire n_2129;
wire n_21291;
wire n_21292;
wire n_21294;
wire n_21295;
wire n_21296;
wire n_21297;
wire n_21298;
wire n_21299;
wire n_213;
wire n_2130;
wire n_21300;
wire n_21301;
wire n_21302;
wire n_21305;
wire n_21306;
wire n_21307;
wire TIMEBOOST_net_1265;
wire n_2131;
wire n_21312;
wire n_21316;
wire n_21317;
wire n_21318;
wire n_2132;
wire n_21322;
wire n_21323;
wire n_21324;
wire n_21326;
wire n_21327;
wire TIMEBOOST_net_2249;
wire n_21329;
wire n_2133;
wire n_21330;
wire n_21331;
wire n_21332;
wire n_21334;
wire n_21335;
wire n_21336;
wire n_21337;
wire n_21338;
wire n_2134;
wire n_21341;
wire n_21342;
wire n_21343;
wire n_21344;
wire n_21345;
wire n_21346;
wire n_21348;
wire n_2135;
wire n_21350;
wire n_21351;
wire n_21353;
wire n_21354;
wire n_21355;
wire n_21356;
wire n_21358;
wire n_21360;
wire n_21361;
wire n_21363;
wire n_21365;
wire n_21366;
wire n_2137;
wire n_21370;
wire n_21371;
wire n_21373;
wire n_21374;
wire n_21375;
wire n_21376;
wire n_21377;
wire n_21378;
wire n_21379;
wire n_21380;
wire n_21381;
wire n_21382;
wire n_21384;
wire n_21385;
wire n_21386;
wire n_21387;
wire TIMEBOOST_net_525;
wire TIMEBOOST_net_2736;
wire n_21390;
wire n_21391;
wire n_21392;
wire n_21393;
wire n_21394;
wire TIMEBOOST_net_2000;
wire n_21397;
wire n_21398;
wire n_21399;
wire n_214;
wire n_2140;
wire n_21402;
wire n_21403;
wire n_21404;
wire n_21405;
wire n_21406;
wire n_21407;
wire n_21408;
wire n_21409;
wire n_2141;
wire n_21410;
wire n_21413;
wire n_21415;
wire n_21416;
wire n_21417;
wire n_21419;
wire n_2142;
wire n_21420;
wire n_21421;
wire n_21422;
wire TIMEBOOST_net_2016;
wire n_21424;
wire n_21425;
wire n_21426;
wire n_21427;
wire n_21428;
wire n_21429;
wire n_2143;
wire n_21430;
wire n_21431;
wire n_21432;
wire n_21433;
wire n_21434;
wire n_21435;
wire TIMEBOOST_net_2694;
wire n_21438;
wire n_2144;
wire TIMEBOOST_net_1324;
wire n_21442;
wire n_21446;
wire n_21447;
wire n_21448;
wire n_21449;
wire n_2145;
wire n_21450;
wire n_21451;
wire n_21452;
wire n_21453;
wire n_21454;
wire n_21455;
wire n_21456;
wire n_21458;
wire n_21459;
wire n_2146;
wire n_21461;
wire n_21462;
wire n_21463;
wire n_21464;
wire n_21466;
wire n_21467;
wire n_2147;
wire n_21470;
wire n_21471;
wire n_21472;
wire n_21473;
wire n_21474;
wire n_21475;
wire n_21476;
wire n_21477;
wire n_21478;
wire n_21479;
wire n_2148;
wire n_21480;
wire n_21481;
wire n_21482;
wire n_21483;
wire n_21484;
wire n_21485;
wire n_21486;
wire n_21487;
wire n_21488;
wire n_21489;
wire n_2149;
wire n_21490;
wire n_21491;
wire n_21492;
wire n_21493;
wire n_21494;
wire n_21495;
wire n_21496;
wire n_21497;
wire n_215;
wire n_21500;
wire n_21501;
wire n_21502;
wire n_21503;
wire n_21504;
wire n_21505;
wire n_21506;
wire n_21507;
wire n_21508;
wire n_21509;
wire n_2151;
wire n_21510;
wire n_21511;
wire n_21514;
wire n_21516;
wire n_21517;
wire n_21518;
wire n_21519;
wire n_2152;
wire n_21520;
wire n_21521;
wire n_21526;
wire n_21527;
wire n_21528;
wire n_21529;
wire n_2153;
wire n_21530;
wire n_21531;
wire n_21533;
wire n_21535;
wire n_21537;
wire n_21538;
wire n_21539;
wire n_2154;
wire n_21540;
wire n_21541;
wire n_21543;
wire n_21544;
wire n_21545;
wire n_21546;
wire n_21547;
wire n_21548;
wire n_2155;
wire n_21552;
wire n_21553;
wire n_21554;
wire n_21556;
wire n_21558;
wire n_2156;
wire n_21560;
wire n_21561;
wire n_21562;
wire n_21563;
wire n_21564;
wire n_21565;
wire n_21566;
wire n_21569;
wire n_2157;
wire n_21571;
wire n_21572;
wire n_21573;
wire n_21574;
wire n_21575;
wire n_21576;
wire n_21578;
wire n_21579;
wire n_2158;
wire n_21580;
wire n_21581;
wire n_21586;
wire n_21587;
wire n_21588;
wire TIMEBOOST_net_959;
wire n_21591;
wire n_21592;
wire n_21593;
wire n_21595;
wire n_21597;
wire n_21598;
wire n_21599;
wire TIMEBOOST_net_36;
wire n_2160;
wire n_21600;
wire n_21601;
wire n_21602;
wire n_21603;
wire n_21604;
wire n_21605;
wire n_21606;
wire n_21609;
wire n_2161;
wire TIMEBOOST_net_1330;
wire n_21611;
wire n_21612;
wire n_21613;
wire n_21615;
wire n_21616;
wire n_21617;
wire n_21618;
wire n_21619;
wire n_21620;
wire n_21621;
wire n_21622;
wire n_21624;
wire n_21625;
wire n_21626;
wire n_21627;
wire n_21628;
wire n_21629;
wire n_2163;
wire n_21630;
wire n_21632;
wire n_21633;
wire n_21634;
wire n_21636;
wire TIMEBOOST_net_2049;
wire n_21639;
wire n_2164;
wire n_21640;
wire n_21641;
wire n_21642;
wire n_21643;
wire n_21644;
wire n_21645;
wire n_21646;
wire n_21647;
wire n_21648;
wire n_2165;
wire n_21654;
wire n_21656;
wire n_21658;
wire n_21659;
wire n_2166;
wire n_21660;
wire n_21661;
wire n_21662;
wire n_21663;
wire n_21664;
wire n_21665;
wire TIMEBOOST_net_2860;
wire n_21668;
wire n_21669;
wire n_2167;
wire n_21670;
wire n_21671;
wire n_21672;
wire TIMEBOOST_net_1403;
wire n_21676;
wire n_21677;
wire n_21678;
wire n_21679;
wire n_21680;
wire n_21682;
wire n_21683;
wire n_21684;
wire n_21685;
wire n_21686;
wire n_21687;
wire n_2169;
wire n_21691;
wire n_21692;
wire n_21693;
wire n_21694;
wire n_21695;
wire n_21696;
wire n_21697;
wire n_21698;
wire n_21699;
wire n_217;
wire n_2170;
wire n_21700;
wire n_21701;
wire n_21702;
wire n_21703;
wire TIMEBOOST_net_599;
wire n_21705;
wire n_21706;
wire n_21707;
wire n_21708;
wire n_21709;
wire n_2171;
wire n_21710;
wire n_21711;
wire TIMEBOOST_net_548;
wire n_21713;
wire n_21714;
wire n_21715;
wire n_21716;
wire n_21718;
wire n_21719;
wire n_2172;
wire n_21720;
wire n_21721;
wire n_21722;
wire n_21723;
wire n_21724;
wire n_21725;
wire n_21726;
wire n_21727;
wire n_21728;
wire n_2173;
wire n_21730;
wire n_21731;
wire n_21732;
wire n_21733;
wire n_21734;
wire n_21735;
wire n_21736;
wire n_21738;
wire n_2174;
wire n_21741;
wire n_21742;
wire n_21743;
wire n_21745;
wire n_21748;
wire n_21749;
wire n_2175;
wire n_21750;
wire n_21751;
wire n_21752;
wire n_21753;
wire n_21754;
wire n_21755;
wire n_21756;
wire n_21757;
wire n_21758;
wire n_21759;
wire n_2176;
wire n_21760;
wire n_21761;
wire n_21762;
wire n_21763;
wire n_21764;
wire TIMEBOOST_net_1332;
wire n_21766;
wire n_21767;
wire n_21768;
wire TIMEBOOST_net_2297;
wire n_2177;
wire n_21772;
wire n_21773;
wire n_21774;
wire n_21775;
wire n_21776;
wire n_21777;
wire n_21778;
wire n_21779;
wire n_2178;
wire n_21780;
wire n_21781;
wire n_21782;
wire n_21783;
wire n_21784;
wire n_21785;
wire n_21786;
wire TIMEBOOST_net_2051;
wire n_21788;
wire n_21789;
wire n_2179;
wire n_21790;
wire n_21791;
wire n_21792;
wire n_21793;
wire n_21794;
wire n_21795;
wire n_21796;
wire n_21797;
wire n_21798;
wire n_21799;
wire n_218;
wire n_2180;
wire n_21800;
wire n_21801;
wire n_21802;
wire n_21803;
wire n_21804;
wire n_21807;
wire n_21808;
wire TIMEBOOST_net_1501;
wire n_2181;
wire n_21810;
wire n_21811;
wire n_21812;
wire n_21813;
wire n_21814;
wire n_21815;
wire n_21816;
wire n_21817;
wire n_21818;
wire n_21819;
wire n_2182;
wire n_21821;
wire n_21822;
wire n_21824;
wire n_21825;
wire n_21826;
wire n_21827;
wire n_21828;
wire n_2183;
wire n_21831;
wire n_21832;
wire n_21833;
wire n_21834;
wire n_21835;
wire n_21836;
wire n_21837;
wire n_21838;
wire n_21839;
wire n_2184;
wire n_21842;
wire n_21843;
wire n_21844;
wire n_21845;
wire n_21847;
wire n_21849;
wire n_2185;
wire n_21851;
wire n_21852;
wire n_21853;
wire n_21854;
wire n_21855;
wire n_21856;
wire n_21857;
wire n_21858;
wire n_21859;
wire n_2186;
wire n_21860;
wire n_21861;
wire n_21862;
wire n_21863;
wire n_21864;
wire n_21865;
wire n_21866;
wire n_21867;
wire n_21868;
wire n_21869;
wire n_2187;
wire n_21870;
wire n_21871;
wire TIMEBOOST_net_608;
wire n_21873;
wire n_21874;
wire n_21875;
wire n_21877;
wire n_21878;
wire n_21879;
wire n_2188;
wire n_21880;
wire n_21881;
wire n_21882;
wire n_21883;
wire n_21884;
wire n_21885;
wire n_21886;
wire n_21887;
wire n_21888;
wire n_21889;
wire n_2189;
wire n_21890;
wire n_21891;
wire n_21892;
wire n_21893;
wire n_21894;
wire n_21895;
wire n_21896;
wire n_21897;
wire n_21898;
wire n_219;
wire n_2190;
wire n_21900;
wire n_21902;
wire n_21903;
wire n_21904;
wire n_21905;
wire n_21906;
wire n_21909;
wire n_2191;
wire n_21910;
wire n_21911;
wire n_21912;
wire n_21913;
wire n_21914;
wire n_21915;
wire n_21916;
wire n_21917;
wire n_21918;
wire n_21919;
wire n_2192;
wire n_21920;
wire n_21921;
wire n_21922;
wire n_21923;
wire n_21924;
wire n_21925;
wire n_21927;
wire n_21929;
wire n_2193;
wire n_21930;
wire n_21931;
wire n_21932;
wire n_21933;
wire n_21936;
wire n_21937;
wire n_21938;
wire n_21939;
wire n_2194;
wire n_21940;
wire n_21941;
wire n_21944;
wire n_21945;
wire n_21946;
wire n_21947;
wire n_2195;
wire n_21950;
wire n_21951;
wire n_21953;
wire n_21954;
wire n_21956;
wire n_21957;
wire n_21958;
wire n_21959;
wire n_2196;
wire n_21960;
wire n_21961;
wire n_21962;
wire n_21963;
wire n_21964;
wire n_21965;
wire n_21966;
wire n_21967;
wire n_21969;
wire n_2197;
wire n_21970;
wire n_21971;
wire n_21972;
wire n_21973;
wire n_21974;
wire n_21975;
wire n_21977;
wire n_21978;
wire n_2198;
wire TIMEBOOST_net_1526;
wire n_21982;
wire n_21983;
wire n_21984;
wire n_21985;
wire n_21987;
wire n_2199;
wire n_21990;
wire n_21994;
wire n_21995;
wire n_21996;
wire n_21997;
wire n_21998;
wire n_21999;
wire n_220;
wire n_2200;
wire n_22002;
wire n_22003;
wire n_22005;
wire n_22008;
wire n_22009;
wire n_2201;
wire n_22010;
wire n_22011;
wire n_22012;
wire n_22014;
wire n_22015;
wire n_22016;
wire n_22018;
wire n_22019;
wire n_2202;
wire n_22020;
wire n_22021;
wire n_22022;
wire n_22027;
wire n_22028;
wire n_22030;
wire n_22031;
wire n_22032;
wire n_22033;
wire n_22034;
wire n_22035;
wire n_22037;
wire n_22038;
wire n_22039;
wire n_2204;
wire n_22041;
wire n_22043;
wire n_22044;
wire n_22045;
wire n_22046;
wire n_22047;
wire n_22048;
wire n_22049;
wire n_2205;
wire n_22052;
wire n_22053;
wire n_22054;
wire n_22055;
wire n_22056;
wire n_22057;
wire n_22058;
wire n_22059;
wire n_2206;
wire n_22060;
wire n_22061;
wire n_22062;
wire n_22063;
wire n_22064;
wire n_22065;
wire n_22066;
wire n_22068;
wire TIMEBOOST_net_1736;
wire n_22078;
wire n_22079;
wire n_2208;
wire n_22080;
wire n_22081;
wire n_22082;
wire n_22083;
wire n_22084;
wire n_22085;
wire n_22086;
wire n_22088;
wire n_22089;
wire n_2209;
wire n_22094;
wire n_22095;
wire n_22098;
wire n_22099;
wire n_221;
wire n_22106;
wire n_22107;
wire n_22108;
wire n_22109;
wire n_2211;
wire n_22110;
wire n_22111;
wire n_22112;
wire n_22113;
wire n_22115;
wire n_22116;
wire n_22117;
wire n_22118;
wire n_22119;
wire n_2212;
wire n_22121;
wire n_22126;
wire TIMEBOOST_net_631;
wire n_22128;
wire n_22129;
wire n_2213;
wire n_22130;
wire n_22131;
wire TIMEBOOST_net_716;
wire n_22134;
wire TIMEBOOST_net_1391;
wire n_22138;
wire n_22139;
wire n_2214;
wire n_22140;
wire n_22144;
wire n_22145;
wire n_22149;
wire n_2215;
wire n_22150;
wire n_22153;
wire n_22154;
wire n_22155;
wire n_22156;
wire n_2216;
wire n_22164;
wire n_22165;
wire n_22167;
wire n_22168;
wire n_22169;
wire n_2217;
wire n_22170;
wire n_22171;
wire n_22172;
wire n_22176;
wire n_22177;
wire n_22178;
wire n_22179;
wire n_2218;
wire n_22180;
wire n_22183;
wire n_22184;
wire n_22185;
wire n_22186;
wire n_22187;
wire n_2219;
wire n_22194;
wire n_22196;
wire TIMEBOOST_net_2316;
wire TIMEBOOST_net_629;
wire n_222;
wire n_22200;
wire n_22201;
wire n_22203;
wire n_22204;
wire n_22205;
wire n_22207;
wire n_22208;
wire n_22209;
wire n_2221;
wire n_22210;
wire n_22212;
wire n_22213;
wire n_22214;
wire n_22216;
wire TIMEBOOST_net_2524;
wire n_2222;
wire n_22220;
wire n_22221;
wire TIMEBOOST_net_630;
wire TIMEBOOST_net_2941;
wire TIMEBOOST_net_2058;
wire n_2223;
wire n_22230;
wire n_22231;
wire n_22232;
wire n_22233;
wire n_22234;
wire n_22235;
wire n_22236;
wire n_22237;
wire n_22238;
wire n_22239;
wire n_2224;
wire n_22242;
wire n_22243;
wire n_22244;
wire n_22245;
wire n_22246;
wire n_22247;
wire n_22248;
wire n_22249;
wire n_2225;
wire n_22253;
wire n_22258;
wire n_22259;
wire n_2226;
wire n_22261;
wire n_22262;
wire n_22263;
wire n_22264;
wire n_22266;
wire n_22267;
wire n_22268;
wire n_22269;
wire n_2227;
wire n_22270;
wire n_22271;
wire n_22272;
wire n_22273;
wire n_22275;
wire n_22279;
wire n_2228;
wire n_22280;
wire n_22284;
wire n_22285;
wire n_22286;
wire n_22287;
wire n_22288;
wire n_2229;
wire n_22291;
wire n_22292;
wire n_22293;
wire n_22294;
wire n_22295;
wire n_22296;
wire n_22299;
wire TIMEBOOST_net_1544;
wire n_2230;
wire n_22300;
wire n_22301;
wire n_22303;
wire n_22304;
wire n_22305;
wire n_22306;
wire n_22307;
wire n_22308;
wire n_22309;
wire n_2231;
wire n_22311;
wire n_22312;
wire n_22313;
wire n_22314;
wire n_22316;
wire n_22317;
wire n_22318;
wire n_22319;
wire n_2232;
wire n_22326;
wire n_22327;
wire n_22328;
wire n_2233;
wire n_22330;
wire n_22332;
wire n_22335;
wire n_22336;
wire n_22337;
wire n_22338;
wire n_22339;
wire n_2234;
wire n_22340;
wire n_22341;
wire n_22342;
wire n_22343;
wire n_22344;
wire n_22345;
wire n_22346;
wire n_22347;
wire n_22349;
wire n_22351;
wire n_22352;
wire TIMEBOOST_net_745;
wire n_22354;
wire n_22355;
wire n_22356;
wire n_22357;
wire n_22358;
wire n_22359;
wire n_22361;
wire n_22362;
wire n_22363;
wire TIMEBOOST_net_626;
wire n_22367;
wire n_22368;
wire n_2237;
wire n_22370;
wire TIMEBOOST_net_2737;
wire n_22374;
wire n_22375;
wire n_22377;
wire n_22378;
wire n_22379;
wire n_2238;
wire n_22380;
wire n_22381;
wire n_22382;
wire n_22383;
wire n_22385;
wire n_22386;
wire n_22387;
wire n_22388;
wire n_22389;
wire n_2239;
wire n_22390;
wire n_22391;
wire n_22392;
wire n_22393;
wire n_22395;
wire n_22396;
wire n_22397;
wire n_22398;
wire n_22399;
wire n_224;
wire n_2240;
wire n_22404;
wire n_22405;
wire n_22406;
wire n_22407;
wire n_2241;
wire TIMEBOOST_net_2320;
wire n_22411;
wire TIMEBOOST_net_2319;
wire n_22413;
wire n_22415;
wire n_22416;
wire n_22417;
wire n_22419;
wire n_22420;
wire n_22421;
wire n_22423;
wire n_22424;
wire n_22425;
wire n_22426;
wire n_22428;
wire n_2243;
wire n_22430;
wire n_22431;
wire n_22432;
wire n_22434;
wire TIMEBOOST_net_1339;
wire n_22436;
wire n_22438;
wire n_22439;
wire n_2244;
wire n_22443;
wire n_22444;
wire n_22445;
wire n_22446;
wire n_22447;
wire n_22448;
wire n_22449;
wire n_2245;
wire n_22450;
wire n_22453;
wire n_22455;
wire n_22456;
wire n_22457;
wire n_22458;
wire n_22459;
wire n_2246;
wire n_22460;
wire n_22461;
wire n_22462;
wire n_22463;
wire n_22464;
wire n_22465;
wire n_22466;
wire n_22468;
wire n_22469;
wire n_2247;
wire n_22470;
wire n_22472;
wire n_22473;
wire n_22474;
wire n_22475;
wire n_22476;
wire n_22479;
wire n_2248;
wire n_22480;
wire n_22481;
wire n_22482;
wire n_22483;
wire n_22484;
wire n_22485;
wire n_22486;
wire n_22487;
wire n_22488;
wire n_22489;
wire n_2249;
wire n_22490;
wire n_22491;
wire n_22492;
wire n_22493;
wire n_22494;
wire n_22495;
wire n_22496;
wire n_22497;
wire n_22498;
wire n_22499;
wire n_225;
wire n_2250;
wire n_22500;
wire n_22501;
wire n_22502;
wire n_22503;
wire n_22504;
wire n_22505;
wire n_22507;
wire n_22508;
wire n_2251;
wire n_22511;
wire n_22513;
wire n_22514;
wire n_22518;
wire n_2252;
wire n_22521;
wire n_22522;
wire n_22523;
wire n_22524;
wire n_22525;
wire n_22526;
wire n_22527;
wire n_22528;
wire n_2253;
wire n_22531;
wire n_22535;
wire n_22536;
wire n_22537;
wire n_22538;
wire TIMEBOOST_net_1435;
wire n_2254;
wire n_22540;
wire n_22542;
wire n_22543;
wire n_22544;
wire n_22545;
wire n_22548;
wire n_22549;
wire n_2255;
wire n_22550;
wire n_22553;
wire n_22554;
wire TIMEBOOST_net_769;
wire n_22556;
wire n_22558;
wire TIMEBOOST_net_789;
wire n_22560;
wire n_22562;
wire n_22564;
wire n_22566;
wire n_22567;
wire n_22568;
wire n_2257;
wire n_22570;
wire n_22573;
wire n_22574;
wire n_22575;
wire n_2258;
wire n_22580;
wire n_22581;
wire n_22584;
wire n_22585;
wire n_22586;
wire n_22587;
wire n_22588;
wire n_22589;
wire n_2259;
wire n_22591;
wire n_22593;
wire n_22594;
wire n_22596;
wire n_22597;
wire n_22598;
wire n_226;
wire n_2260;
wire n_22601;
wire TIMEBOOST_net_736;
wire n_22603;
wire n_22604;
wire n_22606;
wire n_22608;
wire n_2261;
wire n_22611;
wire n_22612;
wire n_22613;
wire n_22614;
wire n_22617;
wire n_22618;
wire n_22619;
wire n_22620;
wire n_22621;
wire n_22622;
wire n_22624;
wire n_22625;
wire n_22629;
wire n_2263;
wire n_22630;
wire n_22631;
wire n_22632;
wire n_22633;
wire n_22634;
wire n_22635;
wire n_22636;
wire n_22637;
wire n_22639;
wire n_2264;
wire n_22640;
wire n_22641;
wire n_22643;
wire n_22644;
wire n_22645;
wire n_22646;
wire n_22647;
wire n_22648;
wire n_22649;
wire n_2265;
wire n_22650;
wire n_22652;
wire n_22653;
wire n_22654;
wire n_22655;
wire n_22656;
wire n_22657;
wire n_22658;
wire n_22659;
wire n_2266;
wire n_22660;
wire n_22661;
wire n_22667;
wire n_22668;
wire n_22669;
wire TIMEBOOST_net_1870;
wire n_22670;
wire n_22671;
wire n_22672;
wire n_22673;
wire n_22674;
wire n_22675;
wire n_22676;
wire n_22677;
wire n_2268;
wire n_22682;
wire n_22684;
wire n_22685;
wire n_22686;
wire n_22687;
wire n_22688;
wire n_22689;
wire n_2269;
wire n_22690;
wire n_22692;
wire n_22693;
wire n_22694;
wire n_22695;
wire n_22697;
wire n_22698;
wire n_22699;
wire n_227;
wire n_2270;
wire n_22700;
wire n_22703;
wire n_22704;
wire n_22705;
wire n_22706;
wire n_22707;
wire n_22708;
wire n_22709;
wire n_2271;
wire n_22710;
wire n_22712;
wire n_22715;
wire n_22716;
wire n_22717;
wire n_22718;
wire n_22719;
wire n_2272;
wire n_22720;
wire n_22721;
wire n_22722;
wire n_22725;
wire n_22726;
wire n_22727;
wire n_22728;
wire n_22729;
wire n_2273;
wire n_22730;
wire n_22731;
wire n_22732;
wire n_22733;
wire n_22734;
wire n_22736;
wire n_22737;
wire n_22738;
wire n_22739;
wire n_2274;
wire n_22742;
wire n_22743;
wire n_22744;
wire n_22745;
wire n_22746;
wire n_22747;
wire n_22748;
wire n_22750;
wire n_22751;
wire n_22752;
wire n_22754;
wire n_22755;
wire n_22756;
wire n_22757;
wire n_22758;
wire n_22759;
wire n_2276;
wire n_22760;
wire n_22761;
wire n_22762;
wire n_22763;
wire n_22765;
wire n_22766;
wire n_22767;
wire n_22769;
wire n_2277;
wire n_22770;
wire n_22771;
wire n_22772;
wire n_22773;
wire n_22774;
wire n_22776;
wire n_22777;
wire n_22778;
wire n_2278;
wire n_22782;
wire n_22783;
wire n_22784;
wire n_22785;
wire n_22786;
wire n_22787;
wire n_22788;
wire n_22789;
wire n_2279;
wire n_22790;
wire n_22792;
wire n_22793;
wire n_22794;
wire n_22795;
wire n_22796;
wire n_228;
wire n_2280;
wire n_22800;
wire n_22801;
wire n_22802;
wire n_22803;
wire n_22804;
wire n_22806;
wire n_22807;
wire n_22808;
wire n_22809;
wire n_22810;
wire n_22811;
wire n_22812;
wire n_22813;
wire n_22814;
wire n_22815;
wire n_22816;
wire n_22817;
wire n_22818;
wire n_22819;
wire n_2282;
wire n_22820;
wire n_22822;
wire n_22823;
wire n_22826;
wire n_22827;
wire n_22828;
wire n_22829;
wire n_22832;
wire n_22833;
wire n_22834;
wire n_22835;
wire n_22839;
wire n_2284;
wire n_22840;
wire n_22841;
wire n_22842;
wire n_22843;
wire n_22844;
wire n_22845;
wire n_22846;
wire n_22847;
wire n_22848;
wire n_22849;
wire n_2285;
wire n_22850;
wire n_22851;
wire n_22852;
wire n_22853;
wire n_22854;
wire n_22855;
wire n_22856;
wire n_22857;
wire n_22858;
wire n_22859;
wire n_2286;
wire n_22861;
wire n_22862;
wire n_22864;
wire TIMEBOOST_net_2155;
wire n_22867;
wire n_22868;
wire n_22869;
wire TIMEBOOST_net_1434;
wire n_22871;
wire n_22872;
wire n_22873;
wire n_22874;
wire n_22875;
wire n_22876;
wire n_22877;
wire n_22878;
wire n_22879;
wire n_2288;
wire n_22880;
wire n_22881;
wire n_22882;
wire n_22883;
wire n_22884;
wire n_22885;
wire TIMEBOOST_net_1572;
wire n_22887;
wire n_22888;
wire n_22889;
wire n_2289;
wire n_22892;
wire n_22893;
wire n_22894;
wire n_22897;
wire n_22898;
wire n_22899;
wire n_229;
wire n_2290;
wire n_22900;
wire n_22901;
wire n_22902;
wire n_22903;
wire n_22907;
wire n_22908;
wire n_22912;
wire n_22913;
wire n_22914;
wire n_22917;
wire n_22918;
wire n_2292;
wire n_22920;
wire n_22921;
wire n_22922;
wire n_22923;
wire n_22924;
wire n_22925;
wire n_22926;
wire n_22927;
wire n_22929;
wire n_2293;
wire n_22930;
wire n_22931;
wire n_22933;
wire n_22934;
wire n_22935;
wire n_22936;
wire n_22937;
wire n_22938;
wire n_22939;
wire n_2294;
wire n_22940;
wire n_22941;
wire n_22942;
wire n_22944;
wire n_22945;
wire n_22947;
wire n_22949;
wire n_2295;
wire n_22950;
wire n_22951;
wire n_22952;
wire n_22953;
wire n_22954;
wire n_22957;
wire TIMEBOOST_net_2172;
wire n_22959;
wire n_2296;
wire n_22960;
wire n_22961;
wire n_22962;
wire n_22963;
wire n_22964;
wire n_22965;
wire n_22966;
wire n_22967;
wire n_22968;
wire n_2297;
wire n_22970;
wire n_22971;
wire n_22972;
wire n_22973;
wire n_22978;
wire n_22979;
wire n_2298;
wire n_22980;
wire n_22981;
wire n_22982;
wire n_22983;
wire n_22984;
wire n_22985;
wire n_22987;
wire TIMEBOOST_net_1471;
wire n_22989;
wire n_2299;
wire n_22990;
wire n_22991;
wire n_22992;
wire n_22993;
wire n_22994;
wire n_22995;
wire n_22996;
wire n_22998;
wire n_230;
wire n_2300;
wire n_23000;
wire n_23002;
wire n_23004;
wire n_23006;
wire n_23007;
wire n_23008;
wire n_23009;
wire n_2301;
wire n_23010;
wire n_23011;
wire n_23012;
wire n_23014;
wire n_23015;
wire n_23017;
wire n_23018;
wire n_23019;
wire n_2302;
wire TIMEBOOST_net_2803;
wire n_23022;
wire n_23023;
wire n_23026;
wire n_23027;
wire TIMEBOOST_net_841;
wire n_23029;
wire n_2303;
wire n_23030;
wire n_23031;
wire n_23032;
wire n_23033;
wire n_23034;
wire n_23035;
wire n_23036;
wire n_23037;
wire n_23038;
wire n_23039;
wire n_2304;
wire n_23040;
wire n_23042;
wire n_23043;
wire n_23044;
wire n_23045;
wire n_23046;
wire n_23047;
wire n_2305;
wire n_23051;
wire n_23052;
wire n_23053;
wire n_23054;
wire n_23055;
wire n_23056;
wire n_23057;
wire n_23058;
wire n_23059;
wire n_2306;
wire n_23060;
wire n_23061;
wire n_23064;
wire n_23066;
wire n_23067;
wire n_23069;
wire n_2307;
wire n_23071;
wire n_23072;
wire n_23073;
wire n_23074;
wire n_23075;
wire n_23077;
wire n_23078;
wire n_23079;
wire n_2308;
wire n_23083;
wire n_23084;
wire n_23085;
wire n_23086;
wire n_23087;
wire n_23088;
wire n_23089;
wire n_23090;
wire n_23091;
wire n_23092;
wire n_23093;
wire n_23094;
wire n_23095;
wire n_23096;
wire n_23097;
wire TIMEBOOST_net_812;
wire n_2310;
wire n_23100;
wire n_23101;
wire n_23105;
wire n_23106;
wire n_23107;
wire n_23108;
wire n_2311;
wire n_23110;
wire n_23111;
wire n_23112;
wire n_23113;
wire n_23114;
wire n_23115;
wire n_23116;
wire n_23117;
wire n_23118;
wire n_23119;
wire n_23120;
wire n_23121;
wire n_23122;
wire n_23123;
wire n_23124;
wire n_23126;
wire n_23127;
wire n_23128;
wire n_23129;
wire n_2313;
wire n_23131;
wire n_23132;
wire n_23133;
wire n_23135;
wire n_23136;
wire n_23137;
wire n_23138;
wire n_2314;
wire n_23140;
wire n_23141;
wire n_23142;
wire n_23143;
wire n_23144;
wire n_23145;
wire n_23148;
wire n_23149;
wire n_23150;
wire n_23151;
wire n_23152;
wire n_23153;
wire n_23154;
wire n_23155;
wire n_23156;
wire n_23157;
wire n_23158;
wire n_23159;
wire n_23160;
wire n_23161;
wire n_23165;
wire n_23166;
wire n_23167;
wire n_23169;
wire n_2317;
wire n_23170;
wire n_23172;
wire n_23173;
wire n_23174;
wire n_23175;
wire n_23176;
wire TIMEBOOST_net_805;
wire n_23178;
wire n_23179;
wire n_2318;
wire n_23181;
wire n_23182;
wire n_23183;
wire n_23184;
wire n_23185;
wire n_23186;
wire n_23187;
wire n_23188;
wire n_23189;
wire n_2319;
wire n_23190;
wire n_23191;
wire n_23192;
wire n_23193;
wire n_23194;
wire n_23195;
wire n_23196;
wire n_23197;
wire n_232;
wire n_2320;
wire n_23201;
wire n_23202;
wire n_23204;
wire n_23205;
wire n_23206;
wire n_23207;
wire n_23208;
wire n_2321;
wire n_23210;
wire n_23211;
wire n_23212;
wire n_23213;
wire n_23214;
wire n_23215;
wire n_23216;
wire n_2322;
wire n_23220;
wire n_23221;
wire n_23222;
wire n_23223;
wire n_23224;
wire n_23225;
wire n_23226;
wire n_23227;
wire n_23228;
wire n_23229;
wire n_2323;
wire TIMEBOOST_net_1568;
wire n_23232;
wire n_23234;
wire n_23235;
wire n_23236;
wire n_23237;
wire TIMEBOOST_net_860;
wire n_2324;
wire n_23242;
wire n_23243;
wire n_23244;
wire n_23245;
wire n_23246;
wire n_23248;
wire n_23249;
wire n_2325;
wire n_23250;
wire n_23251;
wire n_23252;
wire n_23253;
wire n_23254;
wire n_23259;
wire n_2326;
wire n_23260;
wire n_23261;
wire n_23264;
wire n_23265;
wire n_23266;
wire n_23267;
wire n_23269;
wire n_2327;
wire n_23270;
wire n_23271;
wire n_23276;
wire TIMEBOOST_net_55;
wire n_23278;
wire n_23279;
wire n_2328;
wire n_23281;
wire n_23282;
wire n_23283;
wire n_23284;
wire n_23286;
wire n_23287;
wire n_23288;
wire n_23289;
wire n_2329;
wire n_23290;
wire n_23291;
wire n_23294;
wire n_23295;
wire n_23296;
wire n_23297;
wire n_23298;
wire n_23299;
wire n_233;
wire n_2330;
wire n_23300;
wire n_23301;
wire n_23302;
wire n_23303;
wire n_23304;
wire n_23305;
wire n_23307;
wire n_23308;
wire n_23309;
wire n_2331;
wire n_23310;
wire n_23311;
wire n_23312;
wire n_23313;
wire TIMEBOOST_net_2129;
wire n_23315;
wire n_23317;
wire n_23319;
wire n_2332;
wire n_23320;
wire n_23321;
wire n_23322;
wire TIMEBOOST_net_2136;
wire n_23325;
wire n_23326;
wire n_23327;
wire n_23328;
wire n_23329;
wire n_2333;
wire n_23330;
wire n_23331;
wire n_23332;
wire n_23333;
wire n_23334;
wire n_23335;
wire n_23336;
wire n_23339;
wire n_23341;
wire n_23342;
wire n_23343;
wire n_23344;
wire n_23345;
wire n_23346;
wire n_23347;
wire n_23348;
wire n_23349;
wire n_2335;
wire n_23350;
wire n_23353;
wire n_23356;
wire n_23357;
wire n_23358;
wire n_23359;
wire n_2336;
wire n_23360;
wire n_23361;
wire TIMEBOOST_net_2746;
wire n_23363;
wire n_23365;
wire n_23366;
wire n_23367;
wire n_23368;
wire n_23369;
wire TIMEBOOST_net_1084;
wire n_23370;
wire n_23371;
wire n_23373;
wire n_23374;
wire n_23376;
wire n_23377;
wire n_23378;
wire n_2338;
wire n_23380;
wire n_23382;
wire n_23383;
wire n_23384;
wire n_23385;
wire n_23386;
wire n_23387;
wire n_23388;
wire n_23390;
wire n_23391;
wire n_23393;
wire n_23394;
wire n_23395;
wire n_23396;
wire n_23397;
wire n_23398;
wire n_23399;
wire n_234;
wire n_2340;
wire n_23400;
wire n_23403;
wire n_23404;
wire n_23405;
wire n_23407;
wire n_23408;
wire n_23409;
wire n_2341;
wire n_23410;
wire n_23411;
wire n_23412;
wire n_23414;
wire n_23416;
wire n_23417;
wire n_23418;
wire n_23419;
wire n_2342;
wire n_23420;
wire TIMEBOOST_net_2253;
wire n_23422;
wire n_23423;
wire n_23424;
wire TIMEBOOST_net_2795;
wire n_23426;
wire n_23427;
wire n_23428;
wire n_23429;
wire n_2343;
wire n_23430;
wire n_23431;
wire n_23432;
wire n_23437;
wire n_23438;
wire n_23439;
wire n_2344;
wire TIMEBOOST_net_1494;
wire n_23441;
wire n_23443;
wire n_23444;
wire n_23445;
wire n_23447;
wire n_23448;
wire n_23449;
wire n_2345;
wire n_23450;
wire n_23451;
wire n_23452;
wire n_23453;
wire n_23455;
wire n_23456;
wire n_23457;
wire n_23458;
wire n_23459;
wire n_2346;
wire n_23461;
wire n_23462;
wire n_23463;
wire TIMEBOOST_net_1497;
wire n_23466;
wire n_23468;
wire n_23469;
wire n_2347;
wire TIMEBOOST_net_820;
wire n_23471;
wire n_23472;
wire n_23473;
wire n_23474;
wire n_23475;
wire n_23476;
wire TIMEBOOST_net_887;
wire n_23479;
wire n_2348;
wire n_23480;
wire n_23481;
wire n_23482;
wire TIMEBOOST_net_2145;
wire n_23486;
wire n_23488;
wire n_23489;
wire n_2349;
wire n_23490;
wire n_23491;
wire n_23492;
wire n_23493;
wire n_23494;
wire n_23495;
wire n_23496;
wire n_23497;
wire n_23498;
wire n_23499;
wire n_235;
wire n_2350;
wire n_23500;
wire TIMEBOOST_net_925;
wire n_23502;
wire n_23503;
wire n_23504;
wire TIMEBOOST_net_68;
wire n_23506;
wire n_23507;
wire n_23508;
wire n_23509;
wire n_2351;
wire n_23512;
wire n_23513;
wire n_23514;
wire n_23515;
wire n_23516;
wire n_23517;
wire n_23518;
wire n_23519;
wire n_2352;
wire n_23520;
wire n_23521;
wire n_23522;
wire n_23523;
wire n_23524;
wire n_23526;
wire n_23527;
wire n_23528;
wire n_23529;
wire n_2353;
wire n_23530;
wire n_23531;
wire n_23532;
wire n_23533;
wire n_23534;
wire n_23535;
wire TIMEBOOST_net_71;
wire n_23537;
wire n_23538;
wire n_23539;
wire n_2354;
wire n_23540;
wire n_23541;
wire n_23542;
wire n_23543;
wire n_23544;
wire n_23545;
wire n_23546;
wire n_23547;
wire n_23548;
wire n_23549;
wire n_2355;
wire n_23550;
wire n_23551;
wire n_23554;
wire n_23555;
wire n_23556;
wire n_23557;
wire n_23558;
wire n_23559;
wire TIMEBOOST_net_243;
wire n_23560;
wire n_23561;
wire n_23562;
wire n_23563;
wire n_23564;
wire n_23565;
wire n_23566;
wire n_23567;
wire n_23568;
wire n_23569;
wire n_2357;
wire n_23570;
wire n_23571;
wire n_23572;
wire n_23574;
wire n_23576;
wire n_23577;
wire n_23578;
wire n_23579;
wire n_2358;
wire n_23580;
wire n_23581;
wire n_23582;
wire TIMEBOOST_net_2133;
wire n_23584;
wire TIMEBOOST_net_1868;
wire n_23586;
wire n_23587;
wire n_23588;
wire n_2359;
wire n_23590;
wire n_23591;
wire n_23592;
wire n_23593;
wire n_23594;
wire n_23595;
wire n_23596;
wire n_23599;
wire n_236;
wire n_2360;
wire n_23600;
wire n_23601;
wire n_23602;
wire n_23603;
wire n_23604;
wire n_23605;
wire n_23606;
wire TIMEBOOST_net_76;
wire TIMEBOOST_net_2350;
wire n_23609;
wire n_2361;
wire n_23611;
wire n_23613;
wire n_23615;
wire n_23616;
wire TIMEBOOST_net_113;
wire n_23618;
wire n_23619;
wire n_23620;
wire n_23626;
wire n_23627;
wire n_23628;
wire n_23629;
wire n_2363;
wire n_23630;
wire n_23631;
wire n_23632;
wire n_23633;
wire n_23634;
wire n_23635;
wire n_23636;
wire n_23637;
wire n_23638;
wire n_23639;
wire n_2364;
wire n_23640;
wire n_23641;
wire n_23642;
wire n_23643;
wire n_23644;
wire n_23645;
wire n_23646;
wire n_23647;
wire n_23648;
wire n_23649;
wire n_23651;
wire n_23652;
wire n_23653;
wire n_23656;
wire n_23658;
wire n_23659;
wire n_2366;
wire TIMEBOOST_net_2731;
wire n_23661;
wire n_23662;
wire n_23663;
wire n_23664;
wire n_23665;
wire n_23666;
wire n_23668;
wire n_23669;
wire n_2367;
wire n_23670;
wire n_23671;
wire n_23672;
wire n_23675;
wire n_23676;
wire n_23677;
wire n_23679;
wire n_2368;
wire n_23680;
wire n_23681;
wire n_23682;
wire n_23683;
wire n_23684;
wire n_23685;
wire TIMEBOOST_net_916;
wire n_23687;
wire n_23688;
wire n_23689;
wire n_2369;
wire n_23690;
wire n_23691;
wire n_23692;
wire n_23693;
wire n_23694;
wire n_23695;
wire n_23697;
wire n_23698;
wire n_23699;
wire n_237;
wire n_2370;
wire n_23700;
wire n_23701;
wire n_23702;
wire n_23703;
wire n_23704;
wire n_23705;
wire n_23707;
wire n_23708;
wire n_23709;
wire TIMEBOOST_net_1552;
wire n_23711;
wire n_23712;
wire n_23713;
wire n_23714;
wire n_23716;
wire n_23717;
wire n_23718;
wire n_23719;
wire TIMEBOOST_net_1894;
wire n_23720;
wire n_23721;
wire n_23722;
wire n_23723;
wire n_23724;
wire n_2373;
wire n_23731;
wire n_23732;
wire n_23733;
wire n_23734;
wire n_23735;
wire n_23736;
wire n_23737;
wire n_23738;
wire n_23739;
wire n_2374;
wire n_23740;
wire n_23741;
wire n_23742;
wire n_23743;
wire n_23746;
wire n_23747;
wire n_23748;
wire n_23749;
wire n_2375;
wire n_23750;
wire n_23751;
wire n_23752;
wire n_23753;
wire n_23754;
wire n_23757;
wire n_23758;
wire n_23759;
wire n_23760;
wire n_23761;
wire n_23762;
wire n_23763;
wire n_23764;
wire n_23765;
wire n_23766;
wire n_23767;
wire n_23768;
wire n_23769;
wire n_23770;
wire n_23771;
wire n_23772;
wire n_23773;
wire n_23774;
wire n_23775;
wire n_23777;
wire n_23778;
wire n_23779;
wire n_2378;
wire n_23783;
wire n_23786;
wire n_23787;
wire n_23788;
wire n_23789;
wire n_2379;
wire n_23790;
wire n_23791;
wire n_23792;
wire n_23793;
wire n_23794;
wire n_23795;
wire n_23796;
wire n_23797;
wire n_23798;
wire n_238;
wire n_2380;
wire n_23800;
wire n_23801;
wire n_23802;
wire n_23803;
wire n_23804;
wire n_23806;
wire n_23807;
wire n_23808;
wire n_23809;
wire n_2381;
wire n_23810;
wire n_23811;
wire n_23812;
wire n_23813;
wire n_23814;
wire n_23815;
wire n_23817;
wire n_23818;
wire n_23819;
wire n_2382;
wire n_23820;
wire n_23821;
wire n_23822;
wire n_23823;
wire n_23824;
wire n_23825;
wire n_23826;
wire n_23827;
wire n_2383;
wire n_23830;
wire n_23831;
wire n_23832;
wire n_23833;
wire n_23834;
wire n_23836;
wire n_23837;
wire n_23838;
wire n_2384;
wire n_23844;
wire n_23845;
wire n_23846;
wire n_23847;
wire n_23848;
wire n_2385;
wire n_23850;
wire n_23851;
wire n_23853;
wire n_23854;
wire n_23855;
wire n_23856;
wire n_23857;
wire n_23859;
wire n_2386;
wire n_23860;
wire n_23862;
wire n_23863;
wire n_23864;
wire n_23865;
wire n_23866;
wire n_23867;
wire n_23868;
wire n_23869;
wire n_2387;
wire TIMEBOOST_net_953;
wire n_23872;
wire n_23873;
wire n_23874;
wire n_23876;
wire n_23878;
wire n_23879;
wire n_2388;
wire n_23880;
wire n_23881;
wire n_23883;
wire n_23884;
wire n_23885;
wire n_23886;
wire n_23887;
wire n_23888;
wire n_23889;
wire n_2389;
wire n_23890;
wire n_23891;
wire n_23892;
wire n_23894;
wire n_23895;
wire n_23897;
wire n_23898;
wire n_23899;
wire TIMEBOOST_net_2620;
wire n_2390;
wire n_23900;
wire n_23901;
wire n_23903;
wire n_23904;
wire n_23905;
wire n_23906;
wire n_23907;
wire n_23908;
wire n_23909;
wire n_2391;
wire n_23910;
wire n_23911;
wire n_23914;
wire n_23917;
wire n_23918;
wire n_23919;
wire n_2392;
wire n_23920;
wire n_23921;
wire n_23922;
wire n_23923;
wire n_23924;
wire n_23925;
wire n_23926;
wire n_23927;
wire n_23928;
wire n_2393;
wire n_23930;
wire n_23932;
wire n_23933;
wire n_23934;
wire n_23936;
wire n_23937;
wire n_23938;
wire n_23939;
wire n_2394;
wire n_23941;
wire n_23943;
wire n_23944;
wire n_23945;
wire n_23946;
wire n_23947;
wire n_23948;
wire n_23949;
wire TIMEBOOST_net_1106;
wire n_23950;
wire n_23951;
wire n_23952;
wire n_23953;
wire n_23954;
wire n_23955;
wire n_23956;
wire n_23957;
wire n_23958;
wire n_23959;
wire n_2396;
wire n_23962;
wire n_23963;
wire n_23964;
wire n_23965;
wire n_23966;
wire n_23967;
wire n_23968;
wire n_23969;
wire n_2397;
wire n_23970;
wire n_23971;
wire n_23972;
wire n_23973;
wire n_23978;
wire n_23979;
wire n_2398;
wire n_23980;
wire n_23981;
wire n_23984;
wire n_23985;
wire n_23986;
wire n_23987;
wire n_23988;
wire n_23989;
wire n_23990;
wire n_23991;
wire n_23992;
wire n_23993;
wire n_23994;
wire n_23995;
wire n_23996;
wire n_23997;
wire n_23998;
wire n_23999;
wire n_240;
wire n_24000;
wire n_24001;
wire n_24002;
wire n_24003;
wire n_24005;
wire n_24006;
wire n_24007;
wire n_24008;
wire n_24009;
wire TIMEBOOST_net_251;
wire n_24010;
wire n_24011;
wire n_24012;
wire n_24013;
wire n_24014;
wire n_24015;
wire n_24016;
wire n_24017;
wire n_24018;
wire n_24019;
wire n_2402;
wire n_24023;
wire n_24024;
wire n_24025;
wire n_24026;
wire n_24028;
wire n_24029;
wire n_24030;
wire n_24031;
wire n_24032;
wire n_24033;
wire n_24034;
wire n_24035;
wire n_24036;
wire n_24037;
wire n_24039;
wire n_2404;
wire n_24040;
wire n_24041;
wire n_24042;
wire n_24043;
wire n_24044;
wire n_24045;
wire n_24046;
wire n_24047;
wire n_24048;
wire n_24049;
wire n_2405;
wire n_24050;
wire n_24051;
wire n_24052;
wire n_24053;
wire n_24054;
wire n_24055;
wire n_24056;
wire n_24057;
wire TIMEBOOST_net_165;
wire n_24059;
wire n_2406;
wire n_24061;
wire n_24062;
wire n_24063;
wire n_24064;
wire n_24065;
wire n_24066;
wire n_24067;
wire n_24068;
wire TIMEBOOST_net_143;
wire n_2407;
wire n_24070;
wire n_24071;
wire n_24072;
wire n_24074;
wire n_24075;
wire n_24076;
wire n_24077;
wire n_24078;
wire n_24079;
wire n_2408;
wire n_24080;
wire n_24081;
wire TIMEBOOST_net_2192;
wire n_24084;
wire n_24085;
wire n_24086;
wire n_24087;
wire n_24088;
wire n_24090;
wire n_24091;
wire n_24092;
wire n_24093;
wire n_24094;
wire TIMEBOOST_net_982;
wire n_24097;
wire n_24099;
wire n_241;
wire n_2410;
wire n_24100;
wire n_24101;
wire n_24102;
wire n_24105;
wire n_24106;
wire n_24107;
wire TIMEBOOST_net_2744;
wire n_24110;
wire n_24111;
wire n_24112;
wire n_24113;
wire n_24114;
wire n_24115;
wire n_24119;
wire n_2412;
wire n_24121;
wire n_24122;
wire n_24125;
wire n_24127;
wire TIMEBOOST_net_168;
wire n_2413;
wire n_24131;
wire n_24132;
wire n_24137;
wire n_24139;
wire n_24142;
wire n_24143;
wire n_24144;
wire n_24145;
wire n_24146;
wire n_24147;
wire n_24148;
wire n_24149;
wire TIMEBOOST_net_1050;
wire n_24150;
wire n_24151;
wire n_24152;
wire n_24153;
wire n_24154;
wire n_24155;
wire n_24157;
wire n_24158;
wire n_24159;
wire n_2416;
wire n_24160;
wire n_24162;
wire n_24163;
wire n_24164;
wire n_24165;
wire n_24166;
wire n_24169;
wire n_24170;
wire n_24171;
wire n_24172;
wire n_24173;
wire n_24175;
wire TIMEBOOST_net_2555;
wire n_24178;
wire n_24181;
wire n_24182;
wire n_24183;
wire TIMEBOOST_net_221;
wire n_24185;
wire TIMEBOOST_net_220;
wire n_24188;
wire n_24189;
wire n_2419;
wire n_24190;
wire n_24191;
wire n_24192;
wire n_24193;
wire n_24194;
wire n_24195;
wire n_24196;
wire TIMEBOOST_net_2740;
wire n_2420;
wire n_24200;
wire n_24201;
wire TIMEBOOST_net_898;
wire TIMEBOOST_net_2663;
wire n_24204;
wire n_24207;
wire n_24208;
wire n_2421;
wire n_24210;
wire n_24215;
wire n_24217;
wire n_24218;
wire n_24219;
wire n_2422;
wire n_24221;
wire n_24222;
wire n_24224;
wire n_24225;
wire TIMEBOOST_net_1580;
wire n_24229;
wire n_2423;
wire n_24230;
wire n_24231;
wire TIMEBOOST_net_1981;
wire n_24234;
wire n_24235;
wire n_24236;
wire n_24237;
wire n_24238;
wire n_24239;
wire n_2424;
wire n_24240;
wire n_24241;
wire n_24246;
wire TIMEBOOST_net_2821;
wire n_24248;
wire n_24249;
wire n_2425;
wire n_24250;
wire n_24251;
wire n_24254;
wire n_24256;
wire n_24257;
wire n_24258;
wire n_24259;
wire n_2426;
wire n_24262;
wire n_24263;
wire n_24264;
wire n_24265;
wire n_24267;
wire n_24268;
wire n_24269;
wire n_2427;
wire n_24270;
wire n_24272;
wire TIMEBOOST_net_1534;
wire n_24274;
wire n_24275;
wire n_24276;
wire n_24277;
wire n_2428;
wire n_24283;
wire n_24284;
wire n_24285;
wire TIMEBOOST_net_203;
wire n_24288;
wire n_24289;
wire n_2429;
wire n_24290;
wire n_24291;
wire n_24292;
wire n_24293;
wire TIMEBOOST_net_228;
wire TIMEBOOST_net_1975;
wire n_24297;
wire n_24299;
wire n_243;
wire n_2430;
wire n_24300;
wire n_24301;
wire n_24302;
wire n_24305;
wire n_24306;
wire n_24307;
wire n_24308;
wire n_24309;
wire n_2431;
wire n_24310;
wire n_24311;
wire n_24312;
wire TIMEBOOST_net_230;
wire TIMEBOOST_net_229;
wire n_24316;
wire n_24318;
wire n_24319;
wire n_2432;
wire n_24320;
wire n_24321;
wire n_24322;
wire n_24323;
wire n_24325;
wire n_24326;
wire n_24327;
wire n_2433;
wire n_24330;
wire n_24332;
wire n_24336;
wire n_24339;
wire n_2434;
wire n_24340;
wire n_24341;
wire n_24342;
wire n_24343;
wire n_24344;
wire n_24345;
wire n_24346;
wire n_24347;
wire n_24348;
wire TIMEBOOST_net_2551;
wire n_24350;
wire n_24352;
wire n_24354;
wire n_24355;
wire n_24359;
wire n_2436;
wire n_24360;
wire n_24361;
wire n_24362;
wire n_24363;
wire n_24364;
wire n_24366;
wire n_24367;
wire n_24368;
wire n_24369;
wire n_2437;
wire n_24370;
wire n_24372;
wire n_24373;
wire n_24375;
wire n_24379;
wire n_24380;
wire n_24381;
wire n_24382;
wire n_24383;
wire n_24384;
wire n_24386;
wire n_24389;
wire n_2439;
wire n_24390;
wire n_24391;
wire n_24392;
wire n_24393;
wire n_24394;
wire n_24395;
wire n_24396;
wire TIMEBOOST_net_214;
wire n_24398;
wire n_24399;
wire n_244;
wire n_2440;
wire n_24402;
wire TIMEBOOST_net_235;
wire n_24404;
wire n_24405;
wire n_24406;
wire n_24407;
wire n_24408;
wire n_2441;
wire TIMEBOOST_net_2925;
wire TIMEBOOST_net_1983;
wire n_24414;
wire n_24415;
wire n_24416;
wire n_24417;
wire n_24419;
wire n_2442;
wire n_24420;
wire n_24421;
wire n_24422;
wire n_24423;
wire n_24424;
wire n_24425;
wire n_24426;
wire n_24429;
wire n_2443;
wire n_24432;
wire n_24433;
wire TIMEBOOST_net_2060;
wire TIMEBOOST_net_234;
wire n_24436;
wire n_24438;
wire TIMEBOOST_net_2211;
wire n_24441;
wire n_24442;
wire n_24443;
wire n_24444;
wire n_24445;
wire n_24446;
wire n_24447;
wire n_24448;
wire n_24449;
wire n_2445;
wire n_24451;
wire n_24452;
wire n_24453;
wire n_24454;
wire n_24455;
wire n_24456;
wire n_24457;
wire n_24458;
wire n_2446;
wire n_24461;
wire n_24462;
wire n_24463;
wire n_24464;
wire n_24465;
wire n_24466;
wire n_24467;
wire n_24469;
wire n_2447;
wire n_24471;
wire n_24472;
wire n_24473;
wire TIMEBOOST_net_248;
wire n_24476;
wire n_24477;
wire n_24478;
wire n_24479;
wire n_2448;
wire n_24480;
wire n_24481;
wire n_24484;
wire n_24485;
wire n_24486;
wire n_24488;
wire n_24489;
wire n_2449;
wire n_24490;
wire n_24491;
wire n_24492;
wire n_24493;
wire n_24494;
wire TIMEBOOST_net_2219;
wire n_24497;
wire n_24498;
wire n_24499;
wire n_245;
wire n_2450;
wire n_24500;
wire n_24501;
wire n_24502;
wire n_24503;
wire n_24505;
wire n_24506;
wire n_24507;
wire n_24508;
wire n_2451;
wire n_24510;
wire TIMEBOOST_net_2877;
wire n_24513;
wire n_24514;
wire n_24515;
wire n_24518;
wire n_24519;
wire n_2452;
wire n_24520;
wire n_24521;
wire n_24522;
wire TIMEBOOST_net_1892;
wire n_24529;
wire n_2453;
wire n_24531;
wire n_24532;
wire n_24534;
wire n_24535;
wire n_24536;
wire n_24537;
wire n_24539;
wire n_24541;
wire n_24542;
wire n_24543;
wire n_24544;
wire n_24546;
wire n_24547;
wire n_24548;
wire n_24549;
wire n_2455;
wire n_24550;
wire n_24551;
wire TIMEBOOST_net_2411;
wire n_24553;
wire n_24554;
wire n_24555;
wire n_24556;
wire n_2456;
wire n_24560;
wire n_24561;
wire n_24562;
wire n_24563;
wire TIMEBOOST_net_2948;
wire n_24566;
wire n_24568;
wire n_24569;
wire n_2457;
wire n_24570;
wire TIMEBOOST_net_238;
wire n_24573;
wire n_24574;
wire n_24576;
wire n_24577;
wire n_24578;
wire n_24579;
wire n_2458;
wire n_24580;
wire n_24581;
wire n_24582;
wire n_24585;
wire n_24586;
wire n_24587;
wire n_24588;
wire n_24590;
wire n_24591;
wire n_24592;
wire n_24593;
wire TIMEBOOST_net_1583;
wire TIMEBOOST_net_1073;
wire n_24598;
wire n_246;
wire n_2460;
wire TIMEBOOST_net_1893;
wire n_24601;
wire n_24602;
wire TIMEBOOST_net_260;
wire n_24604;
wire n_24605;
wire n_24606;
wire n_24607;
wire n_24608;
wire n_24609;
wire n_2461;
wire n_24610;
wire n_24612;
wire n_24613;
wire n_24614;
wire TIMEBOOST_net_171;
wire TIMEBOOST_net_249;
wire n_24618;
wire TIMEBOOST_net_2321;
wire n_24620;
wire n_24621;
wire TIMEBOOST_net_963;
wire n_24623;
wire n_24624;
wire TIMEBOOST_net_1673;
wire n_24626;
wire n_24627;
wire n_24628;
wire n_24629;
wire n_2463;
wire n_24630;
wire n_24632;
wire n_24633;
wire n_24635;
wire n_24636;
wire n_24637;
wire n_24638;
wire n_24639;
wire n_2464;
wire n_24642;
wire n_24645;
wire n_24646;
wire TIMEBOOST_net_177;
wire n_24648;
wire n_2465;
wire n_24650;
wire TIMEBOOST_net_1081;
wire n_24652;
wire n_24653;
wire n_24655;
wire n_24656;
wire n_24657;
wire n_24659;
wire n_2466;
wire n_24660;
wire n_24661;
wire n_24664;
wire n_24665;
wire n_24666;
wire n_24667;
wire n_24668;
wire n_24669;
wire n_2467;
wire n_24670;
wire n_24671;
wire n_24672;
wire n_24673;
wire n_24674;
wire n_24675;
wire n_24676;
wire n_24677;
wire n_24680;
wire n_24682;
wire n_24683;
wire n_24684;
wire n_24685;
wire TIMEBOOST_net_176;
wire n_24687;
wire n_24688;
wire n_2469;
wire n_24690;
wire n_24691;
wire n_24692;
wire n_24694;
wire n_24695;
wire TIMEBOOST_net_242;
wire TIMEBOOST_net_1683;
wire n_24698;
wire n_24699;
wire n_247;
wire TIMEBOOST_net_2574;
wire TIMEBOOST_net_1203;
wire n_24701;
wire n_24702;
wire n_24703;
wire n_24704;
wire n_24705;
wire n_24706;
wire n_24707;
wire n_24708;
wire n_24711;
wire n_24712;
wire n_24713;
wire n_24714;
wire n_24715;
wire n_24716;
wire n_24717;
wire n_24718;
wire n_24719;
wire n_2472;
wire n_24720;
wire n_24721;
wire n_24722;
wire n_24723;
wire n_24726;
wire TIMEBOOST_net_1995;
wire n_24729;
wire n_2473;
wire n_24733;
wire n_24734;
wire n_24735;
wire n_24736;
wire n_24737;
wire n_24738;
wire n_24739;
wire n_2474;
wire n_24740;
wire n_24741;
wire n_24742;
wire n_24743;
wire n_24746;
wire n_24747;
wire n_24748;
wire n_2475;
wire n_24750;
wire n_24751;
wire n_24752;
wire n_24754;
wire TIMEBOOST_net_1012;
wire n_24756;
wire n_24757;
wire TIMEBOOST_net_1598;
wire n_2476;
wire n_24760;
wire n_24761;
wire n_24762;
wire n_24763;
wire n_24764;
wire n_24765;
wire n_24766;
wire n_24767;
wire n_24768;
wire n_24769;
wire n_2477;
wire n_24770;
wire n_24771;
wire n_24774;
wire n_24775;
wire n_24776;
wire n_24777;
wire n_24778;
wire n_24779;
wire n_2478;
wire n_24780;
wire n_24781;
wire n_24782;
wire n_24783;
wire n_24784;
wire n_24785;
wire n_24787;
wire n_24788;
wire n_2479;
wire n_24791;
wire n_24792;
wire n_24793;
wire n_24794;
wire n_24797;
wire n_24798;
wire n_24799;
wire n_248;
wire n_2480;
wire n_24800;
wire TIMEBOOST_net_233;
wire n_24802;
wire n_24803;
wire n_24804;
wire n_24805;
wire TIMEBOOST_net_2621;
wire n_24808;
wire n_24810;
wire n_24813;
wire n_24815;
wire n_24816;
wire n_24817;
wire TIMEBOOST_net_223;
wire n_24819;
wire n_24820;
wire n_24821;
wire n_24822;
wire n_24823;
wire n_24825;
wire n_24826;
wire n_24828;
wire n_24829;
wire n_2483;
wire n_24830;
wire n_24831;
wire n_24832;
wire n_24833;
wire n_24834;
wire n_24836;
wire n_24837;
wire n_24838;
wire n_24839;
wire n_2484;
wire n_24842;
wire n_24844;
wire n_24845;
wire n_24846;
wire n_24848;
wire n_2485;
wire n_24850;
wire n_24851;
wire n_24852;
wire n_24853;
wire n_24857;
wire TIMEBOOST_net_186;
wire n_24859;
wire n_2486;
wire n_24860;
wire n_24861;
wire n_24862;
wire n_24864;
wire n_24865;
wire n_24867;
wire n_24868;
wire n_24869;
wire n_2487;
wire n_24870;
wire n_24872;
wire n_24873;
wire n_24874;
wire n_24875;
wire n_24876;
wire n_24877;
wire n_24878;
wire n_24879;
wire n_2488;
wire n_24880;
wire n_24881;
wire n_24882;
wire n_24883;
wire n_24884;
wire n_24887;
wire n_2489;
wire n_24891;
wire n_24892;
wire n_24893;
wire n_24894;
wire n_24895;
wire n_24896;
wire n_24897;
wire n_24898;
wire n_24899;
wire n_249;
wire n_24900;
wire n_24901;
wire n_24902;
wire n_24903;
wire n_24904;
wire n_24905;
wire n_24906;
wire n_24907;
wire n_24908;
wire n_24909;
wire n_2491;
wire n_24910;
wire n_24911;
wire n_24912;
wire n_24913;
wire n_24914;
wire n_24915;
wire TIMEBOOST_net_920;
wire n_24918;
wire n_24919;
wire n_2492;
wire n_24920;
wire n_24921;
wire n_24922;
wire n_24923;
wire n_24924;
wire n_24929;
wire TIMEBOOST_net_1046;
wire n_24930;
wire n_24932;
wire n_24933;
wire n_24934;
wire n_24935;
wire n_24936;
wire n_24937;
wire n_24938;
wire n_24939;
wire n_2494;
wire n_24940;
wire n_24941;
wire n_24942;
wire n_24943;
wire n_24944;
wire n_24945;
wire n_24946;
wire n_2495;
wire n_24953;
wire n_24954;
wire n_24955;
wire n_24956;
wire n_24957;
wire n_24958;
wire n_24959;
wire n_2496;
wire TIMEBOOST_net_1927;
wire n_24961;
wire n_24962;
wire n_24963;
wire n_24964;
wire n_24966;
wire n_24967;
wire n_24968;
wire n_24969;
wire n_2497;
wire n_24970;
wire n_24971;
wire n_24972;
wire n_24974;
wire n_24975;
wire n_24976;
wire n_24977;
wire n_24978;
wire n_24979;
wire n_2498;
wire n_24980;
wire n_24981;
wire n_24982;
wire n_24983;
wire n_24984;
wire n_24985;
wire n_24986;
wire n_24987;
wire n_24989;
wire n_2499;
wire n_24990;
wire n_24992;
wire n_24993;
wire n_24994;
wire n_24995;
wire n_24996;
wire n_24997;
wire n_24998;
wire n_24999;
wire n_250;
wire n_2500;
wire n_25000;
wire n_25001;
wire n_25002;
wire n_25003;
wire n_25004;
wire n_25005;
wire n_25006;
wire n_25007;
wire n_25008;
wire n_2501;
wire TIMEBOOST_net_2730;
wire n_25011;
wire n_25013;
wire n_25015;
wire n_25016;
wire n_25017;
wire n_25018;
wire TIMEBOOST_net_1213;
wire n_2502;
wire n_25020;
wire n_25021;
wire n_25022;
wire n_25023;
wire n_25024;
wire n_25025;
wire n_25026;
wire n_25027;
wire n_25028;
wire n_25029;
wire n_2503;
wire n_25030;
wire n_25031;
wire n_25032;
wire n_25033;
wire TIMEBOOST_net_236;
wire n_25035;
wire n_25036;
wire n_25037;
wire n_25038;
wire n_25039;
wire n_2504;
wire n_25040;
wire n_25041;
wire n_25042;
wire TIMEBOOST_net_2833;
wire n_25044;
wire n_25045;
wire n_25046;
wire n_25047;
wire n_25048;
wire n_25049;
wire n_2505;
wire n_25050;
wire n_25052;
wire n_25053;
wire n_25055;
wire n_25056;
wire n_25057;
wire n_25058;
wire n_25059;
wire n_2506;
wire n_25060;
wire n_25061;
wire n_25062;
wire n_25063;
wire n_25064;
wire n_25065;
wire n_25066;
wire n_25067;
wire TIMEBOOST_net_2720;
wire n_25069;
wire TIMEBOOST_net_1108;
wire n_25070;
wire n_25071;
wire n_25072;
wire n_25073;
wire n_25074;
wire n_25075;
wire n_25076;
wire n_25077;
wire n_2508;
wire n_25081;
wire n_25082;
wire n_25083;
wire n_25084;
wire n_25085;
wire n_25086;
wire n_25087;
wire n_25088;
wire n_25089;
wire n_25090;
wire TIMEBOOST_net_2358;
wire n_25092;
wire n_25093;
wire n_25094;
wire n_25095;
wire n_25096;
wire TIMEBOOST_net_2437;
wire n_25098;
wire n_25099;
wire n_251;
wire n_2510;
wire n_25100;
wire n_25101;
wire n_25102;
wire n_25103;
wire n_25104;
wire n_25105;
wire n_25106;
wire n_25107;
wire n_25108;
wire n_25109;
wire n_2511;
wire n_25111;
wire n_25112;
wire n_25113;
wire n_25114;
wire n_25116;
wire n_25117;
wire n_25118;
wire n_25119;
wire n_2512;
wire n_25120;
wire n_25122;
wire n_25124;
wire n_25125;
wire n_25126;
wire n_25127;
wire n_25128;
wire n_25129;
wire n_25130;
wire n_25132;
wire n_25133;
wire n_25134;
wire n_25135;
wire n_25136;
wire n_25138;
wire n_25139;
wire n_2514;
wire n_25140;
wire n_25141;
wire n_25142;
wire n_25143;
wire n_25144;
wire n_25145;
wire n_25146;
wire n_25147;
wire n_25148;
wire n_25149;
wire n_2515;
wire n_25150;
wire n_25151;
wire n_25152;
wire n_25153;
wire n_25154;
wire n_25155;
wire n_25157;
wire n_25158;
wire n_2516;
wire n_25160;
wire n_25161;
wire n_25162;
wire n_25163;
wire n_25164;
wire n_25166;
wire n_25167;
wire n_25168;
wire n_25169;
wire n_2517;
wire TIMEBOOST_net_2747;
wire n_25172;
wire n_25175;
wire n_25176;
wire n_25178;
wire n_25179;
wire n_2518;
wire n_25180;
wire n_25181;
wire n_25182;
wire n_25184;
wire n_25185;
wire n_25186;
wire n_25187;
wire n_25188;
wire n_25189;
wire n_2519;
wire n_25191;
wire n_25192;
wire n_25193;
wire n_25194;
wire n_25195;
wire n_25196;
wire n_25197;
wire n_25198;
wire n_25199;
wire n_252;
wire n_2520;
wire n_25200;
wire n_25203;
wire n_25204;
wire n_25205;
wire n_25206;
wire n_25207;
wire n_25208;
wire n_25209;
wire n_2521;
wire n_25210;
wire n_25211;
wire n_25212;
wire n_25213;
wire n_25216;
wire n_25217;
wire n_25218;
wire n_25219;
wire n_2522;
wire n_25220;
wire n_25221;
wire n_25222;
wire n_25223;
wire n_25224;
wire n_25229;
wire n_2523;
wire n_25231;
wire n_25233;
wire n_25234;
wire n_25239;
wire n_2524;
wire n_25241;
wire n_25242;
wire n_25243;
wire n_25244;
wire n_25245;
wire n_25246;
wire n_25247;
wire n_25248;
wire n_2525;
wire n_25250;
wire n_25251;
wire n_25253;
wire n_25254;
wire n_25256;
wire n_25257;
wire n_25258;
wire n_25259;
wire n_2526;
wire n_25261;
wire n_25262;
wire n_25265;
wire n_25267;
wire n_25268;
wire n_25272;
wire n_25275;
wire n_25276;
wire n_25277;
wire n_25279;
wire n_2528;
wire n_25280;
wire n_25281;
wire n_25282;
wire n_25284;
wire n_25285;
wire n_25286;
wire n_25287;
wire n_25288;
wire TIMEBOOST_net_2180;
wire n_25290;
wire n_25291;
wire n_25292;
wire TIMEBOOST_net_372;
wire n_25295;
wire n_253;
wire n_2530;
wire n_25301;
wire n_25302;
wire n_25303;
wire n_25304;
wire n_25306;
wire n_25307;
wire n_25308;
wire n_25309;
wire n_2531;
wire n_25310;
wire n_25311;
wire n_25312;
wire n_25316;
wire n_25318;
wire n_25319;
wire n_2532;
wire n_25320;
wire n_25321;
wire n_25323;
wire n_25327;
wire n_25328;
wire n_25329;
wire n_2533;
wire n_25331;
wire n_25333;
wire n_25334;
wire n_25335;
wire n_25336;
wire n_25337;
wire n_2534;
wire n_25340;
wire n_25341;
wire n_25342;
wire n_25343;
wire n_25344;
wire n_25345;
wire n_25346;
wire n_25347;
wire n_25348;
wire n_25349;
wire n_2535;
wire n_25350;
wire n_25351;
wire n_25352;
wire n_25353;
wire n_25354;
wire n_25355;
wire n_25356;
wire n_25357;
wire n_25358;
wire n_25359;
wire n_25361;
wire n_25363;
wire n_25365;
wire n_25366;
wire n_25368;
wire n_25369;
wire n_2537;
wire n_25370;
wire n_25371;
wire n_25372;
wire n_25373;
wire n_25375;
wire n_25377;
wire n_25378;
wire n_25379;
wire n_2538;
wire n_25380;
wire n_25381;
wire n_25382;
wire n_25383;
wire n_25385;
wire n_25386;
wire n_25388;
wire n_25389;
wire n_2539;
wire n_25390;
wire TIMEBOOST_net_1873;
wire n_25394;
wire n_25395;
wire n_25396;
wire n_25397;
wire n_25398;
wire n_25399;
wire n_254;
wire n_2540;
wire n_25401;
wire n_25403;
wire n_25404;
wire n_25405;
wire n_25407;
wire n_25408;
wire n_25409;
wire n_2541;
wire n_25410;
wire n_25412;
wire n_25413;
wire n_25414;
wire n_25415;
wire n_25416;
wire n_25418;
wire n_2542;
wire n_25421;
wire n_25422;
wire n_25424;
wire n_25425;
wire n_25426;
wire n_25427;
wire n_25428;
wire n_25429;
wire n_2543;
wire n_25430;
wire n_25431;
wire n_25432;
wire n_25433;
wire n_25436;
wire n_25437;
wire n_25438;
wire n_25439;
wire n_2544;
wire n_25440;
wire n_25441;
wire n_25444;
wire n_25445;
wire n_25446;
wire n_25447;
wire n_2545;
wire n_25451;
wire n_25452;
wire n_25453;
wire n_25454;
wire n_25455;
wire n_25457;
wire n_25458;
wire n_2546;
wire n_25460;
wire n_25461;
wire n_25462;
wire n_25463;
wire n_25464;
wire n_25465;
wire n_25466;
wire n_25467;
wire n_25468;
wire n_25469;
wire n_25470;
wire n_25471;
wire n_25472;
wire n_25473;
wire n_25476;
wire n_25477;
wire n_25478;
wire n_25479;
wire n_2548;
wire n_25482;
wire n_25485;
wire n_25486;
wire n_25487;
wire n_25488;
wire n_2549;
wire n_25493;
wire n_25494;
wire n_25495;
wire n_25499;
wire n_255;
wire n_2550;
wire n_25500;
wire n_25501;
wire n_25502;
wire n_25503;
wire n_25504;
wire n_25505;
wire n_25506;
wire n_25507;
wire n_25509;
wire n_2551;
wire n_25511;
wire n_25513;
wire n_25514;
wire n_25515;
wire n_25516;
wire n_25517;
wire n_25518;
wire n_25519;
wire n_25521;
wire n_25522;
wire n_25524;
wire n_25525;
wire n_25526;
wire n_25527;
wire n_25528;
wire n_25529;
wire n_25531;
wire n_25532;
wire n_25533;
wire n_25534;
wire n_25535;
wire n_25536;
wire n_25537;
wire n_25538;
wire n_2554;
wire n_25540;
wire n_25542;
wire n_25543;
wire n_25544;
wire n_25545;
wire n_25547;
wire n_25548;
wire TIMEBOOST_net_1138;
wire n_2555;
wire n_25551;
wire n_25552;
wire n_25553;
wire n_25554;
wire n_25555;
wire n_2556;
wire n_25561;
wire n_25562;
wire n_25564;
wire n_25565;
wire n_25567;
wire TIMEBOOST_net_2756;
wire n_25570;
wire n_25571;
wire n_25572;
wire n_25573;
wire n_25574;
wire n_25575;
wire n_25576;
wire n_25577;
wire n_25578;
wire n_25579;
wire n_2558;
wire n_25580;
wire n_25581;
wire n_25582;
wire n_25583;
wire n_25584;
wire n_25585;
wire n_25586;
wire n_25588;
wire n_25589;
wire n_2559;
wire n_25591;
wire TIMEBOOST_net_1233;
wire n_25593;
wire n_25594;
wire n_25595;
wire n_25598;
wire n_256;
wire n_25600;
wire n_25601;
wire n_25602;
wire n_25604;
wire n_25605;
wire n_25606;
wire n_25607;
wire n_25608;
wire n_2561;
wire n_25612;
wire n_25613;
wire n_25614;
wire n_25615;
wire n_25616;
wire n_25618;
wire n_25619;
wire n_2562;
wire n_25622;
wire n_25623;
wire n_25624;
wire n_25625;
wire n_25626;
wire n_25627;
wire n_25628;
wire n_25629;
wire n_2563;
wire n_25630;
wire n_25631;
wire n_25632;
wire n_25633;
wire n_25634;
wire n_25635;
wire n_25637;
wire n_25638;
wire n_25639;
wire n_25640;
wire n_25641;
wire n_25642;
wire n_25644;
wire n_25645;
wire n_25647;
wire n_25648;
wire n_2565;
wire n_25650;
wire n_25651;
wire TIMEBOOST_net_2516;
wire n_25653;
wire n_25654;
wire n_25655;
wire n_25656;
wire n_2566;
wire n_25660;
wire n_25661;
wire n_25662;
wire n_25667;
wire n_25668;
wire n_25669;
wire n_2567;
wire n_25670;
wire n_25671;
wire n_25672;
wire n_25673;
wire n_25675;
wire n_25676;
wire n_25677;
wire n_25678;
wire n_25679;
wire n_25680;
wire n_25683;
wire n_25684;
wire n_25685;
wire n_25686;
wire n_25687;
wire n_25688;
wire n_25689;
wire n_2569;
wire n_25690;
wire n_25691;
wire n_25692;
wire n_25693;
wire n_25694;
wire n_25695;
wire n_25696;
wire n_25697;
wire n_257;
wire n_2570;
wire n_25702;
wire n_25704;
wire TIMEBOOST_net_1160;
wire TIMEBOOST_net_375;
wire n_25707;
wire n_25708;
wire n_25709;
wire n_2571;
wire n_25710;
wire n_25711;
wire n_25712;
wire n_25713;
wire n_25714;
wire n_25715;
wire n_25716;
wire n_25717;
wire n_25718;
wire n_25719;
wire n_25720;
wire n_25721;
wire n_25722;
wire n_25723;
wire n_25724;
wire n_25725;
wire n_25726;
wire n_25727;
wire n_25729;
wire n_2573;
wire n_25730;
wire n_25731;
wire n_25732;
wire n_25733;
wire n_25734;
wire n_25735;
wire n_25736;
wire n_25738;
wire n_25739;
wire n_2574;
wire n_25740;
wire n_25741;
wire n_25743;
wire n_25744;
wire n_25745;
wire n_25746;
wire n_25747;
wire n_25748;
wire n_25749;
wire n_2575;
wire n_25750;
wire n_25751;
wire n_25753;
wire n_25757;
wire n_25758;
wire n_25759;
wire n_2576;
wire n_25760;
wire n_25761;
wire n_25762;
wire n_25763;
wire n_25764;
wire TIMEBOOST_net_1161;
wire n_2577;
wire n_25771;
wire n_25772;
wire n_25773;
wire n_25774;
wire n_25775;
wire n_25776;
wire n_25777;
wire TIMEBOOST_net_1189;
wire n_25781;
wire n_25782;
wire n_25783;
wire n_25785;
wire n_25786;
wire n_25788;
wire n_25789;
wire n_2579;
wire TIMEBOOST_net_2003;
wire n_25793;
wire n_25799;
wire n_258;
wire n_25800;
wire n_25801;
wire n_25802;
wire n_25803;
wire n_25804;
wire TIMEBOOST_net_1772;
wire n_25810;
wire n_25812;
wire n_25813;
wire n_25816;
wire n_25817;
wire n_25818;
wire n_25819;
wire n_2582;
wire n_25821;
wire n_25822;
wire n_25823;
wire n_25824;
wire n_25826;
wire n_25828;
wire n_25829;
wire n_2583;
wire TIMEBOOST_net_415;
wire n_25831;
wire n_25832;
wire n_25834;
wire n_25839;
wire n_2584;
wire n_25840;
wire n_25843;
wire n_25845;
wire n_25846;
wire n_25847;
wire n_25849;
wire n_25854;
wire n_25855;
wire n_25856;
wire n_25859;
wire TIMEBOOST_net_2891;
wire n_25867;
wire n_25868;
wire n_25869;
wire n_2587;
wire n_25870;
wire n_25874;
wire n_25875;
wire n_25876;
wire TIMEBOOST_net_1771;
wire n_2588;
wire n_25881;
wire n_25882;
wire n_25883;
wire n_25884;
wire n_25885;
wire n_25889;
wire n_2589;
wire n_25890;
wire n_25891;
wire n_25893;
wire TIMEBOOST_net_459;
wire n_25895;
wire n_25898;
wire n_259;
wire n_2590;
wire n_25900;
wire n_25902;
wire n_25903;
wire n_25904;
wire n_25905;
wire n_25906;
wire n_2591;
wire n_25911;
wire n_25912;
wire n_25914;
wire n_25915;
wire n_25916;
wire n_25917;
wire n_25918;
wire n_25919;
wire n_2592;
wire n_25920;
wire n_25922;
wire n_25923;
wire TIMEBOOST_net_1791;
wire n_25925;
wire n_25928;
wire n_2593;
wire n_25931;
wire n_25932;
wire n_25933;
wire n_25934;
wire n_25935;
wire n_25937;
wire n_25938;
wire n_25939;
wire n_2594;
wire n_25940;
wire TIMEBOOST_net_2283;
wire n_25947;
wire n_25948;
wire n_25949;
wire n_2595;
wire n_25950;
wire n_25951;
wire n_25952;
wire n_25953;
wire n_25954;
wire n_25955;
wire n_25956;
wire n_2596;
wire n_25962;
wire n_25963;
wire n_25964;
wire n_25966;
wire n_25967;
wire n_25968;
wire n_25969;
wire TIMEBOOST_net_2313;
wire n_25971;
wire n_25972;
wire n_25973;
wire n_25974;
wire n_25975;
wire n_25976;
wire n_25977;
wire n_25980;
wire n_25982;
wire n_25983;
wire n_25984;
wire n_25986;
wire TIMEBOOST_net_1668;
wire n_2599;
wire TIMEBOOST_net_2767;
wire TIMEBOOST_net_423;
wire n_25994;
wire n_25997;
wire n_25998;
wire n_25999;
wire n_260;
wire n_2600;
wire n_26000;
wire TIMEBOOST_net_2885;
wire n_26002;
wire n_26003;
wire n_26004;
wire n_26005;
wire n_26006;
wire n_26007;
wire n_26008;
wire n_26009;
wire n_2601;
wire n_26010;
wire n_26011;
wire n_26013;
wire n_26014;
wire n_26015;
wire n_26016;
wire n_26019;
wire n_2602;
wire n_26020;
wire n_26021;
wire n_26022;
wire TIMEBOOST_net_523;
wire n_26025;
wire n_26026;
wire n_26027;
wire n_26028;
wire n_26029;
wire n_2603;
wire TIMEBOOST_net_1209;
wire n_26032;
wire n_26033;
wire TIMEBOOST_net_433;
wire n_26036;
wire n_26037;
wire TIMEBOOST_net_425;
wire n_26039;
wire n_2604;
wire n_26040;
wire n_26041;
wire n_26042;
wire n_26044;
wire n_26045;
wire n_26048;
wire n_26049;
wire n_2605;
wire n_26051;
wire TIMEBOOST_net_1212;
wire n_26054;
wire n_26055;
wire TIMEBOOST_net_2488;
wire n_26057;
wire n_26058;
wire n_26059;
wire n_2606;
wire n_26060;
wire n_26061;
wire n_26062;
wire TIMEBOOST_net_1707;
wire TIMEBOOST_net_1706;
wire TIMEBOOST_net_1314;
wire n_26068;
wire n_26069;
wire n_2607;
wire TIMEBOOST_net_1299;
wire n_26072;
wire n_26073;
wire TIMEBOOST_net_1375;
wire n_26076;
wire n_26077;
wire n_26078;
wire n_26079;
wire n_2608;
wire n_26081;
wire n_26083;
wire n_26084;
wire n_26085;
wire n_26086;
wire n_26087;
wire n_26089;
wire n_2609;
wire n_26090;
wire n_26091;
wire n_26092;
wire TIMEBOOST_net_2085;
wire TIMEBOOST_net_1218;
wire n_26097;
wire n_26098;
wire n_261;
wire n_26100;
wire n_26101;
wire TIMEBOOST_net_1708;
wire n_26104;
wire n_26106;
wire n_26107;
wire n_2611;
wire n_26110;
wire n_26111;
wire n_26112;
wire n_26114;
wire n_26115;
wire n_26116;
wire TIMEBOOST_net_2916;
wire n_26118;
wire TIMEBOOST_net_1709;
wire n_2612;
wire n_26120;
wire n_26121;
wire TIMEBOOST_net_2705;
wire n_26124;
wire n_26125;
wire n_26128;
wire n_26129;
wire n_2613;
wire n_26130;
wire n_26131;
wire n_26132;
wire n_26133;
wire n_26134;
wire n_26135;
wire n_26136;
wire n_26137;
wire n_26138;
wire n_26139;
wire n_2614;
wire n_26140;
wire n_26142;
wire n_26143;
wire n_26144;
wire n_26146;
wire n_26147;
wire n_26149;
wire n_2615;
wire n_26150;
wire n_26152;
wire n_26153;
wire n_26154;
wire TIMEBOOST_net_427;
wire n_26156;
wire n_26157;
wire n_26158;
wire n_2616;
wire n_26160;
wire n_26161;
wire n_26162;
wire n_26163;
wire TIMEBOOST_net_1967;
wire TIMEBOOST_net_1222;
wire n_26167;
wire n_26169;
wire n_2617;
wire n_26171;
wire n_26173;
wire n_26174;
wire n_26175;
wire n_26176;
wire n_26178;
wire n_26179;
wire n_2618;
wire n_26180;
wire n_26181;
wire n_26184;
wire n_26185;
wire n_26186;
wire n_26188;
wire n_2619;
wire n_26190;
wire n_26191;
wire n_26192;
wire n_26193;
wire n_26194;
wire n_26195;
wire n_26196;
wire n_26198;
wire n_262;
wire n_2620;
wire n_26200;
wire n_26201;
wire n_26202;
wire n_26204;
wire TIMEBOOST_net_462;
wire n_26206;
wire n_26207;
wire n_26208;
wire TIMEBOOST_net_272;
wire TIMEBOOST_net_2704;
wire n_26212;
wire n_26213;
wire n_26214;
wire n_26215;
wire n_26216;
wire n_26217;
wire n_26218;
wire n_26219;
wire n_2622;
wire n_26220;
wire n_26221;
wire n_26222;
wire TIMEBOOST_net_1315;
wire n_26224;
wire n_26225;
wire n_26226;
wire n_26227;
wire n_26228;
wire n_2623;
wire n_26230;
wire n_26232;
wire n_26233;
wire n_26234;
wire n_26235;
wire n_26236;
wire n_26237;
wire n_26238;
wire n_26239;
wire n_2624;
wire n_26240;
wire n_26245;
wire n_26246;
wire n_26247;
wire n_26248;
wire n_26249;
wire n_2625;
wire n_26250;
wire n_26251;
wire n_26252;
wire n_26253;
wire n_26254;
wire n_26258;
wire n_2626;
wire TIMEBOOST_net_1319;
wire n_26262;
wire n_26263;
wire n_26264;
wire n_26265;
wire n_26266;
wire n_26267;
wire TIMEBOOST_net_2624;
wire n_2627;
wire n_26271;
wire n_26272;
wire n_26276;
wire n_26277;
wire n_26278;
wire n_26279;
wire n_2628;
wire TIMEBOOST_net_1193;
wire n_26283;
wire TIMEBOOST_net_1807;
wire n_2629;
wire n_26290;
wire n_26291;
wire n_26292;
wire n_26293;
wire n_26294;
wire n_26295;
wire n_26296;
wire n_26297;
wire n_26298;
wire n_26299;
wire n_263;
wire n_2630;
wire n_26300;
wire n_26301;
wire n_26302;
wire n_26303;
wire n_26304;
wire n_26306;
wire n_26307;
wire n_26308;
wire n_2631;
wire n_26310;
wire n_26311;
wire n_26312;
wire n_26313;
wire n_26314;
wire n_26316;
wire n_26318;
wire n_26319;
wire n_26320;
wire n_26322;
wire n_26323;
wire n_26324;
wire n_26325;
wire n_26326;
wire n_26327;
wire n_26328;
wire n_26329;
wire n_2633;
wire n_26330;
wire n_26331;
wire n_26332;
wire n_26333;
wire TIMEBOOST_net_1718;
wire n_26335;
wire TIMEBOOST_net_1225;
wire n_26337;
wire n_26338;
wire n_2634;
wire n_26340;
wire n_26343;
wire n_26345;
wire n_26346;
wire n_26348;
wire n_26349;
wire n_2635;
wire n_26350;
wire n_26351;
wire n_26352;
wire TIMEBOOST_net_2217;
wire n_26354;
wire n_26355;
wire n_26358;
wire n_26359;
wire n_2636;
wire n_26360;
wire n_26361;
wire n_26362;
wire n_26363;
wire n_26364;
wire n_26365;
wire n_26366;
wire n_26367;
wire n_26368;
wire n_26369;
wire n_2637;
wire n_26370;
wire n_26371;
wire n_26372;
wire n_26373;
wire n_26374;
wire TIMEBOOST_net_1378;
wire n_26376;
wire n_26377;
wire n_26378;
wire TIMEBOOST_net_1364;
wire n_2638;
wire n_26381;
wire n_26382;
wire n_26383;
wire n_26384;
wire n_26385;
wire n_26386;
wire n_26387;
wire n_26389;
wire n_2639;
wire n_26390;
wire n_26392;
wire n_26393;
wire n_26394;
wire TIMEBOOST_net_472;
wire n_26398;
wire n_26399;
wire n_264;
wire n_2640;
wire n_26400;
wire n_26401;
wire n_26403;
wire n_26406;
wire n_26407;
wire n_26409;
wire n_2641;
wire n_26410;
wire TIMEBOOST_net_2931;
wire n_26412;
wire n_26413;
wire n_26414;
wire n_26415;
wire n_26416;
wire n_26417;
wire n_26418;
wire n_26419;
wire n_2642;
wire n_26420;
wire n_26421;
wire n_26422;
wire n_26424;
wire n_26425;
wire n_26426;
wire n_26427;
wire n_26428;
wire n_26429;
wire n_2643;
wire n_26434;
wire TIMEBOOST_net_1808;
wire n_26437;
wire n_26439;
wire n_2644;
wire n_26440;
wire n_26442;
wire n_26444;
wire n_26445;
wire n_26447;
wire n_26448;
wire TIMEBOOST_net_532;
wire n_26451;
wire n_26452;
wire n_26453;
wire n_26454;
wire n_26456;
wire n_26458;
wire n_2646;
wire n_26461;
wire n_26462;
wire n_26463;
wire n_26464;
wire n_26465;
wire n_26466;
wire n_26467;
wire n_26468;
wire n_26469;
wire n_2647;
wire n_26471;
wire n_26472;
wire n_26473;
wire n_26477;
wire n_26478;
wire n_26479;
wire n_26480;
wire n_26484;
wire n_26486;
wire n_26487;
wire n_2649;
wire n_26491;
wire n_26493;
wire n_26494;
wire n_26495;
wire n_26496;
wire n_26497;
wire n_26498;
wire n_265;
wire n_2650;
wire n_26500;
wire n_26501;
wire n_26502;
wire n_26503;
wire n_26504;
wire n_26506;
wire n_26507;
wire n_26508;
wire n_26509;
wire n_2651;
wire n_26510;
wire TIMEBOOST_net_440;
wire n_26512;
wire TIMEBOOST_net_2934;
wire n_26514;
wire n_26516;
wire n_26518;
wire n_26519;
wire n_2652;
wire n_26520;
wire n_26521;
wire n_26522;
wire n_26524;
wire n_26525;
wire n_26526;
wire n_26527;
wire n_26528;
wire n_26529;
wire n_26530;
wire n_26531;
wire n_26532;
wire n_26533;
wire n_26536;
wire n_26537;
wire TIMEBOOST_net_1120;
wire n_26539;
wire n_2654;
wire n_26540;
wire n_26541;
wire n_26542;
wire n_26544;
wire n_26546;
wire n_26547;
wire n_26548;
wire n_26549;
wire n_2655;
wire n_26550;
wire n_26551;
wire n_26552;
wire n_26553;
wire n_26555;
wire n_26557;
wire n_26558;
wire n_26559;
wire n_2656;
wire n_26560;
wire n_26563;
wire n_26564;
wire n_26566;
wire n_2657;
wire n_26571;
wire n_26572;
wire n_26573;
wire n_26574;
wire n_26575;
wire TIMEBOOST_net_2887;
wire TIMEBOOST_net_1805;
wire n_26579;
wire n_2658;
wire n_26580;
wire n_26581;
wire n_26582;
wire n_26583;
wire n_26584;
wire n_26586;
wire n_26587;
wire n_26588;
wire n_26589;
wire n_26590;
wire n_26592;
wire n_26594;
wire n_26595;
wire n_26596;
wire n_26597;
wire n_26599;
wire n_266;
wire n_2660;
wire n_26601;
wire n_26602;
wire n_26604;
wire n_26605;
wire n_26606;
wire TIMEBOOST_net_2906;
wire n_26608;
wire n_26609;
wire n_2661;
wire n_26610;
wire n_26611;
wire n_26612;
wire n_26613;
wire n_26614;
wire n_26615;
wire n_26616;
wire n_26617;
wire n_26620;
wire n_26622;
wire n_26623;
wire n_26624;
wire n_26625;
wire n_26626;
wire n_26627;
wire n_26628;
wire n_26629;
wire n_2663;
wire n_26630;
wire n_26633;
wire n_26634;
wire n_26636;
wire n_26637;
wire n_26638;
wire n_26639;
wire n_2664;
wire n_26640;
wire n_26641;
wire n_26642;
wire n_26643;
wire n_26644;
wire n_26645;
wire n_26646;
wire n_26647;
wire n_26648;
wire n_2665;
wire n_26652;
wire n_26653;
wire n_26654;
wire n_26655;
wire n_26656;
wire n_26657;
wire n_26658;
wire n_26659;
wire n_2666;
wire n_26660;
wire n_26661;
wire n_26663;
wire n_26664;
wire TIMEBOOST_net_1323;
wire n_26666;
wire n_26668;
wire n_26669;
wire n_2667;
wire n_26670;
wire n_26671;
wire n_26672;
wire n_26673;
wire n_26674;
wire n_26675;
wire n_26677;
wire n_26679;
wire n_2668;
wire n_26680;
wire n_26681;
wire n_26682;
wire n_26683;
wire n_26684;
wire n_26685;
wire n_26686;
wire n_26687;
wire n_26688;
wire n_26689;
wire n_26690;
wire n_26691;
wire n_26692;
wire n_26693;
wire n_26694;
wire n_26695;
wire n_26696;
wire n_26697;
wire n_26698;
wire n_26699;
wire n_267;
wire n_26700;
wire n_26701;
wire n_26702;
wire n_26703;
wire n_26704;
wire n_26705;
wire n_26707;
wire n_26708;
wire n_26709;
wire n_26710;
wire n_26711;
wire n_26712;
wire n_26713;
wire n_26714;
wire n_26715;
wire n_26716;
wire TIMEBOOST_net_2670;
wire n_26718;
wire n_26719;
wire n_2672;
wire TIMEBOOST_net_534;
wire n_26721;
wire n_26722;
wire n_26723;
wire n_26724;
wire n_26725;
wire n_26726;
wire n_26729;
wire n_2673;
wire TIMEBOOST_net_1379;
wire n_26731;
wire n_26732;
wire n_26734;
wire n_26736;
wire n_26737;
wire n_26738;
wire n_26739;
wire n_2674;
wire n_26740;
wire n_26741;
wire n_26742;
wire n_26743;
wire n_26744;
wire n_26745;
wire n_26747;
wire n_26748;
wire n_26749;
wire n_2675;
wire n_26750;
wire n_26751;
wire n_26752;
wire n_26753;
wire n_26754;
wire n_26755;
wire n_26756;
wire TIMEBOOST_net_1369;
wire n_26758;
wire n_26759;
wire n_26761;
wire n_26762;
wire n_26763;
wire n_26764;
wire n_26765;
wire n_26766;
wire n_26767;
wire n_26768;
wire n_26769;
wire TIMEBOOST_net_2892;
wire n_26770;
wire n_26771;
wire n_26772;
wire n_26773;
wire n_26774;
wire n_26775;
wire n_26776;
wire n_26777;
wire n_26778;
wire TIMEBOOST_net_1059;
wire TIMEBOOST_net_2779;
wire n_26781;
wire n_26783;
wire n_26784;
wire n_26785;
wire n_26786;
wire n_26787;
wire n_26788;
wire n_2679;
wire n_26790;
wire n_26791;
wire n_26792;
wire n_26793;
wire n_26794;
wire n_26795;
wire n_26796;
wire n_26797;
wire n_26799;
wire n_268;
wire n_2680;
wire TIMEBOOST_net_607;
wire n_26801;
wire n_26802;
wire n_26804;
wire n_26805;
wire TIMEBOOST_net_1380;
wire n_26807;
wire n_26808;
wire n_26809;
wire n_2681;
wire n_26810;
wire n_26812;
wire n_26813;
wire n_26814;
wire n_26815;
wire n_26816;
wire n_26817;
wire TIMEBOOST_net_2923;
wire n_26819;
wire n_2682;
wire n_26820;
wire n_26821;
wire n_26822;
wire n_26823;
wire n_26824;
wire n_26826;
wire n_26827;
wire n_26828;
wire n_26829;
wire n_2683;
wire n_26830;
wire n_26831;
wire n_26832;
wire n_26833;
wire n_26834;
wire n_26835;
wire n_26836;
wire n_26837;
wire n_26838;
wire n_26839;
wire n_2684;
wire n_26840;
wire n_26844;
wire n_26846;
wire n_26847;
wire n_26848;
wire n_26849;
wire n_2685;
wire n_26850;
wire n_26851;
wire n_26852;
wire n_26853;
wire n_26855;
wire n_2686;
wire n_26860;
wire n_26861;
wire n_26862;
wire n_26863;
wire n_26864;
wire n_26865;
wire n_26866;
wire n_26868;
wire n_26869;
wire n_2687;
wire n_26870;
wire n_26871;
wire n_26872;
wire n_26873;
wire n_26874;
wire n_26875;
wire n_26876;
wire n_26877;
wire n_26878;
wire n_26879;
wire n_2688;
wire n_26880;
wire n_26881;
wire n_26882;
wire n_26883;
wire n_26884;
wire n_26885;
wire n_26886;
wire n_26887;
wire n_26888;
wire n_26889;
wire n_2689;
wire n_26890;
wire n_26891;
wire n_26892;
wire n_26893;
wire n_26894;
wire n_26895;
wire n_26896;
wire n_26897;
wire n_26898;
wire n_26899;
wire n_269;
wire n_2690;
wire n_26900;
wire n_26901;
wire n_26902;
wire n_26903;
wire n_26904;
wire n_26905;
wire n_26906;
wire n_26907;
wire n_26908;
wire n_26909;
wire n_2691;
wire n_26910;
wire n_26911;
wire n_26912;
wire n_26913;
wire n_26914;
wire n_26915;
wire n_26916;
wire TIMEBOOST_net_2778;
wire n_26918;
wire n_26919;
wire n_2692;
wire n_26920;
wire n_26922;
wire n_26924;
wire n_26925;
wire n_26926;
wire n_26927;
wire n_26928;
wire n_26929;
wire n_2693;
wire n_26930;
wire n_26931;
wire n_26932;
wire n_26933;
wire n_26934;
wire n_26935;
wire n_26936;
wire n_26937;
wire n_26938;
wire n_26939;
wire n_2694;
wire n_26940;
wire n_26941;
wire n_26942;
wire n_26943;
wire n_26944;
wire n_26945;
wire n_26946;
wire n_26947;
wire n_26948;
wire n_26949;
wire n_2695;
wire n_26950;
wire n_26951;
wire n_26952;
wire n_26953;
wire n_26954;
wire n_26955;
wire n_26956;
wire n_26957;
wire n_26958;
wire n_26960;
wire n_26961;
wire n_26962;
wire n_26963;
wire TIMEBOOST_net_2317;
wire n_26966;
wire n_26967;
wire n_26968;
wire n_26969;
wire n_2697;
wire n_26970;
wire n_26971;
wire n_26972;
wire n_26973;
wire n_26974;
wire TIMEBOOST_net_1365;
wire n_26976;
wire n_26977;
wire n_26978;
wire TIMEBOOST_net_1331;
wire n_2698;
wire n_26980;
wire n_26981;
wire n_26982;
wire n_26983;
wire n_26984;
wire n_26985;
wire TIMEBOOST_net_680;
wire n_26987;
wire n_26988;
wire n_26989;
wire n_2699;
wire n_26990;
wire n_26991;
wire n_26992;
wire n_26993;
wire n_26996;
wire n_26997;
wire n_26998;
wire n_26999;
wire n_27;
wire n_270;
wire n_2700;
wire n_27000;
wire n_27001;
wire n_27002;
wire TIMEBOOST_net_1581;
wire n_27004;
wire n_27005;
wire n_27006;
wire n_27007;
wire n_27008;
wire n_27009;
wire n_2701;
wire n_27010;
wire n_27011;
wire n_27012;
wire n_27013;
wire n_27014;
wire n_27015;
wire n_27016;
wire n_27017;
wire n_27018;
wire n_27019;
wire n_2702;
wire n_27020;
wire n_27021;
wire n_27022;
wire n_27023;
wire n_27024;
wire n_27025;
wire n_27026;
wire n_27027;
wire n_27028;
wire n_27029;
wire n_27031;
wire n_27032;
wire n_27033;
wire n_27034;
wire n_27035;
wire n_27036;
wire n_27037;
wire n_27038;
wire n_27039;
wire n_2704;
wire n_27040;
wire n_27041;
wire n_27042;
wire n_27043;
wire n_27044;
wire n_27045;
wire n_27046;
wire n_27047;
wire n_2705;
wire n_27050;
wire n_27051;
wire TIMEBOOST_net_1366;
wire TIMEBOOST_net_1333;
wire n_27055;
wire n_27057;
wire n_27058;
wire n_27059;
wire n_2706;
wire n_27062;
wire n_27063;
wire n_27064;
wire TIMEBOOST_net_659;
wire TIMEBOOST_net_606;
wire n_27067;
wire n_27068;
wire n_27070;
wire n_27071;
wire n_27072;
wire n_27073;
wire n_27075;
wire n_27076;
wire n_27077;
wire n_27079;
wire n_27080;
wire n_27081;
wire n_27082;
wire n_27083;
wire n_27086;
wire n_27088;
wire n_27089;
wire n_2709;
wire n_27090;
wire n_27092;
wire n_27093;
wire n_27094;
wire n_27095;
wire n_27096;
wire n_27097;
wire n_27098;
wire n_27099;
wire n_271;
wire n_2710;
wire n_27100;
wire n_27101;
wire n_27102;
wire n_27103;
wire n_27104;
wire n_27107;
wire n_27108;
wire n_27109;
wire n_2711;
wire n_27110;
wire n_27113;
wire n_27117;
wire n_27119;
wire n_2712;
wire n_27120;
wire n_27121;
wire n_27123;
wire n_27124;
wire n_27125;
wire n_27126;
wire n_27127;
wire n_27128;
wire n_27129;
wire n_27130;
wire n_27131;
wire n_27132;
wire n_27133;
wire n_27134;
wire n_27135;
wire n_2714;
wire TIMEBOOST_net_699;
wire n_27143;
wire n_27144;
wire n_27145;
wire n_27146;
wire n_2715;
wire n_27150;
wire n_27151;
wire n_27152;
wire n_27153;
wire TIMEBOOST_net_2819;
wire TIMEBOOST_net_2845;
wire n_27157;
wire n_27158;
wire n_27159;
wire n_2716;
wire n_27160;
wire n_27161;
wire n_27164;
wire n_27165;
wire n_27167;
wire n_27168;
wire n_2717;
wire n_27170;
wire n_27172;
wire n_27173;
wire n_27175;
wire n_27178;
wire n_2718;
wire n_27183;
wire n_27184;
wire TIMEBOOST_net_2117;
wire n_27188;
wire n_27189;
wire n_2719;
wire n_27190;
wire n_27191;
wire n_27192;
wire n_27193;
wire n_27194;
wire n_27198;
wire n_27199;
wire n_272;
wire n_2720;
wire n_27200;
wire n_27201;
wire n_27202;
wire n_27203;
wire n_27204;
wire n_27206;
wire n_27207;
wire n_27208;
wire n_27210;
wire n_27211;
wire n_27213;
wire n_27214;
wire n_27215;
wire n_27216;
wire n_27217;
wire n_27218;
wire n_27219;
wire n_2722;
wire n_27222;
wire n_27223;
wire n_27224;
wire n_27225;
wire n_27226;
wire n_27227;
wire n_27229;
wire n_27230;
wire n_27232;
wire n_27233;
wire n_27234;
wire TIMEBOOST_net_2734;
wire n_27237;
wire n_27238;
wire n_27239;
wire n_2724;
wire n_27240;
wire n_27241;
wire n_27242;
wire n_27243;
wire n_27244;
wire n_27245;
wire n_27246;
wire n_27247;
wire n_2725;
wire n_27250;
wire n_27254;
wire n_27256;
wire n_2726;
wire n_27263;
wire n_27264;
wire TIMEBOOST_net_2106;
wire n_27267;
wire n_27268;
wire n_27269;
wire n_27270;
wire n_27271;
wire n_27272;
wire n_27273;
wire n_27274;
wire n_27276;
wire n_27277;
wire n_27278;
wire n_27279;
wire n_2728;
wire n_27283;
wire n_27284;
wire n_27285;
wire n_2729;
wire n_27291;
wire n_27292;
wire n_27294;
wire n_27295;
wire n_27296;
wire n_27297;
wire n_27298;
wire n_27299;
wire n_273;
wire n_2730;
wire n_27300;
wire n_27301;
wire n_27302;
wire n_27303;
wire n_27304;
wire n_27305;
wire n_27306;
wire n_27307;
wire n_27308;
wire n_27309;
wire n_2731;
wire n_27310;
wire n_27312;
wire n_27313;
wire n_27314;
wire n_27315;
wire n_27318;
wire n_27319;
wire n_2732;
wire n_27320;
wire n_27321;
wire n_27322;
wire n_27323;
wire n_27326;
wire TIMEBOOST_net_2095;
wire n_27329;
wire n_2733;
wire TIMEBOOST_net_714;
wire n_27334;
wire n_27336;
wire n_27337;
wire n_27338;
wire n_27339;
wire n_2734;
wire n_27340;
wire n_27342;
wire n_27343;
wire TIMEBOOST_net_1479;
wire TIMEBOOST_net_2791;
wire n_27347;
wire n_27348;
wire n_27349;
wire n_2735;
wire n_27351;
wire n_27352;
wire n_27353;
wire n_27354;
wire n_27355;
wire n_27356;
wire n_27357;
wire n_27358;
wire n_27359;
wire n_2736;
wire n_27360;
wire n_27361;
wire n_27362;
wire n_27363;
wire n_27364;
wire n_27365;
wire n_27366;
wire n_27367;
wire n_27368;
wire n_27371;
wire n_27373;
wire n_27375;
wire n_27376;
wire n_27378;
wire n_2738;
wire n_27380;
wire n_27381;
wire n_27382;
wire n_27383;
wire n_27384;
wire n_27386;
wire n_27387;
wire n_27388;
wire n_2739;
wire n_27390;
wire n_27391;
wire n_27392;
wire n_27393;
wire n_27394;
wire n_27395;
wire n_27396;
wire n_27397;
wire n_27398;
wire n_27399;
wire n_274;
wire n_2740;
wire n_27400;
wire n_27401;
wire n_27402;
wire n_27403;
wire n_27404;
wire n_27406;
wire TIMEBOOST_net_1815;
wire n_27410;
wire n_27411;
wire n_27413;
wire n_27414;
wire n_27415;
wire n_27416;
wire n_27418;
wire n_2742;
wire n_27420;
wire n_27421;
wire n_27422;
wire n_27423;
wire n_27424;
wire n_27425;
wire n_27426;
wire n_27427;
wire n_27428;
wire n_27429;
wire n_2743;
wire n_27430;
wire TIMEBOOST_net_1393;
wire n_27433;
wire n_27434;
wire n_27436;
wire n_27437;
wire n_27438;
wire n_27439;
wire n_2744;
wire n_27440;
wire n_27441;
wire n_27442;
wire n_27443;
wire n_27447;
wire n_27448;
wire n_27449;
wire n_2745;
wire n_27450;
wire n_27451;
wire n_27452;
wire n_27453;
wire n_27454;
wire n_27455;
wire n_27456;
wire n_27457;
wire n_27458;
wire n_27459;
wire n_2746;
wire n_27460;
wire n_27461;
wire n_27462;
wire n_27463;
wire n_27464;
wire n_27465;
wire n_27466;
wire n_27467;
wire n_27468;
wire n_27469;
wire n_2747;
wire n_27470;
wire n_27471;
wire n_27472;
wire n_27473;
wire n_27476;
wire n_27479;
wire n_2748;
wire n_27480;
wire n_27481;
wire n_27482;
wire n_27483;
wire n_27484;
wire n_27485;
wire n_27486;
wire n_27487;
wire n_27488;
wire n_27489;
wire n_2749;
wire n_27490;
wire n_27491;
wire n_27492;
wire n_27493;
wire n_27494;
wire n_27496;
wire n_27497;
wire n_27498;
wire n_27499;
wire n_275;
wire n_2750;
wire n_27500;
wire n_27501;
wire n_27502;
wire n_27503;
wire n_27504;
wire n_27506;
wire n_27507;
wire n_27509;
wire n_2751;
wire n_27510;
wire n_27511;
wire n_27512;
wire n_27513;
wire n_27514;
wire n_27518;
wire n_27519;
wire n_2752;
wire n_27520;
wire n_27521;
wire n_27522;
wire n_27523;
wire n_27524;
wire n_27525;
wire n_27526;
wire n_27527;
wire n_27528;
wire n_27529;
wire n_2753;
wire n_27531;
wire n_27532;
wire n_27533;
wire n_27534;
wire n_27535;
wire n_27536;
wire n_27537;
wire n_27538;
wire n_27539;
wire n_2754;
wire n_27540;
wire TIMEBOOST_net_616;
wire n_27542;
wire n_27543;
wire n_27544;
wire n_27545;
wire n_27546;
wire n_27547;
wire n_27548;
wire n_27549;
wire n_2755;
wire n_27550;
wire n_27551;
wire n_27554;
wire n_27555;
wire n_27559;
wire n_2756;
wire n_27560;
wire n_27561;
wire n_27565;
wire n_27566;
wire n_27567;
wire n_27568;
wire n_27569;
wire n_27570;
wire n_27571;
wire n_27572;
wire n_27573;
wire n_27574;
wire n_27575;
wire n_27576;
wire n_27578;
wire n_27579;
wire n_2758;
wire n_27580;
wire n_27582;
wire n_27584;
wire n_27585;
wire n_27586;
wire n_27587;
wire n_27588;
wire n_27589;
wire n_27590;
wire n_27593;
wire n_27595;
wire TIMEBOOST_net_1518;
wire n_27598;
wire n_27599;
wire n_276;
wire n_2760;
wire n_27600;
wire n_27601;
wire n_27602;
wire n_27603;
wire n_27604;
wire n_27605;
wire n_27607;
wire n_27608;
wire TIMEBOOST_net_2182;
wire n_2761;
wire n_27610;
wire n_27611;
wire n_27612;
wire n_27613;
wire n_27614;
wire n_27615;
wire n_27617;
wire TIMEBOOST_net_756;
wire n_27619;
wire n_27620;
wire n_27621;
wire n_27622;
wire n_27623;
wire n_27624;
wire n_27625;
wire n_27626;
wire n_27627;
wire n_2763;
wire n_27632;
wire n_27634;
wire n_27635;
wire n_27637;
wire TIMEBOOST_net_2173;
wire n_27639;
wire n_2764;
wire n_27641;
wire n_27642;
wire n_27643;
wire n_27644;
wire n_27645;
wire n_27646;
wire n_27648;
wire n_27649;
wire n_27652;
wire n_27653;
wire n_27654;
wire n_27655;
wire n_27656;
wire n_27657;
wire n_27659;
wire n_2766;
wire n_27661;
wire n_27662;
wire n_27665;
wire n_27666;
wire n_27667;
wire n_27668;
wire n_27669;
wire n_27670;
wire n_27671;
wire n_27672;
wire n_27673;
wire n_27674;
wire n_27675;
wire n_27676;
wire n_27677;
wire n_27678;
wire n_2768;
wire n_27681;
wire n_27682;
wire n_27683;
wire n_27684;
wire TIMEBOOST_net_759;
wire n_27686;
wire n_27687;
wire n_27688;
wire n_2769;
wire n_27690;
wire n_27691;
wire n_27692;
wire n_27693;
wire n_27695;
wire n_27696;
wire n_27697;
wire n_27698;
wire n_277;
wire n_2770;
wire n_27700;
wire n_27701;
wire n_27702;
wire n_27703;
wire n_27705;
wire n_27706;
wire n_27708;
wire n_27709;
wire n_2771;
wire n_27710;
wire n_27711;
wire n_27712;
wire n_27714;
wire n_27715;
wire n_27717;
wire n_27719;
wire TIMEBOOST_net_2625;
wire n_27720;
wire n_27721;
wire n_27723;
wire n_27725;
wire n_27726;
wire n_27727;
wire n_27728;
wire n_27729;
wire n_27730;
wire n_27731;
wire n_27732;
wire n_27733;
wire n_27736;
wire n_27737;
wire n_27738;
wire n_27739;
wire n_2774;
wire n_27741;
wire n_27743;
wire n_27744;
wire n_27745;
wire n_27748;
wire n_27749;
wire n_2775;
wire n_27750;
wire n_27751;
wire n_27752;
wire n_27755;
wire n_27756;
wire n_27757;
wire n_27758;
wire n_27762;
wire n_27763;
wire n_27764;
wire n_27765;
wire n_27766;
wire n_27767;
wire n_27768;
wire n_2777;
wire n_27771;
wire n_27772;
wire n_27773;
wire n_27776;
wire TIMEBOOST_net_2841;
wire n_27778;
wire n_27779;
wire n_2778;
wire n_27780;
wire n_27781;
wire n_27782;
wire n_27783;
wire n_27784;
wire n_27785;
wire n_27787;
wire n_27788;
wire n_27789;
wire n_27790;
wire n_27791;
wire n_27792;
wire n_27794;
wire n_27795;
wire n_27796;
wire n_27797;
wire n_27799;
wire n_278;
wire n_27800;
wire n_27802;
wire n_27803;
wire n_27804;
wire n_27805;
wire n_27806;
wire n_27807;
wire n_27810;
wire n_27812;
wire n_27813;
wire n_27814;
wire n_27815;
wire n_27818;
wire n_27819;
wire n_2782;
wire n_27822;
wire n_27823;
wire n_27824;
wire n_27825;
wire n_27827;
wire n_27830;
wire n_27831;
wire n_27832;
wire n_27833;
wire n_27834;
wire n_27835;
wire n_27836;
wire n_27838;
wire n_27839;
wire n_2784;
wire n_27843;
wire n_27844;
wire n_27845;
wire n_27846;
wire n_27848;
wire n_2785;
wire n_27851;
wire n_27852;
wire n_27853;
wire n_27854;
wire n_27855;
wire n_27858;
wire n_27859;
wire n_2786;
wire n_27860;
wire n_27862;
wire n_27863;
wire n_27864;
wire n_27865;
wire n_27868;
wire n_27869;
wire n_2787;
wire n_27871;
wire n_27872;
wire n_27875;
wire n_27876;
wire n_27877;
wire n_27878;
wire n_27879;
wire n_27880;
wire n_27881;
wire n_27882;
wire n_27883;
wire n_27884;
wire n_27885;
wire n_27887;
wire n_27888;
wire n_27889;
wire n_2789;
wire TIMEBOOST_net_2134;
wire n_27893;
wire n_27894;
wire n_27895;
wire n_27896;
wire n_27899;
wire n_279;
wire n_2790;
wire n_27901;
wire n_27902;
wire n_27903;
wire n_27905;
wire n_27906;
wire n_27907;
wire n_27908;
wire n_27909;
wire n_2791;
wire n_27910;
wire n_27911;
wire n_27912;
wire n_27914;
wire n_27916;
wire n_27917;
wire n_27918;
wire n_27919;
wire n_2792;
wire n_27920;
wire n_27921;
wire n_27922;
wire n_27923;
wire n_27926;
wire n_27928;
wire n_27929;
wire n_2793;
wire n_27931;
wire n_27932;
wire n_27933;
wire n_27934;
wire n_27936;
wire n_27937;
wire n_27938;
wire n_27939;
wire n_2794;
wire n_27940;
wire n_27941;
wire n_27944;
wire n_27948;
wire n_27949;
wire n_2795;
wire n_27950;
wire n_27951;
wire n_27953;
wire n_27954;
wire n_27955;
wire n_27956;
wire n_27957;
wire n_27958;
wire n_27959;
wire n_2796;
wire n_27960;
wire n_27961;
wire n_27962;
wire n_27964;
wire n_27965;
wire n_27966;
wire n_27968;
wire n_2797;
wire n_27970;
wire n_27971;
wire n_27972;
wire n_27973;
wire TIMEBOOST_net_1629;
wire n_27976;
wire n_2798;
wire n_27986;
wire n_27987;
wire n_27988;
wire n_2799;
wire n_27990;
wire n_27991;
wire n_27992;
wire n_27993;
wire n_27994;
wire n_27995;
wire n_27997;
wire n_27998;
wire n_27999;
wire n_280;
wire n_28001;
wire n_28002;
wire n_28003;
wire TIMEBOOST_net_1466;
wire n_28005;
wire n_28006;
wire n_28008;
wire n_28009;
wire n_28010;
wire n_28011;
wire n_28012;
wire n_28014;
wire n_28015;
wire n_28016;
wire n_28018;
wire n_2802;
wire n_28021;
wire n_28022;
wire n_28023;
wire n_28024;
wire n_28025;
wire n_28027;
wire n_28028;
wire n_28029;
wire n_2803;
wire n_28030;
wire n_28031;
wire n_28032;
wire n_28034;
wire n_28035;
wire n_28036;
wire n_28037;
wire n_28038;
wire n_28039;
wire n_28040;
wire n_28041;
wire n_28042;
wire n_28043;
wire n_28044;
wire n_2805;
wire n_28050;
wire n_28051;
wire n_28052;
wire n_28053;
wire n_28054;
wire n_28055;
wire n_28056;
wire n_28057;
wire n_28058;
wire n_28059;
wire TIMEBOOST_net_2838;
wire n_28060;
wire n_28061;
wire n_28062;
wire n_28063;
wire n_28064;
wire n_28065;
wire n_28066;
wire n_28067;
wire n_28068;
wire n_2807;
wire n_28070;
wire n_28071;
wire n_28072;
wire n_28075;
wire n_28076;
wire n_28077;
wire n_28078;
wire n_28079;
wire n_2808;
wire n_28080;
wire n_28082;
wire n_28083;
wire n_28084;
wire n_28085;
wire n_28086;
wire n_28088;
wire n_28089;
wire n_2809;
wire n_28090;
wire n_28091;
wire n_28092;
wire n_28093;
wire n_28094;
wire n_28096;
wire n_28097;
wire n_28098;
wire n_28099;
wire n_281;
wire n_2810;
wire n_28100;
wire TIMEBOOST_net_874;
wire n_28102;
wire n_28105;
wire n_28106;
wire n_28107;
wire n_28108;
wire n_28109;
wire n_28112;
wire n_28113;
wire n_28114;
wire n_28115;
wire n_28116;
wire n_28117;
wire n_28118;
wire n_28119;
wire n_28120;
wire n_28121;
wire n_28122;
wire n_28123;
wire n_28124;
wire n_28125;
wire TIMEBOOST_net_2824;
wire n_28128;
wire n_28129;
wire n_2813;
wire n_28130;
wire n_28131;
wire n_28132;
wire n_28134;
wire n_28135;
wire n_28136;
wire n_28137;
wire n_28138;
wire n_28139;
wire n_2814;
wire n_28140;
wire n_28142;
wire n_28143;
wire TIMEBOOST_net_1478;
wire n_28146;
wire n_28147;
wire n_28148;
wire n_28149;
wire n_28150;
wire n_28152;
wire n_28154;
wire n_28156;
wire n_28157;
wire n_28158;
wire n_28159;
wire n_2816;
wire n_28160;
wire n_28161;
wire n_28162;
wire n_28163;
wire n_28164;
wire n_28165;
wire n_28166;
wire TIMEBOOST_net_2788;
wire n_2817;
wire n_28173;
wire n_28174;
wire n_28175;
wire n_28176;
wire n_28177;
wire n_28179;
wire n_2818;
wire n_28180;
wire n_28181;
wire n_28182;
wire n_28183;
wire n_28186;
wire n_28187;
wire n_28188;
wire n_28189;
wire n_2819;
wire n_28190;
wire n_28191;
wire n_28192;
wire n_28195;
wire n_28196;
wire n_28198;
wire n_28199;
wire n_282;
wire n_2820;
wire n_28200;
wire n_28201;
wire n_28202;
wire n_28203;
wire n_28204;
wire n_28205;
wire TIMEBOOST_net_2875;
wire n_28207;
wire n_28208;
wire n_28209;
wire n_2821;
wire n_28210;
wire n_28211;
wire n_28212;
wire n_28213;
wire n_28214;
wire n_28216;
wire n_28217;
wire n_28218;
wire n_28219;
wire n_28220;
wire n_28221;
wire n_28222;
wire n_28223;
wire n_28224;
wire n_28225;
wire n_28226;
wire n_28227;
wire n_28228;
wire n_28229;
wire n_2823;
wire n_28230;
wire n_28231;
wire n_28232;
wire n_28233;
wire n_28234;
wire n_28238;
wire n_28239;
wire n_2824;
wire n_28240;
wire n_28241;
wire n_28242;
wire n_28243;
wire n_28244;
wire n_28245;
wire n_28246;
wire n_28247;
wire n_28248;
wire n_28249;
wire n_2825;
wire n_28250;
wire n_28251;
wire n_28252;
wire n_28253;
wire n_28254;
wire n_28255;
wire n_28256;
wire n_28257;
wire n_28259;
wire n_2826;
wire n_28261;
wire n_28262;
wire n_28263;
wire n_28264;
wire n_28265;
wire n_28266;
wire TIMEBOOST_net_2539;
wire n_28268;
wire TIMEBOOST_net_52;
wire n_2827;
wire n_28270;
wire n_28271;
wire n_28273;
wire n_28276;
wire n_28277;
wire n_28278;
wire n_28279;
wire n_28280;
wire TIMEBOOST_net_804;
wire n_28282;
wire n_28283;
wire n_28284;
wire n_28285;
wire n_28286;
wire n_28288;
wire n_28289;
wire n_2829;
wire n_28290;
wire n_28291;
wire n_28292;
wire n_28293;
wire n_28294;
wire n_28295;
wire n_28297;
wire n_28298;
wire n_28299;
wire n_283;
wire n_2830;
wire n_28300;
wire n_28302;
wire n_28303;
wire n_28304;
wire n_28305;
wire n_28306;
wire n_28307;
wire n_28308;
wire n_28309;
wire n_2831;
wire n_28310;
wire n_28311;
wire n_28312;
wire n_28314;
wire n_28315;
wire n_28316;
wire n_28317;
wire n_28318;
wire n_28319;
wire n_2832;
wire n_28320;
wire n_28321;
wire n_28322;
wire n_28326;
wire n_28327;
wire n_28328;
wire n_28329;
wire n_28330;
wire n_28331;
wire n_28332;
wire n_28333;
wire n_28334;
wire n_28335;
wire n_28336;
wire n_28338;
wire n_28339;
wire n_2834;
wire n_28340;
wire n_28341;
wire n_28342;
wire n_28343;
wire n_28344;
wire TIMEBOOST_net_2138;
wire n_28347;
wire n_28348;
wire n_28349;
wire n_2835;
wire n_28350;
wire n_28351;
wire n_28352;
wire n_28353;
wire n_28354;
wire n_28355;
wire n_28356;
wire n_28357;
wire n_28358;
wire n_28359;
wire n_2836;
wire n_28360;
wire n_28361;
wire n_28362;
wire n_28363;
wire n_28364;
wire n_28365;
wire n_28366;
wire n_28367;
wire n_28368;
wire n_28369;
wire n_28370;
wire n_28371;
wire n_28372;
wire n_28373;
wire n_28378;
wire n_28379;
wire n_2838;
wire n_28380;
wire n_28381;
wire TIMEBOOST_net_927;
wire n_28383;
wire n_28384;
wire n_28385;
wire n_28387;
wire n_28388;
wire n_28389;
wire n_28390;
wire n_28391;
wire n_28396;
wire n_28397;
wire n_28398;
wire n_28399;
wire n_284;
wire n_2840;
wire n_28401;
wire n_28402;
wire n_28403;
wire n_28404;
wire n_28405;
wire n_28406;
wire n_28407;
wire n_2841;
wire n_28415;
wire n_28416;
wire n_28417;
wire n_28418;
wire n_28419;
wire n_2842;
wire n_28420;
wire n_28421;
wire n_28422;
wire n_28423;
wire n_28424;
wire n_28425;
wire n_28426;
wire n_28427;
wire n_28428;
wire n_2843;
wire n_28434;
wire n_28435;
wire n_28436;
wire n_28437;
wire n_28438;
wire n_28439;
wire n_2844;
wire n_28440;
wire n_28441;
wire n_28445;
wire n_28446;
wire n_28447;
wire n_28448;
wire n_28449;
wire n_2845;
wire n_28450;
wire n_28451;
wire n_28452;
wire n_28453;
wire n_28454;
wire n_28455;
wire n_28457;
wire n_28458;
wire n_2846;
wire n_28460;
wire n_28463;
wire n_28464;
wire n_28465;
wire n_28466;
wire n_28467;
wire n_28468;
wire n_28469;
wire n_2847;
wire n_28472;
wire n_28473;
wire n_28474;
wire n_28475;
wire n_28476;
wire n_28477;
wire n_28478;
wire n_28479;
wire n_2848;
wire n_28480;
wire n_28484;
wire n_28485;
wire n_28486;
wire n_28487;
wire n_28489;
wire n_2849;
wire n_28490;
wire n_28491;
wire n_28492;
wire n_28493;
wire n_28494;
wire n_28495;
wire n_28496;
wire n_28498;
wire n_28499;
wire n_285;
wire n_2850;
wire n_28501;
wire n_28504;
wire n_28505;
wire n_28507;
wire n_28508;
wire n_28509;
wire n_2851;
wire n_28510;
wire n_28511;
wire n_28512;
wire n_28513;
wire n_28514;
wire n_28515;
wire n_2852;
wire n_28520;
wire n_28521;
wire n_28522;
wire n_28523;
wire n_28525;
wire n_28526;
wire n_28527;
wire n_28528;
wire n_28529;
wire n_2853;
wire n_28530;
wire n_28532;
wire n_28533;
wire n_28534;
wire n_28535;
wire n_28536;
wire n_28538;
wire n_28539;
wire n_2854;
wire n_28541;
wire n_28542;
wire n_28543;
wire n_28544;
wire n_28545;
wire n_28547;
wire n_28548;
wire n_28549;
wire n_2855;
wire n_28550;
wire n_28551;
wire n_28552;
wire n_28555;
wire n_28556;
wire n_28557;
wire n_28558;
wire n_28559;
wire n_2856;
wire n_28560;
wire n_28565;
wire n_28566;
wire n_28567;
wire n_28568;
wire n_28569;
wire n_28570;
wire n_28571;
wire n_28572;
wire n_28573;
wire n_28574;
wire n_28575;
wire n_28577;
wire n_28579;
wire n_2858;
wire n_28582;
wire n_28583;
wire n_28585;
wire n_28586;
wire n_28587;
wire n_28588;
wire n_28589;
wire n_2859;
wire n_28590;
wire n_28591;
wire n_28592;
wire TIMEBOOST_net_1649;
wire n_286;
wire n_2860;
wire n_28600;
wire n_28601;
wire n_28602;
wire n_28603;
wire n_28604;
wire n_28605;
wire n_28606;
wire n_28607;
wire n_28608;
wire n_28609;
wire n_2861;
wire n_28610;
wire n_28611;
wire n_28612;
wire n_28615;
wire n_28616;
wire n_28617;
wire n_28618;
wire n_28619;
wire n_2862;
wire n_28620;
wire n_28621;
wire n_28624;
wire n_28625;
wire n_28626;
wire n_28627;
wire n_28628;
wire n_2863;
wire n_28630;
wire n_28631;
wire n_28632;
wire n_28634;
wire n_28635;
wire n_28636;
wire n_28637;
wire n_28638;
wire n_28639;
wire n_2864;
wire n_28643;
wire n_28644;
wire n_28645;
wire n_28646;
wire n_28647;
wire TIMEBOOST_net_103;
wire n_28649;
wire n_2865;
wire n_28650;
wire n_28651;
wire n_28652;
wire n_28654;
wire n_28655;
wire n_28656;
wire n_28657;
wire n_28658;
wire n_28659;
wire n_2866;
wire n_28660;
wire n_28661;
wire n_28664;
wire n_28665;
wire n_28666;
wire n_28667;
wire n_28668;
wire n_28669;
wire n_2867;
wire n_28672;
wire n_28673;
wire n_28674;
wire n_28675;
wire n_28676;
wire n_28677;
wire n_28678;
wire n_28679;
wire n_28680;
wire n_28681;
wire n_28682;
wire n_28683;
wire n_28684;
wire n_28685;
wire n_28689;
wire n_2869;
wire n_28690;
wire n_28691;
wire n_28692;
wire n_28693;
wire n_28694;
wire n_28698;
wire n_28699;
wire n_287;
wire n_2870;
wire n_28701;
wire n_28703;
wire n_28704;
wire n_28705;
wire n_28707;
wire n_28708;
wire n_28709;
wire n_2871;
wire n_28710;
wire n_28711;
wire n_28712;
wire n_28713;
wire n_28714;
wire n_28715;
wire n_28718;
wire n_28719;
wire n_2872;
wire n_28720;
wire n_28721;
wire n_28722;
wire n_28723;
wire n_28724;
wire n_28725;
wire n_28726;
wire n_28728;
wire n_28729;
wire n_2873;
wire n_28730;
wire n_28732;
wire n_28733;
wire n_28734;
wire n_28735;
wire n_28736;
wire n_28737;
wire n_28739;
wire n_2874;
wire n_28740;
wire n_28741;
wire n_28742;
wire n_28743;
wire n_28744;
wire n_28745;
wire n_28746;
wire n_28747;
wire n_28748;
wire n_28749;
wire n_2875;
wire n_28750;
wire n_28751;
wire n_28752;
wire n_28753;
wire n_28754;
wire n_28755;
wire n_28756;
wire n_28757;
wire n_28758;
wire n_2876;
wire n_28761;
wire n_28762;
wire n_28764;
wire n_28766;
wire n_28767;
wire n_28768;
wire n_28769;
wire n_2877;
wire n_28770;
wire n_28771;
wire n_28773;
wire n_28774;
wire n_28775;
wire n_28777;
wire n_28778;
wire n_28779;
wire n_2878;
wire n_28780;
wire n_28781;
wire n_28784;
wire n_28785;
wire n_28786;
wire n_28787;
wire n_28788;
wire n_28789;
wire n_28790;
wire n_28791;
wire n_28793;
wire n_28795;
wire n_28798;
wire n_28799;
wire n_288;
wire n_2880;
wire n_28801;
wire n_28802;
wire n_28803;
wire n_28804;
wire n_28805;
wire n_28806;
wire n_28807;
wire n_28810;
wire n_28811;
wire n_28812;
wire n_28813;
wire n_28815;
wire n_28816;
wire n_28817;
wire n_2882;
wire n_28820;
wire n_28822;
wire n_28823;
wire n_28824;
wire n_28825;
wire n_28826;
wire n_28828;
wire n_28829;
wire n_28830;
wire n_28832;
wire n_28833;
wire n_28834;
wire n_28835;
wire n_28836;
wire n_28837;
wire n_28838;
wire n_28839;
wire n_2884;
wire n_28840;
wire n_28841;
wire n_28842;
wire n_28843;
wire n_28845;
wire n_28846;
wire n_28847;
wire n_28848;
wire n_28849;
wire n_2885;
wire n_28850;
wire n_28851;
wire n_28852;
wire n_28853;
wire n_28856;
wire n_28858;
wire n_28859;
wire n_2886;
wire n_28860;
wire n_28862;
wire n_28863;
wire n_28864;
wire n_28865;
wire n_28866;
wire n_28867;
wire n_28869;
wire n_2887;
wire n_28870;
wire n_28871;
wire n_28872;
wire n_28877;
wire n_28878;
wire n_28879;
wire n_2888;
wire n_28881;
wire n_28882;
wire n_28883;
wire n_28885;
wire n_28886;
wire n_28887;
wire n_28888;
wire n_28889;
wire n_2889;
wire n_28890;
wire n_28891;
wire n_28892;
wire n_28893;
wire n_28894;
wire n_28897;
wire n_28898;
wire n_28899;
wire n_289;
wire n_2890;
wire n_28901;
wire n_28902;
wire n_28903;
wire n_28904;
wire n_28905;
wire n_28906;
wire n_28907;
wire n_28908;
wire n_28909;
wire n_28910;
wire n_28911;
wire n_28912;
wire n_28913;
wire n_28914;
wire n_28915;
wire n_28919;
wire n_2892;
wire n_28921;
wire n_28922;
wire n_28923;
wire n_28924;
wire n_28925;
wire n_28926;
wire n_28927;
wire n_28928;
wire n_28929;
wire n_28930;
wire n_28931;
wire n_28933;
wire n_28934;
wire n_28935;
wire n_28937;
wire n_28939;
wire n_2894;
wire n_28940;
wire n_28941;
wire n_28942;
wire n_28943;
wire n_28945;
wire n_28946;
wire n_28948;
wire n_28949;
wire n_2895;
wire n_28950;
wire n_28951;
wire n_28952;
wire n_28955;
wire n_28956;
wire n_28957;
wire n_28958;
wire n_28959;
wire n_2896;
wire n_28960;
wire n_28961;
wire n_28962;
wire n_28965;
wire n_28966;
wire n_28967;
wire n_28968;
wire n_2897;
wire n_28970;
wire n_28971;
wire n_28972;
wire n_28973;
wire n_28974;
wire n_28975;
wire n_28976;
wire n_28977;
wire n_28978;
wire n_28979;
wire n_2898;
wire n_28982;
wire n_28984;
wire n_28986;
wire n_28987;
wire n_28988;
wire n_28989;
wire n_2899;
wire n_28990;
wire n_28991;
wire n_28992;
wire n_28993;
wire n_28994;
wire n_28995;
wire n_28996;
wire n_28997;
wire n_28998;
wire n_29;
wire n_290;
wire n_2900;
wire n_29000;
wire n_29001;
wire n_29002;
wire n_29003;
wire n_29004;
wire n_29006;
wire n_29007;
wire n_29008;
wire n_2901;
wire n_29010;
wire n_29011;
wire n_29012;
wire n_29013;
wire n_29014;
wire n_29015;
wire n_29016;
wire n_29017;
wire n_29018;
wire TIMEBOOST_net_971;
wire n_2902;
wire n_29020;
wire n_29023;
wire n_29024;
wire n_29025;
wire n_29026;
wire n_29028;
wire n_29029;
wire n_2903;
wire n_29030;
wire n_29031;
wire n_29033;
wire n_29034;
wire n_29036;
wire TIMEBOOST_net_1520;
wire n_29038;
wire n_29039;
wire n_2904;
wire n_29040;
wire n_29041;
wire n_29042;
wire n_29043;
wire n_29044;
wire n_29045;
wire n_29046;
wire n_29047;
wire n_29048;
wire n_29049;
wire n_2905;
wire n_29050;
wire n_29051;
wire n_29053;
wire n_29054;
wire n_29055;
wire n_29056;
wire n_29057;
wire n_29058;
wire n_29059;
wire n_2906;
wire n_29060;
wire n_29062;
wire n_29063;
wire n_29064;
wire n_29065;
wire n_29067;
wire n_29068;
wire n_29069;
wire n_2907;
wire n_29070;
wire n_29071;
wire n_29072;
wire n_29073;
wire n_29074;
wire n_29076;
wire n_29077;
wire n_29078;
wire n_29079;
wire n_2908;
wire n_29080;
wire n_29081;
wire n_29082;
wire n_29083;
wire n_2909;
wire n_29091;
wire n_29092;
wire n_29094;
wire n_29095;
wire TIMEBOOST_net_132;
wire n_29097;
wire n_29098;
wire n_29099;
wire n_291;
wire n_2910;
wire n_29100;
wire n_29101;
wire n_29102;
wire n_29103;
wire n_29104;
wire n_29105;
wire n_29109;
wire n_2911;
wire n_29110;
wire n_29112;
wire n_29113;
wire TIMEBOOST_net_2836;
wire n_29115;
wire n_29116;
wire n_29117;
wire n_29118;
wire TIMEBOOST_net_2605;
wire n_2912;
wire n_29120;
wire n_29121;
wire n_29122;
wire n_29123;
wire n_29124;
wire n_29125;
wire n_29126;
wire n_29127;
wire n_29128;
wire n_29129;
wire n_2913;
wire n_29130;
wire n_29131;
wire n_29132;
wire n_29135;
wire n_29137;
wire n_29139;
wire n_2914;
wire n_29140;
wire n_29141;
wire n_29143;
wire n_29144;
wire n_29145;
wire n_29148;
wire n_29149;
wire n_2915;
wire n_29150;
wire n_29151;
wire n_29154;
wire n_29155;
wire n_29156;
wire n_29157;
wire n_29158;
wire n_29159;
wire n_29160;
wire n_29161;
wire n_29163;
wire n_29164;
wire n_29165;
wire TIMEBOOST_net_119;
wire n_29167;
wire n_29169;
wire TIMEBOOST_net_2755;
wire n_29170;
wire n_29171;
wire n_29172;
wire n_29174;
wire n_29175;
wire n_29176;
wire n_29177;
wire n_2918;
wire n_29180;
wire TIMEBOOST_net_1904;
wire n_29187;
wire n_29188;
wire n_29189;
wire n_2919;
wire n_29190;
wire n_29192;
wire n_29193;
wire n_29194;
wire TIMEBOOST_net_958;
wire n_29196;
wire TIMEBOOST_net_1029;
wire n_29198;
wire n_292;
wire n_2920;
wire n_29200;
wire n_29201;
wire n_29202;
wire n_29203;
wire n_29204;
wire n_29205;
wire n_2921;
wire n_29210;
wire n_29211;
wire TIMEBOOST_net_2750;
wire n_29215;
wire n_29216;
wire n_29217;
wire n_29218;
wire n_29219;
wire n_2922;
wire TIMEBOOST_net_144;
wire n_29223;
wire n_29224;
wire n_29225;
wire n_29226;
wire n_29227;
wire n_29228;
wire n_29229;
wire n_2923;
wire n_29231;
wire n_29232;
wire n_29233;
wire n_29235;
wire n_29236;
wire n_29239;
wire n_2924;
wire n_29240;
wire n_29241;
wire n_29242;
wire n_29243;
wire n_29245;
wire n_29246;
wire n_29247;
wire n_29248;
wire n_29249;
wire TIMEBOOST_net_1591;
wire n_29250;
wire n_29251;
wire n_29252;
wire n_29253;
wire n_29254;
wire n_29255;
wire n_29256;
wire n_29258;
wire n_29260;
wire n_29262;
wire n_29263;
wire n_29265;
wire n_29266;
wire n_29267;
wire n_29268;
wire n_29269;
wire n_2927;
wire n_29270;
wire n_29271;
wire n_29272;
wire n_29273;
wire TIMEBOOST_net_211;
wire n_29279;
wire TIMEBOOST_net_1110;
wire n_29280;
wire TIMEBOOST_net_986;
wire n_29285;
wire n_29286;
wire n_29287;
wire n_29288;
wire n_2929;
wire n_29290;
wire n_29291;
wire n_29292;
wire n_29298;
wire n_29299;
wire n_293;
wire n_2930;
wire n_29301;
wire n_29302;
wire n_29303;
wire TIMEBOOST_net_861;
wire n_29305;
wire n_29306;
wire n_29308;
wire n_29309;
wire n_29310;
wire n_29311;
wire n_29312;
wire n_29313;
wire n_29316;
wire n_29317;
wire n_29318;
wire n_29319;
wire n_2932;
wire n_29322;
wire TIMEBOOST_net_904;
wire TIMEBOOST_net_1530;
wire TIMEBOOST_net_2588;
wire n_29327;
wire n_29328;
wire n_29329;
wire n_29330;
wire n_29332;
wire n_29333;
wire n_29334;
wire n_29335;
wire n_29336;
wire n_29337;
wire n_29339;
wire n_29340;
wire n_29341;
wire TIMEBOOST_net_2849;
wire n_29343;
wire n_29344;
wire n_29345;
wire n_29347;
wire n_29349;
wire n_2935;
wire n_29352;
wire n_29353;
wire TIMEBOOST_net_216;
wire n_29358;
wire n_29359;
wire n_29360;
wire n_29361;
wire n_29362;
wire n_29363;
wire n_29364;
wire n_29365;
wire n_29368;
wire n_29369;
wire n_2937;
wire n_29371;
wire n_29372;
wire n_29373;
wire n_29374;
wire n_29375;
wire n_29376;
wire n_29378;
wire n_29379;
wire n_2938;
wire n_29380;
wire n_29381;
wire n_29382;
wire n_29383;
wire n_29384;
wire n_29385;
wire n_29386;
wire TIMEBOOST_net_1878;
wire n_29388;
wire n_29389;
wire n_2939;
wire TIMEBOOST_net_1051;
wire n_29391;
wire n_29392;
wire n_29393;
wire n_29395;
wire n_29396;
wire n_29397;
wire n_29398;
wire n_29399;
wire n_294;
wire n_2940;
wire n_29400;
wire n_29401;
wire n_29403;
wire TIMEBOOST_net_2372;
wire n_29405;
wire n_29406;
wire n_29407;
wire n_29408;
wire n_29409;
wire n_29410;
wire n_29411;
wire TIMEBOOST_net_1567;
wire n_29413;
wire n_29414;
wire n_29415;
wire n_29417;
wire n_29418;
wire n_29419;
wire n_29420;
wire n_29421;
wire n_29422;
wire TIMEBOOST_net_1913;
wire n_29424;
wire n_29425;
wire TIMEBOOST_net_2848;
wire n_29428;
wire n_2943;
wire n_29431;
wire n_29432;
wire n_29433;
wire n_29436;
wire n_29437;
wire n_29438;
wire n_29439;
wire n_2944;
wire n_29440;
wire n_29441;
wire n_29442;
wire n_29443;
wire n_29444;
wire n_29445;
wire n_29446;
wire n_29448;
wire n_29450;
wire n_29451;
wire n_29453;
wire n_29454;
wire n_29456;
wire n_29457;
wire n_29458;
wire n_29459;
wire n_2946;
wire n_29460;
wire n_29461;
wire n_29462;
wire n_29463;
wire n_29464;
wire n_29465;
wire n_29466;
wire n_29467;
wire n_2947;
wire n_29470;
wire n_29472;
wire n_29473;
wire n_29475;
wire n_29476;
wire n_29477;
wire n_29479;
wire n_2948;
wire n_29480;
wire n_29481;
wire TIMEBOOST_net_244;
wire TIMEBOOST_net_1072;
wire n_29485;
wire TIMEBOOST_net_127;
wire n_29487;
wire n_29488;
wire n_29489;
wire n_2949;
wire n_29490;
wire n_29491;
wire n_29492;
wire n_29494;
wire n_29495;
wire n_29496;
wire n_29497;
wire n_29498;
wire n_295;
wire n_2950;
wire n_29500;
wire n_29501;
wire n_29502;
wire n_29504;
wire n_29505;
wire n_29507;
wire TIMEBOOST_net_1877;
wire n_29509;
wire n_2951;
wire n_29510;
wire n_29511;
wire n_29512;
wire n_29513;
wire n_29514;
wire n_29515;
wire n_29516;
wire n_29518;
wire n_29523;
wire n_29525;
wire n_29526;
wire n_29527;
wire n_29529;
wire n_2953;
wire n_29530;
wire TIMEBOOST_net_2812;
wire n_29532;
wire n_29533;
wire n_29534;
wire n_29535;
wire n_29536;
wire n_29537;
wire n_29538;
wire n_2954;
wire n_29542;
wire n_29543;
wire n_29544;
wire n_29545;
wire TIMEBOOST_net_261;
wire n_29549;
wire n_29550;
wire n_29551;
wire n_29553;
wire n_29554;
wire n_29555;
wire n_29556;
wire n_29558;
wire n_29559;
wire n_2956;
wire n_29560;
wire n_29561;
wire n_29562;
wire n_29564;
wire n_29565;
wire n_29566;
wire n_29568;
wire n_2957;
wire n_29570;
wire n_29571;
wire n_29572;
wire n_29573;
wire n_29574;
wire n_29576;
wire n_29577;
wire n_29579;
wire n_2958;
wire n_29581;
wire n_29582;
wire n_29583;
wire n_29584;
wire n_29585;
wire n_29586;
wire n_29587;
wire n_29588;
wire n_29589;
wire n_2959;
wire n_29590;
wire n_29591;
wire n_29592;
wire n_29593;
wire n_29594;
wire TIMEBOOST_net_227;
wire n_29596;
wire n_29597;
wire n_29598;
wire n_29599;
wire n_296;
wire n_2960;
wire n_29600;
wire n_29601;
wire n_29602;
wire n_29603;
wire n_29604;
wire n_29605;
wire n_29606;
wire n_29607;
wire n_29608;
wire n_29609;
wire n_2961;
wire n_29610;
wire n_29611;
wire n_29612;
wire n_29613;
wire n_29615;
wire n_29616;
wire n_2962;
wire n_29620;
wire n_29621;
wire n_29622;
wire n_29624;
wire n_29628;
wire n_2963;
wire n_29630;
wire n_29631;
wire n_29632;
wire n_29633;
wire n_29634;
wire n_29635;
wire n_29636;
wire n_29637;
wire n_29638;
wire n_29639;
wire n_2964;
wire n_29640;
wire n_29641;
wire n_29642;
wire n_29643;
wire n_29644;
wire n_29645;
wire TIMEBOOST_net_1075;
wire n_29648;
wire n_29649;
wire n_2965;
wire n_29650;
wire n_29651;
wire n_29652;
wire n_29653;
wire n_29654;
wire n_29655;
wire n_29656;
wire n_29657;
wire n_29658;
wire n_29659;
wire TIMEBOOST_net_2609;
wire n_29660;
wire n_29661;
wire n_29663;
wire n_29666;
wire n_29667;
wire n_29668;
wire n_29669;
wire n_2967;
wire n_29670;
wire n_29671;
wire n_29672;
wire n_29673;
wire n_29674;
wire n_29675;
wire n_29676;
wire n_29677;
wire n_29678;
wire n_2968;
wire n_29681;
wire n_29686;
wire n_29687;
wire TIMEBOOST_net_268;
wire n_29689;
wire n_2969;
wire n_29690;
wire n_29691;
wire n_29692;
wire n_29693;
wire n_29694;
wire n_29696;
wire n_29697;
wire n_29698;
wire n_297;
wire n_2970;
wire n_29700;
wire TIMEBOOST_net_1574;
wire n_29702;
wire n_29703;
wire n_29704;
wire TIMEBOOST_net_2944;
wire n_29706;
wire n_29707;
wire n_29708;
wire n_29709;
wire n_29710;
wire n_29711;
wire n_29712;
wire n_29713;
wire n_29714;
wire n_29715;
wire n_29716;
wire n_29717;
wire n_29718;
wire n_29719;
wire TIMEBOOST_net_1158;
wire n_29720;
wire n_29721;
wire n_29722;
wire n_29723;
wire n_29724;
wire n_29725;
wire n_29727;
wire n_29728;
wire n_29729;
wire n_2973;
wire n_29730;
wire TIMEBOOST_net_283;
wire n_29732;
wire n_29733;
wire n_29734;
wire n_29735;
wire n_29736;
wire n_29737;
wire n_29738;
wire n_29739;
wire n_2974;
wire n_29740;
wire n_29741;
wire n_29742;
wire n_29743;
wire n_29744;
wire TIMEBOOST_net_1132;
wire n_29746;
wire n_29747;
wire n_29748;
wire n_29749;
wire n_2975;
wire TIMEBOOST_net_1077;
wire n_29751;
wire n_29752;
wire n_29753;
wire n_29754;
wire n_29755;
wire n_29756;
wire n_29757;
wire n_29758;
wire n_29759;
wire n_2976;
wire n_29760;
wire n_29761;
wire n_29762;
wire n_29763;
wire n_29764;
wire n_29765;
wire n_29766;
wire n_29767;
wire n_29768;
wire n_29769;
wire n_2977;
wire n_29770;
wire n_29771;
wire n_29773;
wire n_29775;
wire n_29776;
wire n_29777;
wire n_29778;
wire n_29779;
wire n_2978;
wire n_29780;
wire n_29781;
wire n_29783;
wire n_29784;
wire n_29785;
wire n_29786;
wire n_29787;
wire n_29788;
wire n_29789;
wire n_2979;
wire n_29790;
wire n_29791;
wire n_29792;
wire n_29793;
wire n_29794;
wire n_29795;
wire n_29796;
wire n_29797;
wire n_29799;
wire n_298;
wire n_2980;
wire n_29800;
wire n_29801;
wire n_29802;
wire n_29803;
wire n_29804;
wire n_29805;
wire n_29806;
wire n_29807;
wire n_29808;
wire n_29809;
wire n_29810;
wire n_29811;
wire n_29812;
wire n_29813;
wire n_29814;
wire n_29815;
wire n_29816;
wire n_29817;
wire n_29818;
wire n_29819;
wire n_2982;
wire n_29820;
wire n_29821;
wire n_29822;
wire n_29823;
wire n_29824;
wire n_29825;
wire n_29826;
wire n_29827;
wire n_29828;
wire n_2983;
wire n_29831;
wire n_29832;
wire n_29833;
wire n_29834;
wire n_29835;
wire n_29836;
wire n_29837;
wire n_29838;
wire n_29839;
wire n_29841;
wire n_29842;
wire n_29843;
wire n_29844;
wire n_29845;
wire n_29846;
wire n_29847;
wire n_29848;
wire n_2985;
wire n_29850;
wire n_29851;
wire n_29852;
wire n_29853;
wire n_29854;
wire TIMEBOOST_net_1133;
wire n_29856;
wire n_29857;
wire n_29859;
wire n_2986;
wire n_29860;
wire n_29861;
wire n_29862;
wire n_29863;
wire n_29864;
wire n_29865;
wire n_29866;
wire n_29868;
wire n_29869;
wire n_2987;
wire n_29870;
wire n_29871;
wire n_29872;
wire n_29873;
wire n_29874;
wire n_29875;
wire n_29877;
wire n_29878;
wire n_29879;
wire n_2988;
wire n_29880;
wire n_29881;
wire n_29882;
wire n_29883;
wire n_29884;
wire n_29886;
wire n_29887;
wire n_29888;
wire n_29889;
wire n_2989;
wire n_29890;
wire n_29892;
wire n_29893;
wire n_29894;
wire n_29895;
wire n_29896;
wire n_29897;
wire n_29898;
wire n_29899;
wire n_299;
wire n_2990;
wire TIMEBOOST_net_281;
wire n_29901;
wire n_29902;
wire n_29903;
wire n_29904;
wire n_29905;
wire n_29906;
wire n_29907;
wire n_29908;
wire n_29909;
wire n_2991;
wire n_29910;
wire n_29913;
wire n_29915;
wire n_29916;
wire n_29918;
wire n_29919;
wire n_2992;
wire n_29920;
wire n_29922;
wire n_29925;
wire n_29926;
wire TIMEBOOST_net_1086;
wire n_29928;
wire n_29929;
wire n_29930;
wire n_29931;
wire n_29932;
wire n_29935;
wire n_29936;
wire n_29937;
wire n_29938;
wire n_29939;
wire n_29940;
wire n_29942;
wire n_29943;
wire n_29944;
wire n_29945;
wire n_29946;
wire n_29947;
wire n_2995;
wire n_29951;
wire n_29952;
wire n_29953;
wire n_29954;
wire n_29955;
wire n_29956;
wire n_29957;
wire n_29958;
wire n_29959;
wire n_2996;
wire n_29960;
wire n_29961;
wire n_29962;
wire n_29963;
wire n_29964;
wire n_29965;
wire n_29966;
wire n_29967;
wire n_29968;
wire n_29969;
wire n_2997;
wire n_29970;
wire n_29974;
wire n_29975;
wire n_29976;
wire n_29977;
wire n_2998;
wire n_29982;
wire n_29984;
wire n_29985;
wire n_29986;
wire n_29987;
wire n_29988;
wire n_29989;
wire n_2999;
wire n_29990;
wire n_29992;
wire n_29993;
wire n_29995;
wire n_29996;
wire n_29997;
wire n_29998;
wire n_29999;
wire n_300;
wire n_3000;
wire n_30000;
wire n_30001;
wire n_30002;
wire n_30003;
wire n_30004;
wire n_30005;
wire n_30007;
wire n_30010;
wire n_30011;
wire n_30012;
wire n_30013;
wire n_30014;
wire n_30015;
wire n_30016;
wire n_30017;
wire n_30018;
wire n_30019;
wire n_30020;
wire n_30021;
wire n_30022;
wire n_30023;
wire n_30024;
wire n_30025;
wire n_30026;
wire n_30028;
wire n_30029;
wire TIMEBOOST_net_1948;
wire n_30030;
wire n_30033;
wire n_30034;
wire n_30035;
wire n_30036;
wire n_30037;
wire n_30038;
wire n_30039;
wire n_3004;
wire n_30040;
wire n_30046;
wire n_30049;
wire n_3005;
wire n_30050;
wire n_30051;
wire n_30053;
wire n_30054;
wire n_30055;
wire n_30056;
wire n_30057;
wire n_30059;
wire n_3006;
wire n_30060;
wire n_30061;
wire n_30062;
wire n_30063;
wire n_30064;
wire n_30065;
wire n_30066;
wire n_30067;
wire n_30068;
wire TIMEBOOST_net_1128;
wire n_30071;
wire n_30076;
wire n_30077;
wire n_30078;
wire n_30079;
wire n_3008;
wire n_30080;
wire n_30082;
wire n_30083;
wire n_30084;
wire n_30085;
wire n_30086;
wire n_30088;
wire n_30089;
wire n_3009;
wire n_30090;
wire n_30091;
wire n_30092;
wire n_30093;
wire n_30094;
wire n_30095;
wire n_30096;
wire n_30097;
wire n_30098;
wire n_30099;
wire n_301;
wire n_30100;
wire n_30101;
wire n_30102;
wire n_30103;
wire n_30104;
wire n_30105;
wire TIMEBOOST_net_271;
wire n_30108;
wire n_30111;
wire n_30113;
wire n_30114;
wire n_30116;
wire n_30119;
wire n_3012;
wire n_30120;
wire n_30121;
wire n_30124;
wire n_30125;
wire n_30126;
wire n_30127;
wire n_30128;
wire n_30129;
wire n_3013;
wire n_30130;
wire n_30134;
wire n_30136;
wire n_30138;
wire n_30139;
wire n_3014;
wire n_30140;
wire n_30141;
wire n_30142;
wire n_30143;
wire n_30144;
wire n_30145;
wire n_30147;
wire n_30148;
wire n_30149;
wire n_3015;
wire n_30150;
wire n_30151;
wire n_30152;
wire n_30153;
wire n_30154;
wire n_30155;
wire n_30156;
wire n_30157;
wire n_30158;
wire n_30159;
wire n_3016;
wire n_30160;
wire n_30161;
wire n_30162;
wire n_30163;
wire n_30164;
wire n_30165;
wire n_30166;
wire n_30167;
wire n_30168;
wire n_30170;
wire n_30171;
wire n_30172;
wire n_30173;
wire n_30175;
wire n_30176;
wire n_30177;
wire n_30178;
wire n_30179;
wire n_3018;
wire n_30180;
wire n_30182;
wire n_30183;
wire n_30184;
wire n_30185;
wire n_30186;
wire n_3019;
wire n_30191;
wire n_30192;
wire n_30194;
wire n_30195;
wire n_30196;
wire n_30197;
wire n_30198;
wire n_302;
wire n_3020;
wire n_30200;
wire n_30201;
wire n_30202;
wire n_30203;
wire n_30204;
wire n_30207;
wire n_30208;
wire n_3021;
wire n_30210;
wire n_30211;
wire n_30212;
wire n_30213;
wire n_30214;
wire n_30215;
wire n_30216;
wire n_30217;
wire n_30218;
wire n_30219;
wire n_3022;
wire n_30220;
wire n_30221;
wire n_30223;
wire n_30224;
wire n_30225;
wire n_30226;
wire n_30227;
wire n_30229;
wire n_3023;
wire n_30230;
wire n_30231;
wire n_30232;
wire n_30233;
wire n_30234;
wire n_30235;
wire n_30239;
wire n_3024;
wire n_30240;
wire n_30242;
wire n_30243;
wire n_30244;
wire n_30245;
wire n_30246;
wire n_30247;
wire n_30248;
wire n_30249;
wire n_3025;
wire n_30250;
wire n_30253;
wire n_30254;
wire n_30255;
wire n_30256;
wire n_30258;
wire n_30259;
wire n_3026;
wire n_30260;
wire n_30261;
wire n_30262;
wire n_30263;
wire n_30265;
wire n_30266;
wire n_30267;
wire n_3027;
wire n_30272;
wire n_30273;
wire n_30275;
wire n_30276;
wire n_30277;
wire n_30278;
wire n_30279;
wire TIMEBOOST_net_1130;
wire n_30280;
wire n_30281;
wire n_30283;
wire n_30285;
wire n_30286;
wire n_30288;
wire n_30289;
wire n_3029;
wire n_30290;
wire n_30292;
wire n_30294;
wire n_30295;
wire n_30296;
wire n_30297;
wire n_30298;
wire n_30299;
wire n_303;
wire n_3030;
wire n_30300;
wire n_30302;
wire n_30303;
wire n_30304;
wire n_30305;
wire n_30306;
wire n_30307;
wire n_3031;
wire n_30310;
wire n_30316;
wire n_30317;
wire n_30318;
wire n_30319;
wire n_3032;
wire n_30320;
wire n_30321;
wire n_30322;
wire n_30324;
wire n_30326;
wire n_30327;
wire n_30332;
wire n_30333;
wire n_30334;
wire n_30335;
wire n_30336;
wire n_30337;
wire n_30338;
wire n_30339;
wire n_3034;
wire n_30340;
wire n_30341;
wire n_30343;
wire n_30344;
wire n_30345;
wire n_30347;
wire n_30348;
wire n_30349;
wire n_3035;
wire n_30350;
wire n_30354;
wire n_30355;
wire n_30356;
wire TIMEBOOST_net_2862;
wire n_30358;
wire n_30359;
wire n_30360;
wire n_30364;
wire n_30367;
wire n_30368;
wire n_30369;
wire n_3037;
wire n_30371;
wire n_30372;
wire n_30374;
wire n_30375;
wire n_30376;
wire n_30377;
wire n_30378;
wire n_30379;
wire n_3038;
wire n_30380;
wire n_30381;
wire n_30383;
wire n_30384;
wire n_30385;
wire TIMEBOOST_net_2577;
wire n_30388;
wire n_3039;
wire n_30392;
wire n_30393;
wire n_30394;
wire n_30399;
wire n_304;
wire n_3040;
wire n_30401;
wire n_30403;
wire n_30405;
wire n_30406;
wire n_30407;
wire n_30408;
wire n_30409;
wire n_30410;
wire n_30411;
wire n_30412;
wire n_30413;
wire n_30416;
wire n_30417;
wire n_30418;
wire n_30419;
wire TIMEBOOST_net_2883;
wire n_30420;
wire n_30421;
wire n_30422;
wire n_30423;
wire n_30424;
wire n_30425;
wire n_30426;
wire n_30428;
wire n_30429;
wire n_3043;
wire n_30431;
wire n_30432;
wire n_30433;
wire n_30434;
wire n_30436;
wire n_30437;
wire n_30438;
wire n_3044;
wire n_30440;
wire n_30441;
wire n_30442;
wire n_30443;
wire n_30444;
wire n_30445;
wire n_30446;
wire n_30447;
wire n_30448;
wire n_30449;
wire n_3045;
wire n_30451;
wire n_30452;
wire n_30453;
wire n_30454;
wire n_30455;
wire n_30457;
wire n_30458;
wire n_30459;
wire n_3046;
wire n_30460;
wire n_30461;
wire n_30462;
wire n_30465;
wire n_30466;
wire n_30467;
wire n_30468;
wire n_30469;
wire n_3047;
wire n_30470;
wire n_30471;
wire TIMEBOOST_net_1327;
wire n_30474;
wire n_30475;
wire n_30476;
wire n_30477;
wire n_30478;
wire n_30479;
wire n_3048;
wire n_30480;
wire n_30481;
wire n_30482;
wire n_30483;
wire n_30484;
wire n_30485;
wire n_30486;
wire n_30487;
wire n_30488;
wire n_30489;
wire n_3049;
wire n_30490;
wire n_30492;
wire n_30493;
wire n_30494;
wire n_30495;
wire n_30496;
wire n_30497;
wire n_30498;
wire n_305;
wire n_30500;
wire n_30501;
wire n_30502;
wire n_30504;
wire n_30505;
wire n_30506;
wire n_30508;
wire TIMEBOOST_net_2052;
wire n_3051;
wire n_30510;
wire n_30511;
wire n_30512;
wire TIMEBOOST_net_541;
wire n_30514;
wire n_30515;
wire n_30518;
wire n_30519;
wire n_30520;
wire n_30521;
wire n_30522;
wire n_30525;
wire n_30526;
wire n_30527;
wire n_30528;
wire TIMEBOOST_net_1207;
wire n_30530;
wire TIMEBOOST_net_1842;
wire TIMEBOOST_net_1631;
wire n_30534;
wire n_30535;
wire n_30537;
wire TIMEBOOST_net_473;
wire n_30540;
wire n_30541;
wire n_30542;
wire n_30543;
wire n_30544;
wire n_30545;
wire n_30546;
wire n_30548;
wire n_30549;
wire n_3055;
wire n_30550;
wire TIMEBOOST_net_318;
wire n_30552;
wire n_30553;
wire n_30554;
wire n_30557;
wire n_30558;
wire n_30559;
wire n_3056;
wire TIMEBOOST_net_2826;
wire TIMEBOOST_net_399;
wire n_30564;
wire n_30566;
wire n_3057;
wire n_30572;
wire n_30573;
wire n_30575;
wire n_30576;
wire n_30577;
wire n_30578;
wire TIMEBOOST_net_1126;
wire n_3058;
wire n_30580;
wire n_30582;
wire n_30584;
wire n_30585;
wire n_30586;
wire n_30587;
wire n_30588;
wire n_30589;
wire n_3059;
wire n_30590;
wire n_30591;
wire n_30592;
wire n_30593;
wire n_30597;
wire n_30598;
wire n_30599;
wire n_306;
wire n_30601;
wire n_30603;
wire TIMEBOOST_net_2652;
wire n_30605;
wire n_30608;
wire n_30609;
wire n_3061;
wire n_30610;
wire n_30611;
wire n_30612;
wire n_30614;
wire n_30615;
wire n_30616;
wire n_30617;
wire n_30619;
wire TIMEBOOST_net_1747;
wire n_30621;
wire n_30622;
wire n_30623;
wire n_30624;
wire n_30625;
wire n_30629;
wire n_3063;
wire n_30630;
wire n_30633;
wire n_30634;
wire n_30635;
wire n_30636;
wire n_30637;
wire TIMEBOOST_net_1307;
wire n_30640;
wire n_30643;
wire n_30644;
wire n_3065;
wire n_30650;
wire n_30652;
wire n_30653;
wire n_30655;
wire n_30656;
wire n_30657;
wire n_30658;
wire n_30659;
wire n_3066;
wire n_30662;
wire n_30663;
wire n_3067;
wire n_30670;
wire n_30671;
wire n_30672;
wire n_30673;
wire n_30674;
wire n_30675;
wire n_30676;
wire n_30677;
wire n_30678;
wire n_3068;
wire TIMEBOOST_net_1295;
wire n_30683;
wire n_30687;
wire n_30688;
wire n_30689;
wire n_3069;
wire n_30690;
wire n_30691;
wire n_30692;
wire n_30693;
wire n_30697;
wire n_30698;
wire n_3070;
wire n_30701;
wire n_30703;
wire n_30706;
wire TIMEBOOST_net_1739;
wire n_3071;
wire n_30711;
wire TIMEBOOST_net_547;
wire n_30713;
wire n_30714;
wire n_30718;
wire n_30719;
wire n_3072;
wire n_30720;
wire n_30721;
wire n_30722;
wire n_30723;
wire n_30724;
wire n_30727;
wire n_30729;
wire n_3073;
wire n_30731;
wire n_30733;
wire n_30734;
wire n_30735;
wire n_30736;
wire n_30737;
wire n_30739;
wire n_30741;
wire n_30743;
wire n_30744;
wire n_30747;
wire n_30749;
wire n_3075;
wire n_30750;
wire n_30751;
wire n_30756;
wire n_30757;
wire n_30758;
wire n_3076;
wire n_30760;
wire n_30763;
wire n_30765;
wire n_30766;
wire n_30767;
wire n_30769;
wire n_30771;
wire n_30772;
wire n_30773;
wire n_30774;
wire n_30776;
wire n_30783;
wire n_30785;
wire n_30786;
wire n_30787;
wire TIMEBOOST_net_2397;
wire n_30790;
wire n_30791;
wire n_30799;
wire n_308;
wire n_3080;
wire n_30800;
wire n_30801;
wire n_30803;
wire n_30806;
wire n_30807;
wire n_30808;
wire TIMEBOOST_net_2725;
wire n_30811;
wire n_30812;
wire n_30813;
wire n_30814;
wire n_30817;
wire n_30818;
wire n_3082;
wire n_30820;
wire TIMEBOOST_net_1871;
wire n_30823;
wire n_30824;
wire n_30825;
wire n_30828;
wire n_30829;
wire n_3083;
wire n_30830;
wire n_30832;
wire n_30833;
wire n_30834;
wire n_30835;
wire n_30836;
wire n_30837;
wire n_30838;
wire n_30839;
wire n_3084;
wire n_30840;
wire n_30841;
wire n_30842;
wire n_30843;
wire TIMEBOOST_net_1696;
wire TIMEBOOST_net_2713;
wire n_30847;
wire n_30849;
wire n_3085;
wire n_30851;
wire n_30852;
wire n_30855;
wire n_30856;
wire n_30857;
wire n_30858;
wire n_30859;
wire n_3086;
wire n_30860;
wire TIMEBOOST_net_555;
wire n_30862;
wire n_30863;
wire n_30864;
wire n_30865;
wire n_30867;
wire n_30869;
wire n_3087;
wire n_30870;
wire TIMEBOOST_net_1210;
wire n_30875;
wire n_30876;
wire n_30877;
wire n_30878;
wire n_30879;
wire n_3088;
wire TIMEBOOST_net_1745;
wire n_30882;
wire n_30883;
wire TIMEBOOST_net_413;
wire n_30885;
wire n_30887;
wire n_30888;
wire n_30889;
wire n_3089;
wire n_30890;
wire n_30892;
wire n_30893;
wire n_30894;
wire n_30895;
wire n_30896;
wire n_30897;
wire n_30898;
wire n_30899;
wire n_309;
wire n_3090;
wire n_30900;
wire n_30901;
wire n_30902;
wire n_30903;
wire n_30904;
wire n_30905;
wire n_30906;
wire n_30908;
wire n_3091;
wire n_30910;
wire TIMEBOOST_net_2252;
wire n_30912;
wire n_30913;
wire n_30914;
wire n_30915;
wire n_30917;
wire n_30918;
wire n_30919;
wire n_3092;
wire n_30920;
wire n_30921;
wire n_30922;
wire n_30923;
wire TIMEBOOST_net_379;
wire n_30925;
wire n_30926;
wire n_3093;
wire n_30930;
wire n_30933;
wire n_30936;
wire n_30937;
wire n_30938;
wire n_30939;
wire n_30940;
wire n_30942;
wire n_30943;
wire n_30944;
wire n_30945;
wire n_30946;
wire n_30947;
wire n_30948;
wire n_30949;
wire n_30950;
wire n_30951;
wire n_30952;
wire n_30953;
wire n_30954;
wire n_30955;
wire n_30956;
wire n_30958;
wire n_3096;
wire n_30960;
wire n_30961;
wire n_30962;
wire n_30963;
wire n_30965;
wire n_30967;
wire n_30968;
wire n_30969;
wire n_3097;
wire n_30970;
wire n_30971;
wire n_30972;
wire n_30973;
wire n_30974;
wire n_30975;
wire n_30976;
wire n_30977;
wire n_30978;
wire n_30979;
wire n_3098;
wire n_30987;
wire n_30988;
wire n_30989;
wire n_30991;
wire n_30992;
wire TIMEBOOST_net_2867;
wire n_30995;
wire n_30996;
wire n_30997;
wire n_30998;
wire n_310;
wire n_3100;
wire n_31001;
wire n_31003;
wire n_31004;
wire n_31005;
wire n_31007;
wire n_31008;
wire n_3101;
wire n_31010;
wire n_31011;
wire n_31012;
wire n_31013;
wire n_31014;
wire n_31015;
wire n_31016;
wire n_31017;
wire n_31018;
wire n_3102;
wire n_31021;
wire n_31022;
wire n_31023;
wire n_31025;
wire n_31026;
wire n_31027;
wire n_31029;
wire n_3103;
wire n_31030;
wire TIMEBOOST_net_2047;
wire n_31032;
wire n_31034;
wire n_31035;
wire n_31036;
wire TIMEBOOST_net_1388;
wire n_31038;
wire n_31039;
wire n_3104;
wire n_31040;
wire n_31041;
wire n_31042;
wire n_31043;
wire n_31044;
wire n_31045;
wire n_31046;
wire n_31048;
wire n_3105;
wire n_31050;
wire n_31051;
wire n_31053;
wire n_31054;
wire n_31055;
wire n_31056;
wire n_31057;
wire n_31058;
wire n_3106;
wire n_31060;
wire n_31061;
wire n_31062;
wire n_31063;
wire n_31064;
wire n_31065;
wire n_31066;
wire n_31067;
wire n_3107;
wire n_31070;
wire n_31071;
wire n_31073;
wire n_31074;
wire n_31075;
wire n_31076;
wire n_31077;
wire n_31079;
wire n_3108;
wire n_31081;
wire n_31082;
wire n_31083;
wire n_31086;
wire n_31088;
wire n_31089;
wire n_3109;
wire n_31090;
wire n_31091;
wire n_31092;
wire n_31093;
wire n_31094;
wire n_31095;
wire n_31097;
wire n_31099;
wire n_311;
wire n_31100;
wire n_31101;
wire n_31103;
wire n_31105;
wire n_31107;
wire n_31108;
wire n_31109;
wire n_3111;
wire n_31110;
wire n_31111;
wire n_31112;
wire n_31114;
wire n_31115;
wire n_31116;
wire n_31117;
wire n_31118;
wire n_31119;
wire n_3112;
wire n_31120;
wire n_31121;
wire n_31122;
wire n_31123;
wire n_31124;
wire n_31125;
wire n_31126;
wire TIMEBOOST_net_424;
wire n_3113;
wire n_31130;
wire TIMEBOOST_net_2700;
wire n_31132;
wire TIMEBOOST_net_2073;
wire n_31136;
wire TIMEBOOST_net_421;
wire n_31138;
wire n_31139;
wire n_3114;
wire n_31140;
wire n_31141;
wire n_31142;
wire n_31143;
wire n_31144;
wire n_31145;
wire n_31147;
wire n_31148;
wire n_31149;
wire n_3115;
wire n_31150;
wire n_31151;
wire n_31152;
wire n_31153;
wire TIMEBOOST_net_2643;
wire n_31156;
wire n_31158;
wire n_3116;
wire n_31160;
wire n_31161;
wire n_31162;
wire n_31163;
wire n_31164;
wire n_31165;
wire n_31169;
wire n_3117;
wire n_31171;
wire n_31172;
wire n_31174;
wire n_31175;
wire n_31176;
wire n_31177;
wire n_3118;
wire n_31180;
wire n_31182;
wire n_31183;
wire n_31184;
wire n_31185;
wire n_31186;
wire n_31187;
wire n_31189;
wire n_3119;
wire n_31190;
wire n_31191;
wire n_31192;
wire n_31193;
wire n_31194;
wire n_31196;
wire n_31197;
wire n_31198;
wire n_31199;
wire n_312;
wire n_3120;
wire n_31200;
wire n_31201;
wire n_31202;
wire n_31203;
wire n_31204;
wire n_31205;
wire n_31206;
wire n_31207;
wire n_31208;
wire n_31209;
wire n_31210;
wire n_31211;
wire n_31212;
wire n_31213;
wire n_31214;
wire n_31216;
wire n_31219;
wire n_3122;
wire n_31220;
wire n_31221;
wire n_31222;
wire n_31223;
wire n_31224;
wire TIMEBOOST_net_385;
wire n_31226;
wire n_31227;
wire n_31228;
wire n_31229;
wire n_3123;
wire n_31230;
wire n_31231;
wire n_31232;
wire n_31233;
wire n_31234;
wire n_31236;
wire n_31237;
wire n_31239;
wire n_3124;
wire n_31241;
wire n_31242;
wire n_31243;
wire n_31244;
wire n_31245;
wire n_31246;
wire n_31249;
wire n_3125;
wire n_31251;
wire n_31253;
wire n_31254;
wire n_31255;
wire n_31256;
wire n_31257;
wire n_31258;
wire n_31259;
wire n_3126;
wire n_31260;
wire n_31261;
wire n_31262;
wire n_31263;
wire n_31264;
wire n_31265;
wire TIMEBOOST_net_2090;
wire n_31267;
wire n_31268;
wire n_31269;
wire n_3127;
wire n_31270;
wire n_31271;
wire n_31272;
wire n_31273;
wire n_31275;
wire n_31276;
wire n_31277;
wire n_31279;
wire n_3128;
wire n_31280;
wire n_31281;
wire n_31282;
wire n_31283;
wire n_31284;
wire n_31285;
wire n_31286;
wire n_31287;
wire n_31288;
wire n_31289;
wire n_31290;
wire TIMEBOOST_net_1165;
wire n_31292;
wire n_31293;
wire n_31294;
wire n_31295;
wire n_31296;
wire n_31297;
wire n_31298;
wire TIMEBOOST_net_2920;
wire n_313;
wire n_3130;
wire n_31300;
wire n_31301;
wire n_31302;
wire n_31303;
wire n_31304;
wire n_31305;
wire n_31308;
wire n_3131;
wire n_31311;
wire n_31312;
wire n_31313;
wire n_31314;
wire n_31315;
wire n_31316;
wire n_31317;
wire n_31318;
wire n_31319;
wire n_3132;
wire n_31320;
wire n_31321;
wire n_31322;
wire n_31323;
wire n_31324;
wire n_31325;
wire n_31326;
wire n_31327;
wire n_31328;
wire n_31329;
wire n_3133;
wire n_31330;
wire n_31331;
wire n_31332;
wire n_31333;
wire n_31334;
wire n_31335;
wire n_31336;
wire n_31338;
wire n_31339;
wire n_31340;
wire n_31341;
wire n_31342;
wire n_31343;
wire n_31344;
wire n_31345;
wire n_31346;
wire n_31347;
wire n_31348;
wire n_31349;
wire n_3135;
wire n_31350;
wire n_31351;
wire n_31352;
wire n_31353;
wire n_31354;
wire n_31355;
wire n_31356;
wire n_31357;
wire n_31358;
wire n_31359;
wire n_31360;
wire n_31361;
wire n_31363;
wire n_31365;
wire n_31368;
wire n_31369;
wire n_3137;
wire n_31370;
wire n_31371;
wire n_31372;
wire n_31374;
wire n_31375;
wire n_31376;
wire n_31377;
wire n_31379;
wire n_3138;
wire n_31380;
wire n_31381;
wire n_31382;
wire n_31383;
wire TIMEBOOST_net_2715;
wire n_31385;
wire n_31386;
wire n_31387;
wire n_31388;
wire n_31389;
wire n_31390;
wire n_31391;
wire n_31392;
wire n_31393;
wire n_31394;
wire n_31395;
wire n_31396;
wire n_31397;
wire TIMEBOOST_net_1764;
wire n_31399;
wire n_314;
wire n_3140;
wire n_31400;
wire n_31401;
wire n_31402;
wire n_31403;
wire n_31404;
wire n_31405;
wire n_31407;
wire n_31408;
wire n_31409;
wire n_3141;
wire n_31410;
wire n_31411;
wire n_31412;
wire n_31414;
wire n_31415;
wire n_31416;
wire n_31417;
wire n_31418;
wire n_31419;
wire n_3142;
wire n_31420;
wire n_31421;
wire TIMEBOOST_net_572;
wire n_31424;
wire n_31425;
wire n_31426;
wire n_31428;
wire n_31429;
wire n_31430;
wire n_31431;
wire n_31432;
wire n_31433;
wire n_31434;
wire n_31435;
wire n_31437;
wire n_31438;
wire n_31439;
wire n_31440;
wire n_31441;
wire n_31442;
wire n_31443;
wire n_31445;
wire n_31446;
wire n_31447;
wire n_31448;
wire n_31449;
wire TIMEBOOST_net_1096;
wire n_31453;
wire n_31454;
wire n_31455;
wire n_31456;
wire n_31457;
wire n_31458;
wire n_31459;
wire n_31460;
wire n_31461;
wire n_31462;
wire n_31463;
wire n_31465;
wire n_31466;
wire n_31467;
wire n_31468;
wire n_31469;
wire n_3147;
wire n_31470;
wire n_31471;
wire n_31472;
wire n_31473;
wire n_31474;
wire n_31475;
wire n_31476;
wire n_31477;
wire n_3148;
wire n_31481;
wire n_31482;
wire n_31483;
wire n_31484;
wire n_31485;
wire n_31486;
wire n_31487;
wire n_31488;
wire n_31489;
wire n_3149;
wire n_31490;
wire n_31491;
wire n_31492;
wire n_31494;
wire n_31497;
wire n_31498;
wire n_31499;
wire n_315;
wire n_3150;
wire n_31500;
wire n_31501;
wire n_31502;
wire n_31504;
wire TIMEBOOST_net_1396;
wire n_31506;
wire n_31508;
wire n_31509;
wire n_3151;
wire n_31510;
wire n_31511;
wire n_31512;
wire n_31513;
wire n_31514;
wire n_31515;
wire n_31518;
wire n_31519;
wire n_3152;
wire n_31520;
wire n_31521;
wire n_31522;
wire n_31523;
wire n_31524;
wire n_31525;
wire n_31526;
wire n_31527;
wire n_31528;
wire n_31529;
wire n_31530;
wire n_31532;
wire n_31533;
wire n_31534;
wire n_31535;
wire n_31536;
wire n_31537;
wire n_31538;
wire n_3154;
wire n_31540;
wire n_31541;
wire n_31542;
wire n_31543;
wire n_31544;
wire n_31545;
wire n_31546;
wire n_31547;
wire n_31548;
wire n_31549;
wire n_3155;
wire n_31550;
wire n_31551;
wire n_31553;
wire n_31554;
wire TIMEBOOST_net_1508;
wire n_31556;
wire n_31557;
wire n_31558;
wire n_31559;
wire n_3156;
wire n_31560;
wire n_31561;
wire n_31563;
wire n_31564;
wire n_31565;
wire n_31567;
wire n_31568;
wire n_31569;
wire n_3157;
wire n_31570;
wire n_31571;
wire n_31572;
wire n_31573;
wire n_31574;
wire n_31576;
wire n_31577;
wire n_31578;
wire n_31579;
wire n_3158;
wire n_31580;
wire n_31581;
wire n_31582;
wire n_31583;
wire n_31584;
wire n_31585;
wire n_31586;
wire n_31587;
wire n_31588;
wire n_31589;
wire n_3159;
wire n_31591;
wire n_31593;
wire n_31594;
wire n_31599;
wire n_316;
wire n_3160;
wire TIMEBOOST_net_730;
wire n_31605;
wire n_31606;
wire n_31607;
wire n_31608;
wire n_31609;
wire n_3161;
wire n_31610;
wire n_31611;
wire n_31612;
wire n_31613;
wire n_31614;
wire n_31615;
wire n_31616;
wire n_31617;
wire n_31618;
wire n_31619;
wire n_31620;
wire n_31621;
wire n_31622;
wire n_31623;
wire n_31624;
wire n_31625;
wire n_31626;
wire n_31627;
wire n_31628;
wire n_31629;
wire n_3163;
wire n_31630;
wire n_31631;
wire n_31632;
wire n_31633;
wire n_31634;
wire n_31635;
wire n_31636;
wire n_31637;
wire n_31638;
wire n_31639;
wire n_3164;
wire n_31640;
wire n_31641;
wire n_31642;
wire n_31643;
wire n_31644;
wire n_31645;
wire n_31646;
wire n_31647;
wire n_31648;
wire n_31649;
wire n_3165;
wire n_31652;
wire n_31653;
wire n_31655;
wire TIMEBOOST_net_1804;
wire TIMEBOOST_net_266;
wire n_31664;
wire n_31666;
wire n_31667;
wire n_31668;
wire n_31669;
wire n_3167;
wire n_31670;
wire n_31671;
wire n_31672;
wire n_31673;
wire n_31676;
wire n_31677;
wire n_31678;
wire TIMEBOOST_net_741;
wire n_31681;
wire n_31682;
wire n_31683;
wire n_31684;
wire n_31685;
wire n_31686;
wire n_31687;
wire n_31688;
wire n_31689;
wire n_3169;
wire n_31690;
wire n_31691;
wire n_31692;
wire n_31693;
wire n_31697;
wire n_31698;
wire n_31699;
wire n_317;
wire n_3170;
wire n_31700;
wire n_31701;
wire n_31702;
wire n_31703;
wire n_31704;
wire n_31705;
wire n_31706;
wire n_31708;
wire n_31709;
wire n_31713;
wire n_31714;
wire n_31715;
wire n_31716;
wire n_31718;
wire n_31719;
wire n_3172;
wire n_31720;
wire n_31721;
wire n_31725;
wire n_31727;
wire n_31729;
wire n_3173;
wire n_31730;
wire TIMEBOOST_net_740;
wire TIMEBOOST_net_739;
wire n_31735;
wire n_31736;
wire n_31737;
wire n_31738;
wire n_3174;
wire n_31740;
wire TIMEBOOST_net_576;
wire n_31742;
wire n_31743;
wire n_31744;
wire n_31745;
wire n_31746;
wire n_31747;
wire n_31748;
wire n_3175;
wire n_31750;
wire n_31751;
wire n_31752;
wire n_31754;
wire n_31755;
wire n_31756;
wire TIMEBOOST_net_1811;
wire TIMEBOOST_net_1810;
wire n_31759;
wire n_3176;
wire n_31760;
wire TIMEBOOST_net_1809;
wire n_31763;
wire n_31764;
wire n_31765;
wire n_31766;
wire n_31768;
wire n_31769;
wire n_3177;
wire n_31770;
wire TIMEBOOST_net_577;
wire n_31773;
wire n_31774;
wire n_31775;
wire n_31776;
wire n_31777;
wire n_31778;
wire n_31779;
wire n_31780;
wire n_31781;
wire n_31782;
wire n_31783;
wire n_31784;
wire n_31785;
wire TIMEBOOST_net_742;
wire n_31787;
wire n_31788;
wire n_3179;
wire n_31791;
wire n_31793;
wire n_31794;
wire n_31795;
wire n_31796;
wire n_31797;
wire n_31799;
wire n_318;
wire n_31800;
wire n_31801;
wire n_31802;
wire n_31803;
wire n_31804;
wire n_31805;
wire n_31806;
wire n_31807;
wire n_31808;
wire n_31809;
wire n_31810;
wire n_31813;
wire TIMEBOOST_net_737;
wire n_31815;
wire n_31816;
wire n_31819;
wire n_31821;
wire n_31823;
wire n_31824;
wire n_31825;
wire n_31826;
wire n_31827;
wire n_31828;
wire n_31829;
wire n_3183;
wire n_31830;
wire n_31831;
wire n_31832;
wire n_31833;
wire n_31834;
wire n_31835;
wire n_31836;
wire n_31837;
wire n_31838;
wire n_31839;
wire n_3184;
wire n_31840;
wire n_31841;
wire n_31842;
wire n_31843;
wire TIMEBOOST_net_2115;
wire n_31847;
wire n_31848;
wire n_3185;
wire n_31850;
wire n_31851;
wire n_31852;
wire n_31853;
wire n_31854;
wire n_31855;
wire n_31856;
wire TIMEBOOST_net_1219;
wire n_31858;
wire n_31859;
wire n_3186;
wire n_31861;
wire n_31862;
wire n_31863;
wire n_31864;
wire n_31868;
wire n_31869;
wire TIMEBOOST_net_1129;
wire n_31871;
wire n_31872;
wire n_31875;
wire n_31876;
wire n_31877;
wire n_31878;
wire n_31879;
wire n_31880;
wire n_31881;
wire n_31882;
wire n_31883;
wire n_31884;
wire n_31885;
wire n_31886;
wire n_31887;
wire n_31888;
wire n_3189;
wire n_31893;
wire n_31894;
wire n_31895;
wire n_31896;
wire n_31897;
wire n_31898;
wire n_319;
wire n_3190;
wire n_31902;
wire n_31903;
wire TIMEBOOST_net_583;
wire TIMEBOOST_net_2495;
wire TIMEBOOST_net_1779;
wire TIMEBOOST_net_1422;
wire n_31908;
wire n_31909;
wire n_3191;
wire n_31910;
wire n_31911;
wire n_31912;
wire n_31913;
wire n_31914;
wire n_31915;
wire n_31916;
wire n_31919;
wire n_3192;
wire n_31920;
wire n_31929;
wire TIMEBOOST_net_2648;
wire n_31930;
wire n_31931;
wire n_31932;
wire n_31934;
wire n_31935;
wire n_31936;
wire n_31937;
wire n_31938;
wire n_31939;
wire n_3194;
wire n_31940;
wire n_31941;
wire n_31947;
wire n_31948;
wire n_31949;
wire n_3195;
wire n_31951;
wire TIMEBOOST_net_2781;
wire n_31953;
wire n_31954;
wire n_31955;
wire n_31956;
wire n_31958;
wire n_31959;
wire n_3196;
wire n_31960;
wire n_31966;
wire n_31967;
wire n_31968;
wire n_31969;
wire n_31970;
wire n_31971;
wire n_31972;
wire n_31974;
wire n_31975;
wire n_31976;
wire n_31977;
wire n_31978;
wire n_31979;
wire n_3198;
wire n_31980;
wire n_31981;
wire n_31988;
wire n_31989;
wire n_3199;
wire n_31990;
wire n_31991;
wire n_31992;
wire n_31993;
wire n_31994;
wire n_31996;
wire TIMEBOOST_net_667;
wire n_31998;
wire n_31999;
wire n_320;
wire n_3200;
wire n_32000;
wire n_32001;
wire n_32002;
wire n_32003;
wire n_32004;
wire n_32005;
wire n_32006;
wire n_32007;
wire n_32008;
wire TIMEBOOST_net_1782;
wire TIMEBOOST_net_1781;
wire TIMEBOOST_net_2087;
wire n_3202;
wire n_32020;
wire n_32021;
wire n_32024;
wire n_32026;
wire n_32027;
wire n_32028;
wire n_32029;
wire n_32032;
wire n_32033;
wire n_32034;
wire n_32035;
wire n_3204;
wire n_32044;
wire n_32046;
wire TIMEBOOST_net_1353;
wire n_3205;
wire n_32051;
wire n_32052;
wire TIMEBOOST_net_771;
wire n_32055;
wire TIMEBOOST_net_581;
wire n_32057;
wire n_32058;
wire n_32060;
wire n_32061;
wire n_32063;
wire n_32064;
wire n_32065;
wire n_32068;
wire n_3207;
wire n_32070;
wire n_32072;
wire n_32075;
wire n_32076;
wire n_32077;
wire n_32079;
wire n_3208;
wire n_32081;
wire n_32082;
wire n_32083;
wire n_32085;
wire n_32086;
wire n_32087;
wire n_32088;
wire n_32089;
wire n_3209;
wire n_32090;
wire n_32093;
wire n_32094;
wire n_32098;
wire n_32099;
wire n_321;
wire n_3210;
wire n_32100;
wire n_32101;
wire n_32102;
wire n_32103;
wire n_32104;
wire n_32106;
wire n_32107;
wire n_32108;
wire n_32109;
wire n_3211;
wire n_32110;
wire n_32111;
wire n_32112;
wire n_32113;
wire n_32114;
wire n_32115;
wire n_32116;
wire n_32118;
wire n_32119;
wire n_3212;
wire n_32120;
wire n_32122;
wire n_32123;
wire n_32124;
wire n_32125;
wire n_32126;
wire n_32127;
wire n_32128;
wire n_32129;
wire n_3213;
wire n_32130;
wire n_32132;
wire n_32133;
wire n_32134;
wire n_32135;
wire n_32136;
wire n_32137;
wire n_32138;
wire n_32139;
wire n_3214;
wire n_32142;
wire n_32143;
wire n_32145;
wire n_32147;
wire TIMEBOOST_net_753;
wire n_32149;
wire n_3215;
wire n_32150;
wire n_32151;
wire n_32152;
wire n_32154;
wire n_32156;
wire n_32157;
wire n_32158;
wire n_3216;
wire n_32161;
wire n_32162;
wire n_32163;
wire n_32164;
wire n_32168;
wire n_32169;
wire n_3217;
wire n_32170;
wire n_32171;
wire n_32172;
wire n_32173;
wire n_32174;
wire n_32175;
wire n_32176;
wire n_32178;
wire n_3218;
wire n_32180;
wire n_32182;
wire n_32183;
wire n_32184;
wire n_32185;
wire n_32186;
wire n_32187;
wire n_32188;
wire n_32189;
wire n_32190;
wire n_32191;
wire n_32192;
wire n_32195;
wire n_32196;
wire n_32197;
wire n_32198;
wire n_322;
wire n_3220;
wire n_32200;
wire n_32201;
wire n_32202;
wire n_32203;
wire n_32204;
wire n_32205;
wire n_32206;
wire n_32207;
wire n_32208;
wire n_32209;
wire n_32210;
wire n_32211;
wire n_32214;
wire n_32215;
wire n_32216;
wire n_32218;
wire n_32219;
wire n_3222;
wire n_32220;
wire TIMEBOOST_net_755;
wire n_32222;
wire n_32223;
wire n_32224;
wire n_32225;
wire n_32226;
wire n_32227;
wire n_32228;
wire n_32229;
wire TIMEBOOST_net_2383;
wire n_32230;
wire n_32231;
wire n_32232;
wire n_32234;
wire n_32235;
wire n_32236;
wire n_32237;
wire n_32238;
wire n_32239;
wire n_3224;
wire n_32240;
wire n_32241;
wire n_32242;
wire n_32243;
wire n_32244;
wire n_32245;
wire n_32247;
wire n_32248;
wire n_32249;
wire n_3225;
wire n_32250;
wire n_32251;
wire n_32252;
wire n_32254;
wire n_32255;
wire n_32256;
wire n_32257;
wire n_32258;
wire n_32259;
wire n_32260;
wire n_32261;
wire n_32262;
wire n_32263;
wire TIMEBOOST_net_2280;
wire n_32266;
wire n_32269;
wire n_3227;
wire n_32271;
wire n_32272;
wire n_32273;
wire n_32274;
wire n_32275;
wire n_32276;
wire n_32277;
wire n_32278;
wire n_32279;
wire n_3228;
wire n_32280;
wire n_32281;
wire n_32283;
wire n_32285;
wire n_32286;
wire n_32287;
wire n_32288;
wire n_32289;
wire n_3229;
wire n_32290;
wire n_32291;
wire n_32292;
wire n_32293;
wire n_32294;
wire n_32295;
wire n_32296;
wire n_323;
wire n_32300;
wire n_32301;
wire TIMEBOOST_net_710;
wire n_32303;
wire n_32304;
wire n_32305;
wire n_3231;
wire n_32310;
wire n_32311;
wire n_32312;
wire n_32313;
wire n_32314;
wire n_32315;
wire n_32316;
wire n_32318;
wire n_32319;
wire n_3232;
wire n_32324;
wire n_32325;
wire n_32326;
wire n_3233;
wire n_32330;
wire n_32333;
wire n_32334;
wire n_32335;
wire n_32336;
wire n_32337;
wire n_32338;
wire n_32339;
wire n_32340;
wire n_32341;
wire n_32342;
wire n_32343;
wire n_32346;
wire n_32347;
wire n_32348;
wire n_32349;
wire n_32350;
wire n_32352;
wire n_32353;
wire n_32354;
wire n_32355;
wire n_32356;
wire n_32357;
wire n_32358;
wire n_3236;
wire n_32360;
wire n_32362;
wire n_32363;
wire n_32364;
wire n_32365;
wire n_32366;
wire n_32367;
wire TIMEBOOST_net_1638;
wire n_32370;
wire n_32373;
wire n_32374;
wire n_32375;
wire n_32376;
wire n_32377;
wire n_32378;
wire n_32379;
wire n_3238;
wire n_32380;
wire n_32381;
wire n_32382;
wire n_32384;
wire n_32387;
wire n_32388;
wire n_32389;
wire n_3239;
wire n_32390;
wire n_32391;
wire n_32392;
wire n_32394;
wire n_32395;
wire n_32399;
wire n_324;
wire n_3240;
wire n_32402;
wire n_32403;
wire n_32404;
wire n_32405;
wire n_32406;
wire n_32407;
wire n_32408;
wire n_32409;
wire n_3241;
wire n_32410;
wire n_32411;
wire n_32412;
wire n_32413;
wire n_32414;
wire n_32415;
wire n_32416;
wire n_32417;
wire n_32418;
wire n_32419;
wire n_3242;
wire n_32420;
wire n_32421;
wire n_32422;
wire n_32423;
wire n_32424;
wire n_32425;
wire n_32426;
wire n_32427;
wire n_32428;
wire n_3243;
wire n_32431;
wire n_32432;
wire n_32433;
wire TIMEBOOST_net_1433;
wire n_32436;
wire TIMEBOOST_net_795;
wire n_32439;
wire n_3244;
wire n_32440;
wire n_32441;
wire n_32442;
wire n_32443;
wire n_32444;
wire n_32445;
wire n_32446;
wire n_32447;
wire n_32448;
wire n_32449;
wire n_3245;
wire n_32450;
wire n_32451;
wire n_32452;
wire n_32453;
wire n_32454;
wire n_32455;
wire n_32456;
wire n_32457;
wire n_32458;
wire n_32459;
wire n_3246;
wire n_32460;
wire n_32461;
wire n_32462;
wire n_32463;
wire n_32464;
wire n_32466;
wire n_32467;
wire n_32468;
wire n_32469;
wire n_32471;
wire n_32472;
wire n_32473;
wire TIMEBOOST_net_22;
wire n_32479;
wire n_3248;
wire n_32480;
wire n_32481;
wire n_32482;
wire n_32483;
wire n_32484;
wire n_32485;
wire n_32486;
wire n_32487;
wire n_32488;
wire n_32489;
wire n_32490;
wire n_32491;
wire n_32492;
wire n_32493;
wire n_32494;
wire n_32495;
wire n_32496;
wire n_32497;
wire n_32498;
wire n_32499;
wire n_325;
wire n_3250;
wire n_32500;
wire n_32501;
wire n_32502;
wire n_32503;
wire n_32504;
wire n_32505;
wire n_32506;
wire n_32507;
wire n_32508;
wire n_32509;
wire n_32510;
wire n_32511;
wire n_32513;
wire n_32515;
wire n_32516;
wire n_32517;
wire n_32518;
wire n_32519;
wire TIMEBOOST_net_267;
wire n_32520;
wire n_32521;
wire n_32522;
wire n_32523;
wire n_32525;
wire TIMEBOOST_net_1432;
wire n_32529;
wire n_32530;
wire n_32531;
wire n_32532;
wire n_32533;
wire n_32534;
wire n_32535;
wire n_32536;
wire n_32537;
wire n_32538;
wire n_32539;
wire n_3254;
wire n_32540;
wire n_32541;
wire n_32542;
wire n_32543;
wire n_32545;
wire n_32546;
wire n_32547;
wire n_32548;
wire n_32549;
wire n_3255;
wire n_32551;
wire n_32552;
wire n_32553;
wire n_32554;
wire n_32555;
wire n_32556;
wire n_32557;
wire n_32558;
wire n_32559;
wire n_32560;
wire n_32561;
wire n_32562;
wire n_32563;
wire n_32564;
wire n_32565;
wire n_32566;
wire n_32567;
wire n_32568;
wire n_32569;
wire n_3257;
wire n_32571;
wire n_32572;
wire n_32573;
wire n_32574;
wire n_32575;
wire n_32577;
wire n_32578;
wire n_32579;
wire n_3258;
wire n_32582;
wire n_32583;
wire n_32584;
wire n_32585;
wire n_32586;
wire n_32587;
wire n_32588;
wire n_32589;
wire n_3259;
wire n_32590;
wire TIMEBOOST_net_10;
wire n_32594;
wire n_32595;
wire n_32596;
wire n_32597;
wire n_32598;
wire n_32599;
wire n_326;
wire n_3260;
wire n_32600;
wire n_32601;
wire n_32602;
wire n_32603;
wire n_32604;
wire n_32605;
wire n_32606;
wire n_32607;
wire n_32608;
wire TIMEBOOST_net_2639;
wire n_3261;
wire n_32610;
wire n_32611;
wire n_32613;
wire n_32615;
wire n_32616;
wire n_32617;
wire n_32621;
wire n_32622;
wire n_32623;
wire n_32624;
wire n_32625;
wire n_32626;
wire n_32627;
wire n_32628;
wire TIMEBOOST_net_2331;
wire n_3263;
wire n_32630;
wire TIMEBOOST_net_1454;
wire n_32632;
wire n_32634;
wire n_32635;
wire n_32637;
wire n_32638;
wire n_3264;
wire n_32641;
wire n_32643;
wire n_32645;
wire n_32646;
wire n_32647;
wire n_32649;
wire n_3265;
wire n_32651;
wire n_32652;
wire n_32653;
wire n_32654;
wire n_32655;
wire n_32656;
wire n_32657;
wire n_32658;
wire n_32659;
wire n_32660;
wire n_32661;
wire n_32662;
wire n_32663;
wire n_32664;
wire n_32665;
wire n_32666;
wire n_32667;
wire n_32668;
wire n_32669;
wire n_32670;
wire n_32671;
wire n_32672;
wire n_32674;
wire n_32675;
wire n_32676;
wire n_32677;
wire n_32678;
wire n_32679;
wire n_32680;
wire n_32682;
wire n_32683;
wire n_32684;
wire n_32687;
wire n_32688;
wire n_32689;
wire TIMEBOOST_net_360;
wire n_32690;
wire TIMEBOOST_net_807;
wire n_32692;
wire n_32693;
wire n_32694;
wire n_32695;
wire n_32696;
wire n_32697;
wire n_32698;
wire n_32699;
wire n_327;
wire n_3270;
wire n_32701;
wire n_32702;
wire n_32704;
wire n_32706;
wire n_32708;
wire n_32709;
wire n_3271;
wire n_32711;
wire n_32714;
wire n_32715;
wire n_32716;
wire n_32717;
wire n_32718;
wire n_32719;
wire n_3272;
wire n_32720;
wire n_32721;
wire n_32722;
wire n_32723;
wire n_32724;
wire n_32725;
wire n_32726;
wire n_32727;
wire n_32728;
wire n_32729;
wire n_3273;
wire n_32730;
wire n_32731;
wire n_32732;
wire n_32733;
wire n_32734;
wire n_32735;
wire n_32736;
wire n_3274;
wire n_32740;
wire n_32741;
wire TIMEBOOST_net_865;
wire n_32743;
wire TIMEBOOST_net_2896;
wire n_32746;
wire n_32747;
wire n_32748;
wire n_32749;
wire n_3275;
wire n_32750;
wire n_32751;
wire n_32752;
wire n_32754;
wire n_32755;
wire n_32756;
wire n_32757;
wire n_32758;
wire n_32759;
wire TIMEBOOST_net_1639;
wire n_32761;
wire n_32762;
wire n_32763;
wire n_32764;
wire n_32765;
wire n_32766;
wire n_32767;
wire n_32768;
wire n_32769;
wire TIMEBOOST_net_2456;
wire n_32770;
wire n_32772;
wire n_32773;
wire n_32774;
wire n_32775;
wire n_32776;
wire n_32777;
wire n_32778;
wire n_32779;
wire n_32780;
wire n_32781;
wire n_32782;
wire n_32783;
wire n_32784;
wire n_32786;
wire n_32787;
wire n_32788;
wire n_32789;
wire n_3279;
wire n_32791;
wire n_32792;
wire n_32793;
wire n_32794;
wire n_32796;
wire n_32797;
wire n_32798;
wire n_32799;
wire n_328;
wire n_3280;
wire n_32800;
wire n_32801;
wire n_32802;
wire n_32803;
wire n_32804;
wire n_32805;
wire n_32806;
wire n_32807;
wire n_32808;
wire n_32809;
wire n_3281;
wire n_32810;
wire n_32811;
wire n_32812;
wire n_32813;
wire n_32814;
wire n_32815;
wire n_32816;
wire n_32817;
wire n_32818;
wire n_3282;
wire n_32820;
wire n_32821;
wire n_32822;
wire n_32823;
wire n_32824;
wire n_32825;
wire n_32826;
wire n_32827;
wire n_32829;
wire n_32830;
wire n_32831;
wire n_32832;
wire n_32833;
wire n_32834;
wire n_32835;
wire n_32837;
wire n_32838;
wire n_32839;
wire n_32840;
wire n_32841;
wire n_32842;
wire n_32843;
wire TIMEBOOST_net_791;
wire n_32845;
wire n_32846;
wire n_32847;
wire n_32848;
wire n_32849;
wire n_3285;
wire n_32850;
wire n_32851;
wire TIMEBOOST_net_1486;
wire n_32853;
wire n_32854;
wire n_32855;
wire n_32856;
wire n_32857;
wire n_3286;
wire n_32860;
wire n_32861;
wire n_32862;
wire n_32863;
wire n_32864;
wire n_32865;
wire n_32866;
wire n_32867;
wire n_32868;
wire TIMEBOOST_net_2344;
wire n_32870;
wire n_32871;
wire n_32875;
wire n_32876;
wire n_32877;
wire n_32878;
wire n_32879;
wire TIMEBOOST_net_270;
wire TIMEBOOST_net_1480;
wire n_32881;
wire n_32882;
wire n_32883;
wire n_32884;
wire n_32885;
wire n_32886;
wire n_32887;
wire n_32888;
wire n_32889;
wire TIMEBOOST_net_868;
wire n_32893;
wire n_32894;
wire n_32895;
wire n_32897;
wire n_32898;
wire n_32899;
wire n_329;
wire n_32900;
wire n_32901;
wire n_32902;
wire n_32903;
wire n_32904;
wire n_32905;
wire n_32906;
wire TIMEBOOST_net_37;
wire n_32908;
wire n_3291;
wire n_32911;
wire n_32912;
wire n_32914;
wire n_32915;
wire n_32916;
wire n_32918;
wire n_32919;
wire n_32920;
wire TIMEBOOST_net_61;
wire n_32923;
wire n_32924;
wire n_32925;
wire n_32926;
wire n_32927;
wire n_32928;
wire TIMEBOOST_net_2952;
wire n_3293;
wire TIMEBOOST_net_2918;
wire n_32931;
wire n_32934;
wire n_32935;
wire n_32936;
wire n_32939;
wire n_3294;
wire n_32940;
wire n_32941;
wire n_32942;
wire n_32943;
wire n_32944;
wire TIMEBOOST_net_2014;
wire n_32947;
wire n_32948;
wire n_32949;
wire TIMEBOOST_net_2438;
wire n_32951;
wire n_32952;
wire n_32953;
wire n_32954;
wire n_32955;
wire n_32957;
wire n_32959;
wire n_3296;
wire n_32961;
wire n_32962;
wire n_32963;
wire TIMEBOOST_net_905;
wire n_32966;
wire n_32967;
wire n_32968;
wire n_32969;
wire n_3297;
wire n_32970;
wire n_32971;
wire n_32972;
wire n_32973;
wire n_32974;
wire n_32975;
wire n_32976;
wire n_32977;
wire n_32978;
wire n_3298;
wire n_32980;
wire n_32981;
wire n_32982;
wire n_32983;
wire n_32984;
wire n_32985;
wire n_32986;
wire n_32988;
wire n_32989;
wire n_3299;
wire n_32990;
wire n_32991;
wire TIMEBOOST_net_914;
wire n_32994;
wire n_32995;
wire n_32996;
wire n_32997;
wire n_32999;
wire n_330;
wire n_3300;
wire n_33000;
wire n_33001;
wire n_33003;
wire n_33004;
wire n_33005;
wire n_33007;
wire n_33010;
wire n_33011;
wire n_33012;
wire n_33013;
wire n_33014;
wire n_33015;
wire n_33016;
wire n_33017;
wire n_33019;
wire n_3302;
wire n_33020;
wire n_33021;
wire n_33022;
wire n_33023;
wire n_33025;
wire n_33026;
wire n_33027;
wire n_33028;
wire n_33029;
wire n_3303;
wire n_33030;
wire n_33032;
wire n_33033;
wire n_33036;
wire n_33037;
wire n_33038;
wire n_33039;
wire n_3304;
wire n_33040;
wire n_33041;
wire n_33042;
wire n_33043;
wire n_33044;
wire n_33045;
wire n_33046;
wire n_33047;
wire n_33048;
wire n_3305;
wire n_33052;
wire n_33053;
wire n_33055;
wire n_33056;
wire n_33057;
wire n_33058;
wire n_33059;
wire n_3306;
wire n_33060;
wire n_33061;
wire TIMEBOOST_net_2002;
wire n_33063;
wire n_33065;
wire n_33066;
wire n_33067;
wire n_33068;
wire n_33069;
wire n_3307;
wire n_33070;
wire n_33071;
wire n_33072;
wire n_33073;
wire n_33075;
wire n_33077;
wire n_33078;
wire n_33079;
wire n_3308;
wire n_33080;
wire n_33081;
wire n_33082;
wire n_33083;
wire n_33084;
wire n_33085;
wire n_33086;
wire n_33088;
wire n_33089;
wire n_3309;
wire n_33090;
wire n_33091;
wire n_33092;
wire n_33093;
wire n_33097;
wire n_33098;
wire n_33099;
wire n_331;
wire n_3310;
wire n_33100;
wire n_33101;
wire n_33102;
wire n_33103;
wire n_33104;
wire n_33105;
wire n_33106;
wire n_33107;
wire n_33109;
wire n_33110;
wire n_33111;
wire n_33113;
wire n_33114;
wire n_33115;
wire n_33116;
wire n_33117;
wire n_33118;
wire n_33119;
wire n_3312;
wire n_33120;
wire n_33121;
wire n_33122;
wire n_33123;
wire n_33124;
wire n_33125;
wire n_33126;
wire n_33127;
wire n_33128;
wire n_33129;
wire n_3313;
wire n_33130;
wire n_33131;
wire n_33132;
wire n_33135;
wire n_33136;
wire n_33137;
wire n_3314;
wire n_33140;
wire n_33141;
wire n_33143;
wire n_33144;
wire n_33145;
wire n_33146;
wire n_33149;
wire n_3315;
wire n_33150;
wire n_33151;
wire n_33152;
wire n_33155;
wire n_33156;
wire n_33157;
wire n_33158;
wire n_33159;
wire n_3316;
wire n_33160;
wire n_33162;
wire n_33164;
wire n_33166;
wire n_33167;
wire n_33168;
wire n_33169;
wire n_3317;
wire n_33170;
wire n_33171;
wire n_33172;
wire n_33173;
wire n_33178;
wire n_33179;
wire n_3318;
wire n_33181;
wire n_33182;
wire n_33183;
wire n_33184;
wire n_33185;
wire n_33186;
wire n_33188;
wire n_33189;
wire n_3319;
wire n_33190;
wire n_33191;
wire n_33192;
wire n_33193;
wire n_33194;
wire n_33196;
wire n_33198;
wire n_33199;
wire n_332;
wire n_3320;
wire n_33200;
wire n_33201;
wire n_33202;
wire n_33203;
wire n_33204;
wire n_33205;
wire n_33206;
wire n_33207;
wire n_33208;
wire n_3321;
wire n_33210;
wire n_33211;
wire n_33213;
wire n_33215;
wire n_33216;
wire n_33217;
wire n_33218;
wire n_33219;
wire n_3322;
wire n_33220;
wire n_33221;
wire n_33222;
wire n_33223;
wire n_33224;
wire n_33225;
wire n_33227;
wire n_3323;
wire n_33231;
wire n_33233;
wire n_33234;
wire n_33235;
wire n_33236;
wire n_33237;
wire n_33239;
wire n_3324;
wire n_33240;
wire TIMEBOOST_net_66;
wire n_33242;
wire n_33246;
wire n_33247;
wire TIMEBOOST_net_2515;
wire n_33250;
wire n_33251;
wire n_33252;
wire n_33253;
wire n_33254;
wire n_33255;
wire n_33256;
wire TIMEBOOST_net_2160;
wire n_33258;
wire n_33259;
wire n_3326;
wire n_33260;
wire n_33261;
wire n_33262;
wire n_33263;
wire n_33264;
wire n_33265;
wire n_33266;
wire n_33267;
wire n_33268;
wire n_33269;
wire TIMEBOOST_net_2874;
wire n_33270;
wire n_33272;
wire n_33273;
wire n_33274;
wire n_33275;
wire n_33276;
wire TIMEBOOST_net_825;
wire n_33279;
wire n_3328;
wire n_33281;
wire n_33287;
wire n_33288;
wire n_33289;
wire n_3329;
wire n_33290;
wire n_33291;
wire n_33293;
wire n_33294;
wire n_33296;
wire n_33297;
wire n_33298;
wire n_33299;
wire n_333;
wire n_33300;
wire n_33301;
wire n_33302;
wire n_33303;
wire n_33304;
wire n_33305;
wire n_33306;
wire n_33307;
wire n_33308;
wire n_3331;
wire n_33310;
wire n_33311;
wire n_33312;
wire n_33313;
wire n_33314;
wire n_33316;
wire n_33317;
wire TIMEBOOST_net_1841;
wire n_3332;
wire n_33321;
wire n_33322;
wire n_33323;
wire n_33324;
wire n_33325;
wire n_33326;
wire n_33327;
wire n_33328;
wire n_33329;
wire n_3333;
wire n_33330;
wire n_33331;
wire n_33334;
wire n_33335;
wire n_33336;
wire n_33337;
wire n_33338;
wire n_33339;
wire n_3334;
wire n_33340;
wire n_33341;
wire n_33343;
wire n_33344;
wire n_33345;
wire n_33346;
wire n_33347;
wire n_3335;
wire n_33350;
wire n_33351;
wire n_33352;
wire n_33353;
wire n_33354;
wire n_33356;
wire n_33357;
wire n_33358;
wire n_33359;
wire n_3336;
wire n_33360;
wire n_33361;
wire n_33362;
wire n_33363;
wire n_33366;
wire n_33367;
wire n_33368;
wire n_3337;
wire n_33370;
wire n_33371;
wire n_33372;
wire n_33373;
wire n_33374;
wire n_33375;
wire n_33376;
wire n_33377;
wire n_33378;
wire n_33379;
wire n_3338;
wire n_33380;
wire n_33381;
wire n_33382;
wire n_33386;
wire TIMEBOOST_net_112;
wire n_33388;
wire n_3339;
wire n_33390;
wire n_33391;
wire n_33393;
wire n_33394;
wire n_33395;
wire n_33396;
wire n_33397;
wire TIMEBOOST_net_2726;
wire n_334;
wire n_3340;
wire n_33401;
wire n_33402;
wire n_33404;
wire n_33405;
wire n_33406;
wire n_33408;
wire n_33409;
wire n_33410;
wire n_33411;
wire n_33412;
wire n_33413;
wire n_33414;
wire n_33415;
wire n_33416;
wire n_33417;
wire n_33418;
wire n_33419;
wire n_33420;
wire n_33421;
wire n_33423;
wire n_33424;
wire n_33425;
wire n_33426;
wire n_33427;
wire n_33428;
wire n_33429;
wire n_3343;
wire TIMEBOOST_net_2872;
wire n_33434;
wire n_33437;
wire n_33438;
wire n_33440;
wire n_33441;
wire n_33442;
wire n_33443;
wire n_33444;
wire n_33445;
wire n_33446;
wire n_33447;
wire n_33448;
wire n_33449;
wire n_3345;
wire n_33450;
wire n_33451;
wire n_33452;
wire n_33454;
wire n_33455;
wire n_33456;
wire n_33457;
wire n_33458;
wire n_33459;
wire n_3346;
wire n_33461;
wire n_33462;
wire n_33463;
wire n_33464;
wire n_33465;
wire n_33467;
wire n_33468;
wire n_33469;
wire n_3347;
wire n_33470;
wire n_33471;
wire n_33472;
wire TIMEBOOST_net_2943;
wire n_33474;
wire n_33475;
wire n_33476;
wire n_33479;
wire n_33480;
wire n_33481;
wire n_33482;
wire n_33483;
wire n_33484;
wire n_33485;
wire n_33486;
wire n_33487;
wire n_33488;
wire n_33489;
wire n_3349;
wire n_33490;
wire n_33491;
wire n_33492;
wire n_33494;
wire n_33495;
wire n_33496;
wire n_33497;
wire n_33498;
wire n_33499;
wire n_335;
wire TIMEBOOST_net_2254;
wire n_33500;
wire n_33501;
wire n_33503;
wire n_33504;
wire n_33505;
wire n_33506;
wire n_33507;
wire n_33508;
wire n_3351;
wire n_33511;
wire n_33512;
wire n_33513;
wire n_33515;
wire n_33516;
wire n_33517;
wire n_33518;
wire n_33519;
wire n_3352;
wire n_33520;
wire n_33521;
wire n_33524;
wire n_33525;
wire n_33526;
wire n_33527;
wire n_33528;
wire n_33529;
wire n_3353;
wire n_33530;
wire TIMEBOOST_net_2721;
wire n_33532;
wire n_33533;
wire n_33534;
wire n_33535;
wire n_33536;
wire n_33537;
wire n_33539;
wire n_3354;
wire n_33540;
wire n_33541;
wire n_33542;
wire n_33544;
wire n_33545;
wire n_33546;
wire n_33547;
wire n_33549;
wire n_3355;
wire n_33550;
wire n_33552;
wire n_33553;
wire n_33554;
wire n_33556;
wire n_33557;
wire n_33558;
wire n_33559;
wire n_3356;
wire n_33560;
wire n_33561;
wire n_33562;
wire n_33564;
wire n_33567;
wire n_33568;
wire n_3357;
wire TIMEBOOST_net_2823;
wire n_33571;
wire n_33572;
wire n_33573;
wire TIMEBOOST_net_123;
wire n_33576;
wire n_33578;
wire n_33579;
wire n_3358;
wire n_33581;
wire n_33583;
wire n_33584;
wire n_33588;
wire n_33589;
wire TIMEBOOST_net_2221;
wire n_33590;
wire n_33591;
wire n_33592;
wire n_33594;
wire n_33595;
wire n_33596;
wire n_33599;
wire n_336;
wire n_3360;
wire n_33600;
wire n_33601;
wire n_33602;
wire n_33603;
wire n_33604;
wire n_33606;
wire n_33607;
wire n_33608;
wire n_33609;
wire n_3361;
wire n_33610;
wire TIMEBOOST_net_997;
wire n_33613;
wire n_33614;
wire n_33618;
wire n_3362;
wire n_33620;
wire n_33621;
wire n_33622;
wire TIMEBOOST_net_116;
wire n_33624;
wire n_33625;
wire n_33626;
wire n_33627;
wire n_33628;
wire n_33629;
wire n_3363;
wire n_33630;
wire n_33631;
wire n_33632;
wire n_33635;
wire n_33636;
wire n_33637;
wire n_33638;
wire n_33639;
wire n_3364;
wire n_33640;
wire n_33642;
wire n_33643;
wire n_33644;
wire TIMEBOOST_net_995;
wire n_33646;
wire TIMEBOOST_net_183;
wire n_33648;
wire n_3365;
wire n_33651;
wire n_33653;
wire n_33654;
wire n_33655;
wire n_33656;
wire n_33657;
wire n_33660;
wire n_33662;
wire n_33663;
wire n_33664;
wire n_33667;
wire n_33668;
wire n_3367;
wire n_33670;
wire n_33671;
wire n_33672;
wire n_33673;
wire n_33674;
wire n_33675;
wire n_33677;
wire n_3368;
wire n_33680;
wire n_33681;
wire n_33682;
wire n_33683;
wire n_33684;
wire n_33685;
wire n_33686;
wire n_33687;
wire n_33688;
wire n_33689;
wire n_3369;
wire n_33690;
wire n_33691;
wire n_33693;
wire n_33695;
wire n_33697;
wire TIMEBOOST_net_1799;
wire n_33699;
wire n_337;
wire n_3370;
wire n_33700;
wire n_33701;
wire n_33702;
wire n_33703;
wire n_33704;
wire n_33705;
wire n_33706;
wire n_33707;
wire n_33708;
wire TIMEBOOST_net_273;
wire n_33711;
wire n_33714;
wire n_33715;
wire n_33717;
wire n_33718;
wire n_33719;
wire n_3372;
wire n_33720;
wire n_33721;
wire n_33722;
wire n_33723;
wire n_33724;
wire n_33725;
wire n_33728;
wire n_33729;
wire n_3373;
wire n_33730;
wire n_33731;
wire n_33732;
wire n_33733;
wire n_33735;
wire n_33737;
wire n_33738;
wire n_33739;
wire n_33740;
wire n_33741;
wire n_33743;
wire n_33745;
wire n_33746;
wire n_33747;
wire n_33748;
wire n_3375;
wire n_33750;
wire n_33752;
wire n_33753;
wire TIMEBOOST_net_1560;
wire n_33756;
wire n_33757;
wire n_33758;
wire n_33759;
wire n_3376;
wire n_33760;
wire n_33761;
wire n_33762;
wire n_33763;
wire n_33764;
wire n_33765;
wire n_33768;
wire n_33769;
wire n_3377;
wire n_33771;
wire n_33772;
wire n_33773;
wire n_33775;
wire n_33776;
wire n_33777;
wire n_33778;
wire n_33779;
wire n_33780;
wire n_33781;
wire n_33782;
wire n_33784;
wire n_33785;
wire n_33787;
wire n_3379;
wire n_33792;
wire n_33793;
wire n_33794;
wire n_33795;
wire n_33796;
wire n_33797;
wire n_33798;
wire n_33799;
wire n_338;
wire n_3380;
wire n_33800;
wire n_33801;
wire n_33802;
wire n_33803;
wire n_33804;
wire n_33805;
wire TIMEBOOST_net_106;
wire n_33807;
wire n_33809;
wire n_3381;
wire n_33810;
wire n_33812;
wire n_33813;
wire n_33814;
wire n_33815;
wire n_33816;
wire n_33817;
wire TIMEBOOST_net_1859;
wire n_33820;
wire n_33825;
wire n_33826;
wire n_33827;
wire n_33829;
wire n_3383;
wire n_33830;
wire n_33831;
wire n_33832;
wire n_33833;
wire n_33834;
wire n_33835;
wire n_3384;
wire n_33840;
wire n_33841;
wire n_33842;
wire n_33843;
wire n_33844;
wire n_33846;
wire n_33847;
wire n_33849;
wire n_3385;
wire n_33850;
wire n_33851;
wire n_33852;
wire TIMEBOOST_net_1953;
wire n_33855;
wire TIMEBOOST_net_107;
wire TIMEBOOST_net_246;
wire n_3386;
wire n_33862;
wire n_33863;
wire n_33864;
wire n_33865;
wire n_33868;
wire TIMEBOOST_net_846;
wire n_3387;
wire n_33870;
wire n_33871;
wire n_33872;
wire n_33873;
wire n_33874;
wire n_33875;
wire n_33876;
wire n_33877;
wire n_33878;
wire n_33879;
wire n_3388;
wire n_33880;
wire n_33881;
wire n_33882;
wire n_33884;
wire n_33885;
wire n_33887;
wire n_33888;
wire n_33889;
wire n_3389;
wire n_33890;
wire n_33891;
wire n_33892;
wire n_33893;
wire n_33894;
wire n_33895;
wire n_33896;
wire n_33897;
wire n_33898;
wire n_339;
wire n_3390;
wire n_33900;
wire n_33901;
wire n_33903;
wire n_33904;
wire n_33905;
wire n_33906;
wire n_33907;
wire n_33908;
wire n_3391;
wire n_33910;
wire n_33911;
wire n_33912;
wire n_33913;
wire n_33914;
wire n_33917;
wire n_33918;
wire n_33919;
wire TIMEBOOST_net_2832;
wire TIMEBOOST_net_2169;
wire n_33922;
wire n_33923;
wire n_33924;
wire n_33925;
wire n_33926;
wire n_33927;
wire n_33928;
wire n_33929;
wire n_3393;
wire n_33930;
wire n_33931;
wire n_33932;
wire n_33933;
wire n_33934;
wire n_33937;
wire n_33938;
wire n_33939;
wire n_3394;
wire n_33940;
wire n_33942;
wire n_33944;
wire n_33945;
wire n_33946;
wire n_3395;
wire n_33950;
wire n_33951;
wire n_33952;
wire n_33953;
wire n_33954;
wire n_33955;
wire n_33956;
wire n_33957;
wire n_33958;
wire n_33959;
wire n_3396;
wire n_33960;
wire n_33961;
wire n_33962;
wire n_33963;
wire n_33964;
wire n_33965;
wire n_33966;
wire n_33967;
wire n_33968;
wire n_33969;
wire n_3397;
wire n_33970;
wire n_33971;
wire n_33972;
wire n_33974;
wire n_33975;
wire n_33976;
wire n_33977;
wire n_33978;
wire n_33979;
wire n_3398;
wire TIMEBOOST_net_1576;
wire n_33981;
wire n_33983;
wire n_33985;
wire n_33986;
wire n_33989;
wire n_33990;
wire n_33991;
wire n_33992;
wire n_33993;
wire n_33994;
wire n_33995;
wire n_33996;
wire n_33997;
wire n_33998;
wire n_33999;
wire n_340;
wire n_3400;
wire n_34000;
wire n_34001;
wire n_34003;
wire n_34005;
wire n_34006;
wire n_34007;
wire n_34008;
wire n_34009;
wire n_34010;
wire n_34011;
wire n_34013;
wire n_34014;
wire n_34015;
wire n_34016;
wire n_34017;
wire n_34019;
wire n_34020;
wire n_34021;
wire n_34022;
wire n_34023;
wire n_34026;
wire n_3403;
wire n_34030;
wire n_34031;
wire n_34032;
wire TIMEBOOST_net_1577;
wire n_34036;
wire n_34037;
wire n_34039;
wire n_3404;
wire n_34040;
wire n_34041;
wire n_34042;
wire n_34043;
wire n_34044;
wire n_34048;
wire n_34049;
wire n_3405;
wire n_34051;
wire n_34052;
wire n_34053;
wire n_34054;
wire n_34055;
wire n_34056;
wire n_34058;
wire n_34059;
wire n_3406;
wire n_34060;
wire n_34061;
wire n_34062;
wire n_34063;
wire n_34064;
wire n_34065;
wire n_34066;
wire n_34067;
wire n_34068;
wire n_34069;
wire n_3407;
wire n_34070;
wire n_34071;
wire n_34072;
wire n_34073;
wire n_34074;
wire n_34075;
wire n_34076;
wire n_34077;
wire n_34078;
wire n_34079;
wire n_3408;
wire n_34080;
wire n_34081;
wire n_34082;
wire n_34083;
wire n_34084;
wire n_34085;
wire n_34086;
wire n_34087;
wire n_34088;
wire n_34089;
wire n_3409;
wire n_34094;
wire n_34095;
wire n_34096;
wire n_34097;
wire n_34098;
wire n_341;
wire n_3410;
wire n_34100;
wire n_34101;
wire n_34102;
wire n_34103;
wire n_34104;
wire n_34105;
wire n_34106;
wire n_34107;
wire n_34108;
wire n_34109;
wire n_3411;
wire n_34110;
wire n_34111;
wire n_34113;
wire n_34114;
wire n_34115;
wire n_34116;
wire n_34117;
wire n_34118;
wire n_34119;
wire n_3412;
wire n_34120;
wire n_34121;
wire n_34122;
wire n_34123;
wire n_34124;
wire n_34126;
wire n_34127;
wire n_34128;
wire n_3413;
wire n_34130;
wire n_34131;
wire n_34132;
wire n_34134;
wire n_34135;
wire n_34136;
wire n_34137;
wire n_34138;
wire n_34139;
wire n_3414;
wire n_34140;
wire n_34141;
wire n_34143;
wire n_34144;
wire n_34145;
wire n_34146;
wire TIMEBOOST_net_2774;
wire n_34148;
wire n_34149;
wire n_3415;
wire n_34150;
wire n_34151;
wire n_34152;
wire n_34153;
wire n_34154;
wire n_34155;
wire n_34157;
wire n_34158;
wire n_3416;
wire n_34160;
wire n_34161;
wire n_34162;
wire n_34163;
wire n_34164;
wire n_34167;
wire n_34168;
wire n_34169;
wire n_3417;
wire n_34170;
wire n_34171;
wire n_34172;
wire n_34173;
wire n_34174;
wire n_34176;
wire n_34177;
wire n_34178;
wire n_34179;
wire n_3418;
wire n_34180;
wire n_34181;
wire n_34182;
wire n_34183;
wire n_34184;
wire n_34186;
wire n_34187;
wire n_34189;
wire n_3419;
wire n_34190;
wire n_34191;
wire n_34192;
wire n_34193;
wire n_34196;
wire n_34197;
wire n_34198;
wire n_34199;
wire n_342;
wire n_34200;
wire n_34201;
wire TIMEBOOST_net_2828;
wire n_34203;
wire n_34204;
wire n_34206;
wire TIMEBOOST_net_1083;
wire n_34209;
wire n_3421;
wire n_34210;
wire n_34211;
wire n_34212;
wire n_34219;
wire n_34220;
wire n_34221;
wire n_34222;
wire n_34223;
wire n_34224;
wire n_34225;
wire n_34226;
wire n_34227;
wire n_34228;
wire n_34229;
wire n_3423;
wire n_34230;
wire n_34231;
wire n_34232;
wire n_34233;
wire n_34234;
wire n_34238;
wire n_34239;
wire n_3424;
wire n_34241;
wire n_34242;
wire TIMEBOOST_net_302;
wire n_34245;
wire n_34246;
wire n_34247;
wire n_34248;
wire n_34249;
wire n_3425;
wire n_34250;
wire n_34251;
wire n_34252;
wire n_34253;
wire n_34256;
wire n_34258;
wire n_34259;
wire n_3426;
wire n_34261;
wire n_34262;
wire n_34263;
wire n_34264;
wire n_34265;
wire n_34266;
wire n_34267;
wire n_34272;
wire n_34273;
wire n_34274;
wire n_34275;
wire n_34276;
wire TIMEBOOST_net_1041;
wire n_34278;
wire n_3428;
wire n_34281;
wire n_34282;
wire n_34283;
wire n_34284;
wire n_34285;
wire n_34287;
wire n_34288;
wire n_34289;
wire n_3429;
wire n_34290;
wire n_34291;
wire n_34292;
wire n_34293;
wire n_34294;
wire n_34296;
wire n_34297;
wire n_34298;
wire n_34299;
wire n_343;
wire n_34300;
wire TIMEBOOST_net_2835;
wire n_34303;
wire n_34304;
wire n_34305;
wire TIMEBOOST_net_2391;
wire n_34307;
wire n_3431;
wire n_34310;
wire n_34311;
wire n_34313;
wire n_34314;
wire n_34315;
wire n_34316;
wire n_34317;
wire n_34318;
wire n_34319;
wire n_34320;
wire n_34321;
wire n_34322;
wire n_34323;
wire n_34324;
wire n_34325;
wire n_34326;
wire n_34327;
wire n_34328;
wire n_34329;
wire n_3433;
wire n_34330;
wire n_34331;
wire n_34332;
wire n_34333;
wire n_34334;
wire n_34335;
wire TIMEBOOST_net_1965;
wire n_34338;
wire n_34339;
wire n_3434;
wire n_34340;
wire n_34342;
wire n_34343;
wire n_34344;
wire n_34345;
wire n_34347;
wire n_34348;
wire n_34349;
wire n_3435;
wire n_34350;
wire n_34351;
wire n_34353;
wire n_34354;
wire n_34355;
wire n_34356;
wire n_34357;
wire n_34358;
wire n_34359;
wire n_3436;
wire n_34362;
wire n_34363;
wire n_34364;
wire n_34365;
wire n_34366;
wire n_34367;
wire n_34368;
wire n_3437;
wire n_34372;
wire n_34374;
wire n_34375;
wire n_34376;
wire n_34377;
wire n_34378;
wire n_34379;
wire n_34380;
wire n_34381;
wire n_34383;
wire n_34384;
wire n_34385;
wire n_34386;
wire n_34387;
wire n_34388;
wire n_34389;
wire n_3439;
wire n_34390;
wire n_34394;
wire n_34395;
wire n_34396;
wire n_34397;
wire n_34398;
wire n_34399;
wire n_344;
wire n_34401;
wire n_34402;
wire n_34403;
wire n_34404;
wire n_34405;
wire n_34406;
wire n_34409;
wire n_34412;
wire n_34413;
wire n_34414;
wire n_34415;
wire n_34417;
wire n_34418;
wire n_34419;
wire TIMEBOOST_net_1116;
wire n_34420;
wire n_34421;
wire n_34423;
wire n_34424;
wire n_34427;
wire n_34428;
wire n_34429;
wire n_34430;
wire n_34433;
wire n_34434;
wire n_34435;
wire n_34437;
wire n_34438;
wire n_34439;
wire n_3444;
wire n_34440;
wire n_34441;
wire n_34442;
wire n_34443;
wire n_34445;
wire n_34446;
wire n_34447;
wire n_34448;
wire n_34450;
wire n_34451;
wire n_34452;
wire n_34453;
wire n_34454;
wire n_34458;
wire n_34459;
wire n_34460;
wire n_34462;
wire n_34463;
wire n_34464;
wire n_34465;
wire n_34466;
wire n_34467;
wire n_3447;
wire n_34472;
wire n_34473;
wire n_34474;
wire n_34475;
wire n_34477;
wire n_34478;
wire n_34479;
wire n_3448;
wire n_34480;
wire n_34481;
wire n_34484;
wire n_34486;
wire n_34487;
wire n_34488;
wire n_34489;
wire n_3449;
wire n_34490;
wire n_34491;
wire n_34492;
wire n_34493;
wire n_34494;
wire n_34496;
wire n_34497;
wire n_34498;
wire n_34499;
wire n_345;
wire n_3450;
wire n_34500;
wire n_34506;
wire n_34507;
wire n_34509;
wire TIMEBOOST_net_1115;
wire TIMEBOOST_net_1092;
wire n_34511;
wire TIMEBOOST_net_2843;
wire n_34514;
wire n_34516;
wire n_34518;
wire n_34519;
wire n_3452;
wire n_34520;
wire n_34521;
wire n_34522;
wire n_34523;
wire n_34525;
wire n_34526;
wire n_34527;
wire n_34528;
wire n_34529;
wire n_3453;
wire TIMEBOOST_net_2854;
wire n_34532;
wire n_34533;
wire n_34534;
wire n_34535;
wire n_34536;
wire n_34537;
wire n_34538;
wire n_34539;
wire n_3454;
wire n_34540;
wire n_34541;
wire n_34542;
wire n_34544;
wire n_34545;
wire n_34546;
wire n_34547;
wire n_34549;
wire n_3455;
wire n_34550;
wire n_34551;
wire n_34552;
wire n_34553;
wire n_34554;
wire n_34558;
wire n_34559;
wire n_3456;
wire TIMEBOOST_net_1093;
wire n_34562;
wire n_34563;
wire n_34564;
wire n_34565;
wire n_34568;
wire n_34569;
wire n_3457;
wire n_34570;
wire n_34571;
wire n_34572;
wire n_34573;
wire n_34574;
wire n_34575;
wire n_34576;
wire n_34577;
wire n_34579;
wire n_3458;
wire n_34580;
wire n_34581;
wire n_34582;
wire n_34585;
wire n_34586;
wire n_34587;
wire n_3459;
wire n_34590;
wire n_34591;
wire n_34592;
wire n_34593;
wire n_34594;
wire n_34595;
wire n_34596;
wire n_34597;
wire n_34598;
wire TIMEBOOST_net_239;
wire n_346;
wire n_3460;
wire n_34600;
wire n_34601;
wire n_34602;
wire n_34603;
wire n_34604;
wire n_34605;
wire n_34606;
wire n_34607;
wire n_34608;
wire n_34609;
wire n_34610;
wire n_34611;
wire n_34612;
wire n_34613;
wire n_34614;
wire n_34615;
wire n_34616;
wire n_34617;
wire n_34618;
wire TIMEBOOST_net_2279;
wire n_34621;
wire n_34622;
wire n_34623;
wire n_34624;
wire n_34625;
wire n_34627;
wire n_34628;
wire n_34629;
wire n_34630;
wire n_34631;
wire n_34632;
wire n_34634;
wire n_34635;
wire n_34637;
wire n_34638;
wire n_34639;
wire TIMEBOOST_net_1624;
wire n_34640;
wire n_34641;
wire n_34642;
wire n_34643;
wire n_34644;
wire n_34645;
wire n_34646;
wire n_34648;
wire n_34649;
wire n_3465;
wire n_34650;
wire n_34651;
wire n_34652;
wire n_34653;
wire n_34654;
wire n_34655;
wire n_34656;
wire n_34657;
wire n_34658;
wire n_34659;
wire n_3466;
wire n_34660;
wire n_34661;
wire n_34662;
wire n_34663;
wire n_34664;
wire n_34666;
wire n_34667;
wire n_34668;
wire n_34669;
wire n_3467;
wire n_34670;
wire n_34671;
wire n_34674;
wire n_34675;
wire n_34676;
wire n_34677;
wire n_34678;
wire n_3468;
wire n_34682;
wire n_34683;
wire n_34684;
wire n_34685;
wire n_34686;
wire n_34687;
wire TIMEBOOST_net_322;
wire n_34692;
wire n_34693;
wire n_34694;
wire n_34695;
wire n_34696;
wire n_34697;
wire n_34698;
wire n_34699;
wire n_347;
wire n_3470;
wire n_34700;
wire n_34701;
wire n_34702;
wire n_34703;
wire n_34704;
wire n_34705;
wire n_34706;
wire n_34707;
wire n_34709;
wire n_3471;
wire n_34710;
wire n_34711;
wire n_34712;
wire n_34713;
wire n_34714;
wire n_34715;
wire n_34716;
wire n_34717;
wire n_34718;
wire n_3472;
wire n_34721;
wire n_34724;
wire n_34725;
wire n_34726;
wire n_34727;
wire n_34728;
wire n_34729;
wire n_3473;
wire n_34730;
wire n_34733;
wire n_34734;
wire n_34735;
wire n_34738;
wire n_34739;
wire n_3474;
wire n_34740;
wire n_34741;
wire n_34742;
wire n_34743;
wire n_34744;
wire n_34745;
wire n_34746;
wire n_34747;
wire n_34748;
wire n_34749;
wire n_3475;
wire n_34751;
wire n_34752;
wire n_34753;
wire n_34754;
wire TIMEBOOST_net_2610;
wire n_34756;
wire n_34757;
wire n_34758;
wire n_34759;
wire n_34760;
wire n_34762;
wire n_34763;
wire n_34764;
wire n_34765;
wire n_34766;
wire n_34767;
wire n_34768;
wire n_34769;
wire n_3477;
wire TIMEBOOST_net_330;
wire n_34772;
wire n_34774;
wire n_34775;
wire n_34776;
wire n_34777;
wire n_34778;
wire n_34779;
wire n_3478;
wire n_34782;
wire n_34783;
wire n_34784;
wire n_34785;
wire n_34786;
wire n_34788;
wire n_34789;
wire n_3479;
wire n_34790;
wire n_34791;
wire TIMEBOOST_net_334;
wire n_34793;
wire TIMEBOOST_net_327;
wire n_34795;
wire TIMEBOOST_net_1102;
wire n_34797;
wire n_348;
wire TIMEBOOST_net_317;
wire n_34800;
wire n_34801;
wire n_34802;
wire n_34803;
wire n_34804;
wire n_34805;
wire n_34806;
wire n_34807;
wire n_34808;
wire n_34809;
wire n_3481;
wire n_34810;
wire n_34811;
wire n_34812;
wire n_34813;
wire n_34814;
wire n_34815;
wire n_34816;
wire n_34817;
wire n_34818;
wire n_34819;
wire n_3482;
wire n_34820;
wire n_34821;
wire n_34822;
wire n_34823;
wire n_34824;
wire n_34825;
wire TIMEBOOST_net_362;
wire n_34827;
wire n_34828;
wire n_34829;
wire n_3483;
wire n_34830;
wire TIMEBOOST_net_1206;
wire TIMEBOOST_net_1071;
wire n_34835;
wire n_34836;
wire n_34839;
wire n_3484;
wire n_34840;
wire n_34841;
wire n_34842;
wire n_34843;
wire n_34844;
wire n_34845;
wire n_34846;
wire n_34847;
wire n_34848;
wire n_34849;
wire n_3485;
wire n_34850;
wire n_34851;
wire n_34852;
wire TIMEBOOST_net_2430;
wire n_34854;
wire n_34855;
wire n_34856;
wire n_34858;
wire TIMEBOOST_net_363;
wire TIMEBOOST_net_1174;
wire n_34861;
wire n_34864;
wire n_34865;
wire n_34866;
wire n_34867;
wire n_34868;
wire n_34869;
wire n_34870;
wire n_34872;
wire n_34873;
wire n_34874;
wire n_34875;
wire n_34876;
wire n_34877;
wire n_34878;
wire n_3488;
wire n_34880;
wire n_34881;
wire n_34883;
wire n_34885;
wire n_34886;
wire n_34888;
wire n_34889;
wire n_3489;
wire n_34890;
wire n_34891;
wire n_34892;
wire n_34893;
wire n_34894;
wire n_34895;
wire n_34896;
wire n_34897;
wire n_34898;
wire n_34899;
wire n_349;
wire n_3490;
wire n_34900;
wire n_34901;
wire n_34903;
wire n_34905;
wire n_34906;
wire n_34907;
wire n_34908;
wire n_3491;
wire n_34911;
wire n_34912;
wire n_34913;
wire n_34914;
wire n_34915;
wire n_34916;
wire n_34917;
wire n_34918;
wire n_34919;
wire n_3492;
wire n_34921;
wire n_34923;
wire n_34924;
wire n_34925;
wire n_34926;
wire n_34927;
wire TIMEBOOST_net_1979;
wire n_34929;
wire n_3493;
wire n_34930;
wire n_34931;
wire n_34933;
wire n_34934;
wire n_34935;
wire n_34936;
wire n_34938;
wire n_3494;
wire n_34940;
wire n_34941;
wire n_34942;
wire n_34943;
wire n_34944;
wire n_34946;
wire n_34947;
wire n_3495;
wire n_34952;
wire n_34953;
wire n_34954;
wire n_34955;
wire n_34956;
wire n_34957;
wire n_34959;
wire n_3496;
wire n_34960;
wire n_34961;
wire n_34962;
wire n_34963;
wire n_34964;
wire n_34965;
wire n_34966;
wire n_34967;
wire n_34971;
wire n_34972;
wire n_34974;
wire TIMEBOOST_net_1176;
wire TIMEBOOST_net_365;
wire n_34978;
wire n_3498;
wire n_34980;
wire n_34981;
wire n_34982;
wire n_34983;
wire n_34985;
wire n_34988;
wire n_34989;
wire n_3499;
wire n_34990;
wire n_34991;
wire TIMEBOOST_net_1178;
wire n_34993;
wire TIMEBOOST_net_1607;
wire n_34996;
wire n_34999;
wire n_350;
wire n_3500;
wire n_35000;
wire n_35001;
wire n_35003;
wire n_35005;
wire n_35006;
wire n_35008;
wire n_35009;
wire n_3501;
wire TIMEBOOST_net_1045;
wire n_35012;
wire TIMEBOOST_net_338;
wire n_35016;
wire n_35017;
wire n_35018;
wire n_35019;
wire n_3502;
wire n_35020;
wire n_35021;
wire n_35025;
wire n_35026;
wire n_35029;
wire n_3503;
wire n_35030;
wire TIMEBOOST_net_1175;
wire TIMEBOOST_net_2718;
wire n_35034;
wire TIMEBOOST_net_405;
wire n_35037;
wire n_3504;
wire n_35041;
wire n_35042;
wire n_35043;
wire n_35044;
wire n_35045;
wire n_35046;
wire n_35047;
wire n_35048;
wire n_35049;
wire n_3505;
wire n_35053;
wire n_35055;
wire TIMEBOOST_net_1660;
wire n_35057;
wire n_35058;
wire n_35059;
wire n_3506;
wire n_35060;
wire TIMEBOOST_net_1695;
wire n_35063;
wire n_35065;
wire n_35069;
wire n_3507;
wire n_35070;
wire n_35071;
wire n_35072;
wire n_35073;
wire n_35075;
wire n_35077;
wire n_35078;
wire n_3508;
wire TIMEBOOST_net_2830;
wire n_35083;
wire n_35084;
wire n_35086;
wire n_35087;
wire n_35088;
wire n_35089;
wire n_3509;
wire n_35090;
wire n_35092;
wire n_35093;
wire TIMEBOOST_net_368;
wire n_35095;
wire n_35096;
wire n_35097;
wire n_35098;
wire n_35099;
wire n_3510;
wire n_35100;
wire n_35101;
wire n_35102;
wire TIMEBOOST_net_344;
wire n_35106;
wire n_35107;
wire n_35108;
wire n_35109;
wire n_3511;
wire n_35110;
wire n_35111;
wire n_35112;
wire n_35113;
wire TIMEBOOST_net_1671;
wire TIMEBOOST_net_370;
wire n_35118;
wire n_35119;
wire TIMEBOOST_net_1990;
wire n_35121;
wire n_35122;
wire n_35123;
wire n_35125;
wire n_35126;
wire n_35127;
wire n_35128;
wire n_35130;
wire n_35132;
wire n_35133;
wire n_35134;
wire n_35135;
wire n_35136;
wire n_35137;
wire TIMEBOOST_net_1182;
wire n_35139;
wire TIMEBOOST_net_429;
wire n_35140;
wire n_35141;
wire n_35143;
wire n_35145;
wire n_35146;
wire n_35147;
wire n_35148;
wire n_35150;
wire n_35152;
wire n_35154;
wire n_35155;
wire n_35156;
wire n_35157;
wire n_35159;
wire n_35160;
wire n_35161;
wire n_35162;
wire n_35163;
wire n_35164;
wire n_35167;
wire n_35168;
wire n_35169;
wire TIMEBOOST_net_371;
wire n_35171;
wire n_35172;
wire TIMEBOOST_net_1027;
wire n_35174;
wire n_35175;
wire n_35177;
wire n_35178;
wire n_35179;
wire n_3518;
wire n_35180;
wire n_35183;
wire n_35184;
wire TIMEBOOST_net_2777;
wire n_35187;
wire n_35188;
wire n_35189;
wire n_3519;
wire n_35190;
wire n_35191;
wire n_35192;
wire n_35193;
wire n_35194;
wire n_35195;
wire n_35196;
wire n_35197;
wire n_35198;
wire n_35199;
wire n_35200;
wire n_35201;
wire n_35204;
wire n_35205;
wire n_35207;
wire n_3521;
wire n_35210;
wire n_35211;
wire TIMEBOOST_net_2770;
wire n_35213;
wire n_35214;
wire n_35215;
wire n_35216;
wire n_35217;
wire n_35218;
wire n_35219;
wire n_3522;
wire n_35220;
wire n_35221;
wire n_35223;
wire n_35224;
wire n_35225;
wire n_35226;
wire n_35228;
wire n_35229;
wire n_35230;
wire n_35231;
wire n_35234;
wire n_35235;
wire n_35236;
wire n_35237;
wire n_35239;
wire n_35240;
wire n_35241;
wire n_35242;
wire n_35243;
wire n_35244;
wire n_35245;
wire n_35246;
wire n_35247;
wire n_35249;
wire n_3525;
wire n_35250;
wire n_35251;
wire n_35252;
wire n_35253;
wire TIMEBOOST_net_432;
wire n_35256;
wire n_35257;
wire n_35258;
wire n_35259;
wire n_3526;
wire n_35260;
wire n_35262;
wire n_35264;
wire n_35265;
wire n_35266;
wire n_35267;
wire n_35268;
wire n_35269;
wire n_3527;
wire n_35270;
wire n_35271;
wire n_35272;
wire n_35273;
wire n_35274;
wire n_35275;
wire n_35277;
wire n_35278;
wire n_35279;
wire n_3528;
wire n_35280;
wire n_35281;
wire n_35282;
wire n_35283;
wire n_35284;
wire n_35285;
wire n_35287;
wire n_35288;
wire n_35289;
wire n_3529;
wire n_35290;
wire n_35292;
wire n_35293;
wire n_35294;
wire n_35296;
wire n_35298;
wire n_35299;
wire n_353;
wire n_3530;
wire n_35303;
wire n_35305;
wire n_35307;
wire n_35309;
wire n_35310;
wire n_35311;
wire n_35312;
wire n_35313;
wire n_35314;
wire n_35315;
wire n_35316;
wire n_35317;
wire n_35318;
wire n_3532;
wire n_35320;
wire n_35321;
wire n_35322;
wire n_35323;
wire n_35324;
wire n_35325;
wire n_35326;
wire n_35327;
wire n_35328;
wire n_35329;
wire n_3533;
wire n_35330;
wire n_35331;
wire n_35332;
wire n_35333;
wire n_35334;
wire n_35335;
wire n_35336;
wire n_35337;
wire n_35338;
wire n_35339;
wire TIMEBOOST_net_1004;
wire n_35340;
wire n_35341;
wire n_35342;
wire n_35343;
wire n_35344;
wire n_35345;
wire n_35346;
wire n_35347;
wire n_35349;
wire n_3535;
wire n_35350;
wire n_35351;
wire n_35352;
wire n_35353;
wire n_35354;
wire n_35355;
wire n_35356;
wire n_35357;
wire n_35358;
wire n_35359;
wire n_3536;
wire n_35360;
wire n_35361;
wire n_35362;
wire n_35363;
wire n_35364;
wire n_35365;
wire TIMEBOOST_net_468;
wire n_35367;
wire n_35368;
wire TIMEBOOST_net_2811;
wire TIMEBOOST_net_467;
wire n_35371;
wire n_35372;
wire n_35373;
wire n_35374;
wire n_35375;
wire n_35376;
wire n_35377;
wire n_35378;
wire n_35379;
wire n_3538;
wire n_35380;
wire n_35381;
wire n_35382;
wire n_35383;
wire TIMEBOOST_net_470;
wire n_35385;
wire n_35386;
wire n_35387;
wire n_35388;
wire n_35389;
wire n_3539;
wire n_35390;
wire n_35391;
wire n_35392;
wire n_35393;
wire n_35394;
wire n_35396;
wire n_35397;
wire n_35398;
wire n_35399;
wire n_354;
wire n_35401;
wire n_35402;
wire n_35403;
wire n_35404;
wire n_35405;
wire n_35406;
wire n_35407;
wire n_35408;
wire n_35409;
wire n_35410;
wire TIMEBOOST_net_1318;
wire n_35413;
wire n_35414;
wire n_35415;
wire n_35416;
wire n_35417;
wire n_35418;
wire n_35419;
wire n_3542;
wire n_35420;
wire n_35421;
wire n_35423;
wire n_35424;
wire n_35425;
wire n_35426;
wire n_35427;
wire n_35428;
wire n_35429;
wire n_3543;
wire n_35430;
wire n_35431;
wire n_35432;
wire n_35433;
wire n_35434;
wire n_35435;
wire n_35436;
wire n_35437;
wire n_35438;
wire n_35439;
wire n_35440;
wire n_35441;
wire TIMEBOOST_net_483;
wire n_35443;
wire n_35444;
wire TIMEBOOST_net_2490;
wire n_35446;
wire n_35447;
wire TIMEBOOST_net_482;
wire n_35449;
wire n_3545;
wire n_35450;
wire n_35451;
wire n_35452;
wire n_35453;
wire n_35454;
wire n_35455;
wire n_35456;
wire n_35457;
wire TIMEBOOST_net_1734;
wire n_35459;
wire n_3546;
wire n_35460;
wire n_35461;
wire n_35462;
wire n_35463;
wire n_35464;
wire n_35465;
wire n_35466;
wire n_35467;
wire n_35468;
wire n_35469;
wire n_3547;
wire n_35470;
wire n_35471;
wire n_35472;
wire n_35473;
wire n_35474;
wire n_35475;
wire n_35476;
wire n_35477;
wire n_35478;
wire n_35479;
wire n_3548;
wire n_35480;
wire n_35481;
wire n_35482;
wire n_35483;
wire n_35484;
wire n_35485;
wire TIMEBOOST_net_2926;
wire n_35487;
wire n_35488;
wire n_35489;
wire n_3549;
wire n_35490;
wire n_35491;
wire n_35493;
wire n_35494;
wire n_35495;
wire n_35496;
wire n_35499;
wire n_355;
wire n_35500;
wire n_35501;
wire n_35502;
wire n_35503;
wire n_35504;
wire n_35505;
wire n_35506;
wire n_35507;
wire n_35508;
wire n_35509;
wire n_3551;
wire n_35510;
wire n_35511;
wire n_35512;
wire n_35513;
wire n_35515;
wire n_35516;
wire n_35517;
wire n_35518;
wire n_35519;
wire n_35520;
wire n_35521;
wire n_35522;
wire n_35523;
wire n_35524;
wire n_35525;
wire n_35526;
wire n_35529;
wire n_35531;
wire n_35532;
wire n_35533;
wire n_35535;
wire n_35536;
wire n_35537;
wire n_35538;
wire n_35539;
wire n_35540;
wire n_35541;
wire n_35542;
wire n_35543;
wire n_35545;
wire n_35546;
wire n_35547;
wire n_35550;
wire n_35551;
wire n_35552;
wire n_35553;
wire n_35554;
wire n_35555;
wire n_35556;
wire n_35557;
wire n_35559;
wire n_3556;
wire TIMEBOOST_net_2957;
wire n_35561;
wire n_35562;
wire n_35565;
wire n_35566;
wire n_35567;
wire n_35569;
wire n_3557;
wire n_35570;
wire TIMEBOOST_net_475;
wire n_35573;
wire n_35574;
wire n_35575;
wire n_35576;
wire n_35577;
wire n_35578;
wire n_35579;
wire n_3558;
wire n_35581;
wire n_35582;
wire n_35583;
wire n_35584;
wire n_35587;
wire n_35588;
wire n_3559;
wire n_35590;
wire n_35591;
wire n_35592;
wire n_35593;
wire n_35594;
wire n_35595;
wire n_35596;
wire n_35597;
wire n_35598;
wire n_35599;
wire n_3560;
wire n_35602;
wire n_35604;
wire n_35605;
wire n_35606;
wire n_3561;
wire n_35611;
wire n_35612;
wire n_35613;
wire TIMEBOOST_net_1349;
wire n_35615;
wire n_35616;
wire n_35617;
wire n_35619;
wire n_3562;
wire n_35620;
wire n_35621;
wire n_35622;
wire n_35623;
wire n_35624;
wire n_35625;
wire n_35626;
wire n_35627;
wire n_35629;
wire n_3563;
wire n_35630;
wire n_35631;
wire n_35633;
wire n_35634;
wire n_35635;
wire n_35638;
wire n_35639;
wire n_3564;
wire n_35640;
wire n_35641;
wire n_35643;
wire n_35644;
wire n_35645;
wire n_35646;
wire n_35647;
wire n_35648;
wire n_35649;
wire n_3565;
wire n_35650;
wire n_35651;
wire n_35653;
wire n_35654;
wire n_35655;
wire n_35656;
wire n_35657;
wire n_35659;
wire n_3566;
wire n_35663;
wire n_35665;
wire n_35667;
wire n_35669;
wire TIMEBOOST_net_346;
wire n_35670;
wire n_35671;
wire n_35672;
wire n_35673;
wire n_35674;
wire n_35675;
wire n_35678;
wire n_35679;
wire n_3568;
wire n_35680;
wire n_35681;
wire n_35682;
wire n_35683;
wire n_35684;
wire n_35687;
wire TIMEBOOST_net_2086;
wire n_35689;
wire n_3569;
wire n_35690;
wire n_35691;
wire n_35692;
wire n_35693;
wire n_35694;
wire n_35696;
wire n_35697;
wire n_35698;
wire n_35699;
wire n_357;
wire n_3570;
wire n_35700;
wire n_35703;
wire n_35704;
wire n_35705;
wire n_35706;
wire n_35707;
wire n_35708;
wire n_35709;
wire n_3571;
wire n_35710;
wire n_35711;
wire n_35712;
wire n_35713;
wire TIMEBOOST_net_568;
wire n_35715;
wire n_35716;
wire n_35717;
wire n_35718;
wire n_35719;
wire n_3572;
wire n_35720;
wire n_35722;
wire n_35723;
wire n_35724;
wire n_35725;
wire n_35726;
wire n_35729;
wire n_3573;
wire n_35732;
wire n_35736;
wire n_35737;
wire n_35738;
wire n_35739;
wire n_35740;
wire n_35742;
wire n_35744;
wire n_35746;
wire n_35747;
wire n_35748;
wire n_35749;
wire n_3575;
wire n_35750;
wire n_35751;
wire n_35752;
wire n_35754;
wire n_35755;
wire n_35757;
wire n_3576;
wire n_35763;
wire n_35764;
wire n_35765;
wire TIMEBOOST_net_1148;
wire n_35767;
wire n_35768;
wire n_35769;
wire n_3577;
wire n_35770;
wire n_35774;
wire n_35776;
wire n_35778;
wire n_35779;
wire n_3578;
wire n_35780;
wire n_35782;
wire n_35783;
wire n_35784;
wire n_35785;
wire TIMEBOOST_net_2850;
wire n_35787;
wire n_35788;
wire n_3579;
wire n_35791;
wire n_35792;
wire n_35793;
wire n_35794;
wire n_35795;
wire n_35796;
wire n_35797;
wire n_35799;
wire n_358;
wire n_3580;
wire n_35800;
wire TIMEBOOST_net_2377;
wire n_35804;
wire n_35805;
wire n_35806;
wire n_35807;
wire n_35808;
wire n_35809;
wire n_3581;
wire n_35810;
wire n_35814;
wire n_35815;
wire n_35819;
wire n_3582;
wire n_35820;
wire n_35821;
wire n_35822;
wire n_35824;
wire n_35826;
wire n_35827;
wire n_35828;
wire n_35829;
wire n_3583;
wire n_35830;
wire n_35831;
wire n_35832;
wire n_35833;
wire n_35834;
wire n_35835;
wire n_35836;
wire n_35839;
wire n_3584;
wire n_35840;
wire n_35841;
wire n_35842;
wire TIMEBOOST_net_1145;
wire n_35845;
wire n_35847;
wire n_35848;
wire n_35849;
wire n_35850;
wire n_35851;
wire TIMEBOOST_net_1147;
wire n_35853;
wire n_35854;
wire n_35856;
wire n_35857;
wire n_35859;
wire n_3586;
wire n_35860;
wire n_35861;
wire n_35864;
wire n_35865;
wire n_35866;
wire n_35867;
wire n_35868;
wire n_35869;
wire n_35870;
wire n_35872;
wire n_35873;
wire n_35874;
wire n_35876;
wire n_35877;
wire n_35878;
wire TIMEBOOST_net_578;
wire n_35880;
wire n_35882;
wire n_35883;
wire n_35884;
wire n_35886;
wire n_35887;
wire n_35888;
wire n_35889;
wire n_35890;
wire n_35891;
wire TIMEBOOST_net_1149;
wire n_35897;
wire TIMEBOOST_net_1351;
wire n_35899;
wire n_3590;
wire n_35900;
wire n_35901;
wire n_35905;
wire n_35906;
wire n_35909;
wire n_3591;
wire n_35910;
wire n_35911;
wire n_35914;
wire n_35916;
wire n_35917;
wire n_35918;
wire n_35919;
wire n_3592;
wire n_35920;
wire n_35921;
wire n_35922;
wire n_35923;
wire n_35926;
wire n_35927;
wire n_35928;
wire n_35929;
wire n_3593;
wire n_35930;
wire n_35931;
wire n_35932;
wire TIMEBOOST_net_2460;
wire n_35934;
wire n_35935;
wire n_35936;
wire n_35937;
wire n_35938;
wire n_35939;
wire n_3594;
wire n_35940;
wire n_35941;
wire n_35945;
wire n_35947;
wire n_35948;
wire n_3595;
wire TIMEBOOST_net_1227;
wire n_35951;
wire n_35952;
wire n_35953;
wire n_35954;
wire n_35955;
wire n_35956;
wire n_35958;
wire n_35959;
wire n_3596;
wire n_35960;
wire n_35961;
wire n_35962;
wire n_35963;
wire n_35964;
wire n_35965;
wire n_35966;
wire n_35967;
wire n_35968;
wire n_35969;
wire n_3597;
wire n_35970;
wire n_35971;
wire n_35972;
wire n_35974;
wire n_35976;
wire n_35977;
wire n_3598;
wire n_35980;
wire TIMEBOOST_net_1341;
wire n_35984;
wire n_35985;
wire n_35987;
wire n_35988;
wire n_35989;
wire TIMEBOOST_net_2893;
wire n_35990;
wire n_35992;
wire n_35993;
wire n_35994;
wire TIMEBOOST_net_357;
wire n_35996;
wire n_360;
wire n_3600;
wire n_36000;
wire n_36001;
wire n_36004;
wire n_36005;
wire n_36007;
wire n_36008;
wire n_36009;
wire n_3601;
wire n_36010;
wire n_36011;
wire n_36012;
wire n_36013;
wire n_36014;
wire n_36015;
wire n_36018;
wire n_36019;
wire n_3602;
wire n_36021;
wire n_36022;
wire n_36023;
wire n_36024;
wire n_36025;
wire n_36026;
wire n_36030;
wire n_36032;
wire n_36033;
wire n_36034;
wire n_36035;
wire n_36036;
wire n_36037;
wire n_36038;
wire n_36039;
wire n_3604;
wire n_36040;
wire n_36043;
wire n_36045;
wire n_36046;
wire n_36047;
wire n_36049;
wire n_3605;
wire n_36050;
wire n_36052;
wire n_36053;
wire n_36054;
wire n_36055;
wire n_36056;
wire n_36058;
wire n_36059;
wire n_3606;
wire n_36062;
wire n_36063;
wire TIMEBOOST_net_476;
wire n_36065;
wire n_36066;
wire TIMEBOOST_net_1340;
wire n_36069;
wire n_3607;
wire n_36071;
wire n_36072;
wire n_36073;
wire n_36074;
wire n_36075;
wire TIMEBOOST_net_1440;
wire n_36079;
wire n_3608;
wire n_36080;
wire n_36081;
wire n_36082;
wire n_36083;
wire n_36084;
wire n_36086;
wire n_36088;
wire TIMEBOOST_net_2951;
wire n_3609;
wire n_36090;
wire n_36091;
wire n_36093;
wire n_36094;
wire n_36095;
wire n_36096;
wire n_36097;
wire n_36098;
wire n_36099;
wire n_361;
wire n_3610;
wire n_36100;
wire n_36102;
wire n_36103;
wire n_36105;
wire n_36108;
wire n_36109;
wire n_36110;
wire n_36111;
wire n_36112;
wire n_36113;
wire n_36114;
wire n_36117;
wire n_36118;
wire n_36119;
wire n_3612;
wire n_36120;
wire n_36121;
wire n_36122;
wire n_36123;
wire n_36124;
wire n_36125;
wire n_36126;
wire n_36127;
wire n_3613;
wire n_36130;
wire n_36132;
wire n_36133;
wire n_36134;
wire n_36135;
wire n_36136;
wire n_36138;
wire n_36139;
wire n_36140;
wire TIMEBOOST_net_2069;
wire n_36143;
wire TIMEBOOST_net_1338;
wire TIMEBOOST_net_602;
wire n_36147;
wire n_36148;
wire n_3615;
wire n_36151;
wire TIMEBOOST_net_779;
wire n_36154;
wire n_36155;
wire n_36156;
wire n_36157;
wire n_36158;
wire n_36159;
wire n_3616;
wire n_36160;
wire n_36161;
wire n_36162;
wire n_36164;
wire n_36165;
wire n_36167;
wire n_36168;
wire n_36169;
wire n_36170;
wire n_36171;
wire n_36172;
wire n_36173;
wire n_36174;
wire n_36175;
wire n_36176;
wire n_36177;
wire n_36178;
wire n_36179;
wire n_36180;
wire n_36182;
wire n_36183;
wire n_36184;
wire n_36185;
wire n_36186;
wire n_36187;
wire n_36188;
wire n_36190;
wire n_36191;
wire n_36192;
wire n_36193;
wire n_36194;
wire n_36195;
wire n_36196;
wire n_36197;
wire n_36198;
wire n_36199;
wire n_362;
wire n_3620;
wire n_36200;
wire n_36203;
wire n_36204;
wire n_36205;
wire n_36206;
wire n_36207;
wire n_36208;
wire n_36209;
wire n_36210;
wire n_36211;
wire n_36212;
wire n_36213;
wire n_36214;
wire n_36215;
wire n_36216;
wire n_36217;
wire n_36218;
wire n_36219;
wire n_36220;
wire n_36221;
wire n_36222;
wire n_36223;
wire n_36224;
wire n_36225;
wire n_36226;
wire n_36227;
wire n_36228;
wire n_36229;
wire n_3623;
wire n_36230;
wire n_36231;
wire n_36232;
wire n_36233;
wire n_36234;
wire n_36235;
wire n_36236;
wire n_36237;
wire n_36238;
wire n_36239;
wire n_3624;
wire n_36240;
wire n_36241;
wire n_36242;
wire n_36243;
wire n_36245;
wire n_36246;
wire n_36247;
wire n_36248;
wire n_3625;
wire n_36250;
wire n_36251;
wire n_36252;
wire n_36253;
wire n_36254;
wire n_36255;
wire n_36256;
wire n_36257;
wire n_36258;
wire n_36259;
wire n_3626;
wire n_36260;
wire n_36261;
wire n_36262;
wire n_36263;
wire n_36264;
wire n_36265;
wire n_36267;
wire n_36268;
wire n_36269;
wire n_3627;
wire n_36270;
wire n_36271;
wire n_36272;
wire n_36273;
wire n_36274;
wire n_36275;
wire n_36276;
wire n_36277;
wire n_36279;
wire n_36280;
wire n_36281;
wire n_36282;
wire n_36283;
wire n_36284;
wire n_36285;
wire n_36286;
wire n_36287;
wire n_36288;
wire n_36289;
wire n_3629;
wire n_36290;
wire n_36291;
wire n_36292;
wire n_36293;
wire n_36294;
wire n_36295;
wire n_36297;
wire n_36298;
wire n_36299;
wire n_363;
wire n_3630;
wire n_36300;
wire n_36301;
wire n_36302;
wire n_36303;
wire n_36304;
wire n_36305;
wire n_36306;
wire n_36307;
wire TIMEBOOST_net_1363;
wire n_36309;
wire n_3631;
wire n_36310;
wire n_36313;
wire n_36314;
wire n_36315;
wire n_36316;
wire n_36317;
wire n_36318;
wire n_36319;
wire n_3632;
wire n_36320;
wire n_36321;
wire n_36322;
wire n_36323;
wire n_36324;
wire n_36325;
wire n_36326;
wire n_36327;
wire n_36328;
wire n_36329;
wire n_3633;
wire n_36330;
wire n_36331;
wire n_36332;
wire n_36333;
wire n_36334;
wire n_36335;
wire n_36336;
wire n_36337;
wire n_36338;
wire n_36339;
wire TIMEBOOST_net_2269;
wire n_36340;
wire n_36343;
wire n_36344;
wire n_36345;
wire n_36346;
wire n_36347;
wire n_36348;
wire n_36349;
wire n_3635;
wire n_36350;
wire TIMEBOOST_net_1404;
wire n_36352;
wire n_36353;
wire n_36354;
wire n_36355;
wire n_36356;
wire n_36358;
wire n_36359;
wire n_3636;
wire n_36360;
wire n_36361;
wire n_36362;
wire n_36363;
wire n_36364;
wire n_36365;
wire n_36366;
wire n_36367;
wire n_36368;
wire n_36369;
wire n_36370;
wire n_36371;
wire n_36372;
wire n_36373;
wire n_36374;
wire TIMEBOOST_net_1374;
wire n_36376;
wire n_36377;
wire n_36378;
wire n_36379;
wire n_3638;
wire n_36381;
wire n_36382;
wire n_36383;
wire n_36384;
wire n_36385;
wire n_36386;
wire n_36387;
wire n_36388;
wire n_36389;
wire n_3639;
wire n_36390;
wire n_36391;
wire n_36392;
wire n_36393;
wire n_36394;
wire n_36395;
wire n_36396;
wire n_36397;
wire n_36398;
wire n_36399;
wire n_3640;
wire n_36400;
wire n_36402;
wire n_36403;
wire n_36404;
wire n_36405;
wire n_36406;
wire n_36407;
wire n_36408;
wire n_36409;
wire n_3641;
wire n_36410;
wire n_36411;
wire n_36412;
wire n_36413;
wire n_36414;
wire n_36415;
wire n_36416;
wire n_36418;
wire n_36419;
wire n_3642;
wire n_36420;
wire n_36421;
wire n_36422;
wire n_36423;
wire n_36424;
wire n_36425;
wire n_36427;
wire n_36428;
wire n_36429;
wire n_3643;
wire n_36430;
wire n_36431;
wire n_36432;
wire n_36433;
wire n_36434;
wire n_36435;
wire n_36437;
wire n_36438;
wire n_36439;
wire n_36440;
wire n_36441;
wire n_36442;
wire n_36444;
wire n_36445;
wire TIMEBOOST_net_1575;
wire n_36447;
wire n_36449;
wire n_3645;
wire n_36450;
wire n_36451;
wire n_36452;
wire n_36453;
wire n_36454;
wire n_36455;
wire n_36457;
wire n_36458;
wire n_3646;
wire n_36460;
wire n_36461;
wire n_36462;
wire n_36463;
wire n_36464;
wire n_36465;
wire n_36466;
wire n_36467;
wire n_36468;
wire n_36469;
wire n_36470;
wire TIMEBOOST_net_2687;
wire TIMEBOOST_net_598;
wire n_36474;
wire TIMEBOOST_net_772;
wire n_36476;
wire n_36477;
wire n_36478;
wire n_36479;
wire n_3648;
wire n_36480;
wire n_36481;
wire n_36482;
wire n_36483;
wire TIMEBOOST_net_692;
wire n_36486;
wire n_36487;
wire TIMEBOOST_net_1795;
wire n_36489;
wire n_3649;
wire n_36490;
wire n_36492;
wire n_36493;
wire n_36494;
wire n_36495;
wire n_36496;
wire n_36497;
wire n_36498;
wire n_36499;
wire n_365;
wire n_3650;
wire n_36501;
wire TIMEBOOST_net_1409;
wire n_36503;
wire n_36504;
wire n_36505;
wire n_36506;
wire n_36507;
wire n_36508;
wire n_3651;
wire n_36510;
wire n_36513;
wire n_36514;
wire n_36515;
wire n_36516;
wire n_36517;
wire TIMEBOOST_net_601;
wire n_3652;
wire n_36520;
wire n_36521;
wire n_36527;
wire n_36528;
wire n_36529;
wire n_3653;
wire n_36530;
wire n_36531;
wire n_36533;
wire n_36534;
wire n_36535;
wire n_36537;
wire TIMEBOOST_net_1407;
wire TIMEBOOST_net_719;
wire n_3654;
wire n_36540;
wire n_36541;
wire n_36542;
wire n_36543;
wire n_36544;
wire n_36545;
wire n_36546;
wire n_36547;
wire n_36549;
wire n_3655;
wire n_36550;
wire n_36551;
wire n_36552;
wire n_36553;
wire TIMEBOOST_net_2099;
wire n_36555;
wire n_36556;
wire n_36557;
wire n_36558;
wire n_36559;
wire n_3656;
wire n_36560;
wire TIMEBOOST_net_1412;
wire TIMEBOOST_net_712;
wire n_36563;
wire n_36564;
wire n_36565;
wire n_36566;
wire n_36567;
wire n_36568;
wire n_36569;
wire TIMEBOOST_net_1408;
wire n_36571;
wire n_36572;
wire n_36573;
wire n_36574;
wire n_36575;
wire n_36576;
wire n_36577;
wire n_36578;
wire n_36579;
wire TIMEBOOST_net_2783;
wire n_36581;
wire TIMEBOOST_net_1816;
wire n_36583;
wire n_36584;
wire n_36585;
wire n_36586;
wire TIMEBOOST_net_612;
wire n_36588;
wire TIMEBOOST_net_1411;
wire n_3659;
wire n_36590;
wire n_36591;
wire n_36592;
wire n_36593;
wire n_36594;
wire n_36595;
wire n_36596;
wire n_36598;
wire n_36599;
wire n_3660;
wire n_36600;
wire n_36601;
wire n_36603;
wire n_36604;
wire n_36607;
wire n_36608;
wire TIMEBOOST_net_713;
wire n_3661;
wire n_36610;
wire n_36611;
wire n_36612;
wire n_36613;
wire n_36614;
wire n_36615;
wire TIMEBOOST_net_2622;
wire TIMEBOOST_net_723;
wire TIMEBOOST_net_611;
wire n_36619;
wire n_36621;
wire n_36622;
wire n_36623;
wire n_36624;
wire n_36625;
wire n_36626;
wire n_36627;
wire n_36628;
wire n_36629;
wire n_3663;
wire n_36630;
wire n_36631;
wire n_36632;
wire TIMEBOOST_net_2128;
wire TIMEBOOST_net_613;
wire n_36635;
wire n_36636;
wire n_36637;
wire n_36638;
wire n_36639;
wire n_36640;
wire n_36641;
wire n_36642;
wire n_36644;
wire n_36645;
wire n_36646;
wire n_36647;
wire TIMEBOOST_net_1798;
wire TIMEBOOST_net_2678;
wire n_36650;
wire n_36651;
wire n_36652;
wire TIMEBOOST_net_1503;
wire n_36654;
wire n_36655;
wire n_36656;
wire n_36657;
wire n_36658;
wire TIMEBOOST_net_1413;
wire n_3666;
wire n_36660;
wire n_36661;
wire n_36662;
wire n_36663;
wire n_36664;
wire n_36666;
wire n_36667;
wire n_36668;
wire n_36669;
wire TIMEBOOST_net_2116;
wire TIMEBOOST_net_1499;
wire n_36672;
wire n_36673;
wire n_36674;
wire n_36675;
wire n_36676;
wire n_36677;
wire n_36678;
wire n_3668;
wire n_36680;
wire n_36681;
wire n_36682;
wire n_36683;
wire n_36684;
wire n_36685;
wire n_36686;
wire TIMEBOOST_net_717;
wire n_36688;
wire n_36689;
wire n_3669;
wire n_36690;
wire n_36691;
wire n_36692;
wire n_36693;
wire n_36695;
wire n_36698;
wire n_36699;
wire n_367;
wire n_3670;
wire n_36700;
wire n_36701;
wire TIMEBOOST_net_1385;
wire n_36703;
wire n_36704;
wire n_36705;
wire n_36706;
wire n_36708;
wire n_36709;
wire n_3671;
wire n_36710;
wire n_36711;
wire n_36712;
wire n_36713;
wire n_36714;
wire n_36715;
wire n_36716;
wire n_36717;
wire n_36718;
wire n_36719;
wire TIMEBOOST_net_2627;
wire n_36720;
wire n_36721;
wire n_36722;
wire n_36723;
wire n_36724;
wire n_36725;
wire n_36726;
wire n_36727;
wire n_36728;
wire n_36729;
wire n_3673;
wire n_36730;
wire n_36731;
wire n_36732;
wire n_36733;
wire n_36734;
wire n_36735;
wire n_36736;
wire n_36737;
wire n_36738;
wire n_36739;
wire n_3674;
wire n_36740;
wire n_36741;
wire n_36742;
wire n_36743;
wire n_36744;
wire n_36745;
wire n_36746;
wire n_36747;
wire n_36748;
wire n_36749;
wire n_36750;
wire n_36751;
wire TIMEBOOST_net_1387;
wire n_36753;
wire n_36754;
wire n_36755;
wire n_36756;
wire n_36757;
wire n_36758;
wire n_36759;
wire n_36760;
wire n_36761;
wire n_36762;
wire n_36763;
wire n_36764;
wire n_36765;
wire n_36766;
wire n_36767;
wire n_36768;
wire n_36769;
wire n_3677;
wire n_36770;
wire n_36771;
wire n_36772;
wire n_36773;
wire n_36774;
wire n_36775;
wire n_36776;
wire n_36777;
wire n_36778;
wire n_3678;
wire n_36780;
wire n_36782;
wire n_36783;
wire n_36784;
wire n_36785;
wire n_36786;
wire n_36787;
wire n_36788;
wire n_36789;
wire n_3679;
wire n_36790;
wire n_36791;
wire n_36792;
wire n_36793;
wire n_36794;
wire n_36796;
wire n_36797;
wire n_36798;
wire n_368;
wire n_36800;
wire n_36801;
wire n_36802;
wire n_36803;
wire n_36805;
wire n_36808;
wire n_3681;
wire n_36810;
wire n_36811;
wire n_36814;
wire n_36816;
wire n_36818;
wire n_36820;
wire n_36822;
wire n_36824;
wire n_36826;
wire n_36828;
wire n_36829;
wire n_3683;
wire n_36830;
wire n_36831;
wire n_36832;
wire n_36833;
wire n_36838;
wire TIMEBOOST_net_278;
wire n_36841;
wire n_36842;
wire n_36844;
wire n_36845;
wire n_36846;
wire n_36847;
wire n_36849;
wire n_3685;
wire n_36851;
wire n_36852;
wire n_36854;
wire n_36855;
wire n_36859;
wire n_3686;
wire n_36860;
wire n_36861;
wire n_36862;
wire n_36863;
wire n_36864;
wire n_36865;
wire n_36866;
wire n_36867;
wire n_36868;
wire n_36869;
wire n_3687;
wire n_36870;
wire n_36871;
wire n_36872;
wire n_36873;
wire n_36874;
wire n_36875;
wire n_36876;
wire n_36877;
wire n_36878;
wire n_36879;
wire n_36880;
wire n_36881;
wire n_36882;
wire n_36883;
wire n_36884;
wire n_36885;
wire n_36886;
wire n_36887;
wire n_36888;
wire n_36889;
wire n_3689;
wire n_36890;
wire n_36891;
wire n_36894;
wire n_36895;
wire n_36896;
wire n_36897;
wire n_36898;
wire n_36899;
wire n_369;
wire n_36900;
wire n_36901;
wire n_36902;
wire n_36903;
wire n_36904;
wire n_36905;
wire n_36906;
wire n_36907;
wire n_36908;
wire n_36909;
wire TIMEBOOST_net_2664;
wire n_36910;
wire n_36911;
wire n_36912;
wire n_36913;
wire n_36914;
wire n_36915;
wire n_36916;
wire n_36917;
wire n_36918;
wire n_36919;
wire n_3692;
wire n_36920;
wire n_36921;
wire n_36922;
wire n_36923;
wire n_36924;
wire n_36925;
wire n_36927;
wire n_36928;
wire n_36929;
wire n_3693;
wire n_36930;
wire n_36931;
wire n_36932;
wire n_36933;
wire n_36934;
wire n_36935;
wire n_36936;
wire n_36937;
wire n_36941;
wire n_36942;
wire n_36943;
wire n_36944;
wire TIMEBOOST_net_2332;
wire n_36946;
wire n_36947;
wire n_36948;
wire TIMEBOOST_net_3;
wire n_3695;
wire n_36950;
wire n_36952;
wire n_36954;
wire n_36955;
wire n_36956;
wire n_36957;
wire n_36958;
wire n_36959;
wire n_3696;
wire n_36960;
wire n_36961;
wire n_36962;
wire n_36963;
wire n_36964;
wire n_36965;
wire n_36966;
wire n_36967;
wire n_36968;
wire n_36969;
wire n_3697;
wire n_36970;
wire n_36971;
wire n_36972;
wire n_36973;
wire n_36974;
wire n_36975;
wire n_36976;
wire n_36978;
wire n_36979;
wire n_3698;
wire n_36980;
wire n_36981;
wire n_36982;
wire n_36983;
wire n_36984;
wire n_36985;
wire n_36986;
wire n_36987;
wire n_36988;
wire n_36989;
wire n_3699;
wire n_36990;
wire n_36991;
wire n_36992;
wire n_36994;
wire n_36996;
wire n_36997;
wire n_36998;
wire n_36999;
wire n_370;
wire n_3700;
wire n_37000;
wire n_37001;
wire n_37002;
wire n_37003;
wire n_37004;
wire n_37005;
wire n_37006;
wire TIMEBOOST_net_1419;
wire n_37008;
wire n_37009;
wire n_3701;
wire n_37010;
wire n_37011;
wire n_37012;
wire n_37013;
wire n_37014;
wire n_37015;
wire n_37016;
wire n_37017;
wire n_37019;
wire n_37020;
wire n_37021;
wire n_37022;
wire n_37023;
wire n_37025;
wire n_37027;
wire n_37028;
wire n_37029;
wire n_37030;
wire n_37031;
wire n_37032;
wire n_37033;
wire n_37034;
wire n_37036;
wire n_37037;
wire n_37038;
wire n_37039;
wire n_3704;
wire n_37040;
wire n_37041;
wire n_37042;
wire n_37043;
wire n_37044;
wire n_37045;
wire n_37046;
wire n_37047;
wire n_37048;
wire n_37049;
wire n_3705;
wire n_37050;
wire n_37051;
wire n_37052;
wire TIMEBOOST_net_788;
wire n_37054;
wire n_37055;
wire n_37056;
wire n_37057;
wire n_37058;
wire n_37059;
wire n_3706;
wire n_37060;
wire n_37061;
wire n_37062;
wire n_37063;
wire n_37064;
wire n_37065;
wire n_37066;
wire n_37067;
wire n_37068;
wire n_37069;
wire n_37070;
wire n_37071;
wire n_37072;
wire n_37073;
wire n_37074;
wire n_37075;
wire n_37076;
wire n_37077;
wire n_37078;
wire n_37079;
wire n_37080;
wire n_37081;
wire n_37083;
wire n_37084;
wire n_37085;
wire n_37086;
wire n_37087;
wire n_37088;
wire n_37089;
wire n_37090;
wire n_37091;
wire n_37092;
wire n_37093;
wire n_37094;
wire n_37095;
wire n_37097;
wire n_37098;
wire n_37099;
wire n_371;
wire n_3710;
wire n_37100;
wire n_37101;
wire n_37102;
wire n_37103;
wire n_37104;
wire n_37105;
wire n_37106;
wire n_37107;
wire n_37108;
wire n_37109;
wire n_37110;
wire n_37111;
wire n_37112;
wire n_37113;
wire n_37115;
wire n_37116;
wire n_37117;
wire n_37118;
wire n_37119;
wire n_37120;
wire n_37121;
wire n_37122;
wire n_37123;
wire n_37124;
wire n_37125;
wire n_37126;
wire n_37127;
wire n_37128;
wire n_37129;
wire n_37130;
wire n_37131;
wire n_37132;
wire n_37133;
wire n_37135;
wire n_37136;
wire n_37138;
wire TIMEBOOST_net_810;
wire n_3714;
wire n_37140;
wire n_37141;
wire n_37142;
wire n_37143;
wire n_37144;
wire n_37145;
wire n_37146;
wire n_37147;
wire n_37148;
wire n_37149;
wire n_3715;
wire n_37150;
wire n_37151;
wire n_37152;
wire n_37153;
wire n_37154;
wire n_37155;
wire n_37156;
wire n_37157;
wire n_37159;
wire n_37160;
wire n_37161;
wire n_37163;
wire n_37164;
wire n_37165;
wire n_37166;
wire n_37167;
wire n_37168;
wire n_37169;
wire n_3717;
wire n_37171;
wire n_37172;
wire n_37173;
wire n_37174;
wire n_37175;
wire n_37176;
wire n_37177;
wire n_37178;
wire n_37179;
wire n_3718;
wire n_37180;
wire n_37181;
wire n_37183;
wire n_37184;
wire n_37185;
wire n_37186;
wire n_37187;
wire n_37188;
wire n_37189;
wire n_37190;
wire n_37191;
wire n_37193;
wire n_37194;
wire n_37195;
wire n_37196;
wire n_37197;
wire n_37198;
wire n_37199;
wire n_372;
wire n_3720;
wire n_37200;
wire n_37201;
wire n_37202;
wire n_37203;
wire n_37204;
wire n_37205;
wire n_37207;
wire n_37209;
wire n_3721;
wire n_37211;
wire n_37212;
wire n_37213;
wire n_37214;
wire n_37215;
wire n_37217;
wire n_37218;
wire n_37219;
wire n_3722;
wire n_37220;
wire n_37221;
wire n_37222;
wire n_37223;
wire n_37224;
wire n_37225;
wire n_37227;
wire n_37228;
wire n_37229;
wire TIMEBOOST_net_282;
wire n_37230;
wire n_37231;
wire n_37232;
wire n_37233;
wire n_37235;
wire n_37236;
wire n_37237;
wire n_37238;
wire n_3724;
wire n_37240;
wire n_37241;
wire n_37242;
wire n_37243;
wire n_37244;
wire n_37245;
wire n_37246;
wire n_37247;
wire n_37248;
wire n_37249;
wire n_3725;
wire n_37250;
wire n_37251;
wire n_37252;
wire n_37253;
wire n_37254;
wire n_37255;
wire n_37256;
wire n_37258;
wire n_37259;
wire n_3726;
wire n_37260;
wire n_37262;
wire n_37264;
wire n_37265;
wire n_37266;
wire n_37268;
wire n_3727;
wire n_37270;
wire n_37271;
wire n_37272;
wire n_37273;
wire n_37274;
wire n_37275;
wire n_37276;
wire n_37277;
wire n_37278;
wire n_37279;
wire n_3728;
wire n_37281;
wire n_37282;
wire n_37283;
wire n_37284;
wire n_37285;
wire n_37286;
wire n_37287;
wire n_37288;
wire n_37289;
wire n_37290;
wire n_37291;
wire n_37292;
wire n_37293;
wire n_37294;
wire n_37295;
wire n_37296;
wire n_37297;
wire n_37298;
wire n_37299;
wire n_373;
wire n_37301;
wire n_37302;
wire n_37303;
wire n_37304;
wire n_37305;
wire n_37306;
wire n_37307;
wire n_37308;
wire n_37309;
wire n_3731;
wire n_37310;
wire n_37311;
wire n_37312;
wire n_37313;
wire n_37314;
wire n_37315;
wire n_37316;
wire n_37317;
wire n_37319;
wire TIMEBOOST_net_390;
wire n_37320;
wire n_37321;
wire n_37322;
wire n_37323;
wire n_37324;
wire n_37325;
wire n_37326;
wire n_37327;
wire n_37328;
wire n_37329;
wire n_3733;
wire n_37330;
wire n_37331;
wire n_37332;
wire n_37333;
wire n_37334;
wire n_37337;
wire n_37339;
wire n_37340;
wire n_37341;
wire n_37342;
wire n_37343;
wire n_37344;
wire n_37345;
wire n_37346;
wire n_37347;
wire n_37348;
wire n_37349;
wire n_3735;
wire n_37350;
wire n_37351;
wire n_37352;
wire n_37353;
wire n_37354;
wire n_37355;
wire n_37356;
wire n_37357;
wire n_37359;
wire n_3736;
wire n_37361;
wire n_37362;
wire n_37363;
wire n_37364;
wire n_37365;
wire n_37366;
wire n_37368;
wire n_37369;
wire n_3737;
wire TIMEBOOST_net_1447;
wire n_37371;
wire n_37372;
wire n_37373;
wire n_37374;
wire n_37375;
wire n_37376;
wire n_37377;
wire n_37379;
wire n_3738;
wire n_37380;
wire n_37381;
wire n_37382;
wire n_37383;
wire n_37384;
wire n_37385;
wire n_37386;
wire n_37387;
wire n_37388;
wire n_37389;
wire TIMEBOOST_net_1117;
wire TIMEBOOST_net_1453;
wire n_37391;
wire n_37392;
wire n_37393;
wire n_37395;
wire n_37396;
wire n_37397;
wire n_37398;
wire n_37399;
wire n_374;
wire TIMEBOOST_net_908;
wire n_37401;
wire n_37402;
wire n_37403;
wire n_37404;
wire n_37405;
wire n_37407;
wire n_37408;
wire n_37409;
wire TIMEBOOST_net_1662;
wire n_37410;
wire n_37411;
wire n_37412;
wire n_37413;
wire n_37414;
wire n_37415;
wire n_37416;
wire n_37417;
wire n_37418;
wire n_37419;
wire n_37421;
wire n_37423;
wire n_37424;
wire n_37425;
wire n_37426;
wire n_37427;
wire n_37428;
wire n_37429;
wire n_3743;
wire n_37430;
wire n_37431;
wire n_37432;
wire n_37433;
wire n_37434;
wire n_37435;
wire n_37436;
wire n_37437;
wire n_37438;
wire n_37439;
wire n_3744;
wire n_37440;
wire n_37441;
wire n_37442;
wire n_37443;
wire n_37444;
wire n_37445;
wire n_37446;
wire n_37447;
wire TIMEBOOST_net_1461;
wire n_37449;
wire n_37451;
wire n_37452;
wire n_37454;
wire n_37455;
wire n_37456;
wire n_37457;
wire n_37458;
wire n_37459;
wire n_3746;
wire n_37460;
wire n_37461;
wire n_37462;
wire TIMEBOOST_net_2743;
wire n_37464;
wire n_37465;
wire n_37466;
wire n_37467;
wire n_37468;
wire n_37469;
wire n_37470;
wire n_37471;
wire n_37472;
wire n_37473;
wire n_37474;
wire n_37475;
wire n_37477;
wire n_37478;
wire n_37479;
wire TIMEBOOST_net_2029;
wire n_37480;
wire n_37481;
wire n_37482;
wire n_37483;
wire n_37484;
wire n_37485;
wire n_37486;
wire n_37487;
wire n_37488;
wire n_37489;
wire n_3749;
wire n_37490;
wire n_37492;
wire n_37493;
wire n_37494;
wire n_37496;
wire n_37497;
wire n_37498;
wire n_37499;
wire n_375;
wire n_3750;
wire n_37500;
wire n_37501;
wire n_37502;
wire n_37504;
wire n_37505;
wire n_37506;
wire n_37507;
wire n_37508;
wire n_37509;
wire n_3751;
wire n_37511;
wire n_37512;
wire n_37513;
wire n_37514;
wire n_37515;
wire n_37516;
wire n_37517;
wire n_37518;
wire n_37519;
wire n_3752;
wire n_37520;
wire n_37521;
wire n_37522;
wire n_37523;
wire n_37524;
wire n_37525;
wire n_37526;
wire n_37527;
wire n_37529;
wire n_3753;
wire n_37531;
wire TIMEBOOST_net_70;
wire n_37534;
wire n_37535;
wire n_37536;
wire TIMEBOOST_net_1861;
wire n_37538;
wire n_37539;
wire n_3754;
wire n_37540;
wire n_37541;
wire n_37542;
wire n_37543;
wire n_37544;
wire n_37545;
wire n_37546;
wire n_37547;
wire n_37548;
wire n_3755;
wire n_37551;
wire n_37554;
wire n_37555;
wire n_37556;
wire n_37557;
wire n_37558;
wire n_37559;
wire n_3756;
wire n_37560;
wire n_37561;
wire TIMEBOOST_net_921;
wire n_37563;
wire TIMEBOOST_net_80;
wire n_37566;
wire n_37568;
wire n_37569;
wire n_3757;
wire n_37571;
wire n_37572;
wire n_37573;
wire n_37574;
wire n_37575;
wire n_37576;
wire n_37577;
wire n_37578;
wire n_37579;
wire n_3758;
wire TIMEBOOST_net_924;
wire n_37581;
wire n_37583;
wire n_37584;
wire n_37585;
wire n_37586;
wire n_37587;
wire n_37589;
wire n_3759;
wire n_37590;
wire n_37593;
wire n_37594;
wire n_37596;
wire n_37597;
wire n_37598;
wire n_376;
wire n_3760;
wire n_37601;
wire n_37602;
wire n_37604;
wire n_37605;
wire n_37606;
wire n_37607;
wire n_37608;
wire n_37609;
wire n_3761;
wire TIMEBOOST_net_2805;
wire n_37611;
wire n_37612;
wire n_37613;
wire n_37614;
wire n_37617;
wire n_37618;
wire n_37619;
wire n_3762;
wire n_37622;
wire n_37623;
wire n_37624;
wire n_37625;
wire n_37626;
wire TIMEBOOST_net_1505;
wire n_37628;
wire TIMEBOOST_net_2825;
wire n_37631;
wire n_37632;
wire n_37634;
wire n_37635;
wire n_37636;
wire n_37637;
wire n_37638;
wire n_37639;
wire n_3764;
wire TIMEBOOST_net_73;
wire n_37644;
wire n_37645;
wire n_37646;
wire n_37647;
wire n_37648;
wire n_37649;
wire n_3765;
wire TIMEBOOST_net_856;
wire n_37653;
wire n_37654;
wire n_37655;
wire n_37656;
wire n_37657;
wire n_37658;
wire n_37659;
wire n_37661;
wire n_37662;
wire n_37663;
wire n_37664;
wire n_37665;
wire TIMEBOOST_net_1509;
wire n_37667;
wire n_37668;
wire n_3767;
wire n_37670;
wire n_37671;
wire n_37672;
wire n_37673;
wire n_37674;
wire n_37676;
wire n_37678;
wire n_3768;
wire n_37680;
wire n_37681;
wire n_37686;
wire n_37687;
wire n_37688;
wire n_37689;
wire n_3769;
wire n_37690;
wire n_37692;
wire n_37693;
wire n_37694;
wire n_37695;
wire n_37696;
wire n_37697;
wire TIMEBOOST_net_2801;
wire n_37699;
wire n_377;
wire n_3770;
wire n_37700;
wire n_37701;
wire n_37702;
wire n_37703;
wire n_37704;
wire n_37707;
wire n_37708;
wire n_37709;
wire n_3771;
wire TIMEBOOST_net_834;
wire n_37711;
wire n_37712;
wire n_37713;
wire n_37715;
wire n_37716;
wire n_37717;
wire TIMEBOOST_net_1800;
wire n_37720;
wire n_37721;
wire n_37722;
wire n_37723;
wire TIMEBOOST_net_1757;
wire n_37725;
wire n_37726;
wire n_37727;
wire n_37728;
wire n_37729;
wire n_3773;
wire n_37730;
wire n_37731;
wire n_37732;
wire n_37733;
wire n_37734;
wire TIMEBOOST_net_1516;
wire n_37737;
wire n_37738;
wire n_37739;
wire n_3774;
wire n_37740;
wire n_37741;
wire n_37742;
wire TIMEBOOST_net_1515;
wire n_37744;
wire n_37745;
wire n_37746;
wire n_37747;
wire n_37748;
wire n_37749;
wire n_3775;
wire n_37750;
wire n_37751;
wire TIMEBOOST_net_2185;
wire n_37753;
wire n_37755;
wire n_37756;
wire n_37757;
wire n_37758;
wire n_37759;
wire n_3776;
wire n_37760;
wire n_37761;
wire n_37762;
wire n_37763;
wire n_37764;
wire n_37765;
wire n_37766;
wire n_37767;
wire n_37768;
wire n_37769;
wire n_3777;
wire n_37770;
wire n_37771;
wire n_37772;
wire n_37773;
wire TIMEBOOST_net_120;
wire n_37775;
wire n_37776;
wire n_37777;
wire n_37778;
wire n_3778;
wire n_37780;
wire n_37781;
wire n_37782;
wire n_37783;
wire n_37784;
wire n_37785;
wire n_37787;
wire n_37788;
wire n_37789;
wire n_37790;
wire n_37791;
wire n_37792;
wire n_37794;
wire n_37795;
wire n_37796;
wire n_37797;
wire n_37798;
wire n_37799;
wire n_378;
wire n_3780;
wire n_37800;
wire n_37801;
wire n_37803;
wire n_37805;
wire n_37806;
wire n_37807;
wire n_37808;
wire n_37809;
wire n_3781;
wire n_37810;
wire n_37811;
wire TIMEBOOST_net_134;
wire n_37813;
wire n_37814;
wire n_37815;
wire n_37816;
wire n_37817;
wire n_37818;
wire n_37819;
wire n_3782;
wire n_37820;
wire n_37821;
wire n_37822;
wire n_37823;
wire TIMEBOOST_net_1522;
wire n_37825;
wire n_37826;
wire n_37827;
wire n_37828;
wire n_37829;
wire n_37830;
wire n_37831;
wire n_37832;
wire n_37833;
wire n_37834;
wire n_37835;
wire n_37836;
wire n_37837;
wire n_37838;
wire n_37839;
wire n_3784;
wire n_37840;
wire n_37841;
wire n_37842;
wire n_37843;
wire n_37844;
wire n_37845;
wire n_37846;
wire n_37847;
wire n_37848;
wire n_37849;
wire TIMEBOOST_net_321;
wire n_37850;
wire TIMEBOOST_net_91;
wire n_37852;
wire n_37853;
wire n_37854;
wire n_37855;
wire n_37856;
wire n_37857;
wire n_37858;
wire n_3786;
wire n_37861;
wire n_37862;
wire n_37863;
wire n_37864;
wire n_37865;
wire n_37866;
wire n_37867;
wire n_37868;
wire n_37869;
wire TIMEBOOST_net_393;
wire n_37871;
wire TIMEBOOST_net_2533;
wire TIMEBOOST_net_93;
wire n_37875;
wire TIMEBOOST_net_92;
wire n_37877;
wire n_37878;
wire TIMEBOOST_net_2157;
wire n_37881;
wire n_37882;
wire n_37883;
wire n_37884;
wire TIMEBOOST_net_2615;
wire n_37887;
wire n_37888;
wire n_37889;
wire TIMEBOOST_net_436;
wire n_37891;
wire n_37892;
wire n_37893;
wire n_37894;
wire n_37895;
wire n_37896;
wire TIMEBOOST_net_1865;
wire n_37898;
wire n_37899;
wire n_379;
wire n_3790;
wire n_37900;
wire n_37901;
wire TIMEBOOST_net_102;
wire TIMEBOOST_net_2890;
wire n_37904;
wire n_37905;
wire n_37906;
wire n_37907;
wire n_37908;
wire n_37909;
wire n_37910;
wire n_37911;
wire n_37912;
wire n_37913;
wire n_37916;
wire n_37917;
wire n_37918;
wire n_37919;
wire n_3792;
wire n_37920;
wire n_37922;
wire n_37923;
wire TIMEBOOST_net_1813;
wire n_37929;
wire TIMEBOOST_net_984;
wire n_37935;
wire TIMEBOOST_net_98;
wire n_37939;
wire n_37940;
wire n_37941;
wire n_37943;
wire n_37944;
wire n_37945;
wire n_37946;
wire n_37947;
wire n_37948;
wire n_37949;
wire n_3795;
wire n_37950;
wire n_37951;
wire n_37952;
wire n_37954;
wire n_37955;
wire n_37956;
wire n_37958;
wire n_37959;
wire n_37960;
wire n_37965;
wire n_37967;
wire n_37968;
wire n_37969;
wire TIMEBOOST_net_1192;
wire n_37970;
wire n_37972;
wire n_37973;
wire n_37974;
wire n_37975;
wire n_37976;
wire TIMEBOOST_net_1021;
wire n_37979;
wire n_37980;
wire n_37981;
wire n_37983;
wire n_37984;
wire n_37985;
wire n_37987;
wire n_37988;
wire n_37989;
wire n_3799;
wire n_37990;
wire n_37991;
wire n_37992;
wire TIMEBOOST_net_1817;
wire TIMEBOOST_net_994;
wire n_38;
wire n_380;
wire n_38000;
wire n_38001;
wire n_38003;
wire n_38004;
wire n_38005;
wire n_38006;
wire n_38007;
wire n_38008;
wire n_38009;
wire n_38010;
wire n_38011;
wire n_38012;
wire TIMEBOOST_net_160;
wire n_38014;
wire n_38016;
wire n_38019;
wire n_3802;
wire n_38020;
wire n_38021;
wire n_38022;
wire n_38026;
wire n_38028;
wire n_3803;
wire n_38032;
wire n_38033;
wire n_38034;
wire n_38035;
wire n_38036;
wire n_38037;
wire n_38038;
wire n_38039;
wire TIMEBOOST_net_2222;
wire n_38041;
wire n_38042;
wire n_38044;
wire n_38045;
wire n_38047;
wire TIMEBOOST_net_1884;
wire n_3805;
wire n_38050;
wire n_38051;
wire n_38053;
wire n_38055;
wire TIMEBOOST_net_159;
wire n_38057;
wire n_38058;
wire TIMEBOOST_net_2552;
wire n_3806;
wire n_38060;
wire n_38062;
wire n_38063;
wire n_38067;
wire n_38068;
wire n_38069;
wire n_3807;
wire n_38070;
wire n_38071;
wire n_38072;
wire n_38073;
wire n_38074;
wire n_38075;
wire n_38076;
wire n_38078;
wire n_38082;
wire n_38083;
wire n_38084;
wire n_38085;
wire n_38087;
wire n_38088;
wire n_38089;
wire n_3809;
wire n_38090;
wire n_38091;
wire n_38092;
wire n_38093;
wire n_38094;
wire n_381;
wire n_3810;
wire n_38102;
wire TIMEBOOST_net_1000;
wire n_38108;
wire n_38109;
wire n_3811;
wire n_38110;
wire n_38111;
wire n_38112;
wire n_38113;
wire n_38114;
wire n_38115;
wire n_38116;
wire n_38117;
wire n_38118;
wire n_38119;
wire n_3812;
wire n_38120;
wire n_38121;
wire n_38122;
wire n_38124;
wire n_38125;
wire n_38126;
wire n_38127;
wire n_38128;
wire n_38129;
wire n_3813;
wire n_38130;
wire n_38131;
wire n_38134;
wire n_38135;
wire TIMEBOOST_net_1011;
wire TIMEBOOST_net_1010;
wire n_38138;
wire n_38139;
wire n_38140;
wire n_38141;
wire n_38142;
wire n_38143;
wire n_38144;
wire n_38145;
wire n_38146;
wire n_38147;
wire n_3815;
wire n_38153;
wire n_38154;
wire n_38156;
wire n_38157;
wire n_38158;
wire n_38159;
wire n_3816;
wire n_38160;
wire n_38161;
wire TIMEBOOST_net_2158;
wire n_38164;
wire n_38166;
wire n_38167;
wire n_38168;
wire n_38169;
wire n_3817;
wire n_38170;
wire n_38171;
wire n_38172;
wire n_38173;
wire n_38174;
wire n_38179;
wire n_38180;
wire n_38181;
wire n_38182;
wire n_38183;
wire n_38184;
wire n_38185;
wire n_38186;
wire n_38187;
wire n_38188;
wire n_3819;
wire n_38190;
wire n_38191;
wire n_38193;
wire n_38196;
wire n_38197;
wire n_38198;
wire n_38199;
wire n_382;
wire n_38200;
wire n_38201;
wire n_38202;
wire n_38204;
wire n_38205;
wire n_38208;
wire n_38209;
wire n_3821;
wire n_38211;
wire n_38212;
wire n_38213;
wire n_38214;
wire n_38215;
wire n_38216;
wire n_38217;
wire n_38218;
wire n_38219;
wire n_3822;
wire n_38220;
wire n_38221;
wire n_38227;
wire n_38228;
wire n_38229;
wire n_38230;
wire n_38231;
wire n_38232;
wire n_38233;
wire n_38234;
wire n_38235;
wire n_38236;
wire n_38237;
wire n_38238;
wire n_38239;
wire n_3824;
wire n_38240;
wire n_38242;
wire n_38243;
wire n_38244;
wire n_38247;
wire n_38248;
wire n_38249;
wire n_3825;
wire n_38250;
wire n_38251;
wire n_38253;
wire n_38254;
wire n_38255;
wire n_38256;
wire n_38258;
wire n_38259;
wire n_38260;
wire n_38261;
wire n_38262;
wire n_38263;
wire n_38266;
wire n_38267;
wire n_38268;
wire n_38269;
wire n_38270;
wire n_38271;
wire n_38272;
wire n_38273;
wire n_38274;
wire n_38276;
wire n_38277;
wire n_38279;
wire n_3828;
wire n_38281;
wire n_38282;
wire n_38283;
wire n_38284;
wire n_38285;
wire n_38286;
wire n_38287;
wire n_38288;
wire n_38290;
wire n_38291;
wire n_38292;
wire n_38293;
wire n_38295;
wire n_38296;
wire n_38297;
wire n_38298;
wire n_383;
wire n_3830;
wire n_38300;
wire n_38301;
wire n_38302;
wire n_38303;
wire n_38304;
wire n_38306;
wire n_38307;
wire n_38308;
wire n_38309;
wire n_38310;
wire n_38311;
wire n_38312;
wire n_38313;
wire n_38314;
wire n_38315;
wire n_38316;
wire n_38317;
wire n_38319;
wire n_3832;
wire n_38320;
wire n_38321;
wire n_38322;
wire n_38323;
wire n_38324;
wire n_38325;
wire n_38326;
wire n_38327;
wire n_38328;
wire n_38329;
wire n_3833;
wire n_38332;
wire n_38333;
wire n_38334;
wire n_38335;
wire n_38336;
wire n_38337;
wire n_38338;
wire n_38339;
wire TIMEBOOST_net_2402;
wire n_38340;
wire TIMEBOOST_net_1101;
wire n_38342;
wire n_38343;
wire n_38344;
wire n_38347;
wire n_38348;
wire n_38349;
wire n_3835;
wire n_38350;
wire n_38352;
wire n_38353;
wire n_38354;
wire n_38355;
wire n_38356;
wire n_38357;
wire n_38358;
wire n_38359;
wire n_38360;
wire n_38361;
wire n_38362;
wire n_38363;
wire n_38364;
wire n_38365;
wire n_38366;
wire n_38367;
wire n_38368;
wire n_38369;
wire n_3837;
wire n_38371;
wire n_38372;
wire n_38373;
wire n_38374;
wire n_38375;
wire n_38376;
wire n_38377;
wire n_38378;
wire n_38379;
wire n_3838;
wire n_38380;
wire n_38381;
wire n_38382;
wire n_38383;
wire n_38384;
wire n_38385;
wire n_38386;
wire n_38387;
wire n_38388;
wire n_38389;
wire TIMEBOOST_net_381;
wire n_38390;
wire n_38391;
wire n_38392;
wire n_38393;
wire n_38394;
wire n_38395;
wire n_38396;
wire n_38397;
wire n_38398;
wire n_38399;
wire n_384;
wire n_3840;
wire n_38400;
wire n_38401;
wire n_38402;
wire n_38403;
wire n_38404;
wire n_38405;
wire n_38406;
wire n_38407;
wire n_38408;
wire n_38409;
wire n_3841;
wire n_38410;
wire n_38411;
wire n_38412;
wire n_38413;
wire n_38414;
wire n_38415;
wire n_38416;
wire n_38417;
wire n_38418;
wire n_38419;
wire n_38420;
wire n_38421;
wire n_38422;
wire n_38423;
wire n_38424;
wire n_38425;
wire n_38426;
wire n_38427;
wire n_38428;
wire n_38429;
wire n_38430;
wire n_38431;
wire n_38432;
wire n_38433;
wire n_38434;
wire n_38435;
wire n_38436;
wire n_38437;
wire n_38438;
wire n_38439;
wire TIMEBOOST_net_2758;
wire n_38440;
wire n_38441;
wire n_38442;
wire n_38443;
wire n_38444;
wire n_38445;
wire n_38446;
wire n_38447;
wire n_38448;
wire n_38449;
wire n_38450;
wire n_38451;
wire n_38452;
wire n_38454;
wire n_38455;
wire n_38456;
wire n_38457;
wire n_38458;
wire n_3846;
wire n_38460;
wire n_38461;
wire n_38462;
wire n_38463;
wire n_38466;
wire n_38467;
wire n_38468;
wire n_38469;
wire n_3847;
wire n_38470;
wire n_38471;
wire n_38472;
wire n_38473;
wire n_38474;
wire n_38475;
wire n_38476;
wire n_38477;
wire n_38478;
wire n_38479;
wire n_3848;
wire n_38480;
wire n_38481;
wire n_38482;
wire n_38483;
wire n_38484;
wire n_38485;
wire n_38486;
wire n_3849;
wire n_38490;
wire n_38491;
wire n_38492;
wire n_38493;
wire n_38494;
wire n_38495;
wire n_38496;
wire n_38497;
wire n_38498;
wire n_38499;
wire n_385;
wire n_3850;
wire n_38500;
wire n_38501;
wire n_38502;
wire n_38503;
wire n_38504;
wire n_38506;
wire n_38508;
wire n_38509;
wire n_3851;
wire n_38510;
wire n_38511;
wire n_38512;
wire n_38514;
wire n_38515;
wire n_38516;
wire n_38517;
wire n_38518;
wire n_38519;
wire n_3852;
wire n_38521;
wire n_38522;
wire n_38523;
wire TIMEBOOST_net_289;
wire n_38525;
wire n_38526;
wire n_38527;
wire n_3853;
wire n_38530;
wire n_38531;
wire n_38534;
wire TIMEBOOST_net_257;
wire n_38537;
wire n_38538;
wire n_38539;
wire n_3854;
wire n_38540;
wire n_38541;
wire n_38543;
wire n_38545;
wire n_38546;
wire n_38547;
wire n_38548;
wire n_3855;
wire n_38550;
wire TIMEBOOST_net_2775;
wire TIMEBOOST_net_1103;
wire n_38553;
wire n_38554;
wire n_38555;
wire n_38556;
wire n_3856;
wire n_38562;
wire n_38563;
wire n_38564;
wire TIMEBOOST_net_1606;
wire TIMEBOOST_net_2504;
wire n_38569;
wire n_3857;
wire n_38570;
wire n_38571;
wire n_38572;
wire n_38573;
wire n_38574;
wire n_38575;
wire n_38577;
wire n_38579;
wire n_3858;
wire n_38580;
wire n_38583;
wire n_38584;
wire n_38586;
wire n_38587;
wire n_38588;
wire n_38589;
wire n_3859;
wire TIMEBOOST_net_1016;
wire n_38591;
wire n_38592;
wire n_38594;
wire n_38595;
wire n_38596;
wire n_38597;
wire n_38598;
wire n_386;
wire n_3860;
wire n_38601;
wire n_38602;
wire n_38603;
wire n_38604;
wire n_38605;
wire n_38606;
wire n_38608;
wire n_38609;
wire n_38610;
wire n_38612;
wire TIMEBOOST_net_312;
wire TIMEBOOST_net_2440;
wire n_38615;
wire n_38616;
wire TIMEBOOST_net_2161;
wire n_3862;
wire n_38622;
wire n_38623;
wire n_38624;
wire TIMEBOOST_net_1111;
wire n_38626;
wire n_38627;
wire n_38628;
wire n_38629;
wire n_3863;
wire n_38630;
wire TIMEBOOST_net_298;
wire n_38633;
wire n_38635;
wire n_38636;
wire n_38637;
wire n_38639;
wire n_3864;
wire n_38640;
wire n_38641;
wire n_38643;
wire TIMEBOOST_net_315;
wire TIMEBOOST_net_2384;
wire n_38647;
wire n_38648;
wire n_38649;
wire n_38650;
wire n_38651;
wire n_38652;
wire n_38653;
wire n_38654;
wire n_38655;
wire n_38656;
wire n_38657;
wire n_38658;
wire n_38659;
wire n_38660;
wire n_38662;
wire n_38663;
wire n_38664;
wire n_38665;
wire n_38666;
wire n_38667;
wire n_38668;
wire n_38669;
wire n_3867;
wire n_38670;
wire n_38671;
wire n_38673;
wire n_38674;
wire n_38676;
wire n_38677;
wire n_38678;
wire TIMEBOOST_net_1685;
wire n_38680;
wire n_38683;
wire n_38685;
wire n_38686;
wire n_38687;
wire TIMEBOOST_net_1958;
wire n_38689;
wire n_38690;
wire n_38691;
wire n_38692;
wire n_38693;
wire n_38694;
wire n_38695;
wire n_38696;
wire n_38697;
wire n_38698;
wire n_387;
wire n_38703;
wire n_38704;
wire n_38705;
wire n_38706;
wire n_38707;
wire n_38708;
wire n_38709;
wire n_3871;
wire n_38710;
wire n_38711;
wire n_38712;
wire n_38713;
wire n_38714;
wire n_38715;
wire n_38716;
wire n_38717;
wire n_38719;
wire n_3872;
wire n_38720;
wire n_38721;
wire n_38722;
wire TIMEBOOST_net_2146;
wire n_38724;
wire n_38725;
wire n_38726;
wire n_38727;
wire n_38728;
wire n_38729;
wire n_3873;
wire n_38730;
wire n_38731;
wire n_38732;
wire n_38734;
wire n_38735;
wire n_38736;
wire n_38737;
wire n_38738;
wire n_38739;
wire n_3874;
wire n_38740;
wire n_38741;
wire n_38742;
wire n_38743;
wire n_38744;
wire n_38745;
wire n_38746;
wire n_38747;
wire n_38748;
wire n_38749;
wire n_3875;
wire n_38750;
wire n_38752;
wire n_38753;
wire n_38754;
wire n_38755;
wire n_38756;
wire n_38757;
wire n_38758;
wire n_38759;
wire n_38760;
wire n_38761;
wire n_38762;
wire n_38763;
wire n_38764;
wire n_38765;
wire n_38766;
wire n_38767;
wire n_38768;
wire n_38769;
wire n_3877;
wire n_38770;
wire TIMEBOOST_net_1156;
wire n_38772;
wire n_38773;
wire n_38774;
wire n_38775;
wire n_38776;
wire n_38778;
wire n_38779;
wire n_38780;
wire n_38781;
wire n_38782;
wire n_38783;
wire n_38784;
wire n_38785;
wire n_38786;
wire n_38787;
wire n_38788;
wire TIMEBOOST_net_1672;
wire n_3879;
wire n_38790;
wire n_38791;
wire n_38792;
wire n_38793;
wire n_38794;
wire n_38795;
wire n_38796;
wire n_38797;
wire n_38798;
wire n_38799;
wire n_3880;
wire n_38800;
wire n_38801;
wire n_38802;
wire n_38803;
wire n_38804;
wire n_38805;
wire n_38806;
wire n_38807;
wire n_38808;
wire n_38809;
wire n_3881;
wire n_38811;
wire n_38812;
wire n_38813;
wire n_38816;
wire n_38817;
wire n_38818;
wire n_3882;
wire n_38820;
wire n_38821;
wire n_38828;
wire n_38829;
wire n_3883;
wire n_38830;
wire n_38831;
wire n_38832;
wire n_38833;
wire n_38834;
wire n_38835;
wire n_38836;
wire n_38837;
wire n_3884;
wire n_38841;
wire n_38842;
wire n_38843;
wire n_38844;
wire n_38845;
wire n_38847;
wire n_3885;
wire n_38852;
wire n_38853;
wire n_38856;
wire n_38857;
wire n_38858;
wire n_38859;
wire n_3886;
wire n_38860;
wire n_38862;
wire n_38863;
wire n_38864;
wire n_38865;
wire n_38868;
wire n_38869;
wire n_3887;
wire n_38872;
wire n_38873;
wire n_38876;
wire n_38877;
wire n_38879;
wire TIMEBOOST_net_386;
wire n_38880;
wire n_38881;
wire n_38882;
wire n_38883;
wire n_38884;
wire n_38885;
wire n_38886;
wire n_38887;
wire n_38888;
wire n_38889;
wire n_38890;
wire n_38892;
wire n_38893;
wire n_38894;
wire n_38895;
wire n_38896;
wire n_38897;
wire n_389;
wire n_3890;
wire n_38900;
wire n_38901;
wire n_38902;
wire n_38903;
wire n_38904;
wire n_38905;
wire n_38906;
wire n_38907;
wire n_38908;
wire n_38909;
wire n_3891;
wire n_38912;
wire n_38915;
wire n_38916;
wire n_38917;
wire n_38919;
wire n_38921;
wire n_38922;
wire n_38924;
wire n_38925;
wire n_38926;
wire n_38927;
wire n_38928;
wire n_38929;
wire TIMEBOOST_net_1669;
wire n_38930;
wire TIMEBOOST_net_1701;
wire n_38932;
wire TIMEBOOST_net_382;
wire n_38934;
wire n_38937;
wire n_38939;
wire n_3894;
wire n_38940;
wire n_38941;
wire n_38942;
wire n_38943;
wire n_38950;
wire n_38951;
wire n_38952;
wire n_38953;
wire TIMEBOOST_net_2403;
wire n_38955;
wire n_38956;
wire n_38957;
wire n_38958;
wire n_38959;
wire n_3896;
wire n_38960;
wire TIMEBOOST_net_2942;
wire n_38963;
wire n_38964;
wire TIMEBOOST_net_1164;
wire n_38966;
wire n_38967;
wire n_38968;
wire n_38969;
wire n_3897;
wire n_38970;
wire n_38971;
wire n_38973;
wire n_38974;
wire n_38975;
wire n_38976;
wire n_38978;
wire n_38980;
wire n_38981;
wire n_38983;
wire n_38984;
wire n_38985;
wire n_38986;
wire n_38987;
wire n_38988;
wire n_38989;
wire n_3899;
wire n_38990;
wire n_38991;
wire n_38992;
wire n_38993;
wire n_38994;
wire n_38995;
wire n_38996;
wire n_38997;
wire n_38998;
wire n_38999;
wire n_390;
wire n_3900;
wire n_39000;
wire n_39001;
wire n_39002;
wire n_39003;
wire n_39004;
wire n_39005;
wire n_39006;
wire n_39007;
wire n_39008;
wire n_39009;
wire TIMEBOOST_net_1184;
wire n_39010;
wire n_39012;
wire n_39013;
wire TIMEBOOST_net_1163;
wire n_39016;
wire n_3902;
wire n_39021;
wire n_39025;
wire n_39026;
wire n_39027;
wire n_39028;
wire n_3903;
wire n_39030;
wire n_39032;
wire n_39033;
wire n_39034;
wire n_39035;
wire n_39037;
wire TIMEBOOST_net_2220;
wire n_3904;
wire n_39040;
wire n_39041;
wire n_39042;
wire n_39043;
wire n_39044;
wire n_39045;
wire n_39046;
wire n_39047;
wire n_39048;
wire n_39049;
wire n_3905;
wire n_39050;
wire n_39051;
wire n_39053;
wire TIMEBOOST_net_355;
wire n_39055;
wire n_39056;
wire n_39057;
wire n_39058;
wire n_39059;
wire n_39060;
wire n_39061;
wire n_39062;
wire n_39063;
wire n_39064;
wire n_39065;
wire n_39068;
wire n_39069;
wire n_39072;
wire n_39074;
wire n_39075;
wire n_39076;
wire n_39077;
wire n_39078;
wire n_39079;
wire n_39080;
wire n_39081;
wire n_39083;
wire n_39084;
wire n_39085;
wire n_39086;
wire n_39087;
wire n_39088;
wire n_39089;
wire n_3909;
wire TIMEBOOST_net_1195;
wire n_39092;
wire n_39094;
wire n_39095;
wire n_39097;
wire n_39098;
wire n_391;
wire n_39100;
wire n_39103;
wire n_39104;
wire n_39105;
wire n_39106;
wire n_39107;
wire n_39108;
wire n_39109;
wire n_3911;
wire n_39110;
wire n_39111;
wire n_39112;
wire n_39113;
wire n_39114;
wire n_39118;
wire n_39120;
wire n_39121;
wire n_39123;
wire n_39125;
wire n_39126;
wire n_39129;
wire n_3913;
wire n_39130;
wire n_39131;
wire TIMEBOOST_net_2078;
wire n_39133;
wire n_39134;
wire n_39135;
wire n_39137;
wire n_39138;
wire n_39139;
wire n_3914;
wire n_39140;
wire n_39141;
wire n_39142;
wire n_39143;
wire n_39144;
wire n_39145;
wire n_39146;
wire n_39147;
wire n_39148;
wire n_39149;
wire n_3915;
wire n_39150;
wire n_39151;
wire n_39152;
wire n_39154;
wire n_39155;
wire n_39156;
wire n_39157;
wire n_39158;
wire TIMEBOOST_net_1627;
wire n_39161;
wire n_39162;
wire n_39163;
wire n_39164;
wire n_39165;
wire n_39166;
wire n_39167;
wire n_39168;
wire n_3917;
wire n_39173;
wire n_39175;
wire n_39176;
wire n_39177;
wire n_39179;
wire n_3918;
wire TIMEBOOST_net_388;
wire n_39181;
wire n_39183;
wire n_39184;
wire n_39185;
wire n_39186;
wire n_39187;
wire n_39189;
wire n_3919;
wire n_39191;
wire n_39192;
wire n_39193;
wire n_39194;
wire n_39195;
wire TIMEBOOST_net_387;
wire n_39199;
wire n_392;
wire n_3920;
wire n_39200;
wire n_39201;
wire n_39202;
wire n_39203;
wire n_39204;
wire n_39205;
wire n_39206;
wire n_39207;
wire n_39208;
wire n_39209;
wire n_39210;
wire n_39211;
wire n_39212;
wire n_39213;
wire n_39214;
wire n_39215;
wire n_39216;
wire n_39217;
wire n_39218;
wire n_39219;
wire n_3922;
wire n_39220;
wire n_39221;
wire n_39222;
wire n_39223;
wire n_39226;
wire n_39227;
wire n_39228;
wire n_39229;
wire n_39230;
wire n_39232;
wire n_39233;
wire n_39234;
wire TIMEBOOST_net_2502;
wire n_39236;
wire n_39237;
wire n_39239;
wire n_39242;
wire n_39243;
wire n_39244;
wire n_39245;
wire n_39246;
wire n_39247;
wire n_39248;
wire n_39249;
wire n_39250;
wire n_39251;
wire n_39252;
wire n_39253;
wire n_39254;
wire n_39256;
wire n_39257;
wire n_39258;
wire n_39259;
wire n_3926;
wire n_39260;
wire n_39261;
wire TIMEBOOST_net_2147;
wire n_39264;
wire n_39265;
wire n_39267;
wire n_39268;
wire n_39269;
wire TIMEBOOST_net_2034;
wire n_39270;
wire n_39271;
wire n_39272;
wire n_39273;
wire n_39274;
wire n_39275;
wire n_39276;
wire n_39277;
wire n_39278;
wire n_39279;
wire n_3928;
wire n_39280;
wire n_39281;
wire TIMEBOOST_net_389;
wire n_39283;
wire n_39284;
wire n_39285;
wire n_39286;
wire n_39287;
wire n_39288;
wire n_39289;
wire n_3929;
wire n_39290;
wire n_39291;
wire n_39292;
wire n_39293;
wire TIMEBOOST_net_392;
wire TIMEBOOST_net_2879;
wire n_39297;
wire n_39298;
wire n_39299;
wire n_393;
wire n_39300;
wire n_39301;
wire n_39302;
wire n_39303;
wire n_39304;
wire n_39305;
wire n_39306;
wire n_39307;
wire n_39308;
wire n_39309;
wire n_3931;
wire n_39310;
wire n_39311;
wire n_39312;
wire n_39313;
wire n_39314;
wire n_39318;
wire n_39319;
wire TIMEBOOST_net_1259;
wire n_39320;
wire n_39321;
wire n_39322;
wire n_39323;
wire n_39324;
wire n_39326;
wire n_39329;
wire n_3933;
wire n_39330;
wire n_39331;
wire n_39332;
wire n_39333;
wire n_39334;
wire n_39335;
wire n_39336;
wire n_39337;
wire n_39338;
wire n_39339;
wire n_3934;
wire n_39340;
wire n_39341;
wire n_39342;
wire n_39343;
wire n_39345;
wire n_39346;
wire n_39347;
wire n_39349;
wire n_3935;
wire n_39350;
wire n_39351;
wire n_39352;
wire n_39353;
wire n_39354;
wire n_39355;
wire n_39356;
wire TIMEBOOST_net_1628;
wire n_39358;
wire n_39359;
wire n_39360;
wire n_39361;
wire n_39362;
wire n_39363;
wire n_39364;
wire n_39365;
wire n_39366;
wire n_39367;
wire n_39368;
wire n_39369;
wire n_39370;
wire n_39371;
wire n_39373;
wire n_39374;
wire n_39375;
wire n_39376;
wire n_39377;
wire n_39378;
wire n_39379;
wire n_39380;
wire n_39381;
wire n_39382;
wire n_39383;
wire n_39384;
wire n_39385;
wire n_39386;
wire n_39391;
wire n_39393;
wire n_39395;
wire n_39396;
wire n_39397;
wire n_39398;
wire n_39399;
wire n_3940;
wire n_39400;
wire n_39401;
wire n_39402;
wire n_39404;
wire n_39405;
wire n_39406;
wire n_39407;
wire n_39408;
wire n_3941;
wire n_39411;
wire n_39412;
wire n_39413;
wire n_39414;
wire n_39415;
wire n_39416;
wire n_39417;
wire n_3942;
wire n_39421;
wire n_39422;
wire n_39423;
wire n_39424;
wire n_39425;
wire n_39426;
wire n_39427;
wire n_39428;
wire n_39429;
wire n_3943;
wire n_39430;
wire n_39431;
wire n_39433;
wire n_39434;
wire n_39435;
wire n_39436;
wire n_39437;
wire n_39438;
wire n_39439;
wire n_3944;
wire n_39440;
wire n_39441;
wire n_39442;
wire n_39443;
wire n_39444;
wire n_39445;
wire n_39446;
wire n_39448;
wire n_3945;
wire n_39450;
wire n_39451;
wire n_39452;
wire n_39453;
wire n_39454;
wire n_39455;
wire n_39457;
wire n_39458;
wire n_39459;
wire n_39460;
wire n_39461;
wire n_39462;
wire n_39463;
wire n_39464;
wire n_39465;
wire n_39466;
wire n_39467;
wire n_39468;
wire n_39469;
wire n_39470;
wire n_39471;
wire n_39472;
wire n_39473;
wire n_39474;
wire n_39475;
wire n_39476;
wire n_39477;
wire n_39478;
wire n_39479;
wire n_3948;
wire n_39480;
wire n_39481;
wire n_39482;
wire n_39483;
wire n_39484;
wire n_39485;
wire n_39487;
wire n_39488;
wire n_39489;
wire n_3949;
wire n_39490;
wire n_39492;
wire n_39493;
wire n_39494;
wire n_39495;
wire n_39496;
wire n_39497;
wire TIMEBOOST_net_495;
wire TIMEBOOST_net_494;
wire n_395;
wire n_3950;
wire n_39500;
wire n_39501;
wire n_39502;
wire n_39503;
wire n_39504;
wire n_39505;
wire n_39506;
wire n_39508;
wire n_39509;
wire n_39510;
wire n_39511;
wire n_39512;
wire n_39513;
wire n_39514;
wire n_39516;
wire n_39517;
wire n_39518;
wire n_39519;
wire n_39520;
wire n_39523;
wire n_39524;
wire n_39525;
wire n_39526;
wire n_39527;
wire n_39528;
wire n_39529;
wire n_3953;
wire n_39531;
wire n_39532;
wire n_39533;
wire n_39534;
wire n_39535;
wire n_39536;
wire n_39537;
wire n_39538;
wire n_39539;
wire n_3954;
wire n_39540;
wire n_39542;
wire n_39543;
wire n_39544;
wire n_39545;
wire n_39548;
wire n_3955;
wire n_39551;
wire n_39552;
wire n_39553;
wire n_39554;
wire n_39555;
wire n_39556;
wire n_39557;
wire n_39558;
wire n_39559;
wire n_3956;
wire n_39560;
wire n_39561;
wire n_39562;
wire n_39566;
wire n_39567;
wire TIMEBOOST_net_396;
wire n_3957;
wire TIMEBOOST_net_498;
wire n_39571;
wire n_39575;
wire n_39577;
wire n_39578;
wire n_39579;
wire n_3958;
wire n_39580;
wire n_39581;
wire n_39582;
wire n_39584;
wire n_39586;
wire n_39587;
wire TIMEBOOST_net_2761;
wire n_39589;
wire n_3959;
wire n_39590;
wire n_39592;
wire n_39593;
wire n_39594;
wire TIMEBOOST_net_502;
wire n_39596;
wire n_39597;
wire n_39598;
wire n_39599;
wire n_396;
wire n_3960;
wire n_39600;
wire n_39601;
wire n_39602;
wire TIMEBOOST_net_1641;
wire TIMEBOOST_net_410;
wire n_39605;
wire TIMEBOOST_net_2053;
wire n_39607;
wire TIMEBOOST_net_1171;
wire TIMEBOOST_net_2856;
wire TIMEBOOST_net_2230;
wire n_39612;
wire n_39614;
wire TIMEBOOST_net_2076;
wire n_39616;
wire n_39617;
wire TIMEBOOST_net_2004;
wire n_39619;
wire n_39621;
wire n_39625;
wire n_39627;
wire n_39628;
wire n_39629;
wire n_3963;
wire n_39633;
wire n_39634;
wire n_39635;
wire n_39636;
wire n_39637;
wire n_39638;
wire n_39639;
wire n_3964;
wire n_39640;
wire n_39642;
wire n_39643;
wire n_39644;
wire n_39645;
wire n_39647;
wire n_39648;
wire TIMEBOOST_net_2278;
wire n_39652;
wire n_39654;
wire n_39655;
wire n_39656;
wire n_39657;
wire TIMEBOOST_net_1350;
wire n_3966;
wire TIMEBOOST_net_1713;
wire n_39661;
wire n_39662;
wire n_39664;
wire n_39665;
wire n_39667;
wire n_39668;
wire n_3967;
wire n_39672;
wire n_39674;
wire n_39675;
wire n_39676;
wire n_39677;
wire n_39678;
wire n_39679;
wire n_3968;
wire n_39680;
wire n_39681;
wire n_39683;
wire n_39684;
wire n_39685;
wire n_39689;
wire n_3969;
wire n_39690;
wire n_39691;
wire n_39692;
wire n_39693;
wire n_39694;
wire n_39695;
wire n_39697;
wire n_39698;
wire n_39699;
wire n_3970;
wire n_39701;
wire n_39702;
wire TIMEBOOST_net_2118;
wire n_39704;
wire n_39705;
wire n_39708;
wire n_39709;
wire n_3971;
wire n_39710;
wire n_39711;
wire n_39712;
wire TIMEBOOST_net_1737;
wire n_39714;
wire TIMEBOOST_net_2905;
wire n_39716;
wire n_39717;
wire n_39718;
wire n_39719;
wire TIMEBOOST_net_2082;
wire TIMEBOOST_net_970;
wire n_39722;
wire n_39723;
wire n_39724;
wire n_39725;
wire n_39727;
wire n_39728;
wire n_39729;
wire n_3973;
wire n_39730;
wire n_39731;
wire n_39732;
wire n_39733;
wire n_39734;
wire n_39735;
wire n_39736;
wire n_39737;
wire n_39738;
wire n_39739;
wire TIMEBOOST_net_411;
wire n_39740;
wire n_39741;
wire n_39742;
wire n_39743;
wire n_39744;
wire n_39745;
wire n_39746;
wire n_39747;
wire n_39748;
wire n_39749;
wire n_3975;
wire n_39750;
wire n_39751;
wire n_39752;
wire n_39753;
wire n_39754;
wire n_39755;
wire n_39756;
wire n_39757;
wire n_39758;
wire n_39759;
wire n_39760;
wire n_39761;
wire n_39762;
wire n_39763;
wire n_39764;
wire n_39765;
wire n_39766;
wire n_39767;
wire n_39768;
wire n_39769;
wire n_3977;
wire n_39770;
wire n_39771;
wire n_39772;
wire n_39773;
wire n_39774;
wire n_39775;
wire n_39776;
wire n_39777;
wire n_39778;
wire n_39779;
wire TIMEBOOST_net_1281;
wire n_39781;
wire n_39782;
wire n_39783;
wire n_39784;
wire n_39785;
wire n_39786;
wire n_39788;
wire n_39789;
wire n_3979;
wire n_39790;
wire n_39791;
wire n_39792;
wire n_39793;
wire n_39795;
wire n_39796;
wire n_39797;
wire n_39798;
wire n_39799;
wire n_398;
wire n_3980;
wire n_39800;
wire n_39801;
wire n_39802;
wire n_39803;
wire n_39804;
wire n_39805;
wire n_39806;
wire n_39807;
wire n_39808;
wire n_3981;
wire n_39810;
wire n_39811;
wire n_39812;
wire n_39814;
wire n_39815;
wire n_39816;
wire n_39817;
wire n_39818;
wire n_3982;
wire n_39820;
wire n_39822;
wire TIMEBOOST_net_1394;
wire n_39824;
wire n_39829;
wire n_3983;
wire n_39830;
wire n_39832;
wire n_39833;
wire TIMEBOOST_net_1346;
wire n_39838;
wire n_3984;
wire n_39840;
wire n_39841;
wire n_39843;
wire n_39844;
wire n_39845;
wire n_39846;
wire n_39847;
wire n_39848;
wire n_39849;
wire n_3985;
wire n_39851;
wire n_39852;
wire n_39853;
wire n_39854;
wire n_39855;
wire n_39857;
wire n_39858;
wire n_39859;
wire n_3986;
wire n_39860;
wire n_39861;
wire n_39862;
wire n_39864;
wire n_39865;
wire n_39866;
wire n_39867;
wire n_39869;
wire n_3987;
wire n_39870;
wire TIMEBOOST_net_1397;
wire n_39872;
wire n_39873;
wire n_39874;
wire n_39875;
wire n_39876;
wire n_39878;
wire TIMEBOOST_net_2614;
wire n_39881;
wire n_39882;
wire n_39889;
wire n_3989;
wire n_39890;
wire n_39891;
wire n_39892;
wire n_39893;
wire n_39894;
wire n_39895;
wire n_39896;
wire n_39897;
wire n_39898;
wire n_39899;
wire n_399;
wire n_3990;
wire n_39900;
wire n_39902;
wire n_39904;
wire n_39905;
wire TIMEBOOST_net_617;
wire n_39907;
wire n_39908;
wire n_3991;
wire n_39910;
wire TIMEBOOST_net_635;
wire n_39914;
wire n_39915;
wire n_39916;
wire n_39917;
wire n_39918;
wire n_39919;
wire n_3992;
wire n_39920;
wire n_39921;
wire n_39922;
wire n_39923;
wire n_39924;
wire n_39925;
wire n_39927;
wire n_39928;
wire n_39929;
wire n_39931;
wire n_39932;
wire n_39934;
wire n_39937;
wire n_39938;
wire n_39939;
wire n_3994;
wire n_39940;
wire n_39941;
wire TIMEBOOST_net_2303;
wire n_39944;
wire n_39945;
wire n_39947;
wire n_3995;
wire n_39950;
wire TIMEBOOST_net_621;
wire n_39953;
wire n_39954;
wire n_39955;
wire n_39956;
wire n_39958;
wire n_39959;
wire n_3996;
wire n_39960;
wire n_39961;
wire n_39962;
wire n_39964;
wire n_39965;
wire n_39966;
wire n_39967;
wire n_39968;
wire n_39969;
wire n_3997;
wire TIMEBOOST_net_1352;
wire n_39971;
wire n_39972;
wire n_39973;
wire n_39974;
wire n_39975;
wire n_39976;
wire n_39977;
wire n_39978;
wire n_3998;
wire n_39980;
wire n_39981;
wire n_39982;
wire n_39983;
wire n_39984;
wire n_39985;
wire n_39986;
wire n_39989;
wire n_39992;
wire TIMEBOOST_net_2876;
wire n_39994;
wire n_39995;
wire n_39996;
wire n_39997;
wire n_39998;
wire n_40;
wire n_400;
wire n_4000;
wire n_40001;
wire n_40002;
wire n_40003;
wire n_40004;
wire n_40005;
wire n_40006;
wire n_40007;
wire TIMEBOOST_net_2335;
wire n_40009;
wire TIMEBOOST_net_625;
wire n_40011;
wire TIMEBOOST_net_622;
wire n_40013;
wire n_40015;
wire n_40016;
wire n_40017;
wire n_40018;
wire n_40019;
wire n_40020;
wire TIMEBOOST_net_642;
wire n_40022;
wire n_40023;
wire n_40024;
wire n_40028;
wire n_40030;
wire TIMEBOOST_net_1589;
wire n_40032;
wire n_40033;
wire n_40034;
wire n_40036;
wire n_40037;
wire n_40038;
wire n_40039;
wire n_40041;
wire n_40042;
wire n_40043;
wire n_40044;
wire n_40045;
wire n_40046;
wire n_40047;
wire n_40048;
wire n_40049;
wire TIMEBOOST_net_1271;
wire n_40050;
wire n_40051;
wire n_40054;
wire n_40057;
wire n_40058;
wire n_40059;
wire n_4006;
wire n_40060;
wire n_40061;
wire n_40062;
wire n_40063;
wire n_40064;
wire n_40066;
wire n_40067;
wire n_40068;
wire n_40069;
wire n_4007;
wire n_40071;
wire n_40072;
wire n_40073;
wire n_40074;
wire n_40076;
wire n_40077;
wire n_40078;
wire n_40079;
wire n_4008;
wire n_40080;
wire n_40081;
wire n_40083;
wire n_40084;
wire n_40085;
wire n_40086;
wire n_40087;
wire n_40089;
wire n_4009;
wire n_40090;
wire n_40091;
wire n_40092;
wire n_40097;
wire n_40098;
wire TIMEBOOST_net_1783;
wire n_401;
wire n_4010;
wire n_40100;
wire n_40101;
wire n_40102;
wire n_40103;
wire n_40104;
wire n_40106;
wire n_40107;
wire n_4011;
wire n_40110;
wire n_40111;
wire n_40112;
wire n_40113;
wire n_40114;
wire n_40115;
wire n_40116;
wire n_40117;
wire n_40118;
wire n_40119;
wire n_4012;
wire n_40120;
wire n_40121;
wire n_40122;
wire n_40123;
wire n_40124;
wire n_40128;
wire n_40130;
wire n_40131;
wire n_40132;
wire n_40133;
wire n_40134;
wire TIMEBOOST_net_624;
wire n_40136;
wire n_40137;
wire n_40138;
wire n_40139;
wire n_4014;
wire n_40140;
wire n_40141;
wire n_40143;
wire n_40144;
wire n_40145;
wire n_40146;
wire n_40148;
wire n_4015;
wire n_40150;
wire n_40151;
wire n_40152;
wire n_40153;
wire n_40154;
wire TIMEBOOST_net_682;
wire n_40156;
wire n_40157;
wire n_40159;
wire n_4016;
wire n_40161;
wire n_40164;
wire n_40165;
wire n_40166;
wire TIMEBOOST_net_645;
wire n_40169;
wire n_40170;
wire n_40171;
wire n_40172;
wire n_40173;
wire n_40174;
wire TIMEBOOST_net_649;
wire n_40177;
wire n_40178;
wire n_40179;
wire n_4018;
wire n_40180;
wire n_40181;
wire n_40182;
wire n_40183;
wire n_40186;
wire n_40187;
wire n_40188;
wire n_40189;
wire n_4019;
wire n_40191;
wire n_40192;
wire n_40193;
wire n_40194;
wire n_40195;
wire n_40196;
wire n_40197;
wire n_40198;
wire n_40199;
wire n_402;
wire n_4020;
wire n_40200;
wire n_40202;
wire n_40204;
wire n_40205;
wire n_40206;
wire n_40207;
wire n_40210;
wire n_40211;
wire n_40212;
wire n_40213;
wire n_40214;
wire n_40215;
wire n_40217;
wire n_40218;
wire n_40219;
wire n_4022;
wire n_40220;
wire n_40221;
wire n_40222;
wire n_40223;
wire n_40224;
wire n_40225;
wire n_40226;
wire TIMEBOOST_net_1400;
wire n_40228;
wire n_40229;
wire n_4023;
wire n_40230;
wire n_40231;
wire n_40232;
wire n_40233;
wire n_40234;
wire n_40235;
wire n_40238;
wire n_40239;
wire n_4024;
wire n_40240;
wire n_40241;
wire n_40242;
wire n_40243;
wire n_40245;
wire n_40246;
wire n_40247;
wire n_40248;
wire n_40249;
wire n_4025;
wire n_40250;
wire n_40251;
wire TIMEBOOST_net_650;
wire n_40253;
wire n_40254;
wire n_40255;
wire n_40256;
wire n_40257;
wire n_40258;
wire n_4026;
wire n_40260;
wire n_40261;
wire n_40262;
wire n_40263;
wire n_40264;
wire n_40265;
wire n_40266;
wire n_40267;
wire n_40269;
wire n_40270;
wire n_40271;
wire n_40272;
wire n_40273;
wire n_40274;
wire n_40277;
wire n_40278;
wire n_40279;
wire n_4028;
wire n_40280;
wire n_40281;
wire n_40282;
wire n_40283;
wire n_40284;
wire n_40285;
wire n_40286;
wire n_40287;
wire n_40288;
wire n_40289;
wire n_4029;
wire n_40290;
wire n_40291;
wire n_40292;
wire n_40293;
wire n_40294;
wire n_40295;
wire n_40297;
wire n_40298;
wire n_40299;
wire n_403;
wire n_4030;
wire n_40300;
wire n_40301;
wire n_40302;
wire n_40303;
wire n_40304;
wire n_40305;
wire n_40306;
wire n_40308;
wire n_40309;
wire n_4031;
wire n_40310;
wire n_40311;
wire n_40312;
wire n_40313;
wire n_40314;
wire n_40315;
wire n_40316;
wire n_40317;
wire n_40318;
wire n_40319;
wire n_4032;
wire n_40320;
wire n_40321;
wire n_40322;
wire n_40323;
wire n_40324;
wire n_40325;
wire n_40326;
wire n_40327;
wire n_40328;
wire n_40329;
wire n_4033;
wire n_40330;
wire n_40331;
wire n_40332;
wire n_40333;
wire n_40335;
wire n_40336;
wire n_40337;
wire n_40338;
wire n_40339;
wire n_4034;
wire n_40340;
wire n_40341;
wire n_40342;
wire n_40343;
wire n_40344;
wire n_40345;
wire n_40346;
wire n_40347;
wire n_40348;
wire n_4035;
wire n_40350;
wire n_40353;
wire n_40354;
wire n_40355;
wire n_40356;
wire n_40357;
wire n_40358;
wire n_40359;
wire n_4036;
wire n_40360;
wire n_40361;
wire n_40362;
wire n_40363;
wire n_40364;
wire n_40365;
wire n_40366;
wire n_40367;
wire n_40368;
wire n_40369;
wire n_4037;
wire n_40370;
wire n_40371;
wire n_40373;
wire n_40374;
wire n_40375;
wire n_40376;
wire n_40377;
wire n_40378;
wire n_40379;
wire n_40380;
wire n_40381;
wire n_40382;
wire n_40383;
wire n_40385;
wire n_40386;
wire n_40387;
wire n_40388;
wire n_40389;
wire n_4039;
wire n_40390;
wire n_40391;
wire n_40392;
wire n_40393;
wire n_40394;
wire n_40395;
wire n_40396;
wire n_40397;
wire n_40398;
wire n_40399;
wire n_404;
wire n_40400;
wire n_40401;
wire n_40402;
wire n_40403;
wire n_40404;
wire n_40405;
wire n_40406;
wire n_40407;
wire n_40408;
wire n_40409;
wire n_4041;
wire n_40410;
wire n_40411;
wire n_40412;
wire n_40414;
wire n_40415;
wire n_40416;
wire n_40417;
wire n_40418;
wire n_40419;
wire n_4042;
wire n_40420;
wire n_40421;
wire n_40422;
wire n_40423;
wire n_40424;
wire n_40425;
wire n_40426;
wire n_40427;
wire n_40428;
wire n_40429;
wire n_40430;
wire n_40431;
wire n_40432;
wire n_40433;
wire n_40434;
wire n_40435;
wire n_40436;
wire n_40437;
wire n_40438;
wire n_40439;
wire n_4044;
wire n_40440;
wire n_40441;
wire n_40442;
wire n_40443;
wire n_40444;
wire n_40445;
wire n_40446;
wire n_40447;
wire n_40448;
wire n_40449;
wire n_4045;
wire n_40450;
wire n_40451;
wire n_40452;
wire n_40453;
wire n_40454;
wire n_40455;
wire n_40456;
wire n_40457;
wire n_40458;
wire n_40459;
wire n_4046;
wire n_40460;
wire n_40461;
wire n_40462;
wire n_40463;
wire n_40464;
wire n_40465;
wire n_40466;
wire n_40467;
wire n_40468;
wire n_40469;
wire n_40470;
wire n_40471;
wire n_40472;
wire n_40473;
wire n_40474;
wire n_40475;
wire n_40476;
wire n_40477;
wire n_40478;
wire n_40479;
wire n_40480;
wire n_40484;
wire n_40485;
wire n_40486;
wire n_40487;
wire n_40488;
wire n_40489;
wire n_4049;
wire n_40490;
wire n_40491;
wire n_40492;
wire n_40493;
wire n_40494;
wire n_40495;
wire n_40496;
wire n_40497;
wire n_40498;
wire n_40499;
wire n_405;
wire n_4050;
wire n_40500;
wire n_40501;
wire n_40502;
wire n_40503;
wire n_40504;
wire n_40505;
wire n_40506;
wire n_40507;
wire n_40508;
wire n_40509;
wire n_4051;
wire n_40510;
wire n_40511;
wire n_40512;
wire n_40513;
wire n_40514;
wire n_40515;
wire n_40516;
wire n_40517;
wire n_40518;
wire n_40519;
wire n_40520;
wire n_40521;
wire n_40522;
wire n_40523;
wire n_40524;
wire n_40525;
wire n_40526;
wire n_40527;
wire n_40528;
wire n_40529;
wire TIMEBOOST_net_1688;
wire n_40530;
wire n_40531;
wire n_40532;
wire n_40534;
wire n_40535;
wire n_40536;
wire n_40537;
wire n_40538;
wire TIMEBOOST_net_685;
wire n_4054;
wire n_40540;
wire n_40541;
wire TIMEBOOST_net_684;
wire n_40543;
wire n_40544;
wire TIMEBOOST_net_767;
wire TIMEBOOST_net_735;
wire TIMEBOOST_net_734;
wire n_40549;
wire TIMEBOOST_net_2436;
wire n_40550;
wire n_40552;
wire n_40553;
wire n_40554;
wire n_40555;
wire n_40556;
wire n_40557;
wire n_40558;
wire n_40559;
wire TIMEBOOST_net_2907;
wire n_40560;
wire n_40561;
wire n_40563;
wire n_40565;
wire n_40567;
wire n_40568;
wire n_4057;
wire n_40572;
wire n_40573;
wire n_40574;
wire n_40575;
wire n_40576;
wire n_40577;
wire n_40578;
wire n_40579;
wire n_4058;
wire n_40580;
wire n_40581;
wire n_40582;
wire n_40583;
wire n_40584;
wire n_40585;
wire n_40586;
wire n_40587;
wire n_40588;
wire n_40589;
wire n_4059;
wire n_40590;
wire n_40591;
wire n_40592;
wire n_40593;
wire n_40594;
wire n_40597;
wire n_40598;
wire n_40599;
wire n_40600;
wire n_40601;
wire n_40602;
wire n_40604;
wire n_40607;
wire n_40608;
wire n_40609;
wire n_4061;
wire n_40610;
wire n_40611;
wire n_40612;
wire n_40614;
wire n_40615;
wire n_40616;
wire n_40617;
wire n_40619;
wire n_4062;
wire n_40622;
wire n_40624;
wire TIMEBOOST_net_2;
wire n_40627;
wire n_40628;
wire n_40629;
wire n_4063;
wire n_40630;
wire n_40631;
wire n_40633;
wire n_40634;
wire n_40636;
wire n_40637;
wire n_40638;
wire n_40639;
wire TIMEBOOST_net_2501;
wire n_40641;
wire TIMEBOOST_net_1425;
wire n_40643;
wire n_40644;
wire n_40645;
wire n_40646;
wire n_40647;
wire n_40649;
wire n_4065;
wire n_40650;
wire n_40651;
wire n_40652;
wire n_40653;
wire n_40654;
wire n_40655;
wire n_40657;
wire n_40658;
wire n_40659;
wire n_40660;
wire n_40662;
wire n_40663;
wire n_40664;
wire n_40667;
wire n_40668;
wire n_40669;
wire n_40670;
wire n_40672;
wire n_40673;
wire n_40674;
wire TIMEBOOST_net_2786;
wire n_40676;
wire n_40679;
wire n_4068;
wire TIMEBOOST_net_2748;
wire n_40681;
wire n_40684;
wire n_40685;
wire n_40686;
wire n_40687;
wire n_40688;
wire n_40689;
wire n_4069;
wire n_40691;
wire n_40692;
wire n_40693;
wire n_40694;
wire n_40695;
wire n_40696;
wire n_40698;
wire n_40699;
wire n_4070;
wire n_40700;
wire n_40701;
wire n_40702;
wire TIMEBOOST_net_842;
wire n_40704;
wire n_40705;
wire n_40706;
wire n_40707;
wire n_40708;
wire n_40709;
wire n_4071;
wire n_40710;
wire n_40711;
wire n_40712;
wire n_40713;
wire n_40714;
wire n_40715;
wire n_40716;
wire n_40717;
wire n_40718;
wire n_40719;
wire n_4072;
wire n_40720;
wire n_40721;
wire n_40723;
wire n_40724;
wire n_40725;
wire n_40726;
wire n_40727;
wire n_40728;
wire n_40729;
wire n_4073;
wire n_40730;
wire n_40732;
wire n_40734;
wire n_40735;
wire n_40737;
wire n_40738;
wire n_40739;
wire TIMEBOOST_net_323;
wire n_40740;
wire n_40741;
wire n_40742;
wire n_40743;
wire n_40744;
wire TIMEBOOST_net_2634;
wire TIMEBOOST_net_38;
wire TIMEBOOST_net_48;
wire n_40749;
wire n_4075;
wire n_40750;
wire n_40751;
wire n_40753;
wire n_40754;
wire n_40756;
wire n_40757;
wire n_40758;
wire TIMEBOOST_net_1465;
wire n_40761;
wire TIMEBOOST_net_2955;
wire n_40763;
wire n_40765;
wire n_40766;
wire n_40767;
wire n_40768;
wire n_40769;
wire TIMEBOOST_net_2033;
wire n_40770;
wire n_40771;
wire n_40772;
wire n_40773;
wire n_40774;
wire n_40775;
wire n_40776;
wire n_40777;
wire n_4078;
wire n_40780;
wire n_40781;
wire n_40782;
wire n_40783;
wire n_40784;
wire n_40785;
wire n_40786;
wire n_40787;
wire n_40788;
wire n_40789;
wire n_40790;
wire n_40791;
wire n_40792;
wire n_40794;
wire n_40795;
wire n_40796;
wire n_40797;
wire n_40798;
wire n_40799;
wire n_408;
wire n_4080;
wire n_40800;
wire n_40801;
wire n_40802;
wire n_40803;
wire n_40805;
wire n_40806;
wire n_40807;
wire n_40808;
wire n_40809;
wire n_4081;
wire n_40810;
wire n_40811;
wire n_40812;
wire n_40813;
wire n_40814;
wire n_40815;
wire n_40816;
wire TIMEBOOST_net_824;
wire n_4082;
wire n_40820;
wire n_40822;
wire n_40823;
wire n_40824;
wire n_40825;
wire n_40826;
wire n_40827;
wire n_40828;
wire n_40829;
wire n_4083;
wire n_40830;
wire n_40831;
wire n_40832;
wire n_40833;
wire n_40834;
wire n_40837;
wire n_40838;
wire n_4084;
wire n_40840;
wire n_40841;
wire n_40842;
wire n_40843;
wire n_40845;
wire n_40846;
wire n_40847;
wire n_40848;
wire n_40849;
wire n_4085;
wire n_40850;
wire n_40851;
wire n_40852;
wire n_40853;
wire n_40856;
wire n_40857;
wire n_40858;
wire n_40859;
wire n_40860;
wire n_40861;
wire n_40862;
wire n_40863;
wire n_40864;
wire n_40865;
wire n_40866;
wire n_40867;
wire n_40868;
wire n_40869;
wire n_4087;
wire n_40872;
wire n_40873;
wire n_40875;
wire n_40876;
wire n_40877;
wire n_40878;
wire n_4088;
wire n_40881;
wire n_40882;
wire n_40883;
wire n_40884;
wire n_40885;
wire n_40886;
wire n_40887;
wire n_40888;
wire n_40889;
wire n_4089;
wire n_40890;
wire n_40891;
wire n_40892;
wire n_40893;
wire n_40894;
wire n_40895;
wire n_40896;
wire n_40897;
wire n_409;
wire n_4090;
wire n_40900;
wire n_40901;
wire n_40902;
wire n_40903;
wire n_40904;
wire n_40905;
wire n_40906;
wire n_40907;
wire n_40908;
wire n_40909;
wire n_4091;
wire n_40910;
wire n_40911;
wire n_40912;
wire n_40913;
wire n_40914;
wire n_40915;
wire n_40917;
wire n_40918;
wire n_40919;
wire n_4092;
wire n_40921;
wire n_40922;
wire n_40923;
wire n_40924;
wire n_40925;
wire n_40926;
wire n_40928;
wire n_40929;
wire n_4093;
wire n_40930;
wire n_40932;
wire n_40933;
wire n_40934;
wire n_40935;
wire n_40936;
wire n_40938;
wire n_40939;
wire TIMEBOOST_net_1599;
wire n_40940;
wire n_40941;
wire n_40942;
wire n_40943;
wire n_40944;
wire n_40945;
wire TIMEBOOST_net_1986;
wire n_40949;
wire n_4095;
wire n_40950;
wire n_40952;
wire n_40953;
wire n_40954;
wire n_40955;
wire n_40956;
wire n_40957;
wire n_40958;
wire n_40959;
wire n_4096;
wire n_40960;
wire n_40961;
wire n_40962;
wire n_40963;
wire n_40964;
wire n_40969;
wire n_4097;
wire n_40970;
wire n_40971;
wire n_40972;
wire n_40975;
wire n_40976;
wire n_40978;
wire n_40979;
wire n_4098;
wire n_40981;
wire n_40982;
wire n_40983;
wire n_40984;
wire n_40986;
wire n_40988;
wire n_40989;
wire n_4099;
wire n_40990;
wire n_40991;
wire n_40992;
wire n_40993;
wire n_40995;
wire n_40996;
wire n_40997;
wire n_40998;
wire n_40999;
wire n_410;
wire n_4100;
wire n_41000;
wire n_41001;
wire n_41002;
wire n_41003;
wire n_41006;
wire n_41007;
wire n_41008;
wire n_41009;
wire n_4101;
wire n_41010;
wire n_41011;
wire n_41012;
wire n_41013;
wire n_41014;
wire n_41015;
wire n_41016;
wire n_41017;
wire n_41018;
wire n_41022;
wire n_41023;
wire n_41026;
wire n_41027;
wire n_41028;
wire n_41029;
wire n_4103;
wire n_41030;
wire n_41031;
wire n_41032;
wire n_41033;
wire n_41036;
wire n_41037;
wire n_41038;
wire n_41039;
wire n_4104;
wire n_41040;
wire n_41041;
wire n_41042;
wire n_41043;
wire n_41044;
wire n_41045;
wire n_41046;
wire n_41047;
wire n_41048;
wire n_41049;
wire n_41050;
wire n_41051;
wire n_41052;
wire n_41053;
wire n_41054;
wire n_41055;
wire n_41056;
wire n_41057;
wire n_41058;
wire n_41059;
wire n_4106;
wire n_41060;
wire n_41061;
wire n_41062;
wire n_41063;
wire n_41064;
wire n_41065;
wire n_4107;
wire n_41070;
wire n_41071;
wire n_41072;
wire n_41073;
wire n_41074;
wire n_41075;
wire n_41076;
wire n_41077;
wire n_41078;
wire n_41079;
wire n_4108;
wire n_41080;
wire n_41081;
wire n_41082;
wire n_41083;
wire n_41084;
wire n_41085;
wire n_41086;
wire n_41087;
wire n_41088;
wire n_41089;
wire n_41090;
wire n_41091;
wire n_41092;
wire n_41093;
wire n_41094;
wire n_41095;
wire n_41096;
wire n_41097;
wire n_41098;
wire n_41099;
wire n_411;
wire n_4110;
wire n_41100;
wire n_41101;
wire n_41102;
wire n_41103;
wire n_41104;
wire n_41107;
wire n_41108;
wire n_41109;
wire n_4111;
wire n_41110;
wire n_41111;
wire n_41112;
wire n_41113;
wire n_41114;
wire n_41116;
wire n_41117;
wire n_41118;
wire n_41119;
wire n_4112;
wire n_41120;
wire n_41121;
wire n_41123;
wire n_41124;
wire n_41125;
wire n_41126;
wire n_41127;
wire n_41128;
wire n_41129;
wire n_4113;
wire n_41130;
wire n_41131;
wire n_41132;
wire n_41133;
wire n_41134;
wire n_41135;
wire n_41136;
wire n_41137;
wire n_41138;
wire n_41139;
wire n_4114;
wire n_41140;
wire n_41141;
wire n_41142;
wire n_41143;
wire n_41144;
wire n_41145;
wire n_41146;
wire n_41147;
wire n_41148;
wire n_41149;
wire n_4115;
wire n_41150;
wire n_41151;
wire n_41152;
wire n_41153;
wire n_41154;
wire n_41155;
wire n_41156;
wire n_41157;
wire n_41158;
wire n_41159;
wire n_4116;
wire n_41160;
wire n_41161;
wire n_41162;
wire n_41163;
wire n_41164;
wire n_41165;
wire n_41166;
wire n_41167;
wire n_41168;
wire n_41169;
wire n_4117;
wire n_41170;
wire n_41171;
wire TIMEBOOST_net_78;
wire n_41173;
wire n_41174;
wire n_41175;
wire n_41176;
wire n_41177;
wire n_41178;
wire n_41179;
wire n_4118;
wire n_41180;
wire n_41183;
wire n_41184;
wire n_41185;
wire n_41186;
wire n_41187;
wire n_4119;
wire n_41190;
wire n_41191;
wire n_41192;
wire n_41193;
wire n_41194;
wire n_41195;
wire n_41196;
wire TIMEBOOST_net_1513;
wire n_41198;
wire n_41199;
wire n_412;
wire TIMEBOOST_net_1778;
wire n_41201;
wire n_41202;
wire n_41203;
wire n_41204;
wire n_41205;
wire n_41206;
wire n_41207;
wire n_41208;
wire TIMEBOOST_net_1776;
wire n_4121;
wire n_41211;
wire n_41212;
wire n_41213;
wire n_41215;
wire n_41217;
wire n_41218;
wire n_41219;
wire n_4122;
wire n_41220;
wire n_41221;
wire n_41222;
wire n_41223;
wire n_41224;
wire n_41225;
wire n_41226;
wire n_41227;
wire n_41228;
wire n_41229;
wire n_41230;
wire n_41231;
wire n_41232;
wire n_41233;
wire n_41234;
wire n_41235;
wire n_41236;
wire n_41237;
wire n_41238;
wire n_41239;
wire n_41240;
wire n_41241;
wire n_41242;
wire n_41243;
wire n_41244;
wire n_41245;
wire n_41246;
wire n_41247;
wire n_41248;
wire n_41249;
wire n_4125;
wire n_41250;
wire n_41251;
wire n_41252;
wire n_41253;
wire n_41254;
wire n_41255;
wire n_41256;
wire n_41257;
wire n_41258;
wire n_4126;
wire n_41260;
wire n_41261;
wire n_41262;
wire n_41263;
wire n_41264;
wire n_41265;
wire n_41266;
wire n_41267;
wire n_41268;
wire n_41269;
wire n_4127;
wire n_41270;
wire n_41271;
wire n_41272;
wire n_41273;
wire n_41274;
wire n_41275;
wire n_41276;
wire n_41277;
wire n_41278;
wire n_41279;
wire n_4128;
wire n_41280;
wire n_41281;
wire n_41282;
wire n_41283;
wire n_41284;
wire n_41285;
wire n_41286;
wire n_41287;
wire n_41288;
wire n_41289;
wire n_4129;
wire n_41290;
wire n_41291;
wire n_41292;
wire n_41293;
wire n_41294;
wire TIMEBOOST_net_2441;
wire n_41296;
wire n_41297;
wire n_41298;
wire n_41299;
wire n_413;
wire TIMEBOOST_net_1172;
wire n_41300;
wire n_41301;
wire n_41302;
wire n_41303;
wire n_41304;
wire n_41305;
wire n_41306;
wire n_41307;
wire n_41308;
wire n_41309;
wire n_4131;
wire n_41310;
wire n_41311;
wire n_41312;
wire n_41313;
wire n_41314;
wire n_41316;
wire n_41317;
wire n_41319;
wire n_4132;
wire n_41320;
wire n_41321;
wire n_41322;
wire n_41324;
wire n_41325;
wire n_41326;
wire n_41327;
wire n_41328;
wire TIMEBOOST_net_101;
wire n_4133;
wire n_41330;
wire n_41333;
wire n_41337;
wire n_41339;
wire n_4134;
wire n_41341;
wire n_41342;
wire n_41343;
wire n_41344;
wire n_41345;
wire n_41347;
wire n_41348;
wire n_41349;
wire n_41353;
wire n_41355;
wire n_41356;
wire n_41357;
wire n_41358;
wire n_41359;
wire n_4136;
wire n_41360;
wire n_41361;
wire n_41362;
wire n_41364;
wire n_41365;
wire n_41366;
wire n_41367;
wire n_41369;
wire n_41370;
wire n_41371;
wire n_41372;
wire n_41374;
wire n_41375;
wire TIMEBOOST_net_2104;
wire n_41378;
wire n_41379;
wire TIMEBOOST_net_457;
wire n_41380;
wire n_41381;
wire n_41382;
wire n_41383;
wire n_41384;
wire n_41385;
wire n_41386;
wire n_41388;
wire n_41389;
wire n_4139;
wire n_41390;
wire n_41391;
wire n_41392;
wire n_41397;
wire n_41398;
wire n_41399;
wire n_414;
wire n_4140;
wire n_41400;
wire n_41401;
wire n_41402;
wire n_41405;
wire n_41406;
wire n_41407;
wire n_41408;
wire n_41409;
wire n_41410;
wire n_41411;
wire n_41412;
wire n_41414;
wire n_41415;
wire n_41416;
wire n_41418;
wire n_41419;
wire n_4142;
wire n_41420;
wire n_41421;
wire n_41422;
wire n_41423;
wire n_41424;
wire n_41426;
wire n_41427;
wire n_41428;
wire n_4143;
wire n_41430;
wire n_41431;
wire n_41432;
wire n_41433;
wire n_41434;
wire n_41435;
wire n_41438;
wire n_4144;
wire n_41440;
wire n_41443;
wire n_41444;
wire n_41445;
wire n_41446;
wire n_41447;
wire TIMEBOOST_net_996;
wire n_41449;
wire n_4145;
wire n_41450;
wire n_41452;
wire n_41453;
wire n_41454;
wire n_41455;
wire n_41456;
wire n_41457;
wire n_41458;
wire n_4146;
wire n_41460;
wire n_41461;
wire n_41462;
wire n_4147;
wire n_41470;
wire n_41471;
wire n_41472;
wire n_41473;
wire n_41474;
wire n_41475;
wire n_41476;
wire n_41477;
wire n_41478;
wire n_41479;
wire n_4148;
wire n_41480;
wire n_41481;
wire n_41482;
wire n_41483;
wire n_41484;
wire n_41485;
wire n_41486;
wire n_41487;
wire n_41488;
wire n_41489;
wire n_4149;
wire n_41490;
wire n_41491;
wire n_41492;
wire n_41494;
wire n_41499;
wire n_415;
wire n_41500;
wire n_41501;
wire n_41502;
wire TIMEBOOST_net_2817;
wire n_41504;
wire n_41505;
wire n_41506;
wire n_41507;
wire n_41508;
wire n_41509;
wire n_41510;
wire n_41511;
wire n_41512;
wire n_41513;
wire n_41514;
wire n_41515;
wire n_41516;
wire n_41517;
wire n_41518;
wire n_41519;
wire n_4152;
wire n_41520;
wire n_41521;
wire n_41522;
wire n_41523;
wire n_41524;
wire n_41525;
wire n_41526;
wire n_41527;
wire n_41528;
wire n_41529;
wire n_41530;
wire n_41531;
wire n_41532;
wire n_41533;
wire n_41534;
wire n_41535;
wire n_41536;
wire n_4154;
wire n_41540;
wire n_41541;
wire n_41542;
wire n_41543;
wire n_41545;
wire n_41546;
wire n_41547;
wire n_41548;
wire n_41549;
wire n_4155;
wire n_41550;
wire n_41551;
wire n_41552;
wire n_41553;
wire n_41557;
wire n_41558;
wire n_4156;
wire n_41560;
wire n_41561;
wire n_41562;
wire n_41563;
wire n_41566;
wire n_4157;
wire n_41571;
wire n_41572;
wire n_41573;
wire n_41574;
wire n_41576;
wire n_41577;
wire n_41578;
wire n_41579;
wire n_4158;
wire n_41580;
wire n_41581;
wire n_41582;
wire n_41583;
wire n_41585;
wire n_41586;
wire n_41587;
wire n_41588;
wire n_41589;
wire n_41590;
wire n_41592;
wire n_41593;
wire n_41594;
wire n_41595;
wire n_41596;
wire n_41598;
wire n_41599;
wire n_416;
wire n_41600;
wire n_41602;
wire n_41604;
wire n_41605;
wire n_41607;
wire n_41608;
wire n_4161;
wire n_41612;
wire n_41613;
wire n_41614;
wire n_41615;
wire n_41616;
wire n_41617;
wire n_41618;
wire n_41619;
wire n_41620;
wire n_41621;
wire n_41622;
wire n_41623;
wire n_41624;
wire n_41626;
wire n_41628;
wire n_41629;
wire n_4163;
wire n_41630;
wire n_41631;
wire n_41632;
wire n_41633;
wire n_41634;
wire n_41635;
wire n_41636;
wire n_41637;
wire n_41638;
wire n_41639;
wire n_41640;
wire n_41641;
wire n_41642;
wire n_41643;
wire n_41645;
wire n_41646;
wire n_41647;
wire n_41648;
wire n_4165;
wire n_41654;
wire n_41656;
wire n_41657;
wire n_41658;
wire n_4166;
wire n_41660;
wire TIMEBOOST_net_1533;
wire n_41662;
wire n_41663;
wire n_41666;
wire n_41667;
wire n_41668;
wire n_41669;
wire n_4167;
wire n_41670;
wire n_41671;
wire n_41672;
wire n_41673;
wire n_41674;
wire n_41675;
wire n_41676;
wire n_41677;
wire n_41678;
wire n_41679;
wire n_4168;
wire n_41680;
wire n_41683;
wire n_41684;
wire n_41685;
wire n_41686;
wire n_41687;
wire n_41688;
wire TIMEBOOST_net_157;
wire n_4169;
wire n_41690;
wire n_41691;
wire n_41692;
wire n_41693;
wire n_41694;
wire n_41695;
wire n_41696;
wire TIMEBOOST_net_2751;
wire n_41698;
wire n_41699;
wire n_417;
wire n_4170;
wire n_41700;
wire n_41701;
wire TIMEBOOST_net_1557;
wire n_41703;
wire n_41704;
wire n_41705;
wire n_41706;
wire n_41707;
wire n_41708;
wire n_41709;
wire n_4171;
wire n_41710;
wire n_41711;
wire n_41712;
wire n_41713;
wire n_41715;
wire n_41716;
wire n_41717;
wire n_4172;
wire n_41721;
wire n_41722;
wire n_41723;
wire n_41724;
wire n_41725;
wire n_41727;
wire n_41729;
wire n_4173;
wire n_41730;
wire n_41731;
wire n_41732;
wire n_41733;
wire n_41734;
wire n_41735;
wire n_41736;
wire n_41737;
wire n_41738;
wire n_4174;
wire n_41740;
wire n_41741;
wire n_41742;
wire n_41743;
wire n_41744;
wire n_41745;
wire TIMEBOOST_net_1033;
wire n_41748;
wire n_41749;
wire n_4175;
wire n_41751;
wire n_41752;
wire n_41753;
wire n_41754;
wire n_41755;
wire n_41756;
wire n_41757;
wire n_41759;
wire n_4176;
wire n_41760;
wire n_41761;
wire n_41762;
wire n_41763;
wire n_41764;
wire n_41765;
wire n_41766;
wire n_41767;
wire TIMEBOOST_net_1007;
wire n_41769;
wire n_4177;
wire n_41770;
wire n_41771;
wire n_41772;
wire n_41773;
wire n_41774;
wire n_41775;
wire n_41776;
wire n_41777;
wire n_41779;
wire n_4178;
wire n_41780;
wire n_41782;
wire n_41783;
wire n_41784;
wire n_41785;
wire n_41786;
wire n_41787;
wire n_41788;
wire n_41789;
wire n_4179;
wire n_41790;
wire n_41791;
wire n_41792;
wire n_41793;
wire n_41794;
wire TIMEBOOST_net_1039;
wire n_41796;
wire n_41797;
wire n_41798;
wire n_41799;
wire n_4180;
wire n_41800;
wire n_41801;
wire n_41803;
wire n_41804;
wire n_41807;
wire n_41808;
wire n_41809;
wire n_41810;
wire n_41812;
wire n_41813;
wire n_41814;
wire TIMEBOOST_net_2553;
wire n_41816;
wire n_41817;
wire n_41818;
wire n_41819;
wire n_41820;
wire n_41822;
wire n_41823;
wire n_41824;
wire n_41825;
wire n_41826;
wire n_41827;
wire n_41828;
wire n_41830;
wire n_41831;
wire n_41832;
wire n_41833;
wire n_41834;
wire n_41835;
wire n_41836;
wire n_41837;
wire n_41838;
wire n_41839;
wire n_4184;
wire n_41840;
wire n_41841;
wire n_41842;
wire n_41843;
wire n_41844;
wire n_41845;
wire n_41846;
wire n_41847;
wire TIMEBOOST_net_414;
wire n_41850;
wire n_41851;
wire n_41852;
wire n_41853;
wire n_41854;
wire n_41856;
wire n_41857;
wire n_41858;
wire n_41859;
wire n_4186;
wire n_41860;
wire n_41861;
wire n_41862;
wire n_41863;
wire n_41864;
wire n_41865;
wire n_41866;
wire n_41867;
wire n_41868;
wire n_41869;
wire n_41870;
wire n_41871;
wire n_41872;
wire n_41873;
wire n_41874;
wire n_41875;
wire n_41876;
wire n_41877;
wire n_41878;
wire n_41879;
wire n_41881;
wire n_41882;
wire n_41884;
wire n_41885;
wire n_41886;
wire n_41887;
wire n_41888;
wire n_41889;
wire n_41890;
wire n_41891;
wire n_41892;
wire n_41893;
wire n_41894;
wire n_41895;
wire n_41896;
wire TIMEBOOST_net_2587;
wire n_41898;
wire n_41899;
wire n_419;
wire n_4190;
wire n_41900;
wire n_41901;
wire n_41902;
wire n_41903;
wire n_41904;
wire n_41905;
wire n_41906;
wire n_41907;
wire n_41908;
wire n_41909;
wire n_4191;
wire n_41910;
wire n_41911;
wire n_41912;
wire n_41915;
wire n_41916;
wire n_41917;
wire n_41918;
wire n_41919;
wire n_4192;
wire n_41920;
wire n_41921;
wire n_41922;
wire n_41923;
wire n_41924;
wire n_41925;
wire n_41926;
wire n_41927;
wire n_41928;
wire n_41929;
wire n_4193;
wire n_41930;
wire n_41931;
wire n_41932;
wire n_41933;
wire n_41934;
wire n_41936;
wire n_41939;
wire n_4194;
wire n_41940;
wire n_41941;
wire n_41943;
wire n_41944;
wire n_41945;
wire n_41946;
wire n_41947;
wire n_41948;
wire n_41949;
wire n_41952;
wire n_41953;
wire n_41954;
wire n_41955;
wire n_41956;
wire n_41957;
wire n_41958;
wire n_41960;
wire n_41961;
wire n_41962;
wire n_41963;
wire n_41964;
wire n_41965;
wire n_41966;
wire n_41967;
wire n_41968;
wire n_41969;
wire n_4197;
wire n_41970;
wire n_41971;
wire n_41972;
wire n_41973;
wire n_41974;
wire n_41976;
wire n_41977;
wire n_41978;
wire TIMEBOOST_net_182;
wire n_4198;
wire n_41980;
wire n_41981;
wire n_41982;
wire n_41983;
wire n_41984;
wire n_41985;
wire n_41986;
wire n_41987;
wire n_41988;
wire n_41989;
wire n_41990;
wire n_41991;
wire n_41992;
wire n_41993;
wire n_41994;
wire n_41995;
wire n_41996;
wire n_41997;
wire n_41998;
wire n_41999;
wire n_42;
wire n_420;
wire n_4200;
wire n_42000;
wire n_42001;
wire n_42002;
wire n_42003;
wire n_42004;
wire n_42005;
wire n_42006;
wire n_42007;
wire n_42008;
wire n_42009;
wire n_4201;
wire n_42010;
wire n_42011;
wire n_42012;
wire n_42013;
wire n_42014;
wire n_42015;
wire n_42016;
wire n_42017;
wire n_42018;
wire n_42019;
wire n_4202;
wire n_42020;
wire n_42021;
wire n_42022;
wire n_42023;
wire n_42024;
wire n_42025;
wire n_42026;
wire n_42027;
wire n_42028;
wire n_42029;
wire n_4203;
wire n_42030;
wire n_42031;
wire n_42032;
wire n_42033;
wire n_42034;
wire n_42035;
wire n_42036;
wire n_42037;
wire n_42038;
wire n_4204;
wire n_42040;
wire n_42041;
wire n_42042;
wire n_42043;
wire n_42045;
wire n_42046;
wire n_42047;
wire n_42048;
wire n_42049;
wire n_42050;
wire n_42051;
wire n_42052;
wire n_42053;
wire n_42054;
wire n_42055;
wire n_42056;
wire n_42057;
wire n_42058;
wire n_42059;
wire n_42060;
wire n_42061;
wire n_42062;
wire n_42063;
wire n_42064;
wire n_42065;
wire n_42066;
wire n_42067;
wire n_42069;
wire n_4207;
wire n_42070;
wire n_42071;
wire n_42072;
wire n_42073;
wire n_42074;
wire TIMEBOOST_net_256;
wire n_42076;
wire n_42077;
wire n_42078;
wire n_42079;
wire n_4208;
wire n_42080;
wire n_42081;
wire TIMEBOOST_net_254;
wire n_42083;
wire n_42084;
wire n_42085;
wire n_42086;
wire n_42087;
wire n_42088;
wire n_42089;
wire n_4209;
wire n_42090;
wire n_42091;
wire n_42092;
wire n_42093;
wire n_42094;
wire n_42095;
wire n_42096;
wire n_42097;
wire n_42098;
wire n_42099;
wire n_4210;
wire n_42100;
wire n_42101;
wire n_42102;
wire n_42103;
wire n_42104;
wire n_42105;
wire n_42106;
wire n_42107;
wire n_42108;
wire n_42109;
wire n_4211;
wire n_42110;
wire n_42111;
wire n_42112;
wire n_42113;
wire n_42114;
wire n_42115;
wire n_42116;
wire n_42117;
wire n_42118;
wire n_42119;
wire n_4212;
wire n_42120;
wire TIMEBOOST_net_255;
wire n_42122;
wire TIMEBOOST_net_206;
wire n_42124;
wire n_42125;
wire n_42128;
wire n_42129;
wire n_4213;
wire n_42130;
wire n_42131;
wire n_42132;
wire n_42133;
wire n_42134;
wire n_42135;
wire n_42136;
wire n_42137;
wire n_42138;
wire n_42139;
wire TIMEBOOST_net_2263;
wire TIMEBOOST_net_1047;
wire n_42141;
wire n_42142;
wire n_42143;
wire n_42144;
wire n_42145;
wire n_42146;
wire n_42147;
wire n_42148;
wire n_42149;
wire n_4215;
wire n_42150;
wire n_42151;
wire n_42152;
wire n_42153;
wire n_42154;
wire n_42155;
wire n_42156;
wire n_42157;
wire n_42158;
wire n_42159;
wire n_4216;
wire n_42160;
wire TIMEBOOST_net_1566;
wire n_42162;
wire n_42163;
wire n_42164;
wire n_42165;
wire n_42166;
wire n_42167;
wire n_42169;
wire n_4217;
wire n_42172;
wire n_42173;
wire n_42175;
wire n_42176;
wire n_42177;
wire n_42178;
wire n_42179;
wire n_4218;
wire n_42180;
wire n_42181;
wire n_42182;
wire n_42183;
wire n_42187;
wire n_42188;
wire n_42189;
wire n_42191;
wire n_42192;
wire n_42193;
wire n_42194;
wire n_42195;
wire n_42196;
wire n_42197;
wire n_42198;
wire n_42199;
wire n_422;
wire n_4220;
wire n_42201;
wire n_42202;
wire n_42203;
wire n_42204;
wire n_42205;
wire n_42206;
wire n_42207;
wire n_42208;
wire n_42209;
wire n_4221;
wire n_42210;
wire n_42211;
wire n_42212;
wire n_42213;
wire n_42214;
wire n_42215;
wire n_42216;
wire n_42218;
wire n_4222;
wire n_42220;
wire n_42221;
wire n_42222;
wire n_42223;
wire n_42225;
wire n_42226;
wire n_42227;
wire n_42232;
wire n_42233;
wire n_42234;
wire n_42235;
wire n_42236;
wire n_42237;
wire n_42238;
wire n_42239;
wire n_42240;
wire n_42241;
wire n_42242;
wire n_42247;
wire n_42248;
wire n_42249;
wire n_4225;
wire n_42251;
wire n_42252;
wire n_42253;
wire n_42254;
wire n_42258;
wire n_42259;
wire n_4226;
wire n_42260;
wire n_42261;
wire n_42262;
wire n_42263;
wire n_42264;
wire n_42265;
wire n_42266;
wire n_42267;
wire n_42268;
wire n_42270;
wire n_42271;
wire n_42272;
wire n_42274;
wire n_42276;
wire n_42277;
wire n_42279;
wire n_4228;
wire n_42280;
wire n_42283;
wire TIMEBOOST_net_1880;
wire n_42285;
wire n_42286;
wire n_42287;
wire n_42288;
wire n_4229;
wire n_42290;
wire n_42291;
wire n_42293;
wire n_42294;
wire n_42295;
wire n_42296;
wire n_42297;
wire n_42298;
wire n_42299;
wire n_423;
wire n_4230;
wire n_42300;
wire n_42302;
wire n_42303;
wire n_42304;
wire n_42306;
wire n_42307;
wire n_42308;
wire n_42309;
wire n_4231;
wire n_42310;
wire n_42311;
wire n_42312;
wire n_42314;
wire n_42316;
wire n_42317;
wire n_42318;
wire n_42321;
wire n_42323;
wire n_42327;
wire n_42328;
wire n_42329;
wire n_4233;
wire n_42330;
wire n_42332;
wire n_42333;
wire n_42334;
wire n_42335;
wire n_42336;
wire n_42337;
wire n_42339;
wire n_4234;
wire n_42340;
wire n_42341;
wire n_42342;
wire n_42343;
wire n_42344;
wire n_42348;
wire n_42349;
wire n_4235;
wire n_42350;
wire n_42351;
wire n_42352;
wire n_42353;
wire n_42354;
wire n_42355;
wire n_42356;
wire n_42357;
wire n_42358;
wire n_42359;
wire n_4236;
wire n_42360;
wire n_42362;
wire n_42363;
wire n_42364;
wire n_42366;
wire n_42367;
wire n_42368;
wire n_4237;
wire n_42370;
wire n_42372;
wire n_42373;
wire n_42374;
wire n_42375;
wire n_42377;
wire n_42378;
wire n_42379;
wire n_4238;
wire n_42381;
wire n_42383;
wire n_42384;
wire n_42385;
wire n_42386;
wire n_42387;
wire n_42388;
wire n_42389;
wire n_42390;
wire n_42391;
wire n_42392;
wire n_42394;
wire n_42395;
wire n_42396;
wire n_42397;
wire n_42398;
wire n_42399;
wire n_424;
wire n_42400;
wire n_42401;
wire n_42402;
wire n_42403;
wire n_42406;
wire n_42408;
wire n_42409;
wire TIMEBOOST_net_2695;
wire n_42410;
wire n_42412;
wire n_42413;
wire n_42414;
wire n_42416;
wire n_42417;
wire n_42418;
wire n_42419;
wire n_4242;
wire n_42420;
wire n_42421;
wire n_42422;
wire n_42423;
wire n_42425;
wire n_42426;
wire n_42427;
wire n_42428;
wire n_4243;
wire n_42433;
wire n_42434;
wire n_42435;
wire n_42437;
wire n_42440;
wire n_42441;
wire n_42442;
wire n_42443;
wire n_42444;
wire n_42445;
wire n_42446;
wire n_42447;
wire n_42448;
wire n_42449;
wire n_4245;
wire n_42450;
wire n_42451;
wire n_42453;
wire n_42454;
wire n_42455;
wire n_42459;
wire TIMEBOOST_net_1127;
wire n_42461;
wire n_42462;
wire n_42463;
wire n_42464;
wire n_42465;
wire n_42466;
wire n_42467;
wire n_42468;
wire n_42469;
wire n_4247;
wire n_42470;
wire n_42472;
wire n_42473;
wire n_42474;
wire n_42475;
wire n_42478;
wire n_4248;
wire n_42480;
wire n_42481;
wire n_42483;
wire TIMEBOOST_net_2006;
wire n_42486;
wire n_42487;
wire n_42488;
wire n_42489;
wire n_4249;
wire n_42490;
wire n_42491;
wire n_42492;
wire n_42494;
wire n_42495;
wire n_42496;
wire n_42497;
wire n_42498;
wire n_425;
wire n_42500;
wire n_42502;
wire n_42503;
wire n_42504;
wire n_42505;
wire n_42507;
wire n_42508;
wire n_42509;
wire n_42510;
wire n_42511;
wire n_42512;
wire n_42514;
wire n_42515;
wire n_42519;
wire n_4252;
wire n_42520;
wire n_42521;
wire n_42522;
wire TIMEBOOST_net_303;
wire n_42524;
wire n_42525;
wire n_42526;
wire n_42527;
wire n_42528;
wire n_42529;
wire n_4253;
wire n_42530;
wire n_42531;
wire n_42532;
wire n_42533;
wire n_42534;
wire n_42535;
wire n_42536;
wire n_42537;
wire n_42538;
wire n_42539;
wire n_4254;
wire n_42540;
wire n_42541;
wire n_42542;
wire n_42545;
wire n_42546;
wire n_42547;
wire n_42549;
wire n_4255;
wire n_42550;
wire n_42551;
wire n_42552;
wire n_42554;
wire n_42555;
wire n_42556;
wire n_42557;
wire n_42558;
wire n_42559;
wire n_4256;
wire n_42562;
wire n_42563;
wire n_42564;
wire n_42565;
wire n_42566;
wire n_42567;
wire n_42569;
wire TIMEBOOST_net_2698;
wire n_42570;
wire n_42574;
wire n_42575;
wire n_42577;
wire n_42580;
wire n_42581;
wire n_42582;
wire n_42583;
wire n_42584;
wire n_42585;
wire n_42586;
wire n_42587;
wire n_42589;
wire TIMEBOOST_net_1197;
wire n_42590;
wire n_42591;
wire n_42592;
wire n_42593;
wire n_42594;
wire n_42595;
wire n_42596;
wire n_42597;
wire n_42598;
wire n_42599;
wire n_426;
wire n_42600;
wire n_42602;
wire n_42603;
wire n_42604;
wire n_42606;
wire n_42607;
wire n_42608;
wire n_42609;
wire n_4261;
wire n_42610;
wire n_42612;
wire n_42614;
wire n_42615;
wire n_42616;
wire n_42618;
wire n_42619;
wire n_4262;
wire n_42620;
wire n_42621;
wire n_42622;
wire n_42623;
wire n_42624;
wire n_42625;
wire n_42626;
wire n_42627;
wire n_42628;
wire n_42629;
wire n_4263;
wire n_42630;
wire n_42631;
wire n_42632;
wire n_42633;
wire n_42634;
wire n_42635;
wire n_42636;
wire n_42637;
wire n_42638;
wire n_42639;
wire n_4264;
wire n_42641;
wire n_42642;
wire n_42644;
wire n_42645;
wire n_42648;
wire n_42649;
wire n_4265;
wire n_42650;
wire n_42652;
wire n_42653;
wire n_42654;
wire n_42655;
wire n_42656;
wire n_42657;
wire n_42659;
wire n_4266;
wire n_42660;
wire n_42661;
wire n_42662;
wire n_42663;
wire n_42664;
wire n_42665;
wire n_42666;
wire n_42668;
wire n_42669;
wire n_4267;
wire n_42670;
wire n_42671;
wire n_42672;
wire n_42673;
wire n_42677;
wire n_42678;
wire n_42679;
wire n_42680;
wire n_42681;
wire n_42683;
wire n_42684;
wire n_42685;
wire n_42686;
wire n_42687;
wire n_42689;
wire n_4269;
wire n_42690;
wire n_42691;
wire n_42692;
wire n_42693;
wire n_42694;
wire n_42698;
wire n_42699;
wire n_427;
wire n_4270;
wire n_42700;
wire n_42701;
wire n_42702;
wire n_42703;
wire n_42704;
wire n_42705;
wire n_42706;
wire n_42707;
wire n_42708;
wire n_4271;
wire n_42710;
wire n_42712;
wire n_42714;
wire n_42715;
wire n_42716;
wire n_42717;
wire n_42718;
wire n_42719;
wire n_4272;
wire n_42721;
wire n_42722;
wire n_42723;
wire n_42724;
wire n_42725;
wire n_42726;
wire n_42727;
wire n_42728;
wire n_42729;
wire n_4273;
wire n_42730;
wire n_42731;
wire n_42732;
wire n_42733;
wire n_42734;
wire n_42736;
wire n_42738;
wire n_4274;
wire n_42740;
wire n_42742;
wire n_42746;
wire n_42747;
wire n_42748;
wire n_42749;
wire n_4275;
wire n_42750;
wire n_42751;
wire n_42752;
wire n_42753;
wire n_42754;
wire n_42755;
wire n_42756;
wire n_42757;
wire n_42758;
wire n_42759;
wire n_4276;
wire n_42760;
wire n_42762;
wire n_42763;
wire n_42764;
wire n_42765;
wire n_42766;
wire n_42767;
wire n_42768;
wire n_42769;
wire n_4277;
wire n_42770;
wire n_42771;
wire n_42772;
wire n_42773;
wire n_42774;
wire n_42775;
wire n_42778;
wire n_42779;
wire n_42780;
wire n_42781;
wire n_42782;
wire n_42783;
wire TIMEBOOST_net_1546;
wire n_42788;
wire n_42789;
wire n_42790;
wire n_42791;
wire n_42792;
wire n_42794;
wire n_42795;
wire n_42796;
wire n_42797;
wire n_42798;
wire n_42799;
wire n_4280;
wire n_42800;
wire n_42801;
wire n_42802;
wire n_42803;
wire n_42804;
wire n_42805;
wire n_42806;
wire n_42807;
wire n_42808;
wire n_4281;
wire n_42810;
wire n_42811;
wire n_42812;
wire n_42813;
wire n_42814;
wire n_42815;
wire n_42816;
wire n_42817;
wire n_42818;
wire n_42821;
wire n_42822;
wire n_42823;
wire n_42825;
wire n_42826;
wire n_42828;
wire n_42829;
wire n_4283;
wire n_42830;
wire n_42831;
wire n_42832;
wire n_42833;
wire n_42834;
wire n_42837;
wire n_42838;
wire n_42839;
wire n_42840;
wire n_42841;
wire n_42842;
wire n_42843;
wire n_42844;
wire n_42845;
wire n_42846;
wire n_42847;
wire n_42848;
wire n_4285;
wire n_42850;
wire n_42851;
wire n_42852;
wire n_42854;
wire n_42855;
wire n_42856;
wire n_42857;
wire TIMEBOOST_net_2429;
wire n_42859;
wire n_4286;
wire n_42860;
wire n_42861;
wire n_42862;
wire n_42864;
wire n_42867;
wire n_42868;
wire n_42869;
wire n_4287;
wire n_42871;
wire n_42873;
wire n_42874;
wire n_42875;
wire n_42876;
wire n_42878;
wire n_42879;
wire n_42881;
wire n_42883;
wire n_42885;
wire n_42886;
wire n_42887;
wire n_42888;
wire n_42889;
wire n_42890;
wire n_42891;
wire n_42894;
wire n_42895;
wire n_42896;
wire n_42897;
wire n_42898;
wire n_42899;
wire n_429;
wire n_42900;
wire n_42902;
wire n_42904;
wire n_42905;
wire n_42906;
wire n_42907;
wire n_42908;
wire n_42909;
wire n_42910;
wire n_42911;
wire n_42912;
wire n_42913;
wire n_42914;
wire n_42916;
wire n_42918;
wire n_42919;
wire n_4292;
wire n_42920;
wire n_42922;
wire n_42923;
wire n_42924;
wire n_42925;
wire n_42926;
wire n_42927;
wire n_42928;
wire TIMEBOOST_net_458;
wire n_42930;
wire n_42931;
wire n_42932;
wire n_42933;
wire n_42934;
wire n_42935;
wire n_42936;
wire n_42938;
wire n_4294;
wire n_42940;
wire n_42941;
wire n_42942;
wire n_42945;
wire n_42946;
wire n_42947;
wire n_42948;
wire n_42949;
wire n_42950;
wire n_42953;
wire n_42954;
wire n_42955;
wire n_42956;
wire n_42957;
wire n_42959;
wire n_4296;
wire n_42961;
wire n_42962;
wire n_42964;
wire n_42965;
wire n_42967;
wire n_42968;
wire n_42969;
wire n_4297;
wire n_42970;
wire n_42971;
wire n_42972;
wire n_42973;
wire n_42974;
wire n_42975;
wire n_42976;
wire n_42977;
wire n_42978;
wire n_4298;
wire n_42980;
wire n_42982;
wire n_42983;
wire n_42984;
wire n_42985;
wire n_42988;
wire n_42989;
wire n_42990;
wire n_42991;
wire n_42992;
wire n_42993;
wire n_42994;
wire TIMEBOOST_net_2668;
wire n_42996;
wire n_42997;
wire n_42998;
wire n_43;
wire n_430;
wire n_4300;
wire n_43000;
wire n_43001;
wire n_43002;
wire n_43003;
wire TIMEBOOST_net_2070;
wire n_43005;
wire n_43006;
wire n_43007;
wire n_43010;
wire n_43011;
wire n_43012;
wire n_43013;
wire n_43014;
wire n_43015;
wire n_43016;
wire n_43018;
wire n_43019;
wire n_4302;
wire n_43020;
wire n_43021;
wire n_43022;
wire n_43023;
wire n_43024;
wire n_43025;
wire n_43026;
wire n_43027;
wire n_43028;
wire n_43029;
wire n_4303;
wire n_43030;
wire n_43031;
wire n_43032;
wire n_43033;
wire n_43034;
wire n_43035;
wire n_43036;
wire n_43037;
wire n_43039;
wire n_4304;
wire n_43040;
wire n_43041;
wire n_43042;
wire n_43043;
wire n_43045;
wire n_43046;
wire n_43048;
wire n_4305;
wire n_43050;
wire n_43051;
wire n_43052;
wire n_43053;
wire n_43054;
wire n_43055;
wire n_43056;
wire n_4306;
wire n_43061;
wire n_43062;
wire n_43064;
wire n_43065;
wire n_43066;
wire n_43067;
wire n_43068;
wire n_43069;
wire n_4307;
wire n_43070;
wire n_43071;
wire n_43072;
wire n_43073;
wire n_43074;
wire n_43075;
wire TIMEBOOST_net_314;
wire n_43083;
wire n_43084;
wire n_43085;
wire n_43087;
wire n_43089;
wire TIMEBOOST_net_1999;
wire n_43090;
wire n_43091;
wire n_43092;
wire TIMEBOOST_net_2260;
wire n_43094;
wire n_43095;
wire n_43096;
wire n_4310;
wire n_43102;
wire n_43103;
wire n_43104;
wire n_43106;
wire n_43108;
wire n_43110;
wire n_43111;
wire TIMEBOOST_net_1258;
wire n_43113;
wire n_43114;
wire n_43115;
wire n_43116;
wire n_43117;
wire n_43118;
wire n_43121;
wire n_43123;
wire n_43125;
wire n_43126;
wire n_43127;
wire n_43128;
wire n_43129;
wire n_4313;
wire n_43130;
wire n_43132;
wire n_43133;
wire n_43134;
wire n_43135;
wire n_43136;
wire n_43138;
wire n_43139;
wire n_4314;
wire n_43140;
wire TIMEBOOST_net_1242;
wire n_43142;
wire n_43143;
wire n_43144;
wire n_43145;
wire n_43146;
wire n_43147;
wire TIMEBOOST_net_2869;
wire n_43149;
wire TIMEBOOST_net_2757;
wire n_43150;
wire n_43151;
wire n_43152;
wire n_43153;
wire n_43154;
wire n_43155;
wire n_43156;
wire n_43157;
wire n_43158;
wire n_43159;
wire n_4316;
wire n_43162;
wire n_43164;
wire n_43165;
wire n_43166;
wire n_43168;
wire n_4317;
wire n_43170;
wire n_43171;
wire n_43172;
wire n_43174;
wire n_43177;
wire n_43178;
wire n_43179;
wire n_4318;
wire TIMEBOOST_net_489;
wire n_43181;
wire n_43182;
wire n_43183;
wire n_43184;
wire n_43185;
wire n_43186;
wire n_43187;
wire n_43188;
wire n_43189;
wire n_4319;
wire n_43190;
wire n_43191;
wire n_43192;
wire n_43193;
wire TIMEBOOST_net_1190;
wire n_43197;
wire n_43199;
wire n_432;
wire n_4320;
wire n_43200;
wire n_43202;
wire n_43203;
wire n_43204;
wire n_43205;
wire n_43206;
wire n_43208;
wire n_4321;
wire n_43211;
wire n_43213;
wire n_43214;
wire n_43215;
wire n_43216;
wire n_43217;
wire TIMEBOOST_net_514;
wire n_4322;
wire n_43220;
wire n_43221;
wire n_43222;
wire n_43223;
wire n_43224;
wire n_43225;
wire n_43226;
wire n_43227;
wire n_43228;
wire n_43229;
wire n_4323;
wire TIMEBOOST_net_2898;
wire n_43233;
wire n_43234;
wire n_43235;
wire n_43236;
wire n_43237;
wire n_43238;
wire n_43239;
wire n_4324;
wire n_43240;
wire n_43241;
wire n_43243;
wire n_43245;
wire n_43247;
wire n_43248;
wire n_4325;
wire n_43250;
wire n_43251;
wire n_43254;
wire n_43255;
wire n_43256;
wire n_43258;
wire n_43259;
wire n_43260;
wire n_43261;
wire n_43262;
wire n_43263;
wire n_43264;
wire n_43265;
wire n_43266;
wire TIMEBOOST_net_493;
wire TIMEBOOST_net_2444;
wire n_43269;
wire n_4327;
wire n_43270;
wire n_43271;
wire n_43272;
wire n_43273;
wire n_43274;
wire n_43275;
wire n_43276;
wire n_43277;
wire n_43278;
wire TIMEBOOST_net_1121;
wire n_43280;
wire n_43281;
wire n_43282;
wire n_43283;
wire n_43284;
wire n_43285;
wire n_43286;
wire n_43287;
wire n_43288;
wire n_4329;
wire n_43291;
wire n_43292;
wire n_43293;
wire n_43297;
wire n_43298;
wire n_43299;
wire n_433;
wire n_4330;
wire n_43300;
wire n_43303;
wire n_43304;
wire n_43305;
wire n_43306;
wire n_43307;
wire n_43309;
wire n_4331;
wire n_43310;
wire n_43311;
wire n_43313;
wire n_43314;
wire n_43315;
wire n_43316;
wire TIMEBOOST_net_511;
wire n_43318;
wire n_43319;
wire n_4332;
wire n_43320;
wire n_43321;
wire n_43322;
wire n_43323;
wire n_43324;
wire n_43325;
wire n_43326;
wire n_43327;
wire n_43328;
wire n_43329;
wire n_4333;
wire n_43330;
wire n_43331;
wire n_43332;
wire n_43333;
wire n_43334;
wire n_43335;
wire n_43337;
wire n_43339;
wire n_4334;
wire n_43341;
wire n_43342;
wire n_43343;
wire n_43344;
wire n_43345;
wire n_43346;
wire n_43347;
wire n_43348;
wire n_43349;
wire n_4335;
wire n_43350;
wire n_43351;
wire n_43352;
wire n_43353;
wire n_43354;
wire n_43355;
wire n_43356;
wire n_43357;
wire n_43358;
wire n_43359;
wire n_4336;
wire n_43360;
wire n_43361;
wire n_43362;
wire n_43363;
wire n_43364;
wire n_43365;
wire n_43366;
wire n_43367;
wire n_43368;
wire n_43369;
wire n_43370;
wire TIMEBOOST_net_1467;
wire n_43372;
wire n_43373;
wire n_43374;
wire n_43375;
wire n_43376;
wire n_43377;
wire n_43378;
wire n_43379;
wire n_4338;
wire n_43381;
wire n_43383;
wire n_43384;
wire n_43385;
wire n_43387;
wire n_43388;
wire n_43389;
wire n_4339;
wire n_43390;
wire n_43391;
wire TIMEBOOST_net_512;
wire n_43393;
wire n_43394;
wire n_43395;
wire n_43396;
wire n_43397;
wire n_43398;
wire n_434;
wire n_4340;
wire n_43400;
wire n_43401;
wire n_43404;
wire n_43405;
wire n_43406;
wire n_43407;
wire n_43408;
wire n_43409;
wire TIMEBOOST_net_1177;
wire n_43411;
wire n_43412;
wire n_43413;
wire n_43414;
wire n_43417;
wire n_43418;
wire n_43420;
wire n_43422;
wire n_43424;
wire n_43425;
wire n_43426;
wire n_43427;
wire n_43428;
wire n_43429;
wire n_4343;
wire n_43430;
wire n_43431;
wire n_43432;
wire n_43433;
wire n_43434;
wire n_43435;
wire n_43437;
wire n_43440;
wire n_43441;
wire n_43442;
wire n_43443;
wire n_43444;
wire n_43446;
wire n_43447;
wire n_43449;
wire n_4345;
wire n_43450;
wire n_43451;
wire n_43452;
wire n_43453;
wire n_43454;
wire n_43455;
wire n_43456;
wire n_43458;
wire n_4346;
wire n_43460;
wire n_43461;
wire n_43462;
wire n_43463;
wire n_43464;
wire n_43465;
wire n_43466;
wire n_43467;
wire n_43468;
wire n_43469;
wire n_4347;
wire n_43470;
wire n_43471;
wire n_43472;
wire n_43473;
wire n_43474;
wire n_43475;
wire n_43477;
wire n_43478;
wire n_43479;
wire n_4348;
wire n_43480;
wire TIMEBOOST_net_2273;
wire n_43482;
wire n_43483;
wire n_43484;
wire n_43485;
wire n_43486;
wire n_43488;
wire n_43489;
wire n_43490;
wire n_43492;
wire n_43493;
wire n_43494;
wire n_43495;
wire n_43497;
wire n_43499;
wire n_435;
wire n_4350;
wire n_43500;
wire n_43501;
wire TIMEBOOST_net_2583;
wire TIMEBOOST_net_1728;
wire n_43504;
wire n_43505;
wire n_43507;
wire n_43508;
wire n_4351;
wire n_43511;
wire n_43514;
wire n_43515;
wire n_43516;
wire n_43517;
wire n_43518;
wire n_43519;
wire n_4352;
wire n_43520;
wire n_43521;
wire n_43522;
wire n_43523;
wire n_43525;
wire n_43526;
wire n_43527;
wire n_43528;
wire n_43529;
wire n_4353;
wire n_43530;
wire TIMEBOOST_net_430;
wire n_43532;
wire n_43533;
wire n_43534;
wire n_43536;
wire n_43537;
wire n_43538;
wire n_43539;
wire n_43540;
wire n_43541;
wire n_43542;
wire n_43543;
wire n_43544;
wire n_43545;
wire n_43546;
wire n_43547;
wire n_43548;
wire n_43549;
wire n_4355;
wire n_43550;
wire n_43551;
wire n_43552;
wire n_43553;
wire n_43554;
wire n_43555;
wire n_43556;
wire n_43557;
wire n_43558;
wire n_43559;
wire n_43560;
wire n_43561;
wire n_43562;
wire n_43563;
wire n_43564;
wire n_43565;
wire n_43566;
wire n_43567;
wire n_43568;
wire n_43569;
wire TIMEBOOST_net_1294;
wire n_43570;
wire n_43571;
wire n_43572;
wire n_43573;
wire n_43574;
wire n_43577;
wire n_43578;
wire n_43579;
wire n_4358;
wire n_43580;
wire n_43581;
wire n_43582;
wire n_43583;
wire n_43584;
wire n_43585;
wire n_43586;
wire n_43587;
wire n_43588;
wire n_43589;
wire n_43590;
wire n_43591;
wire n_43592;
wire n_43593;
wire n_43594;
wire n_43595;
wire n_43596;
wire n_43597;
wire n_43598;
wire n_43599;
wire n_4360;
wire n_43600;
wire n_43601;
wire n_43602;
wire n_43603;
wire n_43604;
wire n_43605;
wire n_43606;
wire n_43607;
wire n_43608;
wire n_43609;
wire n_4361;
wire n_43610;
wire n_43611;
wire n_43612;
wire n_43613;
wire n_43614;
wire n_43615;
wire n_43616;
wire n_43617;
wire n_43618;
wire n_43619;
wire n_4362;
wire n_43620;
wire n_43621;
wire n_43622;
wire n_43623;
wire n_43624;
wire n_43625;
wire n_43626;
wire n_43627;
wire n_43628;
wire n_43629;
wire n_4363;
wire n_43630;
wire n_43631;
wire n_43632;
wire n_43633;
wire n_43634;
wire n_43635;
wire n_43636;
wire n_43637;
wire n_43638;
wire n_43639;
wire n_43640;
wire n_43641;
wire n_43642;
wire n_43644;
wire n_43645;
wire n_43646;
wire n_43648;
wire n_43649;
wire n_4365;
wire n_43650;
wire n_43651;
wire n_43652;
wire n_43653;
wire n_43654;
wire n_43655;
wire n_43656;
wire n_43657;
wire n_43658;
wire n_43659;
wire n_4366;
wire n_43660;
wire n_43661;
wire n_43662;
wire n_43663;
wire n_43664;
wire n_43665;
wire n_43670;
wire n_43672;
wire n_43675;
wire n_43676;
wire n_43677;
wire n_43678;
wire n_4368;
wire n_43680;
wire n_43681;
wire n_43682;
wire n_43683;
wire n_43684;
wire n_43685;
wire n_43686;
wire n_43687;
wire n_43688;
wire n_43689;
wire n_4369;
wire n_43690;
wire n_43691;
wire n_43692;
wire n_43693;
wire n_43694;
wire n_43695;
wire n_43696;
wire n_43697;
wire n_43699;
wire n_437;
wire n_43700;
wire n_43701;
wire n_43702;
wire n_43703;
wire n_43704;
wire TIMEBOOST_net_2198;
wire n_43707;
wire n_43708;
wire n_43709;
wire n_4371;
wire n_43710;
wire n_43711;
wire n_43712;
wire n_43713;
wire n_43714;
wire n_43715;
wire n_43716;
wire n_43717;
wire n_43718;
wire n_43719;
wire n_43720;
wire n_43721;
wire n_43722;
wire n_43723;
wire n_43724;
wire n_43726;
wire n_43727;
wire n_43728;
wire n_43729;
wire n_43730;
wire n_43731;
wire n_43732;
wire n_43735;
wire n_43737;
wire n_43738;
wire n_43739;
wire n_4374;
wire n_43740;
wire n_43741;
wire n_43742;
wire n_43744;
wire n_43745;
wire n_43746;
wire n_43747;
wire n_43748;
wire n_43749;
wire n_43750;
wire n_43751;
wire n_43752;
wire n_43753;
wire n_43754;
wire n_43755;
wire n_43757;
wire n_43758;
wire n_43759;
wire n_4376;
wire n_43760;
wire n_43761;
wire n_43762;
wire n_43763;
wire n_43764;
wire n_43765;
wire n_43766;
wire n_43767;
wire n_43768;
wire n_43770;
wire n_43771;
wire n_43772;
wire n_43773;
wire n_43774;
wire n_43775;
wire n_43776;
wire n_43777;
wire n_43779;
wire n_4378;
wire n_43780;
wire n_43781;
wire n_43782;
wire n_43783;
wire n_43784;
wire n_43785;
wire n_43788;
wire n_43789;
wire n_43790;
wire n_43791;
wire n_43792;
wire n_43793;
wire n_43794;
wire n_43795;
wire n_43796;
wire n_43797;
wire n_43798;
wire n_43799;
wire n_438;
wire n_4380;
wire n_43800;
wire n_43801;
wire n_43802;
wire n_43803;
wire n_43804;
wire n_43805;
wire n_43807;
wire n_43808;
wire n_43809;
wire TIMEBOOST_net_2901;
wire n_43811;
wire n_43813;
wire n_43815;
wire TIMEBOOST_net_2154;
wire n_43817;
wire n_43818;
wire n_43819;
wire n_4382;
wire n_43820;
wire n_43821;
wire n_43822;
wire n_43823;
wire n_43824;
wire n_43827;
wire n_43828;
wire n_43829;
wire n_4383;
wire n_43831;
wire n_43832;
wire n_43833;
wire n_43834;
wire n_43835;
wire n_43836;
wire n_43838;
wire n_43839;
wire n_43840;
wire n_43841;
wire n_43842;
wire n_43844;
wire n_43845;
wire n_43846;
wire n_43847;
wire n_43848;
wire n_43849;
wire n_4385;
wire n_43850;
wire n_43851;
wire n_43852;
wire n_43853;
wire n_43854;
wire n_43855;
wire n_43857;
wire n_43858;
wire n_43859;
wire n_4386;
wire n_43860;
wire n_43861;
wire n_43862;
wire n_43863;
wire n_43864;
wire n_43865;
wire n_43866;
wire n_43867;
wire n_43868;
wire n_43869;
wire n_4387;
wire n_43870;
wire n_43871;
wire n_43872;
wire n_43873;
wire n_43874;
wire n_43875;
wire n_43876;
wire n_43877;
wire n_43878;
wire n_43879;
wire n_4388;
wire n_43880;
wire n_43882;
wire n_43884;
wire n_43885;
wire n_43886;
wire n_43887;
wire n_43888;
wire n_43889;
wire n_4389;
wire n_43890;
wire n_43891;
wire n_43892;
wire n_43893;
wire n_43894;
wire n_43895;
wire n_43896;
wire n_43897;
wire n_43898;
wire n_43899;
wire n_439;
wire n_43900;
wire n_43901;
wire n_43902;
wire n_43903;
wire n_43904;
wire n_43905;
wire n_43906;
wire n_43907;
wire n_43908;
wire n_43909;
wire n_4391;
wire n_43910;
wire n_43911;
wire n_43912;
wire n_43913;
wire n_43914;
wire n_43915;
wire n_43916;
wire n_43917;
wire n_43918;
wire n_43919;
wire n_4392;
wire n_43920;
wire n_4393;
wire n_4394;
wire n_4395;
wire n_4396;
wire n_4397;
wire n_4398;
wire n_4399;
wire n_44;
wire n_4400;
wire n_4401;
wire n_4402;
wire n_44021;
wire n_44026;
wire n_44027;
wire n_44028;
wire n_44029;
wire n_4403;
wire n_44030;
wire n_44032;
wire n_44033;
wire n_44034;
wire n_44035;
wire n_44036;
wire n_44037;
wire n_44038;
wire n_44039;
wire n_4404;
wire n_44040;
wire n_44042;
wire n_44045;
wire n_44046;
wire n_4405;
wire n_44051;
wire n_44052;
wire n_44053;
wire n_44054;
wire n_44055;
wire n_44057;
wire n_44058;
wire n_44059;
wire n_44060;
wire n_44061;
wire n_4407;
wire n_44083;
wire n_441;
wire n_44100;
wire n_44102;
wire n_4411;
wire TIMEBOOST_net_1282;
wire n_44139;
wire n_44147;
wire n_44153;
wire n_44155;
wire n_44158;
wire n_4416;
wire n_44160;
wire n_44162;
wire n_44163;
wire n_44165;
wire n_44166;
wire n_44168;
wire n_4419;
wire n_442;
wire n_4420;
wire TIMEBOOST_net_2267;
wire n_44213;
wire n_44216;
wire n_44218;
wire n_44219;
wire n_4422;
wire n_44222;
wire n_4423;
wire n_4424;
wire n_4425;
wire n_44256;
wire n_44259;
wire n_4426;
wire n_44262;
wire n_44265;
wire n_44267;
wire n_44275;
wire n_44277;
wire n_4428;
wire n_44287;
wire n_44288;
wire n_4429;
wire n_44296;
wire n_443;
wire n_4430;
wire n_44309;
wire n_4431;
wire n_44311;
wire n_44312;
wire n_4432;
wire n_44327;
wire n_44329;
wire n_4433;
wire n_44334;
wire n_4434;
wire n_44344;
wire n_44346;
wire n_44347;
wire n_4435;
wire n_44352;
wire n_44354;
wire n_44355;
wire n_44356;
wire n_4436;
wire n_44360;
wire n_44364;
wire n_44365;
wire n_4437;
wire n_4438;
wire n_4439;
wire n_444;
wire n_4441;
wire n_4442;
wire n_44420;
wire n_44422;
wire n_44423;
wire n_44425;
wire n_44426;
wire n_44428;
wire n_44429;
wire n_4443;
wire n_44430;
wire n_44432;
wire n_44434;
wire n_44437;
wire n_44438;
wire n_44439;
wire n_44441;
wire n_44443;
wire n_44445;
wire n_44447;
wire TIMEBOOST_net_1179;
wire n_44450;
wire n_44451;
wire n_44453;
wire n_44454;
wire n_4446;
wire n_4447;
wire TIMEBOOST_net_2701;
wire n_4449;
wire n_44490;
wire n_44492;
wire n_44498;
wire n_445;
wire n_4451;
wire n_44511;
wire n_44516;
wire n_4452;
wire TIMEBOOST_net_460;
wire n_4454;
wire n_4457;
wire n_44570;
wire n_44575;
wire n_44576;
wire n_44579;
wire n_4458;
wire n_4459;
wire n_44592;
wire n_44594;
wire n_446;
wire n_4460;
wire n_44610;
wire n_4462;
wire n_44621;
wire n_44623;
wire n_44624;
wire n_44626;
wire n_4463;
wire n_44636;
wire n_44637;
wire n_4464;
wire n_4465;
wire n_44650;
wire n_44652;
wire n_44659;
wire n_4466;
wire n_44661;
wire n_4467;
wire n_44672;
wire n_4468;
wire n_44687;
wire n_44690;
wire n_44692;
wire n_44695;
wire n_44696;
wire n_447;
wire n_44710;
wire n_44711;
wire n_44713;
wire n_44717;
wire n_44718;
wire n_4472;
wire n_44720;
wire n_44721;
wire n_44722;
wire n_44723;
wire n_4473;
wire n_4474;
wire n_4475;
wire n_44759;
wire n_4476;
wire n_44761;
wire n_4477;
wire n_44775;
wire n_44776;
wire n_4479;
wire n_44798;
wire n_448;
wire n_4480;
wire n_44804;
wire n_44809;
wire n_4481;
wire n_44811;
wire n_44812;
wire n_44814;
wire n_44815;
wire n_4482;
wire n_44821;
wire n_44823;
wire n_44825;
wire n_44826;
wire n_44827;
wire n_44828;
wire n_44829;
wire n_4483;
wire n_44831;
wire n_44835;
wire n_4484;
wire n_44847;
wire n_44849;
wire n_4485;
wire n_44850;
wire n_44852;
wire n_44853;
wire n_44855;
wire n_4486;
wire n_44866;
wire n_44867;
wire n_44869;
wire n_4487;
wire n_44871;
wire n_44872;
wire n_44875;
wire n_44877;
wire n_4488;
wire n_44887;
wire TIMEBOOST_net_97;
wire n_4490;
wire n_4491;
wire n_4492;
wire n_44920;
wire n_44921;
wire n_44925;
wire n_44926;
wire n_4493;
wire n_4494;
wire n_44944;
wire n_44946;
wire n_4495;
wire n_44954;
wire n_44955;
wire n_44958;
wire n_4496;
wire n_44962;
wire n_4497;
wire n_4498;
wire n_4499;
wire n_44995;
wire n_44996;
wire n_45;
wire n_4500;
wire n_45002;
wire n_45003;
wire n_45008;
wire n_4501;
wire n_45010;
wire n_45012;
wire n_45013;
wire n_4502;
wire n_45023;
wire n_45024;
wire n_45026;
wire n_4503;
wire n_45032;
wire n_4504;
wire n_4505;
wire n_45050;
wire n_4506;
wire n_45060;
wire n_45065;
wire n_45066;
wire n_45067;
wire n_45069;
wire n_4507;
wire n_45070;
wire n_45072;
wire n_45073;
wire n_4508;
wire n_45080;
wire n_45081;
wire TIMEBOOST_net_2840;
wire n_45091;
wire n_451;
wire n_45101;
wire n_4511;
wire n_45118;
wire n_45120;
wire n_45132;
wire n_45134;
wire n_45135;
wire n_45139;
wire n_45145;
wire n_45146;
wire n_45149;
wire n_4515;
wire n_45153;
wire n_45155;
wire n_4516;
wire n_4517;
wire n_4518;
wire n_45180;
wire n_45181;
wire n_45185;
wire n_45186;
wire n_45188;
wire n_4519;
wire n_45190;
wire n_45192;
wire n_45194;
wire n_45198;
wire n_452;
wire n_4520;
wire n_45200;
wire n_45202;
wire n_45204;
wire n_45209;
wire TIMEBOOST_net_348;
wire n_45212;
wire n_45213;
wire n_45214;
wire n_45216;
wire n_45217;
wire n_45224;
wire TIMEBOOST_net_1699;
wire n_4524;
wire n_4525;
wire n_4526;
wire n_4528;
wire n_4529;
wire n_453;
wire n_4530;
wire n_45300;
wire n_45301;
wire n_45304;
wire n_45306;
wire n_45309;
wire n_4531;
wire n_45311;
wire n_45317;
wire n_45319;
wire n_4532;
wire n_45321;
wire n_45322;
wire n_45323;
wire n_45327;
wire n_45329;
wire n_4533;
wire n_45331;
wire n_45332;
wire TIMEBOOST_net_454;
wire n_4535;
wire n_4536;
wire n_4537;
wire n_4538;
wire n_4539;
wire n_454;
wire n_4542;
wire n_4543;
wire n_4544;
wire n_4546;
wire n_45462;
wire n_45463;
wire n_4547;
wire n_45474;
wire n_45475;
wire n_45479;
wire n_4548;
wire n_45484;
wire n_45487;
wire n_45488;
wire n_45489;
wire n_4549;
wire n_45496;
wire n_45497;
wire n_45498;
wire n_45499;
wire n_455;
wire n_4550;
wire n_45501;
wire n_45502;
wire n_45503;
wire n_45505;
wire n_45506;
wire n_45507;
wire n_45508;
wire n_45511;
wire n_45512;
wire n_45513;
wire n_45514;
wire n_45516;
wire n_45517;
wire n_45518;
wire TIMEBOOST_net_1650;
wire n_4552;
wire n_45520;
wire n_45521;
wire n_45523;
wire n_45524;
wire n_45525;
wire n_45527;
wire n_45528;
wire n_45529;
wire n_4553;
wire n_45530;
wire n_45532;
wire n_45533;
wire n_4554;
wire n_4555;
wire n_4556;
wire n_4557;
wire n_4558;
wire n_4559;
wire n_456;
wire n_4560;
wire n_4561;
wire n_45616;
wire n_45617;
wire n_45619;
wire n_4562;
wire n_45622;
wire n_45623;
wire n_45625;
wire n_45627;
wire n_4563;
wire n_45630;
wire n_45631;
wire n_45633;
wire n_4565;
wire n_4568;
wire n_45685;
wire n_45697;
wire n_457;
wire TIMEBOOST_net_1202;
wire TIMEBOOST_net_466;
wire n_45716;
wire n_45717;
wire n_45718;
wire n_4572;
wire n_4573;
wire n_45738;
wire n_45739;
wire n_4574;
wire n_45740;
wire n_45741;
wire n_45744;
wire n_45745;
wire n_45747;
wire n_45748;
wire n_4575;
wire n_45753;
wire n_45754;
wire n_45755;
wire n_45758;
wire n_4576;
wire n_4577;
wire n_4578;
wire n_4579;
wire n_458;
wire TIMEBOOST_net_2286;
wire n_45808;
wire n_45809;
wire n_4581;
wire n_45812;
wire n_45813;
wire n_45814;
wire n_45815;
wire n_45816;
wire n_45817;
wire n_45818;
wire n_45819;
wire n_4582;
wire n_45820;
wire n_45821;
wire n_45824;
wire n_45825;
wire n_45826;
wire n_45827;
wire n_45828;
wire n_4583;
wire n_45840;
wire n_45843;
wire n_45844;
wire n_45845;
wire n_45846;
wire n_4585;
wire n_45858;
wire n_45861;
wire n_45863;
wire n_45864;
wire n_45865;
wire n_45866;
wire n_4587;
wire n_45871;
wire n_45872;
wire n_45873;
wire n_45874;
wire n_45875;
wire n_45878;
wire n_45879;
wire n_4588;
wire n_45880;
wire n_45884;
wire n_45887;
wire n_45889;
wire n_4589;
wire n_45890;
wire n_45891;
wire n_45894;
wire n_45895;
wire n_45896;
wire n_45897;
wire n_45898;
wire n_45899;
wire n_4590;
wire n_45903;
wire n_4591;
wire n_4592;
wire TIMEBOOST_net_2045;
wire n_4594;
wire n_4595;
wire n_4596;
wire n_4597;
wire n_4598;
wire n_4599;
wire n_46;
wire n_460;
wire n_4600;
wire n_4601;
wire n_4602;
wire n_4603;
wire n_4604;
wire n_4605;
wire n_46055;
wire n_4606;
wire n_4608;
wire n_4609;
wire n_461;
wire n_46107;
wire n_4611;
wire n_4612;
wire n_4613;
wire n_46137;
wire n_4614;
wire n_46141;
wire n_46143;
wire n_46145;
wire n_46146;
wire n_46147;
wire n_46148;
wire n_46149;
wire n_4615;
wire n_46150;
wire n_46151;
wire n_46152;
wire n_46153;
wire n_46154;
wire n_46155;
wire n_46156;
wire n_46157;
wire n_46158;
wire n_46159;
wire n_4616;
wire n_46160;
wire n_46161;
wire n_46162;
wire n_46163;
wire n_46164;
wire n_46165;
wire n_46166;
wire n_46167;
wire n_46168;
wire n_46169;
wire n_4617;
wire n_46170;
wire n_46171;
wire n_46172;
wire n_46173;
wire n_46174;
wire n_46175;
wire n_46176;
wire n_46177;
wire n_46178;
wire n_46179;
wire n_46180;
wire n_46181;
wire n_46182;
wire n_46183;
wire n_46184;
wire n_46185;
wire n_46186;
wire n_46187;
wire n_46188;
wire n_46189;
wire n_4619;
wire n_46190;
wire n_46191;
wire n_46192;
wire n_46193;
wire n_46194;
wire n_46195;
wire n_46197;
wire n_462;
wire n_4620;
wire n_46200;
wire n_46202;
wire n_46203;
wire n_46204;
wire n_46205;
wire n_46206;
wire n_46208;
wire n_46209;
wire n_46210;
wire n_46211;
wire n_46212;
wire n_46213;
wire n_46214;
wire n_46215;
wire n_46216;
wire n_46217;
wire n_46218;
wire n_46219;
wire n_4622;
wire n_46220;
wire n_46221;
wire n_46222;
wire n_46223;
wire n_46224;
wire n_46225;
wire n_46226;
wire n_46227;
wire n_46228;
wire n_46229;
wire n_4623;
wire n_46230;
wire n_46231;
wire n_46232;
wire n_46233;
wire n_46234;
wire n_46235;
wire n_46236;
wire n_46237;
wire n_46238;
wire n_46239;
wire n_4624;
wire n_46240;
wire n_46241;
wire n_46242;
wire n_46243;
wire n_46244;
wire n_46245;
wire n_46246;
wire n_46247;
wire n_46248;
wire n_46249;
wire n_4625;
wire n_46250;
wire n_46251;
wire n_46252;
wire n_46253;
wire n_46254;
wire n_4626;
wire n_46285;
wire n_463;
wire n_4630;
wire n_4631;
wire n_4632;
wire n_46337;
wire n_4634;
wire n_46340;
wire n_46342;
wire n_46344;
wire n_46345;
wire n_46347;
wire n_46348;
wire n_46349;
wire n_4635;
wire n_46350;
wire n_46351;
wire n_46352;
wire n_46353;
wire n_46354;
wire n_46355;
wire n_46356;
wire n_46357;
wire n_46358;
wire n_46359;
wire n_4636;
wire n_46360;
wire n_46361;
wire n_46362;
wire n_46363;
wire n_46364;
wire n_46365;
wire n_46366;
wire n_46367;
wire n_46368;
wire n_46369;
wire n_46370;
wire n_46371;
wire n_46372;
wire n_46373;
wire n_46374;
wire n_46375;
wire n_46376;
wire n_46377;
wire n_46378;
wire n_46379;
wire TIMEBOOST_net_1181;
wire n_46380;
wire n_46381;
wire n_46382;
wire n_46383;
wire n_46384;
wire n_46385;
wire n_46386;
wire n_46387;
wire n_46388;
wire n_4639;
wire n_464;
wire n_4641;
wire n_46413;
wire n_46414;
wire n_46415;
wire n_46416;
wire n_46417;
wire n_46418;
wire n_46419;
wire n_4642;
wire n_46420;
wire n_46421;
wire n_46422;
wire n_46423;
wire n_46424;
wire n_46426;
wire n_46427;
wire n_4643;
wire n_4644;
wire n_4646;
wire n_4647;
wire n_4649;
wire n_465;
wire n_4650;
wire n_4652;
wire n_4653;
wire n_4654;
wire n_4656;
wire n_4657;
wire n_4658;
wire n_4659;
wire n_466;
wire n_4660;
wire n_4661;
wire n_4662;
wire n_4664;
wire n_4665;
wire n_4666;
wire n_4667;
wire n_4668;
wire n_4669;
wire n_467;
wire n_4671;
wire n_4672;
wire n_4673;
wire n_4674;
wire n_4675;
wire n_4676;
wire TIMEBOOST_net_1292;
wire n_4679;
wire n_468;
wire n_4680;
wire n_4681;
wire n_4683;
wire n_4685;
wire n_4686;
wire n_4688;
wire n_4689;
wire n_469;
wire n_4690;
wire n_4692;
wire n_4693;
wire n_46933;
wire n_46934;
wire n_46935;
wire n_46936;
wire n_46937;
wire n_46938;
wire n_46939;
wire n_46940;
wire n_46941;
wire n_46942;
wire n_46943;
wire n_46944;
wire n_46947;
wire n_46948;
wire n_46949;
wire n_4695;
wire n_46950;
wire n_46951;
wire n_46952;
wire n_46953;
wire n_46956;
wire n_46957;
wire n_46958;
wire n_46959;
wire n_4696;
wire n_46960;
wire n_46961;
wire n_46962;
wire n_46963;
wire n_46964;
wire n_46965;
wire n_46966;
wire TIMEBOOST_net_1322;
wire n_46968;
wire n_46969;
wire n_4697;
wire n_46972;
wire n_46973;
wire n_46974;
wire n_46975;
wire n_46976;
wire n_46977;
wire n_46978;
wire n_46979;
wire TIMEBOOST_net_1183;
wire n_46980;
wire n_46981;
wire n_46982;
wire n_46984;
wire n_46985;
wire n_46986;
wire n_46987;
wire n_46988;
wire n_46989;
wire n_46990;
wire n_46991;
wire n_46992;
wire n_46993;
wire n_46994;
wire n_46995;
wire n_46996;
wire n_46997;
wire n_46998;
wire n_46999;
wire n_47;
wire n_470;
wire n_4700;
wire n_47000;
wire n_47001;
wire n_47002;
wire n_47003;
wire n_47004;
wire n_47005;
wire n_47006;
wire n_47007;
wire n_47008;
wire n_47009;
wire n_47010;
wire n_47011;
wire n_47012;
wire n_47013;
wire n_47014;
wire n_47015;
wire n_47016;
wire n_47017;
wire n_47018;
wire n_47019;
wire n_4702;
wire n_47020;
wire n_47021;
wire n_47022;
wire n_47023;
wire n_47024;
wire n_47025;
wire n_47026;
wire n_47027;
wire n_4703;
wire n_4704;
wire n_4708;
wire n_4709;
wire n_471;
wire n_4710;
wire n_4713;
wire n_4714;
wire n_4715;
wire n_4716;
wire n_4717;
wire n_47174;
wire n_47175;
wire n_47176;
wire n_47177;
wire n_47179;
wire n_47180;
wire n_47181;
wire n_47182;
wire n_47183;
wire n_47184;
wire n_47185;
wire n_47186;
wire n_47187;
wire n_4719;
wire n_47195;
wire n_47197;
wire n_47199;
wire n_472;
wire n_4720;
wire n_47200;
wire n_47203;
wire n_47207;
wire n_4721;
wire n_47210;
wire n_47211;
wire n_47212;
wire n_47213;
wire n_4722;
wire n_4723;
wire n_47233;
wire n_47235;
wire n_47240;
wire n_47241;
wire n_47242;
wire n_47243;
wire n_47244;
wire n_47245;
wire n_47246;
wire n_47247;
wire n_47248;
wire n_47249;
wire n_47250;
wire n_47251;
wire n_47252;
wire n_47253;
wire n_47254;
wire n_47255;
wire n_47256;
wire n_47257;
wire n_47258;
wire n_47259;
wire n_4726;
wire n_47260;
wire n_47261;
wire n_47262;
wire n_47263;
wire n_47264;
wire n_47265;
wire n_47266;
wire n_47267;
wire n_47268;
wire n_47269;
wire n_4727;
wire n_47270;
wire n_47271;
wire n_47272;
wire n_47273;
wire n_47274;
wire n_47278;
wire n_47279;
wire n_4729;
wire n_4730;
wire n_4731;
wire n_4732;
wire TIMEBOOST_net_2880;
wire n_47332;
wire n_47333;
wire n_47334;
wire n_47335;
wire n_47336;
wire n_47337;
wire n_47340;
wire n_47341;
wire n_4735;
wire n_4736;
wire n_4739;
wire n_4740;
wire n_4741;
wire n_4742;
wire n_4743;
wire n_4745;
wire n_4746;
wire TIMEBOOST_net_1216;
wire n_475;
wire n_4750;
wire n_4751;
wire TIMEBOOST_net_557;
wire n_4753;
wire n_4754;
wire n_4756;
wire n_4757;
wire n_4759;
wire n_476;
wire n_4760;
wire n_4761;
wire n_4762;
wire n_4763;
wire n_4765;
wire n_4766;
wire n_4767;
wire TIMEBOOST_net_1704;
wire n_477;
wire n_4771;
wire TIMEBOOST_net_1200;
wire n_4773;
wire n_4774;
wire n_4775;
wire n_4776;
wire n_4777;
wire n_4779;
wire n_478;
wire n_4780;
wire n_4781;
wire n_4782;
wire n_4783;
wire n_4784;
wire n_4786;
wire n_4787;
wire n_4788;
wire n_4789;
wire n_479;
wire n_4790;
wire n_4792;
wire n_4793;
wire n_4795;
wire n_4796;
wire n_4797;
wire TIMEBOOST_net_2464;
wire n_4799;
wire n_48;
wire n_480;
wire n_4800;
wire n_4802;
wire n_4804;
wire n_4806;
wire n_4807;
wire n_4808;
wire n_4809;
wire n_481;
wire n_4810;
wire n_4811;
wire n_4812;
wire n_4814;
wire n_4815;
wire n_4816;
wire n_4817;
wire n_4818;
wire n_4819;
wire n_482;
wire n_4820;
wire n_4821;
wire n_4823;
wire n_4824;
wire n_4825;
wire n_4826;
wire n_4827;
wire n_4828;
wire n_4830;
wire n_4831;
wire n_4833;
wire n_4834;
wire n_4837;
wire n_4838;
wire n_484;
wire n_4840;
wire n_4841;
wire n_4842;
wire n_4843;
wire n_4844;
wire n_4846;
wire n_4847;
wire n_4848;
wire n_4849;
wire n_485;
wire n_4850;
wire n_4851;
wire n_4852;
wire n_4853;
wire n_4855;
wire n_4856;
wire n_4857;
wire n_4858;
wire n_4860;
wire n_4861;
wire n_4862;
wire n_4863;
wire n_4864;
wire TIMEBOOST_net_537;
wire n_4867;
wire n_4868;
wire n_4871;
wire n_4872;
wire n_4873;
wire n_4874;
wire n_4875;
wire n_4876;
wire n_4878;
wire n_4879;
wire n_488;
wire n_4880;
wire n_4881;
wire n_4884;
wire n_4885;
wire n_4886;
wire n_4887;
wire TIMEBOOST_net_2275;
wire n_489;
wire n_4890;
wire n_4891;
wire n_4892;
wire n_4894;
wire n_4895;
wire n_4898;
wire n_49;
wire n_490;
wire n_4900;
wire n_4901;
wire TIMEBOOST_net_418;
wire n_4904;
wire n_4905;
wire n_4906;
wire n_4907;
wire n_4908;
wire n_491;
wire n_4910;
wire n_4911;
wire n_4912;
wire TIMEBOOST_net_2911;
wire TIMEBOOST_net_560;
wire n_4915;
wire n_4916;
wire n_4917;
wire n_4918;
wire n_4919;
wire n_492;
wire n_4920;
wire n_4921;
wire n_4922;
wire n_4923;
wire n_4925;
wire n_4927;
wire n_4928;
wire n_4929;
wire n_493;
wire n_4930;
wire n_4931;
wire n_4932;
wire n_4933;
wire n_4935;
wire n_4936;
wire TIMEBOOST_net_2282;
wire n_4938;
wire n_4939;
wire n_4940;
wire n_4941;
wire n_4942;
wire TIMEBOOST_net_1786;
wire n_4946;
wire TIMEBOOST_net_2474;
wire n_4948;
wire n_4949;
wire n_495;
wire n_4950;
wire n_4951;
wire TIMEBOOST_net_1237;
wire n_4953;
wire n_4954;
wire n_4956;
wire n_4957;
wire n_4958;
wire n_4959;
wire n_496;
wire n_4962;
wire n_4963;
wire n_4964;
wire n_4965;
wire n_4966;
wire n_4968;
wire n_4969;
wire n_497;
wire n_4970;
wire n_4972;
wire n_4973;
wire n_4974;
wire n_4975;
wire n_4976;
wire n_4978;
wire n_4979;
wire n_498;
wire n_4980;
wire n_4981;
wire n_4986;
wire n_4987;
wire n_4989;
wire n_499;
wire n_4990;
wire TIMEBOOST_net_2287;
wire n_4992;
wire n_4994;
wire n_4995;
wire n_4997;
wire n_4998;
wire n_4999;
wire n_50;
wire n_5000;
wire n_5001;
wire n_5002;
wire n_5003;
wire n_5005;
wire n_5006;
wire n_5009;
wire n_501;
wire TIMEBOOST_net_1283;
wire n_5011;
wire n_5012;
wire n_5013;
wire n_5015;
wire n_5016;
wire n_5017;
wire n_5018;
wire n_5020;
wire n_5021;
wire n_5023;
wire n_5024;
wire n_5025;
wire n_5026;
wire n_5028;
wire n_5030;
wire n_5031;
wire n_5032;
wire n_5035;
wire n_5036;
wire n_504;
wire n_5041;
wire n_5045;
wire TIMEBOOST_net_2676;
wire n_5048;
wire n_5049;
wire n_505;
wire n_5050;
wire n_5051;
wire n_5052;
wire n_5053;
wire n_5054;
wire n_5055;
wire n_5056;
wire n_5057;
wire n_5058;
wire n_5059;
wire n_506;
wire n_5060;
wire n_5061;
wire n_5062;
wire n_5063;
wire n_5064;
wire n_5065;
wire n_5066;
wire n_5067;
wire n_5069;
wire TIMEBOOST_net_2505;
wire n_5071;
wire n_5072;
wire n_5076;
wire n_5077;
wire TIMEBOOST_net_544;
wire n_5079;
wire n_508;
wire n_5080;
wire n_5081;
wire n_5082;
wire n_5083;
wire n_5084;
wire n_5085;
wire n_5087;
wire TIMEBOOST_net_1712;
wire n_509;
wire n_5090;
wire n_5091;
wire TIMEBOOST_net_2762;
wire n_5093;
wire n_5094;
wire n_5095;
wire n_5096;
wire TIMEBOOST_net_2459;
wire n_5098;
wire n_5099;
wire n_51;
wire n_510;
wire n_5101;
wire TIMEBOOST_net_2766;
wire n_5104;
wire n_5105;
wire n_5106;
wire n_5107;
wire n_5108;
wire n_5109;
wire n_511;
wire n_5110;
wire n_5111;
wire n_5112;
wire n_5113;
wire n_5114;
wire n_5115;
wire n_5116;
wire n_5117;
wire n_5121;
wire n_5123;
wire n_5125;
wire n_5127;
wire n_5128;
wire n_5129;
wire n_513;
wire n_5130;
wire n_5131;
wire n_5132;
wire n_5134;
wire n_5136;
wire n_5137;
wire n_5138;
wire n_5139;
wire n_514;
wire n_5140;
wire n_5141;
wire n_5142;
wire n_5143;
wire n_5144;
wire n_5145;
wire n_5146;
wire n_5147;
wire TIMEBOOST_net_1667;
wire n_5149;
wire n_515;
wire n_5150;
wire n_5151;
wire n_5152;
wire n_5153;
wire n_5154;
wire n_5156;
wire n_5157;
wire n_5158;
wire n_5159;
wire n_516;
wire n_5160;
wire n_5161;
wire n_5163;
wire TIMEBOOST_net_2949;
wire n_5165;
wire n_5166;
wire n_5168;
wire n_5169;
wire n_5170;
wire n_5171;
wire n_5172;
wire TIMEBOOST_net_1231;
wire n_5174;
wire n_5175;
wire n_5176;
wire n_5177;
wire n_5178;
wire n_518;
wire n_5181;
wire n_5184;
wire n_5185;
wire n_5186;
wire n_5187;
wire n_5188;
wire n_5189;
wire n_519;
wire TIMEBOOST_net_1716;
wire n_5191;
wire n_5192;
wire n_5193;
wire n_5194;
wire n_5195;
wire n_5196;
wire n_5197;
wire n_5198;
wire n_5199;
wire n_52;
wire n_520;
wire n_5200;
wire n_5203;
wire n_5204;
wire n_5206;
wire n_5207;
wire n_5208;
wire n_5209;
wire n_521;
wire n_5210;
wire n_5211;
wire n_5212;
wire n_5213;
wire n_5215;
wire n_5216;
wire n_5217;
wire n_5218;
wire n_522;
wire n_5221;
wire n_5224;
wire n_5225;
wire n_5226;
wire n_5227;
wire n_5228;
wire n_5229;
wire n_523;
wire n_5230;
wire n_5231;
wire n_5232;
wire n_5233;
wire n_5234;
wire n_5235;
wire n_5236;
wire n_524;
wire n_5240;
wire n_5241;
wire n_5242;
wire n_5243;
wire n_5244;
wire n_5247;
wire n_5248;
wire n_5249;
wire n_5250;
wire n_5251;
wire n_5253;
wire n_5255;
wire TIMEBOOST_net_1243;
wire n_5258;
wire n_5259;
wire TIMEBOOST_net_2186;
wire n_5260;
wire n_5261;
wire n_5262;
wire n_5263;
wire n_5265;
wire n_5266;
wire n_5267;
wire n_527;
wire n_5272;
wire n_5273;
wire n_5274;
wire n_5275;
wire n_5276;
wire n_5277;
wire n_5279;
wire n_528;
wire n_5280;
wire n_5283;
wire n_5284;
wire n_5285;
wire n_5286;
wire n_5287;
wire n_5288;
wire n_5289;
wire n_529;
wire n_5290;
wire n_5291;
wire TIMEBOOST_net_2153;
wire n_5294;
wire n_5295;
wire n_5297;
wire n_5298;
wire n_5299;
wire n_53;
wire n_530;
wire n_5300;
wire n_5301;
wire n_5304;
wire n_5305;
wire TIMEBOOST_net_1710;
wire n_5307;
wire n_5308;
wire n_531;
wire n_5310;
wire n_5312;
wire n_5313;
wire n_5314;
wire n_5315;
wire n_5316;
wire TIMEBOOST_net_564;
wire TIMEBOOST_net_565;
wire TIMEBOOST_net_1511;
wire n_5320;
wire n_5321;
wire n_5322;
wire n_5323;
wire n_5324;
wire n_5325;
wire n_5328;
wire n_5329;
wire n_533;
wire n_5330;
wire n_5331;
wire n_5332;
wire n_5333;
wire n_5334;
wire n_5335;
wire n_5336;
wire n_5339;
wire n_534;
wire n_5340;
wire n_5341;
wire n_5342;
wire n_5343;
wire n_5344;
wire n_5345;
wire n_5346;
wire n_5348;
wire n_5349;
wire n_535;
wire n_5350;
wire n_5351;
wire TIMEBOOST_net_1719;
wire n_5353;
wire TIMEBOOST_net_2763;
wire n_5355;
wire n_5356;
wire n_5357;
wire n_5358;
wire n_5359;
wire n_536;
wire n_5361;
wire n_5362;
wire n_5363;
wire n_5364;
wire n_5365;
wire n_5367;
wire n_5368;
wire TIMEBOOST_net_1261;
wire n_5371;
wire n_5372;
wire n_5373;
wire n_5374;
wire n_5375;
wire n_5377;
wire n_5378;
wire n_5379;
wire n_5380;
wire n_5381;
wire n_5382;
wire n_5384;
wire n_5385;
wire n_5386;
wire n_5387;
wire TIMEBOOST_net_2054;
wire n_5389;
wire n_539;
wire n_5393;
wire n_5394;
wire n_5395;
wire n_5397;
wire n_5399;
wire n_54;
wire n_540;
wire n_5400;
wire n_5402;
wire n_5403;
wire n_5404;
wire n_5405;
wire n_5406;
wire TIMEBOOST_net_2067;
wire n_5408;
wire n_5409;
wire n_541;
wire n_5410;
wire n_5411;
wire n_5412;
wire n_5413;
wire n_5414;
wire n_5415;
wire n_5416;
wire n_5417;
wire n_5418;
wire n_542;
wire n_5420;
wire n_5421;
wire n_5422;
wire n_5423;
wire n_5424;
wire n_5425;
wire n_5426;
wire n_5428;
wire n_5429;
wire n_543;
wire n_5430;
wire n_5431;
wire n_5432;
wire n_5433;
wire n_5434;
wire TIMEBOOST_net_551;
wire n_5436;
wire n_5437;
wire n_5439;
wire n_544;
wire n_5440;
wire n_5441;
wire n_5442;
wire n_5443;
wire n_5444;
wire n_5446;
wire n_5447;
wire TIMEBOOST_net_2946;
wire n_545;
wire n_5450;
wire n_5451;
wire n_5452;
wire n_5454;
wire n_5455;
wire n_5456;
wire n_5457;
wire n_5458;
wire n_5459;
wire n_546;
wire n_5460;
wire n_5461;
wire n_5462;
wire n_5463;
wire n_5464;
wire n_5465;
wire n_5468;
wire n_547;
wire n_5471;
wire n_5472;
wire n_5473;
wire n_5475;
wire n_5476;
wire n_5477;
wire n_5478;
wire n_548;
wire n_5480;
wire n_5481;
wire n_5482;
wire n_5483;
wire n_5484;
wire n_5485;
wire n_5486;
wire n_5487;
wire n_5488;
wire n_5489;
wire n_549;
wire n_5490;
wire n_5491;
wire n_5493;
wire n_5494;
wire n_5495;
wire n_5496;
wire n_5497;
wire n_5498;
wire n_5499;
wire n_55;
wire n_550;
wire n_5500;
wire n_5501;
wire n_5502;
wire n_5503;
wire n_5504;
wire n_5505;
wire n_5506;
wire n_5508;
wire n_5509;
wire n_5510;
wire n_5511;
wire n_5512;
wire n_5516;
wire n_5517;
wire n_5518;
wire n_5520;
wire n_5521;
wire TIMEBOOST_net_1260;
wire n_5523;
wire n_5524;
wire n_5526;
wire n_5527;
wire n_5528;
wire n_5529;
wire n_553;
wire n_5530;
wire n_5531;
wire n_5532;
wire n_5534;
wire n_5535;
wire TIMEBOOST_net_2930;
wire n_5538;
wire n_5539;
wire n_554;
wire n_5540;
wire n_5541;
wire n_5543;
wire TIMEBOOST_net_1262;
wire n_5545;
wire n_5546;
wire n_5547;
wire n_5548;
wire n_5549;
wire n_5550;
wire n_5551;
wire n_5552;
wire n_5553;
wire n_5554;
wire n_5555;
wire n_5556;
wire n_5557;
wire n_5558;
wire n_5559;
wire n_556;
wire n_5561;
wire n_5562;
wire n_5563;
wire n_5564;
wire n_5565;
wire n_5566;
wire n_5567;
wire n_5568;
wire n_5569;
wire n_557;
wire TIMEBOOST_net_556;
wire n_5571;
wire n_5572;
wire TIMEBOOST_net_2921;
wire TIMEBOOST_net_520;
wire TIMEBOOST_net_1762;
wire n_5577;
wire n_5578;
wire n_5579;
wire n_558;
wire n_5580;
wire n_5581;
wire n_5582;
wire n_5583;
wire n_5584;
wire n_5586;
wire n_5587;
wire n_5589;
wire n_559;
wire n_5590;
wire TIMEBOOST_net_2919;
wire n_5592;
wire n_5593;
wire n_5594;
wire n_5595;
wire n_5596;
wire n_5598;
wire n_5599;
wire n_56;
wire n_560;
wire TIMEBOOST_net_1784;
wire n_5601;
wire n_5603;
wire n_5605;
wire n_5606;
wire n_5607;
wire n_5608;
wire n_5609;
wire n_561;
wire n_5610;
wire n_5611;
wire n_5612;
wire n_5613;
wire n_5614;
wire n_5616;
wire n_5617;
wire n_5618;
wire n_5619;
wire n_5620;
wire n_5621;
wire n_5622;
wire n_5624;
wire n_5626;
wire n_5627;
wire n_5628;
wire n_5629;
wire n_563;
wire n_5632;
wire TIMEBOOST_net_1761;
wire n_5636;
wire n_5637;
wire n_5638;
wire n_5639;
wire n_564;
wire n_5641;
wire n_5642;
wire n_5644;
wire n_5645;
wire n_5648;
wire n_565;
wire n_5650;
wire n_5651;
wire TIMEBOOST_net_2235;
wire n_5654;
wire n_5655;
wire n_5656;
wire n_5657;
wire n_5658;
wire n_5659;
wire n_566;
wire n_5660;
wire n_5661;
wire n_5662;
wire n_5663;
wire n_5664;
wire n_5665;
wire n_5666;
wire n_5667;
wire TIMEBOOST_net_1267;
wire n_5669;
wire n_567;
wire TIMEBOOST_net_2043;
wire n_5671;
wire n_5672;
wire n_5673;
wire n_5674;
wire n_5675;
wire n_5676;
wire n_5677;
wire n_5679;
wire n_568;
wire n_5680;
wire n_5681;
wire n_5684;
wire n_5685;
wire n_5688;
wire n_5689;
wire n_569;
wire n_5690;
wire n_5691;
wire n_5692;
wire n_5693;
wire n_5695;
wire n_5696;
wire n_5697;
wire n_5698;
wire n_57;
wire n_570;
wire n_5700;
wire n_5701;
wire n_5702;
wire n_5703;
wire n_5706;
wire n_5707;
wire n_5708;
wire n_5709;
wire n_571;
wire n_5710;
wire n_5711;
wire n_5712;
wire TIMEBOOST_net_2940;
wire n_5714;
wire n_5716;
wire n_5717;
wire n_5718;
wire n_5719;
wire n_572;
wire n_5720;
wire n_5721;
wire n_5723;
wire n_5724;
wire n_5725;
wire n_5726;
wire n_5727;
wire n_5728;
wire n_5730;
wire TIMEBOOST_net_1272;
wire n_5732;
wire TIMEBOOST_net_501;
wire n_5735;
wire n_5736;
wire n_5739;
wire n_5740;
wire n_5741;
wire n_5742;
wire n_5743;
wire n_5746;
wire n_5748;
wire n_5750;
wire n_5751;
wire n_5753;
wire n_5754;
wire n_5755;
wire n_5756;
wire n_5757;
wire n_5759;
wire n_576;
wire TIMEBOOST_net_1300;
wire n_5761;
wire n_5763;
wire n_5765;
wire n_5766;
wire n_5767;
wire n_5768;
wire n_5769;
wire n_5770;
wire n_5771;
wire TIMEBOOST_net_1801;
wire n_5773;
wire n_5774;
wire n_5775;
wire n_5776;
wire n_5777;
wire n_5778;
wire n_5779;
wire n_578;
wire n_5780;
wire n_5782;
wire n_5783;
wire n_5784;
wire n_5785;
wire n_5786;
wire n_5787;
wire n_5788;
wire n_5789;
wire n_579;
wire n_5791;
wire n_5792;
wire n_5793;
wire n_5795;
wire n_5796;
wire n_5797;
wire n_5798;
wire TIMEBOOST_net_2318;
wire n_58;
wire n_580;
wire n_5800;
wire n_5801;
wire n_5802;
wire n_5805;
wire n_5806;
wire n_5807;
wire n_5808;
wire n_581;
wire n_5810;
wire n_5811;
wire n_5812;
wire n_5813;
wire n_5814;
wire n_5815;
wire n_5816;
wire n_5818;
wire TIMEBOOST_net_588;
wire n_582;
wire n_5820;
wire n_5821;
wire n_5823;
wire n_5824;
wire n_5825;
wire TIMEBOOST_net_658;
wire n_5830;
wire TIMEBOOST_net_528;
wire n_5832;
wire n_5833;
wire TIMEBOOST_net_653;
wire n_5835;
wire n_5836;
wire n_5837;
wire n_5838;
wire n_5839;
wire n_584;
wire n_5840;
wire n_5841;
wire n_5842;
wire n_5844;
wire n_5845;
wire n_5852;
wire n_5853;
wire TIMEBOOST_net_664;
wire n_5857;
wire n_5858;
wire n_5859;
wire n_5860;
wire n_5861;
wire n_5862;
wire n_5863;
wire n_5864;
wire n_5866;
wire n_5867;
wire n_5868;
wire n_587;
wire n_5870;
wire n_5871;
wire n_5873;
wire n_5874;
wire n_5875;
wire n_5876;
wire n_5877;
wire n_5878;
wire n_5879;
wire n_588;
wire n_5880;
wire n_5881;
wire n_5882;
wire n_5883;
wire n_5884;
wire TIMEBOOST_net_2768;
wire n_5886;
wire n_5887;
wire n_5888;
wire n_5889;
wire n_589;
wire n_5893;
wire n_5894;
wire n_5895;
wire n_5896;
wire n_5897;
wire n_5898;
wire n_5899;
wire n_59;
wire n_590;
wire n_5900;
wire n_5901;
wire n_5902;
wire n_5904;
wire n_5905;
wire n_5906;
wire n_5907;
wire n_5909;
wire n_591;
wire n_5910;
wire n_5911;
wire n_5913;
wire TIMEBOOST_net_656;
wire n_5915;
wire n_5916;
wire n_5917;
wire n_5918;
wire n_5919;
wire TIMEBOOST_net_561;
wire n_5921;
wire n_5922;
wire n_5923;
wire n_5924;
wire n_5925;
wire n_5926;
wire n_5927;
wire n_5928;
wire n_5929;
wire n_593;
wire n_5930;
wire n_5933;
wire n_5935;
wire n_5937;
wire n_5938;
wire n_5939;
wire n_594;
wire n_5940;
wire n_5941;
wire n_5943;
wire n_5944;
wire TIMEBOOST_net_480;
wire n_5946;
wire n_5947;
wire n_5948;
wire n_5949;
wire n_595;
wire n_5950;
wire n_5951;
wire n_5952;
wire n_5953;
wire n_5955;
wire n_5957;
wire n_5958;
wire n_5959;
wire n_596;
wire n_5961;
wire n_5962;
wire n_5963;
wire n_5964;
wire n_5965;
wire n_5966;
wire n_5967;
wire n_5968;
wire n_5969;
wire n_597;
wire n_5970;
wire n_5971;
wire n_5972;
wire TIMEBOOST_net_530;
wire n_5974;
wire n_5976;
wire n_5977;
wire TIMEBOOST_net_639;
wire n_5979;
wire n_598;
wire n_5980;
wire n_5981;
wire n_5982;
wire n_5983;
wire n_5984;
wire n_5986;
wire n_5987;
wire n_5989;
wire n_599;
wire n_5990;
wire n_5991;
wire n_5992;
wire n_5994;
wire TIMEBOOST_net_2458;
wire n_5996;
wire n_5997;
wire n_5998;
wire n_5999;
wire n_60;
wire n_600;
wire n_6001;
wire n_6002;
wire n_6003;
wire n_6004;
wire n_6005;
wire n_6006;
wire n_6007;
wire n_6008;
wire n_6009;
wire n_601;
wire n_6010;
wire n_6011;
wire n_6012;
wire n_6013;
wire TIMEBOOST_net_671;
wire n_6015;
wire n_6017;
wire n_6019;
wire n_602;
wire n_6020;
wire n_6021;
wire n_6023;
wire n_6024;
wire n_6025;
wire n_6026;
wire n_6028;
wire n_603;
wire n_6032;
wire n_6033;
wire n_6034;
wire n_6036;
wire n_6037;
wire n_6038;
wire n_6039;
wire n_604;
wire n_6040;
wire n_6041;
wire n_6042;
wire n_6043;
wire n_6044;
wire n_6047;
wire n_6048;
wire TIMEBOOST_net_640;
wire n_605;
wire n_6051;
wire n_6052;
wire n_6053;
wire n_6054;
wire n_6055;
wire TIMEBOOST_net_663;
wire n_6059;
wire n_606;
wire n_6061;
wire n_6062;
wire n_6063;
wire n_6064;
wire n_6065;
wire n_6066;
wire n_6067;
wire n_6068;
wire n_6069;
wire n_607;
wire TIMEBOOST_net_492;
wire n_6071;
wire n_6074;
wire n_6076;
wire n_6077;
wire n_608;
wire n_6080;
wire n_6081;
wire n_6082;
wire n_6083;
wire TIMEBOOST_net_1796;
wire n_6085;
wire n_6086;
wire n_6087;
wire n_6089;
wire n_609;
wire n_6090;
wire n_6092;
wire n_6094;
wire n_6096;
wire n_6097;
wire n_6098;
wire n_61;
wire n_610;
wire n_6100;
wire n_6101;
wire n_6102;
wire TIMEBOOST_net_2719;
wire n_6104;
wire n_6105;
wire n_6106;
wire n_6107;
wire n_6108;
wire n_6109;
wire n_611;
wire n_6110;
wire TIMEBOOST_net_2752;
wire n_6112;
wire n_6113;
wire n_6114;
wire n_6115;
wire n_6116;
wire n_6117;
wire n_6118;
wire n_6119;
wire n_612;
wire n_6121;
wire n_6122;
wire n_6123;
wire n_6124;
wire n_6125;
wire n_6127;
wire n_6128;
wire TIMEBOOST_net_670;
wire n_613;
wire n_6130;
wire n_6132;
wire n_6133;
wire n_6135;
wire n_6136;
wire n_6137;
wire n_6138;
wire n_6139;
wire n_614;
wire n_6140;
wire n_6141;
wire n_6142;
wire n_6143;
wire n_6144;
wire n_6145;
wire n_6146;
wire n_6147;
wire n_6148;
wire n_6149;
wire n_615;
wire n_6150;
wire n_6151;
wire TIMEBOOST_net_2591;
wire n_6153;
wire n_6154;
wire TIMEBOOST_net_694;
wire n_6156;
wire n_6157;
wire n_6158;
wire n_6159;
wire n_616;
wire n_6160;
wire TIMEBOOST_net_496;
wire n_6162;
wire n_6163;
wire n_6165;
wire TIMEBOOST_net_1828;
wire n_6167;
wire TIMEBOOST_net_681;
wire n_6169;
wire n_617;
wire n_6170;
wire n_6171;
wire n_6172;
wire n_6173;
wire n_6175;
wire n_6176;
wire n_6177;
wire n_6178;
wire n_6179;
wire TIMEBOOST_net_853;
wire n_6180;
wire n_6181;
wire n_6182;
wire n_6183;
wire n_6184;
wire n_6185;
wire n_6186;
wire n_6187;
wire n_6188;
wire n_6189;
wire n_619;
wire n_6190;
wire n_6191;
wire n_6192;
wire TIMEBOOST_net_698;
wire n_6196;
wire n_6197;
wire n_6198;
wire n_62;
wire n_620;
wire n_6201;
wire TIMEBOOST_net_738;
wire n_6203;
wire n_6204;
wire n_6205;
wire n_6206;
wire n_6207;
wire n_6208;
wire n_6209;
wire n_621;
wire n_6210;
wire n_6212;
wire n_6213;
wire n_6214;
wire n_6215;
wire n_6217;
wire n_6218;
wire n_6219;
wire n_622;
wire n_6220;
wire n_6222;
wire n_6223;
wire n_6224;
wire n_6225;
wire n_6226;
wire n_6228;
wire n_6229;
wire n_623;
wire n_6230;
wire n_6231;
wire n_6233;
wire n_6234;
wire n_6235;
wire n_6237;
wire n_6238;
wire n_6239;
wire n_624;
wire n_6240;
wire n_6241;
wire n_6243;
wire n_6244;
wire n_6245;
wire n_6248;
wire n_625;
wire n_6250;
wire TIMEBOOST_net_1384;
wire n_6253;
wire n_6254;
wire n_6257;
wire n_6259;
wire n_626;
wire n_6260;
wire n_6261;
wire n_6262;
wire n_6263;
wire n_6265;
wire n_6266;
wire n_6267;
wire n_6268;
wire n_6269;
wire n_627;
wire n_6270;
wire TIMEBOOST_net_744;
wire n_6272;
wire n_6276;
wire n_6277;
wire n_6279;
wire n_628;
wire n_6280;
wire n_6281;
wire n_6282;
wire n_6285;
wire n_6286;
wire n_6287;
wire n_6288;
wire n_629;
wire n_6290;
wire n_6291;
wire TIMEBOOST_net_1372;
wire n_6294;
wire n_6295;
wire n_6297;
wire n_6298;
wire n_6299;
wire n_63;
wire n_630;
wire n_6301;
wire TIMEBOOST_net_708;
wire TIMEBOOST_net_750;
wire n_6304;
wire TIMEBOOST_net_1285;
wire n_6308;
wire n_6309;
wire n_631;
wire n_6310;
wire n_6311;
wire n_6312;
wire n_6313;
wire n_6315;
wire n_6316;
wire n_6317;
wire n_6318;
wire n_6319;
wire n_632;
wire n_6320;
wire n_6321;
wire n_6323;
wire n_6324;
wire n_6325;
wire n_6326;
wire n_6327;
wire n_6328;
wire n_6329;
wire n_633;
wire n_6330;
wire TIMEBOOST_net_574;
wire n_6332;
wire n_6334;
wire n_6335;
wire n_6338;
wire n_634;
wire n_6340;
wire n_6341;
wire n_6342;
wire n_6343;
wire TIMEBOOST_net_707;
wire n_6345;
wire n_6346;
wire n_6347;
wire n_6348;
wire TIMEBOOST_net_746;
wire n_635;
wire n_6350;
wire n_6351;
wire n_6352;
wire n_6353;
wire n_6354;
wire n_6355;
wire n_6356;
wire n_6357;
wire n_6358;
wire n_6359;
wire n_636;
wire n_6360;
wire n_6362;
wire n_6363;
wire TIMEBOOST_net_2074;
wire n_6365;
wire TIMEBOOST_net_2091;
wire n_6368;
wire n_6369;
wire n_637;
wire n_6370;
wire n_6371;
wire n_6373;
wire TIMEBOOST_net_2797;
wire TIMEBOOST_net_711;
wire n_6376;
wire n_6379;
wire n_638;
wire n_6380;
wire n_6382;
wire n_6383;
wire n_6384;
wire TIMEBOOST_net_2498;
wire n_6386;
wire n_6387;
wire n_6388;
wire n_6389;
wire n_639;
wire n_6390;
wire n_6391;
wire n_6392;
wire n_6393;
wire n_6394;
wire n_6395;
wire n_6396;
wire TIMEBOOST_net_1373;
wire n_6398;
wire n_6399;
wire n_64;
wire n_640;
wire n_6404;
wire n_6405;
wire n_6407;
wire n_6408;
wire n_6409;
wire n_641;
wire n_6412;
wire n_6413;
wire n_6414;
wire n_6415;
wire n_6416;
wire TIMEBOOST_net_2080;
wire n_6418;
wire n_6419;
wire n_642;
wire n_6425;
wire n_643;
wire n_6435;
wire n_6436;
wire n_6438;
wire n_644;
wire n_6442;
wire n_6443;
wire n_6447;
wire n_6448;
wire n_645;
wire n_6453;
wire n_6454;
wire n_6456;
wire n_646;
wire n_6463;
wire n_6465;
wire n_6466;
wire n_647;
wire n_6471;
wire n_6473;
wire n_6476;
wire n_6477;
wire n_6479;
wire n_648;
wire n_6485;
wire n_6486;
wire n_6487;
wire n_6488;
wire n_6489;
wire n_649;
wire n_6490;
wire n_6491;
wire n_6493;
wire n_6496;
wire n_6499;
wire n_65;
wire n_650;
wire n_6500;
wire n_6502;
wire n_6503;
wire n_6504;
wire n_6505;
wire n_6506;
wire n_6507;
wire n_6509;
wire n_651;
wire n_6510;
wire n_6512;
wire n_6513;
wire n_6517;
wire n_6519;
wire n_652;
wire n_6521;
wire n_6523;
wire n_6524;
wire n_6528;
wire n_6529;
wire n_653;
wire n_6531;
wire n_6535;
wire n_6539;
wire n_654;
wire n_6540;
wire n_6541;
wire n_6542;
wire TIMEBOOST_net_2416;
wire TIMEBOOST_net_2164;
wire n_6546;
wire n_6547;
wire n_655;
wire TIMEBOOST_net_1421;
wire n_6551;
wire n_6552;
wire n_6554;
wire n_6555;
wire n_6556;
wire n_6557;
wire n_6558;
wire n_656;
wire n_6560;
wire n_6561;
wire n_6562;
wire n_6563;
wire n_6564;
wire n_6565;
wire n_6567;
wire n_6569;
wire n_657;
wire n_6570;
wire n_6571;
wire n_6572;
wire n_6574;
wire n_6576;
wire n_6577;
wire n_6578;
wire n_6579;
wire n_658;
wire n_6580;
wire n_6581;
wire n_6582;
wire n_6583;
wire n_6585;
wire n_6586;
wire n_6587;
wire n_6589;
wire n_659;
wire n_6590;
wire n_6591;
wire n_6592;
wire n_6593;
wire n_6594;
wire n_6595;
wire n_6596;
wire n_6597;
wire n_6598;
wire n_6599;
wire n_66;
wire n_660;
wire n_6600;
wire n_6601;
wire n_6607;
wire n_6609;
wire n_661;
wire n_6610;
wire n_6612;
wire n_6613;
wire n_6616;
wire n_6617;
wire n_6618;
wire n_6619;
wire n_662;
wire n_6620;
wire n_6621;
wire n_6624;
wire n_6625;
wire n_6626;
wire n_6627;
wire n_6628;
wire n_663;
wire n_6630;
wire n_6631;
wire n_6633;
wire n_6634;
wire n_6635;
wire n_6637;
wire n_6638;
wire n_6639;
wire n_664;
wire n_6640;
wire n_6641;
wire n_6642;
wire n_6643;
wire n_6644;
wire n_6645;
wire n_6646;
wire n_6648;
wire n_6649;
wire n_665;
wire n_6651;
wire n_6652;
wire n_6653;
wire n_6654;
wire n_6655;
wire n_6656;
wire n_6658;
wire n_666;
wire n_6660;
wire n_6661;
wire n_6664;
wire n_6665;
wire n_6666;
wire n_6667;
wire n_6668;
wire n_6669;
wire n_667;
wire n_6670;
wire n_6671;
wire n_6672;
wire n_6673;
wire n_6674;
wire n_6675;
wire n_6676;
wire n_6679;
wire n_6680;
wire n_6681;
wire n_6683;
wire n_6684;
wire n_6687;
wire n_6688;
wire n_6689;
wire n_669;
wire n_6690;
wire n_6695;
wire n_6696;
wire n_6697;
wire n_6698;
wire n_67;
wire n_670;
wire n_6700;
wire n_6701;
wire n_6703;
wire n_6704;
wire n_6705;
wire n_6706;
wire n_6707;
wire n_6708;
wire n_671;
wire n_6710;
wire n_6711;
wire n_6715;
wire n_6716;
wire n_6717;
wire n_6718;
wire n_6719;
wire n_672;
wire n_6720;
wire n_6721;
wire n_6722;
wire n_6723;
wire n_6724;
wire n_6725;
wire n_6729;
wire TIMEBOOST_net_200;
wire n_6730;
wire n_6731;
wire n_6732;
wire n_6733;
wire n_6734;
wire n_6737;
wire n_6739;
wire n_674;
wire n_6741;
wire n_6742;
wire n_6743;
wire n_6745;
wire n_6746;
wire n_6747;
wire n_6748;
wire n_6749;
wire n_675;
wire n_6752;
wire n_6753;
wire n_6754;
wire n_6755;
wire n_6756;
wire n_6758;
wire n_6759;
wire n_676;
wire n_6760;
wire n_6761;
wire n_6762;
wire n_6763;
wire n_6764;
wire n_6765;
wire n_6767;
wire n_6769;
wire n_677;
wire n_6770;
wire n_6771;
wire n_6772;
wire n_6773;
wire n_6774;
wire n_6775;
wire n_6776;
wire TIMEBOOST_net_2728;
wire n_678;
wire n_6780;
wire n_6782;
wire n_6783;
wire n_6784;
wire n_6789;
wire n_679;
wire n_6790;
wire TIMEBOOST_net_790;
wire n_6798;
wire n_68;
wire TIMEBOOST_net_1418;
wire n_6801;
wire n_6802;
wire n_6803;
wire n_6804;
wire n_6806;
wire n_6809;
wire n_6813;
wire n_6815;
wire n_6816;
wire n_6817;
wire n_6818;
wire n_6819;
wire n_682;
wire n_6822;
wire n_6824;
wire n_6825;
wire n_6826;
wire n_6828;
wire n_6829;
wire n_6830;
wire n_6831;
wire n_6832;
wire n_6833;
wire n_6834;
wire n_6835;
wire n_6836;
wire n_684;
wire TIMEBOOST_net_1468;
wire TIMEBOOST_net_2339;
wire n_6842;
wire n_6843;
wire n_6844;
wire n_6845;
wire n_6847;
wire n_6848;
wire n_6849;
wire n_685;
wire n_6850;
wire n_6851;
wire n_6852;
wire n_6853;
wire n_6854;
wire n_6855;
wire n_6856;
wire n_6857;
wire n_6858;
wire n_6859;
wire n_686;
wire n_6860;
wire n_6861;
wire n_6862;
wire n_6863;
wire n_6864;
wire n_6865;
wire n_6866;
wire n_6867;
wire n_6868;
wire n_6869;
wire n_687;
wire n_6870;
wire n_6871;
wire n_6872;
wire n_6873;
wire n_6874;
wire n_6875;
wire n_6876;
wire n_6877;
wire n_6878;
wire n_6879;
wire n_688;
wire n_6880;
wire n_6881;
wire n_6882;
wire n_6883;
wire n_6884;
wire n_6885;
wire n_6887;
wire n_6889;
wire n_689;
wire n_6890;
wire n_6891;
wire n_6892;
wire n_6893;
wire n_6895;
wire n_6896;
wire n_6897;
wire n_6898;
wire n_6899;
wire n_69;
wire n_690;
wire n_6900;
wire n_6901;
wire n_6903;
wire n_6904;
wire n_6907;
wire n_6908;
wire n_6909;
wire n_691;
wire n_6910;
wire TIMEBOOST_net_1476;
wire n_6914;
wire n_6915;
wire n_6916;
wire n_6918;
wire n_6919;
wire n_692;
wire n_6920;
wire n_6921;
wire n_6922;
wire n_6923;
wire n_6924;
wire n_6925;
wire n_6926;
wire n_6927;
wire n_6928;
wire n_6929;
wire n_693;
wire n_6930;
wire n_6931;
wire n_6932;
wire TIMEBOOST_net_2201;
wire n_6934;
wire n_6935;
wire n_6936;
wire n_6937;
wire n_6938;
wire n_6939;
wire n_694;
wire n_6940;
wire n_6941;
wire n_6942;
wire n_6943;
wire n_6944;
wire n_6945;
wire n_6946;
wire n_6947;
wire n_6948;
wire n_6949;
wire n_695;
wire n_6950;
wire n_6951;
wire n_6952;
wire n_6953;
wire n_6956;
wire n_6957;
wire n_6958;
wire n_6959;
wire n_6960;
wire n_6961;
wire n_6962;
wire n_6963;
wire n_6964;
wire n_6965;
wire n_6966;
wire n_6967;
wire n_6968;
wire n_6969;
wire n_697;
wire n_6970;
wire n_6971;
wire n_6973;
wire n_6974;
wire n_6975;
wire n_6976;
wire n_6977;
wire n_6979;
wire n_698;
wire n_6980;
wire n_6981;
wire n_6984;
wire n_6985;
wire n_6986;
wire n_6987;
wire n_6988;
wire n_6989;
wire n_6990;
wire n_6991;
wire n_6992;
wire n_6993;
wire n_6994;
wire n_6995;
wire n_6996;
wire n_6997;
wire n_6998;
wire n_6999;
wire n_7;
wire n_70;
wire n_700;
wire n_7000;
wire n_7002;
wire n_7003;
wire n_7004;
wire n_7006;
wire n_7007;
wire n_7008;
wire n_7009;
wire n_701;
wire n_7010;
wire n_7011;
wire n_7012;
wire n_7013;
wire n_7014;
wire n_7015;
wire n_7016;
wire n_7017;
wire n_7020;
wire n_7021;
wire n_7022;
wire n_7023;
wire n_7024;
wire n_7025;
wire n_7026;
wire n_7027;
wire n_7028;
wire n_7029;
wire n_703;
wire n_7030;
wire n_7031;
wire n_7033;
wire n_7034;
wire n_7035;
wire n_7036;
wire n_7037;
wire n_704;
wire n_7040;
wire n_7041;
wire n_7042;
wire n_7043;
wire n_7044;
wire n_7045;
wire n_7046;
wire n_7048;
wire n_7049;
wire n_705;
wire n_7050;
wire n_7051;
wire n_7052;
wire n_7053;
wire n_7054;
wire n_7055;
wire n_7056;
wire n_7057;
wire n_7058;
wire n_7059;
wire n_706;
wire n_7060;
wire TIMEBOOST_net_867;
wire n_7062;
wire n_7063;
wire n_7064;
wire n_7065;
wire n_7066;
wire n_7067;
wire n_7068;
wire n_7069;
wire n_707;
wire n_7070;
wire n_7071;
wire n_7072;
wire n_7073;
wire n_7077;
wire n_7078;
wire n_7079;
wire n_708;
wire n_7080;
wire n_7081;
wire n_7082;
wire n_7083;
wire n_7084;
wire n_7085;
wire n_7086;
wire n_7087;
wire n_7088;
wire n_7089;
wire n_709;
wire n_7090;
wire n_7091;
wire n_7092;
wire n_7093;
wire n_7094;
wire n_7095;
wire n_7097;
wire n_7098;
wire n_7099;
wire n_71;
wire n_710;
wire n_7100;
wire n_7101;
wire n_7102;
wire n_7103;
wire n_7105;
wire n_7106;
wire n_7107;
wire n_7108;
wire n_7109;
wire n_711;
wire n_7110;
wire n_7111;
wire n_7112;
wire n_7113;
wire n_7114;
wire n_7116;
wire n_7117;
wire n_7118;
wire n_7119;
wire n_712;
wire n_7120;
wire n_7121;
wire n_7122;
wire n_7123;
wire n_7124;
wire TIMEBOOST_net_878;
wire n_7126;
wire n_7127;
wire n_7128;
wire n_7129;
wire n_713;
wire n_7131;
wire n_7132;
wire n_7134;
wire n_7135;
wire n_7136;
wire n_7137;
wire n_7138;
wire n_7139;
wire n_714;
wire n_7141;
wire n_7143;
wire n_7144;
wire TIMEBOOST_net_1490;
wire n_7146;
wire n_7147;
wire n_715;
wire n_7150;
wire n_7153;
wire n_7154;
wire n_7155;
wire n_7156;
wire n_7157;
wire n_7158;
wire n_7159;
wire n_716;
wire n_7160;
wire n_7161;
wire n_7162;
wire n_7163;
wire n_7164;
wire n_7165;
wire n_7166;
wire n_7167;
wire n_7168;
wire n_7169;
wire n_717;
wire n_7170;
wire n_7171;
wire n_7172;
wire n_7173;
wire n_7177;
wire n_7178;
wire n_7179;
wire n_718;
wire n_7180;
wire n_7181;
wire n_7182;
wire TIMEBOOST_net_884;
wire n_7187;
wire n_7188;
wire n_7189;
wire n_719;
wire n_7190;
wire n_7191;
wire n_7193;
wire n_7194;
wire n_7195;
wire n_7196;
wire n_7197;
wire n_7198;
wire n_7199;
wire n_72;
wire TIMEBOOST_net_901;
wire n_7201;
wire n_7202;
wire n_7203;
wire n_7204;
wire n_7206;
wire n_7207;
wire n_7208;
wire n_7209;
wire n_7210;
wire n_7211;
wire n_7212;
wire n_7215;
wire n_7217;
wire n_7218;
wire n_7219;
wire n_7221;
wire n_7222;
wire n_7223;
wire n_7224;
wire n_7225;
wire n_7226;
wire n_7227;
wire n_7228;
wire n_7229;
wire n_7230;
wire n_7231;
wire TIMEBOOST_net_881;
wire n_7233;
wire n_7234;
wire n_7235;
wire n_7236;
wire n_7237;
wire n_7238;
wire n_7239;
wire n_724;
wire n_7240;
wire n_7241;
wire n_7242;
wire n_7243;
wire n_7244;
wire n_7245;
wire n_7246;
wire n_7247;
wire n_725;
wire n_7250;
wire n_7251;
wire n_7252;
wire n_7254;
wire n_7255;
wire n_7256;
wire n_7257;
wire n_7258;
wire n_726;
wire n_7260;
wire n_7261;
wire n_7262;
wire n_7263;
wire n_7264;
wire n_7265;
wire n_7266;
wire n_7267;
wire n_7268;
wire n_7269;
wire n_727;
wire n_7270;
wire n_7271;
wire n_7272;
wire n_7273;
wire n_7276;
wire n_7277;
wire n_7278;
wire n_7279;
wire n_7280;
wire n_7281;
wire n_7282;
wire n_7283;
wire n_7284;
wire n_7285;
wire n_7286;
wire n_7287;
wire n_7288;
wire n_7289;
wire n_729;
wire n_7290;
wire n_7291;
wire n_7292;
wire n_7294;
wire n_7295;
wire n_7296;
wire n_7297;
wire n_7298;
wire n_7299;
wire n_73;
wire n_730;
wire n_7300;
wire n_7301;
wire n_7302;
wire n_7303;
wire n_7304;
wire n_7305;
wire n_7306;
wire n_7307;
wire n_7308;
wire n_7309;
wire n_731;
wire n_7310;
wire n_7311;
wire n_7313;
wire n_7314;
wire n_7315;
wire n_7316;
wire n_7317;
wire n_7318;
wire n_732;
wire n_7320;
wire n_7321;
wire n_7322;
wire n_7323;
wire n_7324;
wire n_7326;
wire n_7327;
wire n_7328;
wire n_7329;
wire n_733;
wire n_7330;
wire n_7331;
wire n_7332;
wire n_7333;
wire n_7334;
wire n_7335;
wire n_7337;
wire n_7338;
wire n_734;
wire n_7341;
wire n_7342;
wire n_7343;
wire n_7344;
wire n_7345;
wire n_7346;
wire n_7347;
wire n_7348;
wire n_7349;
wire n_7351;
wire n_7352;
wire n_7353;
wire n_7354;
wire n_7355;
wire n_7356;
wire n_7357;
wire n_7358;
wire n_7359;
wire n_736;
wire n_7360;
wire n_7361;
wire n_7362;
wire n_7363;
wire n_7364;
wire n_7365;
wire n_7366;
wire n_7368;
wire n_7369;
wire TIMEBOOST_net_893;
wire n_7371;
wire n_7372;
wire n_7373;
wire n_7374;
wire n_7375;
wire n_7376;
wire n_7377;
wire n_7378;
wire n_7379;
wire n_738;
wire n_7380;
wire n_7381;
wire n_7382;
wire TIMEBOOST_net_2012;
wire n_7384;
wire n_7385;
wire n_7386;
wire n_7387;
wire n_7388;
wire n_7389;
wire n_739;
wire n_7392;
wire n_7393;
wire n_7394;
wire n_7395;
wire n_7396;
wire n_7399;
wire n_74;
wire n_740;
wire n_7400;
wire n_7401;
wire n_7402;
wire n_7403;
wire n_7404;
wire n_7405;
wire n_7406;
wire n_7407;
wire n_7408;
wire n_7409;
wire n_7410;
wire n_7411;
wire n_7412;
wire n_7413;
wire n_7414;
wire n_7415;
wire n_7416;
wire n_7417;
wire n_7418;
wire n_7419;
wire n_742;
wire n_7420;
wire n_7421;
wire n_7422;
wire n_7423;
wire n_7424;
wire n_7425;
wire n_7426;
wire n_7427;
wire n_7428;
wire n_7429;
wire n_743;
wire n_7430;
wire n_7431;
wire n_7432;
wire n_7434;
wire n_7435;
wire n_7436;
wire n_7437;
wire n_7438;
wire n_7439;
wire n_744;
wire n_7440;
wire n_7441;
wire n_7442;
wire n_7443;
wire n_7444;
wire n_7445;
wire n_7446;
wire n_7447;
wire n_7448;
wire n_7449;
wire n_745;
wire n_7450;
wire n_7451;
wire n_7452;
wire n_7453;
wire n_7455;
wire n_7456;
wire n_7457;
wire n_7458;
wire n_746;
wire n_7460;
wire n_7461;
wire n_7462;
wire n_7464;
wire n_7465;
wire n_7466;
wire n_7467;
wire n_7468;
wire n_7469;
wire n_747;
wire n_7470;
wire n_7471;
wire n_7472;
wire n_7473;
wire n_7474;
wire n_7475;
wire n_7476;
wire n_7477;
wire n_7478;
wire n_748;
wire n_7480;
wire n_7481;
wire n_7483;
wire n_7484;
wire n_7486;
wire n_7487;
wire n_7488;
wire n_7489;
wire n_749;
wire n_7490;
wire n_7491;
wire n_7492;
wire n_7493;
wire n_7494;
wire n_7495;
wire n_7496;
wire n_7497;
wire n_7498;
wire n_7499;
wire n_75;
wire n_750;
wire n_7500;
wire n_7501;
wire n_7502;
wire n_7503;
wire n_7505;
wire n_7506;
wire n_7507;
wire n_7509;
wire n_751;
wire n_7510;
wire n_7511;
wire n_7512;
wire n_7513;
wire n_7514;
wire n_7515;
wire n_7516;
wire n_7518;
wire n_7519;
wire n_752;
wire n_7520;
wire n_7521;
wire n_7522;
wire n_7523;
wire n_7524;
wire n_7525;
wire n_7526;
wire n_7527;
wire n_7528;
wire TIMEBOOST_net_130;
wire n_753;
wire n_7530;
wire n_7531;
wire n_7532;
wire TIMEBOOST_net_2617;
wire n_7534;
wire n_7535;
wire n_7536;
wire n_7537;
wire n_7538;
wire n_7539;
wire n_754;
wire n_7540;
wire n_7541;
wire n_7542;
wire n_7543;
wire n_7544;
wire n_7545;
wire n_7546;
wire n_7547;
wire n_7548;
wire n_7549;
wire n_755;
wire n_7550;
wire n_7551;
wire n_7552;
wire n_7554;
wire n_7555;
wire n_7556;
wire n_7557;
wire n_7558;
wire n_7559;
wire n_756;
wire n_7560;
wire TIMEBOOST_net_1037;
wire n_7562;
wire n_7563;
wire n_7564;
wire n_7565;
wire n_7566;
wire n_7567;
wire n_7568;
wire n_7569;
wire n_757;
wire n_7570;
wire n_7571;
wire n_7572;
wire n_7573;
wire n_7574;
wire n_7575;
wire n_7577;
wire n_7578;
wire n_7579;
wire n_7580;
wire n_7581;
wire n_7582;
wire n_7583;
wire n_7584;
wire n_7585;
wire n_7586;
wire n_7587;
wire n_7588;
wire n_7589;
wire n_759;
wire n_7590;
wire n_7591;
wire n_7592;
wire n_7593;
wire n_7594;
wire n_7595;
wire n_7596;
wire n_7597;
wire n_7598;
wire n_7599;
wire n_76;
wire n_7600;
wire n_7601;
wire n_7602;
wire n_7603;
wire n_7604;
wire n_7605;
wire n_7606;
wire n_7608;
wire n_7609;
wire n_761;
wire n_7610;
wire n_7611;
wire n_7612;
wire TIMEBOOST_net_849;
wire n_7614;
wire n_7615;
wire n_7617;
wire n_762;
wire n_7621;
wire n_7622;
wire n_7623;
wire n_7624;
wire n_7625;
wire n_7626;
wire n_7627;
wire n_7628;
wire n_7629;
wire n_763;
wire n_7630;
wire n_7631;
wire n_7632;
wire n_7633;
wire n_7634;
wire n_7636;
wire TIMEBOOST_net_79;
wire n_7639;
wire n_764;
wire n_7640;
wire n_7641;
wire n_7644;
wire n_7646;
wire n_7647;
wire n_765;
wire n_7650;
wire n_7651;
wire n_7654;
wire n_7656;
wire n_7657;
wire n_7658;
wire n_7659;
wire n_766;
wire n_7660;
wire n_7661;
wire n_7662;
wire n_7663;
wire n_7665;
wire n_7667;
wire n_7668;
wire n_7669;
wire n_767;
wire n_7670;
wire n_7671;
wire n_7672;
wire n_7673;
wire n_7674;
wire n_7675;
wire n_7676;
wire n_7677;
wire n_7678;
wire n_7679;
wire n_768;
wire n_7680;
wire n_7681;
wire n_7682;
wire n_7683;
wire TIMEBOOST_net_152;
wire n_7685;
wire n_7686;
wire n_7687;
wire n_7689;
wire n_769;
wire n_7690;
wire n_7691;
wire n_7692;
wire n_7693;
wire n_7695;
wire n_7696;
wire n_7697;
wire n_7698;
wire n_7699;
wire n_77;
wire n_770;
wire n_7700;
wire n_7701;
wire n_7702;
wire n_7703;
wire n_7704;
wire n_7706;
wire n_7707;
wire n_7708;
wire n_7709;
wire n_771;
wire n_7710;
wire n_7711;
wire n_7712;
wire n_7713;
wire n_7714;
wire n_7715;
wire n_7716;
wire n_7717;
wire n_7718;
wire n_7720;
wire n_7722;
wire n_7723;
wire n_7724;
wire n_7725;
wire n_7726;
wire n_7727;
wire n_7728;
wire TIMEBOOST_net_1545;
wire n_773;
wire n_7730;
wire n_7731;
wire n_7732;
wire n_7733;
wire n_7735;
wire n_7736;
wire n_7737;
wire n_7738;
wire n_7739;
wire n_7740;
wire n_7741;
wire n_7742;
wire n_7744;
wire n_7745;
wire TIMEBOOST_net_1909;
wire n_7747;
wire n_7748;
wire n_7749;
wire n_7750;
wire n_7751;
wire n_7752;
wire n_7753;
wire n_7754;
wire n_7756;
wire n_7757;
wire n_7759;
wire n_776;
wire n_7760;
wire n_7761;
wire n_7762;
wire n_7763;
wire n_7764;
wire n_7765;
wire n_7766;
wire n_7767;
wire n_7768;
wire n_7769;
wire n_7771;
wire n_7773;
wire TIMEBOOST_net_2789;
wire n_7775;
wire n_7777;
wire n_778;
wire n_7782;
wire n_7783;
wire n_7784;
wire n_7785;
wire n_7786;
wire n_7787;
wire n_7788;
wire n_7789;
wire n_779;
wire n_7790;
wire TIMEBOOST_net_2248;
wire TIMEBOOST_net_1048;
wire n_7794;
wire n_7795;
wire n_7796;
wire n_7797;
wire n_7798;
wire n_7799;
wire n_78;
wire n_780;
wire n_7801;
wire n_7803;
wire n_7804;
wire n_7805;
wire n_7806;
wire n_7807;
wire n_7809;
wire n_781;
wire n_7810;
wire n_7811;
wire n_7812;
wire n_7813;
wire n_7814;
wire n_7815;
wire n_7816;
wire n_7818;
wire n_7819;
wire n_782;
wire n_7820;
wire n_7821;
wire n_7824;
wire n_7825;
wire n_7827;
wire n_7828;
wire n_7829;
wire n_783;
wire n_7830;
wire n_7831;
wire n_7832;
wire n_7834;
wire n_7835;
wire n_7836;
wire n_7839;
wire n_784;
wire n_7840;
wire n_7841;
wire n_7843;
wire n_7844;
wire n_7846;
wire n_7847;
wire n_7848;
wire n_7849;
wire TIMEBOOST_net_2672;
wire n_7850;
wire n_7852;
wire n_7853;
wire n_7854;
wire n_7855;
wire n_7857;
wire n_7858;
wire n_7859;
wire n_786;
wire n_7860;
wire n_7861;
wire n_7862;
wire n_7863;
wire n_7864;
wire n_7865;
wire n_7866;
wire n_7868;
wire n_7869;
wire n_787;
wire n_7870;
wire n_7871;
wire n_7874;
wire n_7875;
wire n_7877;
wire n_788;
wire n_7880;
wire n_7881;
wire TIMEBOOST_net_1049;
wire n_7883;
wire n_7884;
wire n_7885;
wire n_7887;
wire n_7888;
wire n_7889;
wire n_789;
wire n_7891;
wire n_7894;
wire n_7895;
wire n_7896;
wire n_7897;
wire n_7898;
wire n_79;
wire n_790;
wire n_7900;
wire TIMEBOOST_net_1032;
wire n_7902;
wire TIMEBOOST_net_164;
wire n_7905;
wire n_7908;
wire n_7909;
wire n_791;
wire n_7910;
wire n_7912;
wire n_7913;
wire n_7914;
wire n_7915;
wire n_7916;
wire n_7917;
wire n_7918;
wire n_7919;
wire n_792;
wire n_7920;
wire n_7921;
wire n_7922;
wire n_7923;
wire n_7924;
wire n_7925;
wire TIMEBOOST_net_217;
wire n_7927;
wire n_7928;
wire n_7929;
wire n_793;
wire n_7931;
wire n_7932;
wire n_7933;
wire n_7934;
wire n_7935;
wire n_7936;
wire n_7937;
wire n_7938;
wire n_7939;
wire n_794;
wire n_7940;
wire n_7941;
wire TIMEBOOST_net_2007;
wire n_7943;
wire n_7945;
wire n_7948;
wire n_7949;
wire n_795;
wire n_7950;
wire n_7951;
wire n_7952;
wire n_7953;
wire n_7954;
wire n_7955;
wire n_7957;
wire TIMEBOOST_net_316;
wire n_7959;
wire n_796;
wire n_7960;
wire n_7961;
wire n_7962;
wire n_7963;
wire n_7964;
wire n_7965;
wire n_7966;
wire n_7967;
wire n_7968;
wire n_7969;
wire n_797;
wire n_7970;
wire TIMEBOOST_net_161;
wire n_7973;
wire n_7974;
wire n_7975;
wire n_7976;
wire n_7977;
wire n_7978;
wire n_7979;
wire n_798;
wire n_7980;
wire n_7982;
wire n_7984;
wire n_7985;
wire n_7986;
wire n_7987;
wire n_7988;
wire n_7989;
wire n_799;
wire n_7990;
wire n_7991;
wire n_7992;
wire n_7993;
wire n_7995;
wire n_7996;
wire n_7997;
wire n_7998;
wire n_7999;
wire n_80;
wire n_800;
wire n_8001;
wire n_8002;
wire n_8003;
wire n_8004;
wire n_8005;
wire n_8006;
wire n_8007;
wire n_8008;
wire n_8009;
wire n_801;
wire n_8010;
wire n_8011;
wire n_8012;
wire n_8014;
wire n_8015;
wire n_8016;
wire n_8017;
wire n_8018;
wire n_8019;
wire n_802;
wire n_8021;
wire n_8022;
wire TIMEBOOST_net_1584;
wire n_8024;
wire n_8025;
wire n_8027;
wire n_8028;
wire n_803;
wire n_8030;
wire n_8031;
wire n_8032;
wire TIMEBOOST_net_1625;
wire n_8036;
wire n_8037;
wire n_8038;
wire n_8039;
wire n_804;
wire n_8040;
wire n_8041;
wire n_8042;
wire n_8043;
wire n_8044;
wire n_8045;
wire n_8046;
wire n_8047;
wire n_8048;
wire n_805;
wire n_8050;
wire n_8051;
wire n_8052;
wire n_8053;
wire n_8054;
wire n_8057;
wire n_8058;
wire n_8059;
wire n_806;
wire n_8061;
wire n_8062;
wire n_8063;
wire n_8064;
wire n_8065;
wire n_8066;
wire n_8067;
wire n_8068;
wire n_8069;
wire n_807;
wire TIMEBOOST_net_1604;
wire n_8073;
wire n_8074;
wire n_8075;
wire n_8077;
wire n_8078;
wire n_808;
wire n_8081;
wire n_8082;
wire n_8084;
wire n_8085;
wire n_8086;
wire n_8087;
wire n_809;
wire n_8091;
wire n_8093;
wire n_8094;
wire n_8095;
wire n_8096;
wire n_8097;
wire n_8098;
wire n_8099;
wire n_81;
wire n_8100;
wire n_8101;
wire n_8102;
wire n_8103;
wire n_8104;
wire n_8105;
wire n_8106;
wire n_8107;
wire n_8108;
wire n_8109;
wire n_811;
wire n_8110;
wire n_8111;
wire n_8113;
wire n_8114;
wire n_8115;
wire n_8118;
wire n_8119;
wire n_812;
wire n_8121;
wire n_8122;
wire n_8123;
wire n_8124;
wire n_8125;
wire n_8126;
wire n_8127;
wire n_8128;
wire n_813;
wire TIMEBOOST_net_1536;
wire n_8133;
wire n_8134;
wire n_8135;
wire n_8136;
wire n_8138;
wire n_814;
wire n_8140;
wire n_8141;
wire n_8142;
wire n_8143;
wire n_8144;
wire n_8145;
wire TIMEBOOST_net_2554;
wire n_815;
wire n_8150;
wire n_8151;
wire n_8153;
wire n_8154;
wire n_8155;
wire TIMEBOOST_net_1006;
wire n_8158;
wire n_8159;
wire n_816;
wire n_8160;
wire n_8161;
wire n_8162;
wire n_8163;
wire TIMEBOOST_net_2594;
wire n_8166;
wire n_8167;
wire n_8169;
wire n_817;
wire n_8170;
wire n_8172;
wire n_8173;
wire n_8174;
wire n_8175;
wire n_8176;
wire n_8177;
wire TIMEBOOST_net_1105;
wire TIMEBOOST_net_1941;
wire n_818;
wire n_8180;
wire n_8181;
wire n_8182;
wire n_8183;
wire TIMEBOOST_net_1015;
wire n_8186;
wire n_8187;
wire n_8189;
wire n_819;
wire n_8191;
wire n_8192;
wire n_8193;
wire n_8195;
wire n_8196;
wire n_8197;
wire n_8199;
wire n_82;
wire n_820;
wire n_8200;
wire TIMEBOOST_net_1590;
wire n_8204;
wire TIMEBOOST_net_1537;
wire n_8206;
wire n_8207;
wire n_8208;
wire n_821;
wire n_8211;
wire n_8212;
wire n_8213;
wire n_8215;
wire n_8216;
wire TIMEBOOST_net_1078;
wire n_8219;
wire n_822;
wire n_8220;
wire n_8221;
wire n_8224;
wire n_8225;
wire n_8226;
wire n_8227;
wire n_8229;
wire n_823;
wire n_8230;
wire n_8231;
wire n_8232;
wire n_8234;
wire n_8235;
wire n_8236;
wire n_8237;
wire n_8238;
wire n_8239;
wire n_824;
wire n_8240;
wire n_8242;
wire n_8243;
wire n_8245;
wire n_8246;
wire n_8248;
wire n_825;
wire n_8250;
wire n_8251;
wire n_8252;
wire n_8255;
wire n_8256;
wire n_8258;
wire n_8259;
wire n_826;
wire n_8261;
wire n_8263;
wire n_8264;
wire n_8266;
wire TIMEBOOST_net_1556;
wire n_8268;
wire n_8269;
wire n_827;
wire n_8270;
wire n_8271;
wire n_8273;
wire n_8274;
wire n_8275;
wire n_8277;
wire n_828;
wire n_8281;
wire n_8282;
wire n_8283;
wire n_8284;
wire n_8285;
wire n_8288;
wire n_8289;
wire n_829;
wire n_8291;
wire n_8292;
wire n_8293;
wire n_8294;
wire n_8295;
wire n_8296;
wire TIMEBOOST_net_2834;
wire n_83;
wire n_8300;
wire n_8302;
wire n_8303;
wire n_8304;
wire n_8305;
wire n_8306;
wire n_8307;
wire n_8309;
wire n_831;
wire n_8313;
wire n_8315;
wire n_8316;
wire n_8318;
wire n_8319;
wire n_832;
wire n_8320;
wire n_8321;
wire n_8322;
wire n_8324;
wire TIMEBOOST_net_1124;
wire n_8326;
wire n_8327;
wire n_833;
wire n_8332;
wire n_8335;
wire n_8336;
wire n_8337;
wire n_834;
wire n_8340;
wire n_8342;
wire TIMEBOOST_net_1630;
wire n_8344;
wire n_8345;
wire n_8346;
wire n_8348;
wire n_835;
wire TIMEBOOST_net_1632;
wire n_8351;
wire n_8352;
wire n_8353;
wire n_8354;
wire n_8355;
wire n_8358;
wire n_8359;
wire n_836;
wire n_8360;
wire n_8362;
wire n_8364;
wire n_8365;
wire n_8366;
wire n_8367;
wire n_8368;
wire n_8369;
wire n_837;
wire n_8370;
wire n_8371;
wire n_8372;
wire n_8373;
wire n_8374;
wire n_8375;
wire n_8376;
wire n_8378;
wire n_8379;
wire n_8380;
wire n_8381;
wire n_8382;
wire n_8385;
wire n_8386;
wire n_8387;
wire n_8388;
wire n_8389;
wire n_839;
wire n_8390;
wire n_8392;
wire n_8393;
wire n_8394;
wire n_8395;
wire n_8396;
wire n_8398;
wire n_84;
wire n_840;
wire n_8400;
wire n_8401;
wire n_8402;
wire n_8403;
wire n_8404;
wire n_8405;
wire n_8406;
wire n_8407;
wire n_8409;
wire n_841;
wire n_8410;
wire n_8411;
wire n_8413;
wire n_8414;
wire n_8415;
wire TIMEBOOST_net_2165;
wire n_8419;
wire n_842;
wire n_8420;
wire n_8421;
wire n_8423;
wire n_8424;
wire n_8425;
wire n_8426;
wire n_8427;
wire n_8428;
wire n_8429;
wire n_843;
wire n_8430;
wire n_8431;
wire n_8432;
wire n_8433;
wire n_8434;
wire n_8435;
wire n_8437;
wire n_8439;
wire n_844;
wire n_8440;
wire n_8441;
wire n_8443;
wire n_8444;
wire n_8445;
wire n_8448;
wire n_845;
wire n_8450;
wire n_8453;
wire n_8454;
wire n_8455;
wire n_8456;
wire n_8457;
wire n_846;
wire n_8460;
wire n_8461;
wire n_8462;
wire TIMEBOOST_net_1144;
wire n_8464;
wire n_8465;
wire n_8466;
wire n_8468;
wire n_8469;
wire n_847;
wire n_8470;
wire n_8471;
wire n_8474;
wire n_8476;
wire n_8477;
wire n_8478;
wire n_8479;
wire n_848;
wire n_8480;
wire n_8481;
wire n_8482;
wire n_8483;
wire n_8484;
wire n_8487;
wire n_8488;
wire n_8489;
wire n_849;
wire n_8490;
wire n_8491;
wire n_8492;
wire n_8493;
wire n_8494;
wire n_8495;
wire n_8496;
wire n_8497;
wire n_8498;
wire n_8499;
wire n_85;
wire n_850;
wire n_8503;
wire n_8504;
wire n_8506;
wire n_8507;
wire n_8508;
wire n_8509;
wire n_851;
wire n_8511;
wire n_8512;
wire n_8514;
wire n_8515;
wire n_8517;
wire n_8518;
wire n_8519;
wire n_8520;
wire n_8521;
wire n_8522;
wire n_8523;
wire n_8525;
wire n_8526;
wire n_8528;
wire TIMEBOOST_net_290;
wire n_853;
wire n_8530;
wire n_8531;
wire n_8532;
wire n_8533;
wire n_8534;
wire n_8535;
wire n_8536;
wire n_8539;
wire n_854;
wire n_8540;
wire n_8542;
wire TIMEBOOST_net_2866;
wire n_8545;
wire n_8546;
wire n_8547;
wire n_8548;
wire n_855;
wire n_8550;
wire n_8553;
wire n_8554;
wire n_8555;
wire n_8556;
wire n_8557;
wire n_8558;
wire n_856;
wire n_8560;
wire n_8561;
wire n_8562;
wire n_8566;
wire n_8567;
wire n_8568;
wire n_8569;
wire n_8570;
wire n_8571;
wire n_8572;
wire n_8573;
wire n_8574;
wire n_8575;
wire n_8576;
wire n_8578;
wire TIMEBOOST_net_2776;
wire n_858;
wire n_8580;
wire n_8584;
wire n_8585;
wire n_8587;
wire n_8588;
wire n_8589;
wire n_859;
wire n_8590;
wire n_8591;
wire n_8594;
wire n_8595;
wire n_8596;
wire n_8597;
wire n_8599;
wire n_86;
wire n_860;
wire n_8601;
wire n_8602;
wire n_8603;
wire n_8604;
wire n_8605;
wire n_8606;
wire n_8607;
wire n_8608;
wire n_8609;
wire n_861;
wire n_8610;
wire n_8613;
wire n_8617;
wire n_8619;
wire n_8620;
wire n_8621;
wire n_8622;
wire n_8626;
wire n_8627;
wire n_8628;
wire n_8629;
wire n_863;
wire TIMEBOOST_net_1098;
wire n_8632;
wire n_8633;
wire n_8634;
wire n_8635;
wire n_8637;
wire n_8638;
wire n_8639;
wire n_864;
wire n_8640;
wire n_8641;
wire n_8642;
wire n_8644;
wire n_8645;
wire n_8646;
wire n_8647;
wire n_8648;
wire n_8649;
wire n_865;
wire n_8650;
wire n_8651;
wire n_8653;
wire n_8654;
wire n_8656;
wire n_8657;
wire n_8659;
wire n_866;
wire n_8660;
wire n_8661;
wire TIMEBOOST_net_1095;
wire n_8664;
wire n_8666;
wire n_8667;
wire n_8668;
wire n_867;
wire n_8670;
wire n_8671;
wire n_8676;
wire n_8677;
wire n_8678;
wire n_868;
wire n_8680;
wire n_8681;
wire n_8682;
wire n_8684;
wire n_8685;
wire n_8687;
wire n_8688;
wire n_8689;
wire n_869;
wire n_8690;
wire n_8692;
wire n_8694;
wire n_8696;
wire TIMEBOOST_net_237;
wire n_8698;
wire n_8699;
wire n_87;
wire n_870;
wire n_8700;
wire TIMEBOOST_net_258;
wire n_8703;
wire n_8704;
wire n_8706;
wire n_8707;
wire n_8708;
wire n_8711;
wire n_8714;
wire n_8716;
wire n_8717;
wire n_8718;
wire n_8719;
wire n_872;
wire n_8721;
wire n_8722;
wire n_8723;
wire n_8724;
wire n_8725;
wire n_8726;
wire n_8727;
wire n_8728;
wire n_8729;
wire n_873;
wire n_8730;
wire n_8732;
wire n_8733;
wire n_8734;
wire n_8735;
wire n_8736;
wire n_8737;
wire n_8739;
wire n_874;
wire n_8741;
wire n_8742;
wire TIMEBOOST_net_292;
wire n_8746;
wire n_8747;
wire n_8748;
wire TIMEBOOST_net_293;
wire n_875;
wire n_8750;
wire n_8751;
wire n_8753;
wire n_8755;
wire TIMEBOOST_net_1064;
wire n_876;
wire n_8760;
wire n_8761;
wire n_8762;
wire n_8764;
wire n_8765;
wire n_8766;
wire n_8767;
wire n_8769;
wire n_877;
wire n_8770;
wire n_8771;
wire n_8772;
wire n_8773;
wire n_8774;
wire n_8775;
wire n_8776;
wire n_878;
wire n_8781;
wire n_8782;
wire n_8783;
wire n_8784;
wire n_8786;
wire n_8787;
wire n_8788;
wire n_879;
wire n_8790;
wire n_8791;
wire n_8793;
wire n_8794;
wire n_8795;
wire n_8798;
wire n_8799;
wire n_88;
wire n_8800;
wire n_8803;
wire n_8805;
wire n_8806;
wire n_8809;
wire n_881;
wire n_8810;
wire n_8811;
wire n_8812;
wire n_8813;
wire n_8815;
wire n_8817;
wire n_8819;
wire n_882;
wire n_8820;
wire n_8821;
wire n_8822;
wire n_8824;
wire n_8825;
wire n_8828;
wire n_883;
wire n_8831;
wire n_8832;
wire n_8835;
wire n_8836;
wire n_8838;
wire n_8839;
wire n_884;
wire n_8840;
wire TIMEBOOST_net_296;
wire n_8842;
wire TIMEBOOST_net_1916;
wire TIMEBOOST_net_264;
wire n_8846;
wire TIMEBOOST_net_1527;
wire n_8848;
wire n_8849;
wire n_885;
wire n_8850;
wire n_8852;
wire n_8857;
wire n_8858;
wire n_8859;
wire n_886;
wire n_8860;
wire n_8861;
wire n_8862;
wire n_8863;
wire n_8864;
wire n_8865;
wire n_8867;
wire n_8868;
wire n_8869;
wire n_887;
wire n_8870;
wire n_8872;
wire n_8875;
wire n_8876;
wire n_8879;
wire n_888;
wire n_8880;
wire n_8881;
wire n_8885;
wire TIMEBOOST_net_300;
wire n_8887;
wire n_8889;
wire n_889;
wire n_8891;
wire n_8895;
wire n_8898;
wire n_8899;
wire n_89;
wire n_890;
wire n_8900;
wire n_8902;
wire n_8904;
wire n_8905;
wire n_8908;
wire n_891;
wire n_8910;
wire n_8911;
wire TIMEBOOST_net_1198;
wire n_8914;
wire n_8915;
wire n_8916;
wire n_8919;
wire n_892;
wire n_8920;
wire n_8921;
wire n_8922;
wire n_8923;
wire n_8925;
wire n_8927;
wire n_8929;
wire n_893;
wire n_8930;
wire n_8931;
wire n_8932;
wire n_8933;
wire n_8934;
wire n_8936;
wire n_8937;
wire TIMEBOOST_net_2842;
wire n_8939;
wire n_894;
wire n_8941;
wire n_8942;
wire n_8943;
wire n_8944;
wire n_895;
wire n_8950;
wire n_8951;
wire n_8952;
wire n_8953;
wire n_8955;
wire TIMEBOOST_net_383;
wire n_896;
wire n_8961;
wire n_8962;
wire n_8963;
wire n_8964;
wire n_8965;
wire n_8966;
wire n_8967;
wire n_8968;
wire n_8969;
wire n_897;
wire n_8970;
wire n_8971;
wire n_8972;
wire n_8973;
wire n_8974;
wire n_898;
wire n_8980;
wire n_8981;
wire n_8983;
wire n_8985;
wire n_8986;
wire n_8988;
wire n_8989;
wire n_899;
wire n_8990;
wire n_8992;
wire n_8995;
wire n_8998;
wire n_8999;
wire n_90;
wire n_900;
wire n_9001;
wire n_9002;
wire n_9003;
wire n_9004;
wire n_9005;
wire n_9006;
wire n_9007;
wire n_9009;
wire n_901;
wire n_9010;
wire n_9011;
wire n_9012;
wire TIMEBOOST_net_1615;
wire n_9014;
wire TIMEBOOST_net_1136;
wire n_9017;
wire n_9019;
wire n_902;
wire n_9020;
wire n_9021;
wire n_9025;
wire n_9026;
wire n_9027;
wire n_9028;
wire n_9029;
wire n_903;
wire n_9030;
wire n_9032;
wire n_9034;
wire n_9035;
wire n_9036;
wire n_904;
wire TIMEBOOST_net_2858;
wire n_9041;
wire n_9042;
wire n_9044;
wire n_9046;
wire n_9047;
wire TIMEBOOST_net_1636;
wire TIMEBOOST_net_2696;
wire n_905;
wire n_9050;
wire n_9051;
wire n_9053;
wire n_9057;
wire n_9058;
wire n_906;
wire n_9061;
wire n_9065;
wire n_9066;
wire n_907;
wire n_9070;
wire n_9074;
wire n_9075;
wire n_9076;
wire n_9077;
wire n_9078;
wire n_9079;
wire n_908;
wire n_9080;
wire n_9082;
wire n_9083;
wire n_9084;
wire n_9086;
wire n_9087;
wire n_9088;
wire n_9089;
wire n_909;
wire n_9090;
wire n_9091;
wire n_9092;
wire n_9093;
wire n_9095;
wire n_9097;
wire n_9099;
wire n_91;
wire n_910;
wire n_9101;
wire n_9102;
wire n_9105;
wire n_9108;
wire n_911;
wire n_9110;
wire n_9111;
wire n_9112;
wire n_9113;
wire n_9114;
wire n_9115;
wire n_9116;
wire TIMEBOOST_net_2914;
wire n_9119;
wire n_912;
wire n_9121;
wire n_9124;
wire n_9125;
wire n_9127;
wire n_9128;
wire TIMEBOOST_net_361;
wire n_913;
wire n_9130;
wire n_9132;
wire n_9134;
wire n_9135;
wire n_9136;
wire n_9137;
wire n_9138;
wire n_914;
wire n_9140;
wire TIMEBOOST_net_1066;
wire n_9144;
wire n_9145;
wire n_9146;
wire n_9148;
wire n_915;
wire n_9150;
wire n_9151;
wire n_9152;
wire n_9153;
wire n_9157;
wire TIMEBOOST_net_2315;
wire n_916;
wire n_9161;
wire n_9162;
wire n_9163;
wire n_9165;
wire n_9166;
wire n_9167;
wire n_9168;
wire n_9169;
wire n_9170;
wire n_9172;
wire n_9173;
wire n_9177;
wire n_9178;
wire n_918;
wire n_9180;
wire n_9182;
wire n_9185;
wire n_9188;
wire n_9189;
wire n_919;
wire n_9190;
wire n_9191;
wire n_9194;
wire n_9195;
wire TIMEBOOST_net_2412;
wire n_9197;
wire n_9198;
wire n_92;
wire n_920;
wire n_9200;
wire n_9201;
wire n_9202;
wire n_9203;
wire n_9204;
wire n_9205;
wire n_9206;
wire n_9207;
wire n_9208;
wire n_921;
wire n_9210;
wire n_9212;
wire n_9213;
wire n_9214;
wire n_9215;
wire n_9218;
wire n_9219;
wire n_922;
wire n_9220;
wire n_9223;
wire n_9225;
wire n_9226;
wire n_9228;
wire n_9229;
wire n_923;
wire n_9230;
wire n_9232;
wire n_9234;
wire n_9235;
wire n_9236;
wire n_9237;
wire n_9238;
wire n_9239;
wire n_924;
wire n_9240;
wire n_9241;
wire n_9242;
wire n_9243;
wire n_9245;
wire n_9246;
wire n_9247;
wire n_925;
wire n_9253;
wire n_9254;
wire TIMEBOOST_net_269;
wire n_926;
wire n_9260;
wire n_9261;
wire TIMEBOOST_net_336;
wire n_9263;
wire n_9264;
wire n_9265;
wire n_9266;
wire n_9267;
wire n_9268;
wire n_9269;
wire n_927;
wire n_9271;
wire n_9274;
wire n_9275;
wire n_9276;
wire n_928;
wire n_9281;
wire n_9282;
wire n_9283;
wire n_9284;
wire n_9286;
wire n_9288;
wire n_9289;
wire n_929;
wire n_9290;
wire n_9291;
wire n_9292;
wire n_9293;
wire n_9294;
wire TIMEBOOST_net_306;
wire n_9297;
wire n_9298;
wire n_9299;
wire n_93;
wire n_930;
wire n_9302;
wire n_9304;
wire n_9305;
wire n_9306;
wire n_9308;
wire n_9309;
wire n_931;
wire n_9310;
wire n_9311;
wire n_9313;
wire n_9314;
wire n_9317;
wire n_9318;
wire n_9321;
wire n_9322;
wire n_9323;
wire n_9324;
wire n_9325;
wire n_9326;
wire n_9327;
wire n_9328;
wire n_9330;
wire n_9331;
wire n_9332;
wire n_9333;
wire TIMEBOOST_net_2903;
wire n_9335;
wire n_9337;
wire TIMEBOOST_net_2904;
wire n_934;
wire n_9340;
wire n_9341;
wire n_9342;
wire n_9344;
wire n_9345;
wire n_9346;
wire n_9347;
wire n_9348;
wire n_935;
wire n_9350;
wire n_9351;
wire n_9353;
wire n_9354;
wire n_9355;
wire n_9356;
wire n_9357;
wire TIMEBOOST_net_2929;
wire n_9359;
wire n_936;
wire n_9360;
wire n_9362;
wire n_9363;
wire n_9365;
wire n_9366;
wire n_9367;
wire n_9368;
wire n_9369;
wire n_937;
wire n_9370;
wire n_9371;
wire n_9372;
wire n_9374;
wire n_9376;
wire n_9377;
wire n_9378;
wire n_9379;
wire n_938;
wire n_9380;
wire n_9381;
wire n_9385;
wire n_9386;
wire n_9387;
wire n_9389;
wire n_9390;
wire n_9391;
wire n_9392;
wire n_9393;
wire n_9396;
wire n_9397;
wire n_9398;
wire n_9399;
wire n_94;
wire n_9400;
wire n_9401;
wire n_9402;
wire n_9403;
wire n_9404;
wire n_9405;
wire n_9406;
wire n_9407;
wire n_9408;
wire n_9409;
wire n_941;
wire n_9410;
wire n_9411;
wire n_9413;
wire n_9415;
wire TIMEBOOST_net_1689;
wire n_9417;
wire n_9419;
wire n_942;
wire n_9420;
wire n_9422;
wire n_9424;
wire n_9425;
wire n_9428;
wire n_9429;
wire n_943;
wire n_9430;
wire n_9431;
wire n_9432;
wire n_9433;
wire n_9434;
wire n_9435;
wire n_9436;
wire n_9437;
wire n_9438;
wire n_9439;
wire n_944;
wire n_9440;
wire n_9441;
wire n_9442;
wire TIMEBOOST_net_1664;
wire n_9446;
wire n_9447;
wire n_945;
wire n_9450;
wire n_9452;
wire TIMEBOOST_net_1732;
wire n_9456;
wire n_9457;
wire n_946;
wire n_9461;
wire n_9462;
wire n_9463;
wire n_9464;
wire n_9465;
wire n_9468;
wire n_947;
wire n_9474;
wire n_9475;
wire n_9476;
wire n_9478;
wire n_948;
wire n_9480;
wire n_9481;
wire n_9482;
wire n_9485;
wire n_9486;
wire n_9489;
wire n_949;
wire TIMEBOOST_net_1735;
wire n_9492;
wire n_9493;
wire n_9494;
wire n_9495;
wire n_9496;
wire n_95;
wire n_950;
wire n_9502;
wire n_9503;
wire n_9504;
wire n_9505;
wire n_9506;
wire n_9507;
wire n_9509;
wire n_951;
wire n_9510;
wire n_9513;
wire n_9514;
wire n_9515;
wire n_9516;
wire n_9517;
wire n_9518;
wire n_9519;
wire n_9520;
wire n_9521;
wire n_9523;
wire n_9524;
wire n_9525;
wire n_9526;
wire n_9527;
wire n_9528;
wire n_9531;
wire n_9532;
wire n_9535;
wire n_9538;
wire n_954;
wire n_9541;
wire n_9542;
wire n_9543;
wire n_9544;
wire n_9546;
wire n_9547;
wire n_9548;
wire n_9549;
wire n_955;
wire n_9550;
wire n_9551;
wire n_9552;
wire n_9553;
wire n_9554;
wire n_9555;
wire n_9556;
wire n_9558;
wire n_9559;
wire n_956;
wire n_9560;
wire n_9561;
wire n_9562;
wire n_9563;
wire n_9564;
wire n_9565;
wire n_9567;
wire n_9568;
wire n_9569;
wire n_957;
wire n_9570;
wire n_9571;
wire n_9572;
wire n_9573;
wire n_9574;
wire n_9578;
wire n_9579;
wire n_958;
wire n_9580;
wire TIMEBOOST_net_2224;
wire n_9582;
wire n_9583;
wire n_9584;
wire n_9586;
wire n_9587;
wire n_9588;
wire n_959;
wire n_9591;
wire n_9592;
wire n_9593;
wire n_9594;
wire n_9595;
wire n_9596;
wire n_9598;
wire n_96;
wire n_960;
wire n_9601;
wire n_9602;
wire n_9603;
wire n_9604;
wire n_9605;
wire n_9606;
wire n_9607;
wire TIMEBOOST_net_2592;
wire n_9609;
wire n_961;
wire TIMEBOOST_net_2667;
wire n_9611;
wire n_9613;
wire n_9615;
wire n_9616;
wire n_9617;
wire n_9618;
wire n_962;
wire n_9620;
wire n_9621;
wire n_9623;
wire n_9624;
wire n_9625;
wire n_9626;
wire n_9627;
wire n_9628;
wire n_9629;
wire n_963;
wire TIMEBOOST_net_342;
wire n_9631;
wire n_9633;
wire n_9634;
wire n_9635;
wire n_9637;
wire n_9638;
wire n_9639;
wire n_964;
wire n_9640;
wire n_9641;
wire n_9642;
wire n_9643;
wire n_9644;
wire n_9647;
wire n_9648;
wire n_9649;
wire n_965;
wire n_9650;
wire n_9651;
wire n_9653;
wire n_9654;
wire n_9655;
wire n_9656;
wire n_9657;
wire n_9658;
wire n_9659;
wire n_966;
wire n_9660;
wire n_9663;
wire n_9664;
wire n_9665;
wire n_9666;
wire n_9667;
wire n_9668;
wire n_967;
wire n_9670;
wire n_9671;
wire n_9672;
wire TIMEBOOST_net_343;
wire n_9674;
wire n_9675;
wire n_9676;
wire n_9681;
wire n_9682;
wire n_9685;
wire n_9686;
wire n_9687;
wire n_9688;
wire n_9689;
wire n_969;
wire n_9692;
wire n_9693;
wire n_9694;
wire n_9695;
wire n_9696;
wire n_9698;
wire n_9699;
wire n_97;
wire n_970;
wire n_9701;
wire TIMEBOOST_net_2346;
wire n_9703;
wire n_9704;
wire n_9706;
wire n_9707;
wire n_9712;
wire n_9713;
wire n_9714;
wire n_9716;
wire n_9717;
wire n_9718;
wire n_9719;
wire n_972;
wire n_9720;
wire n_9721;
wire n_9722;
wire n_9723;
wire n_9724;
wire n_9726;
wire n_9727;
wire n_9728;
wire n_9729;
wire n_973;
wire n_9730;
wire n_9733;
wire n_9734;
wire n_9735;
wire n_9737;
wire n_9738;
wire TIMEBOOST_net_2580;
wire n_974;
wire n_9740;
wire n_9741;
wire n_9742;
wire n_9743;
wire n_9744;
wire n_9745;
wire n_9746;
wire n_9747;
wire n_9748;
wire n_9749;
wire n_975;
wire n_9750;
wire TIMEBOOST_net_1230;
wire n_9754;
wire n_9755;
wire n_9757;
wire n_9758;
wire TIMEBOOST_net_1702;
wire n_976;
wire n_9760;
wire n_9761;
wire n_9762;
wire n_9763;
wire n_9764;
wire n_9767;
wire n_9768;
wire n_977;
wire n_9770;
wire n_9771;
wire n_9772;
wire n_9773;
wire n_9774;
wire n_9775;
wire n_9776;
wire n_9777;
wire n_978;
wire n_9780;
wire n_9781;
wire n_9782;
wire n_9783;
wire n_9784;
wire n_9785;
wire n_9786;
wire n_9787;
wire n_9788;
wire n_9789;
wire n_979;
wire n_9790;
wire n_9791;
wire TIMEBOOST_net_2020;
wire n_9794;
wire n_9795;
wire n_98;
wire n_980;
wire n_9800;
wire n_9801;
wire TIMEBOOST_net_1738;
wire n_9804;
wire n_9806;
wire n_9807;
wire n_9808;
wire n_9809;
wire n_981;
wire n_9811;
wire n_9813;
wire n_9814;
wire n_9815;
wire n_9816;
wire TIMEBOOST_net_2947;
wire n_9819;
wire n_982;
wire n_9820;
wire n_9822;
wire n_9824;
wire n_9825;
wire n_9826;
wire n_9827;
wire n_9828;
wire n_9829;
wire n_983;
wire n_9830;
wire n_9831;
wire n_9832;
wire n_9833;
wire n_9834;
wire n_9835;
wire n_9836;
wire n_9837;
wire n_9838;
wire n_9839;
wire n_984;
wire n_9840;
wire n_9841;
wire n_9842;
wire n_9843;
wire n_9844;
wire n_9845;
wire TIMEBOOST_net_2001;
wire TIMEBOOST_net_2924;
wire n_9849;
wire n_985;
wire n_9850;
wire n_9851;
wire n_9852;
wire n_9853;
wire n_9854;
wire n_9855;
wire n_9856;
wire TIMEBOOST_net_444;
wire n_9859;
wire n_986;
wire n_9860;
wire n_9861;
wire n_9862;
wire n_9864;
wire n_9866;
wire n_9867;
wire n_9868;
wire n_9869;
wire n_987;
wire n_9870;
wire n_9873;
wire n_9874;
wire n_9875;
wire n_9876;
wire n_9877;
wire n_9878;
wire TIMEBOOST_net_1277;
wire n_988;
wire n_9880;
wire n_9881;
wire n_9882;
wire n_9883;
wire n_9884;
wire n_9885;
wire n_9886;
wire TIMEBOOST_net_1220;
wire n_9888;
wire n_989;
wire n_9890;
wire n_9892;
wire n_9893;
wire n_9895;
wire n_9896;
wire n_9897;
wire n_9898;
wire n_9899;
wire n_99;
wire n_990;
wire n_9900;
wire n_9901;
wire n_9904;
wire n_9905;
wire n_9906;
wire n_9907;
wire n_9908;
wire n_9909;
wire n_991;
wire n_9910;
wire n_9913;
wire n_9915;
wire n_9916;
wire n_9917;
wire n_9918;
wire n_9919;
wire n_992;
wire n_9921;
wire n_9923;
wire n_9924;
wire n_9925;
wire n_9926;
wire n_9927;
wire n_9928;
wire TIMEBOOST_net_450;
wire n_993;
wire n_9930;
wire n_9931;
wire n_9932;
wire n_9934;
wire n_9935;
wire n_9936;
wire n_9937;
wire n_9939;
wire n_9941;
wire n_9942;
wire n_9944;
wire n_9946;
wire n_9947;
wire n_995;
wire n_9951;
wire n_9952;
wire n_9953;
wire n_9954;
wire n_9955;
wire n_9956;
wire n_9957;
wire n_9958;
wire n_9959;
wire n_9960;
wire n_9961;
wire n_9962;
wire n_9963;
wire n_9964;
wire n_9965;
wire n_9966;
wire TIMEBOOST_net_2908;
wire n_9968;
wire n_997;
wire n_9970;
wire n_9971;
wire n_9974;
wire n_9975;
wire n_9978;
wire n_9979;
wire n_998;
wire n_9980;
wire n_9982;
wire n_9983;
wire TIMEBOOST_net_2658;
wire n_9987;
wire n_9988;
wire n_9989;
wire n_999;
wire n_9991;
wire n_9992;
wire TIMEBOOST_net_774;
wire n_9994;
wire n_9999;
wire state_cordic_1_;

// Start cells
in01s01 FE_OCPC1043_n_42367 ( .a(n_42367), .o(FE_OCPN1043_n_42367) );
in01s02 FE_OCPC1044_n_42367 ( .a(FE_OCPN1043_n_42367), .o(FE_OCPN1044_n_42367) );
in01s03 FE_OCPC1047_n_23581 ( .a(n_23581), .o(FE_OCPN1047_n_23581) );
in01m06 FE_OCPC1048_n_23581 ( .a(n_23581), .o(FE_OCPN1048_n_23581) );
in01s06 FE_OCPC1049_n_23581 ( .a(FE_OCPN1047_n_23581), .o(FE_OCPN1049_n_23581) );
in01m08 FE_OCPC1050_n_23581 ( .a(FE_OCPN1048_n_23581), .o(FE_OCPN1050_n_23581) );
in01s01 FE_OCPC1051_n_2702 ( .a(n_2702), .o(FE_OCPN1051_n_2702) );
in01s01 FE_OCPC1052_n_2702 ( .a(FE_OCPN1051_n_2702), .o(FE_OCPN1052_n_2702) );
in01s01 FE_OCPC1055_n_38087 ( .a(n_38087), .o(FE_OCPN1055_n_38087) );
in01s02 FE_OCPC1056_n_38087 ( .a(FE_OCPN1055_n_38087), .o(FE_OCPN1056_n_38087) );
in01s02 FE_OCPC1061_n_44460 ( .a(FE_OCP_RBN4288_n_44563), .o(FE_OCPN1061_n_44460) );
in01s01 FE_OCPC1063_n_44461 ( .a(FE_OCP_RBN6740_n_44563), .o(FE_OCPN1063_n_44461) );
in01s01 FE_OCPC1064_n_44461 ( .a(FE_OCP_RBN6740_n_44563), .o(FE_OCPN1064_n_44461) );
in01s01 FE_OCPC1065_n_44461 ( .a(FE_OCPN1064_n_44461), .o(FE_OCPN1065_n_44461) );
in01s01 FE_OCPC1066_n_44461 ( .a(FE_OCPN1065_n_44461), .o(FE_OCPN1066_n_44461) );
in01s01 FE_OCPC1067_n_44461 ( .a(FE_OCPN1065_n_44461), .o(FE_OCPN1067_n_44461) );
in01s02 FE_OCPC1068_n_21973 ( .a(n_21973), .o(FE_OCPN1068_n_21973) );
in01s01 FE_OCPC1070_n_44267 ( .a(FE_OCP_RBN6185_n_44267), .o(FE_OCPN1070_n_44267) );
in01s02 FE_OCPC1071_n_44267 ( .a(FE_OCPN1070_n_44267), .o(FE_OCPN1071_n_44267) );
in01f02 FE_OCPC1072_n_12638 ( .a(n_12638), .o(FE_OCPN1072_n_12638) );
in01f02 FE_OCPC1073_n_12638 ( .a(FE_OCPN1072_n_12638), .o(FE_OCPN1073_n_12638) );
in01s06 FE_OCPC1077_n_13831 ( .a(FE_OCP_RBN6650_n_13818), .o(FE_OCPN1077_n_13831) );
in01s01 FE_OCPC1078_n_8915 ( .a(n_8915), .o(FE_OCPN1078_n_8915) );
in01s01 FE_OCPC1079_n_8915 ( .a(FE_OCPN1078_n_8915), .o(FE_OCPN1079_n_8915) );
in01s01 FE_OCPC1080_n_24819 ( .a(n_24819), .o(FE_OCPN1080_n_24819) );
in01s01 FE_OCPC1081_n_24819 ( .a(FE_OCPN1080_n_24819), .o(FE_OCPN1081_n_24819) );
in01s01 FE_OCPC1082_n_8388 ( .a(n_8388), .o(FE_OCPN1082_n_8388) );
in01s01 FE_OCPC1083_n_8388 ( .a(FE_OCPN1082_n_8388), .o(FE_OCPN1083_n_8388) );
in01s01 FE_OCPC1084_n_8388 ( .a(FE_OCPN1082_n_8388), .o(FE_OCPN1084_n_8388) );
in01s01 FE_OCPC1085_n_8499 ( .a(n_8499), .o(FE_OCPN1085_n_8499) );
in01s01 FE_OCPC1086_n_8499 ( .a(FE_OCPN1085_n_8499), .o(FE_OCPN1086_n_8499) );
in01s01 FE_OCPC1087_n_25481 ( .a(FE_OCP_RBN6797_n_25211), .o(FE_OCPN1087_n_25481) );
in01s01 FE_OCPC1088_n_25481 ( .a(FE_OCPN1087_n_25481), .o(FE_OCPN1088_n_25481) );
in01s01 FE_OCPC1089_n_39089 ( .a(n_39089), .o(FE_OCPN1089_n_39089) );
in01s02 FE_OCPC1090_n_39089 ( .a(FE_OCPN1089_n_39089), .o(FE_OCPN1090_n_39089) );
in01s01 FE_OCPC1091_n_9014 ( .a(FE_OCP_RBN6721_FE_OCP_DRV_N6264_n_9014), .o(FE_OCPN1091_n_9014) );
in01s01 FE_OCPC1092_n_9014 ( .a(FE_OCPN1091_n_9014), .o(FE_OCPN1092_n_9014) );
in01s01 FE_OCPC1093_n_4459 ( .a(n_4459), .o(FE_OCPN1093_n_4459) );
in01s01 FE_OCPC1094_n_4459 ( .a(FE_OCPN1093_n_4459), .o(FE_OCPN1094_n_4459) );
in01s01 FE_OCPC1095_n_25318 ( .a(n_25318), .o(FE_OCPN1095_n_25318) );
in01s01 FE_OCPC1096_n_25318 ( .a(FE_OCPN1095_n_25318), .o(FE_OCPN1096_n_25318) );
in01s06 FE_OCPC1201_n_45450 ( .a(FE_OCP_RBN5513_n_44365), .o(FE_OCPN1201_n_45450) );
in01s20 FE_OCPC1202_n_45450 ( .a(FE_OCPN1201_n_45450), .o(FE_OCPN1202_n_45450) );
in01s01 FE_OCPC1203_n_7663 ( .a(n_7663), .o(FE_OCPN1203_n_7663) );
in01s01 FE_OCPC1204_n_7663 ( .a(FE_OCPN1203_n_7663), .o(FE_OCPN1204_n_7663) );
in01s02 FE_OCPC1205_n_46990 ( .a(n_46990), .o(FE_OCPN1205_n_46990) );
in01s02 FE_OCPC1206_n_46990 ( .a(FE_OCPN1205_n_46990), .o(FE_OCPN1206_n_46990) );
in01s01 FE_OCPC1207_n_8185 ( .a(FE_OCP_RBN2678_n_8163), .o(FE_OCPN1207_n_8185) );
in01s01 FE_OCPC1208_n_8185 ( .a(FE_OCPN1207_n_8185), .o(FE_OCPN1208_n_8185) );
in01s01 FE_OCPC1209_n_8846 ( .a(n_8846), .o(FE_OCPN1209_n_8846) );
in01s01 FE_OCPC1210_n_8846 ( .a(FE_OCPN1209_n_8846), .o(FE_OCPN1210_n_8846) );
in01s01 FE_OCPC1212_n_19354 ( .a(FE_OCP_DRV_N1447_n_19354), .o(FE_OCPN1212_n_19354) );
in01s01 FE_OCPC1213_n_21166 ( .a(n_21166), .o(FE_OCPN1213_n_21166) );
in01s01 FE_OCPC1214_n_21166 ( .a(FE_OCPN1213_n_21166), .o(FE_OCPN1214_n_21166) );
in01m02 FE_OCPC1215_n_21946 ( .a(n_21946), .o(FE_OCPN1215_n_21946) );
in01m06 FE_OCPC1216_n_21946 ( .a(FE_OCPN1215_n_21946), .o(FE_OCPN1216_n_21946) );
in01s01 FE_OCPC1217_n_11012 ( .a(n_11012), .o(FE_OCPN1217_n_11012) );
in01s01 FE_OCPC1218_n_11012 ( .a(FE_OCPN1217_n_11012), .o(FE_OCPN1218_n_11012) );
in01s01 FE_OCPC1219_n_40863 ( .a(n_40863), .o(FE_OCPN1219_n_40863) );
in01s01 FE_OCPC1220_n_40863 ( .a(FE_OCPN1219_n_40863), .o(FE_OCPN1220_n_40863) );
in01s01 FE_OCPC1221_n_41211 ( .a(n_41211), .o(FE_OCPN1221_n_41211) );
in01s01 FE_OCPC1222_n_41211 ( .a(FE_OCPN1221_n_41211), .o(FE_OCPN1222_n_41211) );
in01s01 FE_OCPC1223_n_43521 ( .a(n_43521), .o(FE_OCPN1223_n_43521) );
in01s01 FE_OCPC1224_n_43521 ( .a(FE_OCPN1223_n_43521), .o(FE_OCPN1224_n_43521) );
in01s01 FE_OCPC1226_n_43357 ( .a(n_43341), .o(FE_OCPN1226_n_43357) );
in01s01 FE_OCPC1227_n_43605 ( .a(n_43605), .o(FE_OCPN1227_n_43605) );
in01s01 FE_OCPC1228_n_43605 ( .a(FE_OCPN1227_n_43605), .o(FE_OCPN1228_n_43605) );
in01s01 FE_OCPC1229_n_43601 ( .a(n_43601), .o(FE_OCPN1229_n_43601) );
in01s01 FE_OCPC1230_n_43601 ( .a(FE_OCPN1229_n_43601), .o(FE_OCPN1230_n_43601) );
in01s01 FE_OCPC1233_n_33341 ( .a(n_33341), .o(FE_OCPN1233_n_33341) );
in01s01 FE_OCPC1234_n_33341 ( .a(FE_OCPN1233_n_33341), .o(FE_OCPN1234_n_33341) );
in01f06 FE_OCPC1235_n_27207 ( .a(n_27207), .o(FE_OCPN1235_n_27207) );
in01m04 FE_OCPC1236_n_27207 ( .a(FE_OCPN1235_n_27207), .o(FE_OCPN1236_n_27207) );
in01s01 FE_OCPC1237_n_30470 ( .a(n_30470), .o(FE_OCPN1237_n_30470) );
in01s01 FE_OCPC1238_n_30470 ( .a(FE_OCPN1237_n_30470), .o(FE_OCPN1238_n_30470) );
in01m01 FE_OCPC1239_n_13412 ( .a(n_13412), .o(FE_OCPN1239_n_13412) );
in01s02 FE_OCPC1240_n_13412 ( .a(FE_OCPN1239_n_13412), .o(FE_OCPN1240_n_13412) );
in01s01 FE_OCPC1241_n_12633 ( .a(n_12633), .o(FE_OCPN1241_n_12633) );
in01s02 FE_OCPC1242_n_12633 ( .a(FE_OCPN1241_n_12633), .o(FE_OCPN1242_n_12633) );
in01s01 FE_OCPC1243_n_13992 ( .a(FE_OCP_RBN5039_n_13927), .o(FE_OCPN1243_n_13992) );
in01s01 FE_OCPC1244_n_13992 ( .a(FE_OCPN1243_n_13992), .o(FE_OCPN1244_n_13992) );
in01s01 FE_OCPC1245_n_19645 ( .a(n_19645), .o(FE_OCPN1245_n_19645) );
in01s01 FE_OCPC1246_n_19645 ( .a(FE_OCPN1245_n_19645), .o(FE_OCPN1246_n_19645) );
in01s01 FE_OCPC1247_n_22291 ( .a(n_22291), .o(FE_OCPN1247_n_22291) );
in01s01 FE_OCPC1248_n_22291 ( .a(FE_OCPN1247_n_22291), .o(FE_OCPN1248_n_22291) );
in01s01 FE_OCPC1249_n_13882 ( .a(n_13882), .o(FE_OCPN1249_n_13882) );
in01s02 FE_OCPC1250_n_13882 ( .a(FE_OCPN1249_n_13882), .o(FE_OCPN1250_n_13882) );
in01s01 FE_OCPC1251_n_19314 ( .a(FE_OCP_DRV_N1446_n_19314), .o(FE_OCPN1251_n_19314) );
in01s01 FE_OCPC1252_n_19314 ( .a(FE_OCPN1251_n_19314), .o(FE_OCPN1252_n_19314) );
in01m01 FE_OCPC1253_n_23815 ( .a(n_23815), .o(FE_OCPN1253_n_23815) );
in01s01 FE_OCPC1256_n_28656 ( .a(FE_OCPUNCON3473_n_28656), .o(FE_OCPN1256_n_28656) );
in01s01 FE_OCPC1257_n_18854 ( .a(n_18854), .o(FE_OCPN1257_n_18854) );
in01s01 FE_OCPC1258_n_18854 ( .a(FE_OCPN1257_n_18854), .o(FE_OCPN1258_n_18854) );
in01s02 FE_OCPC1263_n_20971 ( .a(FE_OCP_RBN3003_n_20432), .o(FE_OCPN1263_n_20971) );
in01s01 FE_OCPC1267_n_29155 ( .a(n_29155), .o(FE_OCPN1267_n_29155) );
in01s01 FE_OCPC1268_n_29155 ( .a(FE_OCPN1267_n_29155), .o(FE_OCPN1268_n_29155) );
in01s01 FE_OCPC1269_n_30577 ( .a(n_30577), .o(FE_OCPN1269_n_30577) );
in01s01 FE_OCPC1270_n_30577 ( .a(FE_OCPN1269_n_30577), .o(FE_OCPN1270_n_30577) );
in01s01 FE_OCPC1271_n_31403 ( .a(FE_OFN4731_n_31403), .o(FE_OCPN1271_n_31403) );
in01s01 FE_OCPC1272_n_31403 ( .a(FE_OCPN1271_n_31403), .o(FE_OCPN1272_n_31403) );
in01s01 FE_OCPC1274_n_15708 ( .a(n_15762), .o(FE_OCPN1274_n_15708) );
in01s01 FE_OCPC1275_n_31773 ( .a(n_31773), .o(FE_OCPN1275_n_31773) );
in01s01 FE_OCPC1276_n_31773 ( .a(FE_OCPN1275_n_31773), .o(FE_OCPN1276_n_31773) );
in01s01 FE_OCPC1277_n_15656 ( .a(n_15656), .o(FE_OCPN1277_n_15656) );
in01s01 FE_OCPC1278_n_15656 ( .a(FE_OCPN1277_n_15656), .o(FE_OCPN1278_n_15656) );
in01s01 FE_OCPC1279_n_30823 ( .a(n_30823), .o(FE_OCPN1279_n_30823) );
in01s01 FE_OCPC1280_n_30823 ( .a(FE_OCPN1279_n_30823), .o(FE_OCPN1280_n_30823) );
in01s01 FE_OCPC1281_n_21007 ( .a(n_21007), .o(FE_OCPN1281_n_21007) );
in01s01 FE_OCPC1287_n_29375 ( .a(FE_OCPUNCON1743_n_29375), .o(FE_OCPN1287_n_29375) );
in01s01 FE_OCPC1288_n_29375 ( .a(FE_OCPN1287_n_29375), .o(FE_OCPN1288_n_29375) );
in01s01 FE_OCPC1289_n_19384 ( .a(FE_OFN4804_n_19384), .o(FE_OCPN1289_n_19384) );
in01s01 FE_OCPC1290_n_19384 ( .a(FE_OCPN1289_n_19384), .o(FE_OCPN1290_n_19384) );
in01s01 FE_OCPC1291_n_29439 ( .a(n_29439), .o(FE_OCPN1291_n_29439) );
in01s01 FE_OCPC1293_n_26296 ( .a(FE_OCP_DRV_N1482_n_26296), .o(FE_OCPN1293_n_26296) );
in01s01 FE_OCPC1294_n_26296 ( .a(FE_OCPN1293_n_26296), .o(FE_OCPN1294_n_26296) );
in01s06 FE_OCPC1295_n_45450 ( .a(FE_OCP_RBN5513_n_44365), .o(FE_OCPN1295_n_45450) );
in01m06 FE_OCPC1296_n_45450 ( .a(FE_OCPN1295_n_45450), .o(FE_OCPN1296_n_45450) );
in01s01 FE_OCPC1297_n_30134 ( .a(n_30134), .o(FE_OCPN1297_n_30134) );
in01s02 FE_OCPC1298_n_30134 ( .a(FE_OCPN1297_n_30134), .o(FE_OCPN1298_n_30134) );
in01s01 FE_OCPC1299_n_30136 ( .a(n_30136), .o(FE_OCPN1299_n_30136) );
in01s01 FE_OCPC1300_n_30136 ( .a(FE_OCPN1299_n_30136), .o(FE_OCPN1300_n_30136) );
in01s01 FE_OCPC1302_n_23771 ( .a(n_23772), .o(FE_OCPN1302_n_23771) );
in01s01 FE_OCPC1303_n_35945 ( .a(n_35945), .o(FE_OCPN1303_n_35945) );
in01s02 FE_OCPC1304_n_35945 ( .a(FE_OCPN1303_n_35945), .o(FE_OCPN1304_n_35945) );
in01s01 FE_OCPC1306_n_13721 ( .a(FE_OCPN1696_n_13721), .o(FE_OCPN1306_n_13721) );
in01s01 FE_OCPC1307_n_23677 ( .a(n_23677), .o(FE_OCPN1307_n_23677) );
in01m04 FE_OCPC1309_n_25431 ( .a(n_25431), .o(FE_OCPN1309_n_25431) );
in01f04 FE_OCPC1310_n_25431 ( .a(FE_OCPN1309_n_25431), .o(FE_OCPN1310_n_25431) );
in01s01 FE_OCPC1311_FE_OCP_RBN1024_n_24125 ( .a(FE_OCP_RBN1024_n_24125), .o(FE_OCPN1311_FE_OCP_RBN1024_n_24125) );
in01s02 FE_OCPC1312_FE_OCP_RBN1024_n_24125 ( .a(FE_OCPN1311_FE_OCP_RBN1024_n_24125), .o(FE_OCPN1312_FE_OCP_RBN1024_n_24125) );
in01s01 FE_OCPC1313_n_25126 ( .a(n_25126), .o(FE_OCPN1313_n_25126) );
in01s01 FE_OCPC1314_n_25126 ( .a(FE_OCPN1313_n_25126), .o(FE_OCPN1314_n_25126) );
in01s02 FE_OCPC1316_n_20265 ( .a(n_20266), .o(FE_OCPN1316_n_20265) );
in01s01 FE_OCPC1317_n_24682 ( .a(n_24682), .o(FE_OCPN1317_n_24682) );
in01s01 FE_OCPC1318_n_24682 ( .a(FE_OCPN1317_n_24682), .o(FE_OCPN1318_n_24682) );
in01s01 FE_OCPC1319_n_31403 ( .a(FE_OFN4731_n_31403), .o(FE_OCPN1319_n_31403) );
in01s01 FE_OCPC1320_n_31403 ( .a(FE_OCPN1319_n_31403), .o(FE_OCPN1320_n_31403) );
in01s01 FE_OCPC1321_n_33714 ( .a(n_33714), .o(FE_OCPN1321_n_33714) );
in01s01 FE_OCPC1324_n_14577 ( .a(FE_OCP_RBN2081_n_14554), .o(FE_OCPN1324_n_14577) );
in01s01 FE_OCPC1325_n_45050 ( .a(n_45050), .o(FE_OCPN1325_n_45050) );
in01s01 FE_OCPC1326_n_45050 ( .a(FE_OCPN1325_n_45050), .o(FE_OCPN1326_n_45050) );
in01s01 FE_OCPC1327_n_16192 ( .a(n_16192), .o(FE_OCPN1327_n_16192) );
in01s01 FE_OCPC1329_FE_OFN1196_n_27014 ( .a(FE_OFN1196_n_27014), .o(FE_OCPN1329_FE_OFN1196_n_27014) );
in01s01 FE_OCPC1330_FE_OFN1196_n_27014 ( .a(FE_OCPN1329_FE_OFN1196_n_27014), .o(FE_OCPN1330_FE_OFN1196_n_27014) );
in01s01 FE_OCPC1331_n_30281 ( .a(n_30281), .o(FE_OCPN1331_n_30281) );
in01s01 FE_OCPC1332_n_30281 ( .a(FE_OCPN1331_n_30281), .o(FE_OCPN1332_n_30281) );
in01s01 FE_OCPC1333_n_23467 ( .a(FE_RN_1116_0), .o(FE_OCPN1333_n_23467) );
in01s01 FE_OCPC1334_n_23467 ( .a(FE_OCPN1333_n_23467), .o(FE_RN_1641_0) );
in01s01 FE_OCPC1335_n_25673 ( .a(n_25673), .o(FE_OCPN1335_n_25673) );
in01s01 FE_OCPC1336_n_25673 ( .a(FE_OCPN1335_n_25673), .o(FE_OCPN1336_n_25673) );
in01s01 FE_OCPC1337_n_25775 ( .a(n_25775), .o(FE_OCPN1337_n_25775) );
in01s01 FE_OCPC1338_n_25775 ( .a(FE_OCPN1337_n_25775), .o(FE_OCPN1338_n_25775) );
in01s03 FE_OCPC1340_n_27246 ( .a(n_27366), .o(FE_OCPN1340_n_27246) );
in01s10 FE_OCPC1341_n_11927 ( .a(n_11927), .o(FE_OCPN1341_n_11927) );
in01s20 FE_OCPC1342_n_11927 ( .a(FE_OCPN1341_n_11927), .o(FE_OCPN1342_n_11927) );
in01s02 FE_OCPC1343_n_12313 ( .a(n_12313), .o(FE_OCPN1343_n_12313) );
in01s06 FE_OCPC1344_n_12313 ( .a(FE_OCPN1343_n_12313), .o(FE_OCPN1344_n_12313) );
in01s01 FE_OCPC1345_n_24142 ( .a(n_24142), .o(FE_OCPN1345_n_24142) );
in01s01 FE_OCPC1346_n_24142 ( .a(FE_OCPN1345_n_24142), .o(FE_OCPN1346_n_24142) );
in01s01 FE_OCPC1350_n_35312 ( .a(FE_OCP_DRV_N1427_n_35312), .o(FE_OCPN1350_n_35312) );
in01s01 FE_OCPC1351_n_26530 ( .a(n_26530), .o(FE_OCPN1351_n_26530) );
in01s01 FE_OCPC1352_n_26530 ( .a(FE_OCPN1351_n_26530), .o(FE_OCPN1352_n_26530) );
in01s01 FE_OCPC1353_n_22484 ( .a(n_22484), .o(FE_OCPN1353_n_22484) );
in01s02 FE_OCPC1354_n_22484 ( .a(FE_OCPN1353_n_22484), .o(FE_OCPN1354_n_22484) );
in01s01 FE_OCPC1355_n_23335 ( .a(n_23335), .o(FE_OCPN1355_n_23335) );
in01s02 FE_OCPC1356_n_23335 ( .a(FE_OCPN1355_n_23335), .o(FE_OCPN1356_n_23335) );
in01m01 FE_OCPC1357_n_17778 ( .a(n_17778), .o(FE_OCPN1357_n_17778) );
in01s01 FE_OCPC1358_n_17778 ( .a(FE_OCPN1357_n_17778), .o(FE_OCPN1358_n_17778) );
in01s06 FE_OCPC1359_n_12370 ( .a(n_12370), .o(FE_OCPN1359_n_12370) );
in01m03 FE_OCPC1360_n_12370 ( .a(FE_OCPN1359_n_12370), .o(FE_OCPN1360_n_12370) );
in01s02 FE_OCPC1361_n_23684 ( .a(n_23684), .o(FE_OCPN1361_n_23684) );
in01m04 FE_OCPC1362_n_23684 ( .a(FE_OCPN1361_n_23684), .o(FE_OCPN1362_n_23684) );
in01s02 FE_OCPC1363_n_29615 ( .a(n_29615), .o(FE_OCPN1363_n_29615) );
in01s04 FE_OCPC1364_n_29615 ( .a(FE_OCPN1363_n_29615), .o(FE_OCPN1364_n_29615) );
in01s01 FE_OCPC1365_n_29573 ( .a(FE_OCP_DRV_N1892_n_29573), .o(FE_OCPN1365_n_29573) );
in01s01 FE_OCPC1366_n_29573 ( .a(FE_OCPN1365_n_29573), .o(FE_OCPN1366_n_29573) );
in01s01 FE_OCPC1367_n_23923 ( .a(n_23923), .o(FE_OCPN1367_n_23923) );
in01s01 FE_OCPC1368_n_23923 ( .a(FE_OCPN1367_n_23923), .o(FE_OCPN1368_n_23923) );
in01s01 FE_OCPC1369_n_34288 ( .a(n_34288), .o(FE_OCPN1369_n_34288) );
in01s01 FE_OCPC1370_n_34288 ( .a(FE_OCPN1369_n_34288), .o(FE_OCPN1370_n_34288) );
in01s01 FE_OCPC1371_n_13510 ( .a(n_13510), .o(FE_OCPN1371_n_13510) );
in01s01 FE_OCPC1372_n_13510 ( .a(FE_OCPN1371_n_13510), .o(FE_OCPN1372_n_13510) );
in01s01 FE_OCPC1373_n_34051 ( .a(n_34051), .o(FE_OCPN1373_n_34051) );
in01s01 FE_OCPC1375_n_30612 ( .a(n_30612), .o(FE_OCPN1375_n_30612) );
in01s01 FE_OCPC1376_n_30612 ( .a(FE_OCPN1375_n_30612), .o(FE_OCPN1376_n_30612) );
in01s01 FE_OCPC1377_n_17836 ( .a(FE_OCPUNCON5302_n_17836), .o(FE_OCPN1377_n_17836) );
in01s01 FE_OCPC1379_n_33640 ( .a(n_33640), .o(FE_OCPN1379_n_33640) );
in01s01 FE_OCPC1380_n_33640 ( .a(FE_OCPN1379_n_33640), .o(FE_OCPN1380_n_33640) );
in01s01 FE_OCPC1381_n_45026 ( .a(n_45026), .o(FE_OCPN1381_n_45026) );
in01s06 FE_OCPC1382_n_45026 ( .a(FE_OCPN1381_n_45026), .o(FE_OCPN1382_n_45026) );
in01s01 FE_OCPC1383_n_21896 ( .a(n_21896), .o(FE_OCPN1383_n_21896) );
in01s01 FE_OCPC1384_n_21896 ( .a(FE_OCPN1383_n_21896), .o(FE_OCPN1384_n_21896) );
in01s01 FE_OCPC1385_n_21199 ( .a(n_21199), .o(FE_OCPN1385_n_21199) );
in01s01 FE_OCPC1386_n_21199 ( .a(FE_OCPN1385_n_21199), .o(FE_OCPN1386_n_21199) );
in01s01 FE_OCPC1387_n_20555 ( .a(n_20555), .o(FE_OCPN1387_n_20555) );
in01s01 FE_OCPC1388_n_20555 ( .a(FE_OCPN1387_n_20555), .o(FE_OCPN1388_n_20555) );
in01s01 FE_OCPC1389_n_26054 ( .a(n_26054), .o(FE_OCPN1389_n_26054) );
in01s01 FE_OCPC1390_n_26054 ( .a(FE_OCPN1389_n_26054), .o(FE_OCPN1390_n_26054) );
in01s01 FE_OCPC1391_n_15462 ( .a(n_15462), .o(FE_OCPN1391_n_15462) );
in01s01 FE_OCPC1393_n_22801 ( .a(n_22801), .o(FE_OCPN1393_n_22801) );
in01s02 FE_OCPC1394_n_22801 ( .a(FE_OCPN1393_n_22801), .o(FE_OCPN1394_n_22801) );
in01s01 FE_OCPC1395_n_27211 ( .a(n_27211), .o(FE_OCPN1395_n_27211) );
in01s01 FE_OCPC1396_n_27211 ( .a(FE_OCPN1395_n_27211), .o(FE_OCPN1396_n_27211) );
in01s01 FE_OCPC1397_n_14742 ( .a(n_14742), .o(FE_OCPN1397_n_14742) );
in01s01 FE_OCPC1398_n_14742 ( .a(FE_OCPN1397_n_14742), .o(FE_OCPN1398_n_14742) );
in01m20 FE_OCPC1400_n_28095 ( .a(n_27911), .o(FE_OCPN1400_n_28095) );
in01s01 FE_OCPC1401_FE_OFN1196_n_27014 ( .a(FE_OCPN1330_FE_OFN1196_n_27014), .o(FE_OCPN1401_FE_OFN1196_n_27014) );
in01s06 FE_OCPC1402_FE_OFN1196_n_27014 ( .a(FE_OCPN1401_FE_OFN1196_n_27014), .o(FE_OCPN1402_FE_OFN1196_n_27014) );
in01s01 FE_OCPC1403_n_30823 ( .a(FE_OCPN1280_n_30823), .o(FE_OCPN1403_n_30823) );
in01s02 FE_OCPC1404_n_30823 ( .a(FE_OCPN1403_n_30823), .o(FE_OCPN1404_n_30823) );
in01s01 FE_OCPC1435_n_21278 ( .a(n_21278), .o(FE_OCPN1435_n_21278) );
in01s06 FE_OCPC1605_n_45697 ( .a(n_45697), .o(FE_OCPN1605_n_45697) );
in01s20 FE_OCPC1606_n_45697 ( .a(FE_OCPN1605_n_45697), .o(FE_OCPN1606_n_45697) );
in01s04 FE_OCPC1607_n_18176 ( .a(n_18176), .o(FE_OCPN1607_n_18176) );
in01s04 FE_OCPC1608_n_18176 ( .a(FE_OCPN1607_n_18176), .o(FE_OCPN1608_n_18176) );
in01s01 FE_OCPC1609_n_23503 ( .a(n_23503), .o(FE_OCPN1609_n_23503) );
in01s01 FE_OCPC1610_n_23503 ( .a(FE_OCPN1609_n_23503), .o(FE_OCPN1610_n_23503) );
in01s01 FE_OCPC1611_n_44174 ( .a(FE_OCP_RBN3171_n_44211), .o(FE_OCPN1611_n_44174) );
in01s01 FE_OCPC1612_n_44174 ( .a(FE_OCPN1611_n_44174), .o(FE_OCPN1612_n_44174) );
in01s01 FE_OCPC1613_n_7630 ( .a(n_7630), .o(FE_OCPN1613_n_7630) );
in01s01 FE_OCPC1614_n_7630 ( .a(FE_OCPN1613_n_7630), .o(FE_OCPN1614_n_7630) );
in01s01 FE_OCPC1615_n_12371 ( .a(n_12371), .o(FE_OCPN1615_n_12371) );
in01s02 FE_OCPC1616_n_12371 ( .a(FE_OCPN1615_n_12371), .o(FE_OCPN1616_n_12371) );
in01s01 FE_OCPC1617_n_8444 ( .a(n_8444), .o(FE_OCPN1617_n_8444) );
in01s01 FE_OCPC1618_n_8444 ( .a(FE_OCPN1617_n_8444), .o(FE_OCPN1618_n_8444) );
in01m01 FE_OCPC1619_n_3361 ( .a(n_3361), .o(FE_OCPN1619_n_3361) );
in01s02 FE_OCPC1620_n_3361 ( .a(FE_OCPN1619_n_3361), .o(FE_OCPN1620_n_3361) );
in01s01 FE_OCPC1621_n_36947 ( .a(n_36947), .o(FE_OCPN1621_n_36947) );
in01s01 FE_OCPC1622_n_36947 ( .a(FE_OCPN1621_n_36947), .o(FE_OCPN1622_n_36947) );
in01s01 FE_OCPC1623_n_37661 ( .a(n_37661), .o(FE_OCPN1623_n_37661) );
in01s01 FE_OCPC1624_n_37661 ( .a(FE_OCPN1623_n_37661), .o(FE_OCPN1624_n_37661) );
in01s01 FE_OCPC1625_n_38135 ( .a(n_38135), .o(FE_OCPN1625_n_38135) );
in01s01 FE_OCPC1626_n_38135 ( .a(FE_OCPN1625_n_38135), .o(FE_OCPN1626_n_38135) );
in01s01 FE_OCPC1627_n_34452 ( .a(n_34452), .o(FE_OCPN1627_n_34452) );
in01s01 FE_OCPC1628_n_34452 ( .a(FE_OCPN1627_n_34452), .o(FE_OCPN1628_n_34452) );
in01s01 FE_OCPC1629_n_33196 ( .a(n_33196), .o(FE_OCPN1629_n_33196) );
in01s01 FE_OCPC1630_n_33196 ( .a(FE_OCPN1629_n_33196), .o(FE_OCPN1630_n_33196) );
in01s01 FE_OCPC1632_n_1835 ( .a(n_1836), .o(FE_OCPN1632_n_1835) );
in01s01 FE_OCPC1633_n_33588 ( .a(n_33588), .o(FE_OCPN1633_n_33588) );
in01s01 FE_OCPC1634_n_33588 ( .a(FE_OCPN1633_n_33588), .o(FE_OCPN1634_n_33588) );
in01s01 FE_OCPC1635_n_18860 ( .a(FE_OCP_DRV_N5354_n_18860), .o(FE_OCPN1635_n_18860) );
in01s01 FE_OCPC1636_n_18860 ( .a(FE_OCPN1635_n_18860), .o(FE_OCPN1636_n_18860) );
in01s01 FE_OCPC1637_n_45081 ( .a(n_45081), .o(FE_OCPN1637_n_45081) );
in01s01 FE_OCPC1638_n_45081 ( .a(FE_OCPN1637_n_45081), .o(FE_OCPN1638_n_45081) );
in01s01 FE_OCPC1639_n_35367 ( .a(n_35367), .o(FE_OCPN1639_n_35367) );
in01s01 FE_OCPC1641_FE_OCP_RBN1596_n_14823 ( .a(FE_OCP_RBN1596_n_14823), .o(FE_OCPN1641_FE_OCP_RBN1596_n_14823) );
in01s01 FE_OCPC1642_FE_OCP_RBN1596_n_14823 ( .a(FE_OCPN1641_FE_OCP_RBN1596_n_14823), .o(FE_OCPN1642_FE_OCP_RBN1596_n_14823) );
in01s01 FE_OCPC1643_n_16866 ( .a(n_16866), .o(FE_OCPN1643_n_16866) );
in01s01 FE_OCPC1644_n_16866 ( .a(FE_OCPN1643_n_16866), .o(FE_OCPN1644_n_16866) );
in01s01 FE_OCPC1645_n_18860 ( .a(FE_OCP_DRV_N5354_n_18860), .o(FE_OCPN1645_n_18860) );
in01s01 FE_OCPC1646_n_18860 ( .a(FE_OCPN1645_n_18860), .o(FE_OCPN1646_n_18860) );
in01s06 FE_OCPC1649_n_44734 ( .a(FE_OCP_RBN2412_n_44722), .o(FE_OCPN1649_n_44734) );
in01s06 FE_OCPC1650_n_11918 ( .a(n_11918), .o(FE_OCPN1650_n_11918) );
in01m06 FE_OCPC1651_n_11918 ( .a(FE_OCPN1650_n_11918), .o(FE_OCPN1651_n_11918) );
in01s10 FE_OCPC1652_n_23078 ( .a(n_23078), .o(FE_OCPN1652_n_23078) );
in01s10 FE_OCPC1653_n_23078 ( .a(FE_OCPN1652_n_23078), .o(FE_OCPN1653_n_23078) );
in01s01 FE_OCPC1655_n_12488 ( .a(FE_OCPN1658_n_12488), .o(FE_OCPN1655_n_12488) );
in01s02 FE_OCPC1656_n_12368 ( .a(n_12368), .o(FE_OCPN1656_n_12368) );
in01s06 FE_OCPC1657_n_12368 ( .a(FE_OCPN1656_n_12368), .o(FE_OCPN1657_n_12368) );
in01s02 FE_OCPC1658_n_12488 ( .a(n_12488), .o(FE_OCPN1658_n_12488) );
in01s02 FE_OCPC1659_n_12488 ( .a(FE_OCPN1658_n_12488), .o(FE_OCPN1659_n_12488) );
in01s01 FE_OCPC1660_n_37661 ( .a(n_37661), .o(FE_OCPN1660_n_37661) );
in01s01 FE_OCPC1661_n_37661 ( .a(FE_OCPN1660_n_37661), .o(FE_OCPN1661_n_37661) );
in01s01 FE_OCPC1662_n_4556 ( .a(n_4556), .o(FE_OCPN1662_n_4556) );
in01s02 FE_OCPC1663_n_4556 ( .a(FE_OCPN1662_n_4556), .o(FE_OCPN1663_n_4556) );
in01s01 FE_OCPC1664_FE_OCP_RBN1138_n_19270 ( .a(FE_OCP_RBN1138_n_19270), .o(FE_OCPN1664_FE_OCP_RBN1138_n_19270) );
in01s02 FE_OCPC1665_FE_OCP_RBN1138_n_19270 ( .a(FE_OCPN1664_FE_OCP_RBN1138_n_19270), .o(FE_OCPN1665_FE_OCP_RBN1138_n_19270) );
in01s01 FE_OCPC1666_n_39207 ( .a(n_39207), .o(FE_OCPN1666_n_39207) );
in01s01 FE_OCPC1667_n_39207 ( .a(FE_OCPN1666_n_39207), .o(FE_OCPN1667_n_39207) );
in01s02 FE_OCPC1668_n_23941 ( .a(n_23941), .o(FE_OCPN1668_n_23941) );
in01s01 FE_OCPC1669_n_23941 ( .a(FE_OCPN1668_n_23941), .o(FE_OCPN1669_n_23941) );
in01s01 FE_OCPC1670_n_39371 ( .a(n_39371), .o(FE_OCPN1670_n_39371) );
in01s01 FE_OCPC1671_n_39371 ( .a(FE_OCPN1670_n_39371), .o(FE_OCPN1671_n_39371) );
in01s01 FE_OCPC1672_n_14055 ( .a(n_14055), .o(FE_OCPN1672_n_14055) );
in01s01 FE_OCPC1674_n_25721 ( .a(n_25721), .o(FE_OCPN1674_n_25721) );
in01s01 FE_OCPC1675_n_25721 ( .a(FE_OCPN1674_n_25721), .o(FE_OCPN1675_n_25721) );
in01s01 FE_OCPC1676_n_27062 ( .a(n_27062), .o(FE_OCPN1676_n_27062) );
in01s01 FE_OCPC1677_n_27062 ( .a(FE_OCPN1676_n_27062), .o(FE_OCPN1677_n_27062) );
in01s01 FE_OCPC1679_n_27315 ( .a(FE_OCPN1762_n_30708), .o(FE_OCPN1679_n_27315) );
in01s01 FE_OCPC1680_n_30614 ( .a(n_30614), .o(FE_OCPN1680_n_30614) );
in01s02 FE_OCPC1681_n_30614 ( .a(FE_OCPN1680_n_30614), .o(FE_OCPN1681_n_30614) );
in01s01 FE_OCPC1682_n_27210 ( .a(n_27210), .o(FE_OCPN1682_n_27210) );
in01s01 FE_OCPC1683_n_27210 ( .a(FE_OCPN1682_n_27210), .o(FE_OCPN1683_n_27210) );
in01s01 FE_OCPC1684_n_14555 ( .a(n_14555), .o(FE_OCPN1684_n_14555) );
in01s01 FE_OCPC1685_n_14555 ( .a(FE_OCPN1684_n_14555), .o(FE_OCPN1685_n_14555) );
in01s06 FE_OCPC1686_n_23097 ( .a(n_23097), .o(FE_OCPN1686_n_23097) );
in01s06 FE_OCPC1687_n_23097 ( .a(FE_OCPN1686_n_23097), .o(FE_OCPN1687_n_23097) );
in01s06 FE_OCPC1688_n_23167 ( .a(n_23167), .o(FE_OCPN1688_n_23167) );
in01s06 FE_OCPC1689_n_23167 ( .a(FE_OCPN1688_n_23167), .o(FE_OCPN1689_n_23167) );
in01s01 FE_OCPC1690_n_10105 ( .a(n_10105), .o(FE_OCPN1690_n_10105) );
in01s01 FE_OCPC1692_n_33140 ( .a(n_33140), .o(FE_OCPN1692_n_33140) );
in01s01 FE_OCPC1693_n_33140 ( .a(FE_OCPN1692_n_33140), .o(FE_OCPN1693_n_33140) );
in01s01 FE_OCPC1694_n_12836 ( .a(n_12836), .o(FE_OCPN1694_n_12836) );
in01s02 FE_OCPC1695_n_12836 ( .a(FE_OCPN1694_n_12836), .o(FE_OCPN1695_n_12836) );
in01s01 FE_OCPC1696_n_13721 ( .a(n_13721), .o(FE_OCPN1696_n_13721) );
in01s01 FE_OCPC1698_n_34118 ( .a(n_34118), .o(FE_OCPN1698_n_34118) );
in01s01 FE_OCPC1699_n_34118 ( .a(FE_OCPN1698_n_34118), .o(FE_OCPN1699_n_34118) );
in01s01 FE_OCPC1700_n_33544 ( .a(n_33544), .o(FE_OCPN1700_n_33544) );
in01s01 FE_OCPC1701_n_33544 ( .a(FE_OCPN1700_n_33544), .o(FE_OCPN1701_n_33544) );
in01s01 FE_OCPC1702_n_14210 ( .a(FE_OCP_RBN5801_n_13962), .o(FE_OCPN1702_n_14210) );
in01s01 FE_OCPC1703_n_14210 ( .a(FE_OCPN1702_n_14210), .o(FE_OCPN1703_n_14210) );
in01m01 FE_OCPC1704_n_14730 ( .a(n_14730), .o(FE_OCPN1704_n_14730) );
in01s06 FE_OCPC1705_n_14730 ( .a(FE_OCPN1704_n_14730), .o(FE_OCPN1705_n_14730) );
in01s01 FE_OCPC1706_n_21229 ( .a(n_21229), .o(FE_OCPN1706_n_21229) );
in01s01 FE_OCPC1707_n_21229 ( .a(FE_OCPN1706_n_21229), .o(FE_OCPN1707_n_21229) );
in01s01 FE_OCPC1708_FE_OFN739_n_17093 ( .a(FE_OFN739_n_17093), .o(FE_OCPN1708_FE_OFN739_n_17093) );
in01s01 FE_OCPC1709_FE_OFN739_n_17093 ( .a(FE_OCPN1708_FE_OFN739_n_17093), .o(FE_OCPN1709_FE_OFN739_n_17093) );
in01s01 FE_OCPC1710_n_45073 ( .a(n_45073), .o(FE_OCPN1710_n_45073) );
in01s01 FE_OCPC1711_n_45073 ( .a(FE_OCPN1710_n_45073), .o(FE_OCPN1711_n_45073) );
in01s01 FE_OCPC1712_n_42306 ( .a(n_42306), .o(FE_OCPN1712_n_42306) );
in01s01 FE_OCPC1713_n_42306 ( .a(FE_OCPN1712_n_42306), .o(FE_OCPN1713_n_42306) );
in01s02 FE_OCPC1714_n_43449 ( .a(n_43449), .o(FE_OCPN1714_n_43449) );
in01s02 FE_OCPC1715_n_43449 ( .a(FE_OCPN1714_n_43449), .o(FE_OCPN1715_n_43449) );
in01m01 FE_OCPC1716_n_12311 ( .a(n_12311), .o(FE_OCPN1716_n_12311) );
in01m03 FE_OCPC1717_n_12311 ( .a(FE_OCPN1716_n_12311), .o(FE_OCPN1717_n_12311) );
in01s08 FE_OCPC1718_n_28065 ( .a(n_28065), .o(FE_OCPN1718_n_28065) );
in01s01 FE_OCPC1721_n_23818 ( .a(n_23819), .o(FE_OCPN1721_n_23818) );
in01s01 FE_OCPC1722_n_29060 ( .a(n_29060), .o(FE_OCPN1722_n_29060) );
in01s01 FE_OCPC1725_n_33136 ( .a(n_33137), .o(FE_OCPN1725_n_33136) );
in01s01 FE_OCPC1726_n_18099 ( .a(n_18099), .o(FE_OCPN1726_n_18099) );
in01s01 FE_OCPC1727_n_18099 ( .a(FE_OCPN1726_n_18099), .o(FE_OCPN1727_n_18099) );
in01s01 FE_OCPC1728_n_34096 ( .a(FE_OCP_DRV_N6907_n_34096), .o(FE_OCPN1728_n_34096) );
in01s02 FE_OCPC1732_n_14524 ( .a(n_14524), .o(FE_OCPN1732_n_14524) );
in01s06 FE_OCPC1733_n_14524 ( .a(FE_OCPN1732_n_14524), .o(FE_OCPN1733_n_14524) );
in01s01 FE_OCPC1736_n_27009 ( .a(n_27009), .o(FE_OCPN1736_n_27009) );
in01s01 FE_OCPC1737_n_27009 ( .a(FE_OCPN1736_n_27009), .o(FE_OCPN1737_n_27009) );
in01s01 FE_OCPC1738_n_33968 ( .a(n_33968), .o(FE_OCPN1738_n_33968) );
in01s01 FE_OCPC1739_n_33968 ( .a(FE_OCPN1738_n_33968), .o(FE_OCPN1739_n_33968) );
in01s01 FE_OCPC1740_n_18591 ( .a(n_18591), .o(FE_OCPN1740_n_18591) );
in01s01 FE_OCPC1741_n_18591 ( .a(FE_OCPN1740_n_18591), .o(FE_OCPN1741_n_18591) );
in01s01 FE_OCPC1762_n_30708 ( .a(n_27315), .o(FE_OCPN1762_n_30708) );
in01s01 FE_OCPC1763_n_30708 ( .a(FE_OCPN1762_n_30708), .o(FE_OCPN1763_n_30708) );
in01s10 FE_OCPC1902_n_32712 ( .a(FE_OCP_RBN6520_n_32706), .o(FE_OCPN1902_n_32712) );
in01s01 FE_OCPC1903_n_32554 ( .a(n_32554), .o(FE_OCPN1903_n_32554) );
in01s01 FE_OCPC1904_n_32554 ( .a(FE_OCPN1903_n_32554), .o(FE_OCPN1904_n_32554) );
in01s10 FE_OCPC1905_n_23322 ( .a(n_23322), .o(FE_OCPN1905_n_23322) );
in01s10 FE_OCPC1906_n_23322 ( .a(FE_OCPN1905_n_23322), .o(FE_OCPN1906_n_23322) );
in01s01 FE_OCPC1907_n_17921 ( .a(n_17921), .o(FE_OCPN1907_n_17921) );
in01s01 FE_OCPC1908_n_17921 ( .a(FE_OCPN1907_n_17921), .o(FE_OCPN1908_n_17921) );
in01s01 FE_OCPC1909_n_40921 ( .a(n_40921), .o(FE_OCPN1909_n_40921) );
in01s01 FE_OCPC1910_n_40921 ( .a(FE_OCPN1909_n_40921), .o(FE_OCPN1910_n_40921) );
in01s01 FE_OCPC1911_n_33907 ( .a(n_33907), .o(FE_OCPN1911_n_33907) );
in01s01 FE_OCPC1912_n_33907 ( .a(FE_OCPN1911_n_33907), .o(FE_OCPN1912_n_33907) );
in01s01 FE_OCPC1915_n_22111 ( .a(n_22111), .o(FE_OCPN1915_n_22111) );
in01s06 FE_OCPC1916_n_22111 ( .a(FE_OCPN1915_n_22111), .o(FE_OCPN1916_n_22111) );
in01s01 FE_OCPC1917_n_29571 ( .a(n_29571), .o(FE_OCPN1917_n_29571) );
in01s01 FE_OCPC1918_n_29571 ( .a(FE_OCPN1917_n_29571), .o(FE_OCPN1918_n_29571) );
in01s01 FE_OCPC1919_n_22393 ( .a(n_22393), .o(FE_OCPN1919_n_22393) );
in01s06 FE_OCPC1920_n_22393 ( .a(FE_OCPN1919_n_22393), .o(FE_OCPN1920_n_22393) );
in01s01 FE_OCPC1921_n_24962 ( .a(FE_OCPUNCON3472_n_24962), .o(FE_OCPN1921_n_24962) );
in01s01 FE_OCPC1922_n_24962 ( .a(FE_OCPN1921_n_24962), .o(FE_OCPN1922_n_24962) );
in01s01 FE_OCPC1923_n_20430 ( .a(n_20430), .o(FE_OCPN1923_n_20430) );
in01s01 FE_OCPC1924_n_20430 ( .a(FE_OCPN1923_n_20430), .o(FE_OCPN1924_n_20430) );
in01s01 FE_OCPC1925_n_34516 ( .a(n_34516), .o(FE_OCPN1925_n_34516) );
in01s01 FE_OCPC1926_n_34516 ( .a(FE_OCPN1925_n_34516), .o(FE_OCPN1926_n_34516) );
in01s01 FE_OCPC1927_n_30385 ( .a(n_30385), .o(FE_OCPN1927_n_30385) );
in01s01 FE_OCPC1928_n_30385 ( .a(FE_OCPN1927_n_30385), .o(FE_OCPN1928_n_30385) );
in01s01 FE_OCPC1932_n_9114 ( .a(n_9197), .o(FE_OCPN1932_n_9114) );
in01s01 FE_OCPC1933_n_26801 ( .a(FE_OCP_DRV_N5159_n_26801), .o(FE_OCPN1933_n_26801) );
in01s01 FE_OCPC1934_n_26801 ( .a(FE_OCPN1933_n_26801), .o(FE_OCPN1934_n_26801) );
in01s01 FE_OCPC1935_n_31676 ( .a(n_31676), .o(FE_OCPN1935_n_31676) );
in01s01 FE_OCPC1936_n_31676 ( .a(FE_OCPN1935_n_31676), .o(FE_OCPN1936_n_31676) );
in01s01 FE_OCPC1937_n_31719 ( .a(n_31719), .o(FE_OCPN1937_n_31719) );
in01s01 FE_OCPC1938_n_31719 ( .a(FE_OCPN1937_n_31719), .o(FE_OCPN1938_n_31719) );
in01s01 FE_OCPC1939_delay_sub_ln23_0_unr23_stage8_stallmux_q ( .a(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(FE_OCPN1939_delay_sub_ln23_0_unr23_stage8_stallmux_q) );
in01s01 FE_OCPC1940_delay_sub_ln23_0_unr23_stage8_stallmux_q ( .a(FE_OCPN1939_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(FE_OCPN1940_delay_sub_ln23_0_unr23_stage8_stallmux_q) );
in01s01 FE_OCPC1941_n_20723 ( .a(n_20723), .o(FE_OCPN1941_n_20723) );
in01s01 FE_OCPC1942_n_20723 ( .a(FE_OCPN1941_n_20723), .o(FE_OCPN1942_n_20723) );
in01s01 FE_OCPC1946_delay_sub_ln23_0_unr23_stage8_stallmux_q ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(FE_OCPN1946_delay_sub_ln23_0_unr23_stage8_stallmux_q) );
in01s01 FE_OCPC1947_delay_sub_ln23_0_unr23_stage8_stallmux_q ( .a(FE_OCPN1946_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(FE_OCPN1947_delay_sub_ln23_0_unr23_stage8_stallmux_q) );
in01s01 FE_OCPC1949_delay_sub_ln23_0_unr23_stage8_stallmux_q ( .a(FE_OCPN1947_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(FE_OCPN1949_delay_sub_ln23_0_unr23_stage8_stallmux_q) );
in01s01 FE_OCPC1950_delay_sub_ln23_0_unr23_stage8_stallmux_q ( .a(FE_OCPN1949_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(FE_OCPN1950_delay_sub_ln23_0_unr23_stage8_stallmux_q) );
in01s06 FE_OCPC1951_delay_sub_ln23_0_unr23_stage8_stallmux_q ( .a(FE_OCPN1949_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q) );
in01s01 FE_OCPC1952_n_36121 ( .a(n_36121), .o(FE_OCPN1952_n_36121) );
in01s01 FE_OCPC1953_n_36121 ( .a(FE_OCPN1952_n_36121), .o(FE_OCPN1953_n_36121) );
in01s01 FE_OCPC1955_n_36050 ( .a(n_36119), .o(FE_OCPN1955_n_36050) );
in01s01 FE_OCPC3529_n_28829 ( .a(FE_OCP_DRV_N6884_n_28829), .o(FE_OCPN3529_n_28829) );
in01s01 FE_OCPC3531_n_26468 ( .a(n_26468), .o(FE_OCPN3531_n_26468) );
in01s03 FE_OCPC3541_n_32436 ( .a(n_32436), .o(FE_OCPN3541_n_32436) );
in01m03 FE_OCPC3542_n_32436 ( .a(FE_OCPN3541_n_32436), .o(FE_OCPN3542_n_32436) );
in01s01 FE_OCPC3543_n_1448 ( .a(n_1448), .o(FE_OCPN3543_n_1448) );
in01s01 FE_OCPC3544_n_1448 ( .a(FE_OCPN3543_n_1448), .o(FE_OCPN3544_n_1448) );
in01s02 FE_OCPC3545_n_1705 ( .a(n_1705), .o(FE_OCPN3545_n_1705) );
in01s02 FE_OCPC3546_n_1705 ( .a(FE_OCPN3545_n_1705), .o(FE_OCPN3546_n_1705) );
in01s06 FE_OCPC3547_n_28043 ( .a(n_28043), .o(FE_OCPN3547_n_28043) );
in01s06 FE_OCPC3548_n_28043 ( .a(FE_OCPN3547_n_28043), .o(FE_OCPN3548_n_28043) );
in01m08 FE_OCPC3549_n_28381 ( .a(n_28381), .o(FE_OCPN3549_n_28381) );
in01m10 FE_OCPC3550_n_28381 ( .a(FE_OCPN3549_n_28381), .o(FE_OCPN3550_n_28381) );
in01s02 FE_OCPC3551_n_33225 ( .a(n_33225), .o(FE_OCPN3551_n_33225) );
in01s04 FE_OCPC3552_n_33225 ( .a(FE_OCPN3551_n_33225), .o(FE_OCPN3552_n_33225) );
in01s01 FE_OCPC3553_n_12671 ( .a(n_12671), .o(FE_OCPN3553_n_12671) );
in01s02 FE_OCPC3554_n_12671 ( .a(FE_OCPN3553_n_12671), .o(FE_OCPN3554_n_12671) );
in01s01 FE_OCPC3555_n_40986 ( .a(n_40986), .o(FE_OCPN3555_n_40986) );
in01s01 FE_OCPC3556_n_40986 ( .a(FE_OCPN3555_n_40986), .o(FE_OCPN3556_n_40986) );
in01s01 FE_OCPC3557_n_7673 ( .a(n_7673), .o(FE_OCPN3557_n_7673) );
in01s01 FE_OCPC3559_n_2386 ( .a(n_2386), .o(FE_OCPN3559_n_2386) );
in01s01 FE_OCPC3560_n_2386 ( .a(FE_OCPN3559_n_2386), .o(FE_OCPN3560_n_2386) );
in01s01 FE_OCPC3561_n_3317 ( .a(n_3317), .o(FE_OCPN3561_n_3317) );
in01s01 FE_OCPC3562_n_3317 ( .a(FE_OCPN3561_n_3317), .o(FE_OCPN3562_n_3317) );
in01s01 FE_OCPC3563_n_38731 ( .a(n_38731), .o(FE_OCPN3563_n_38731) );
in01s01 FE_OCPC3564_n_38731 ( .a(FE_OCPN3563_n_38731), .o(FE_OCPN3564_n_38731) );
in01s01 FE_OCPC3565_n_10214 ( .a(n_10214), .o(FE_OCPN3565_n_10214) );
in01s01 FE_OCPC3567_n_8348 ( .a(n_8348), .o(FE_OCPN3567_n_8348) );
in01s01 FE_OCPC3568_n_8348 ( .a(FE_OCPN3567_n_8348), .o(FE_OCPN3568_n_8348) );
in01s01 FE_OCPC3569_n_19303 ( .a(FE_OCP_RBN3714_n_19241), .o(FE_OCPN3569_n_19303) );
in01s01 FE_OCPC3570_n_19303 ( .a(FE_OCPN3569_n_19303), .o(FE_OCPN3570_n_19303) );
in01s02 FE_OCPC3571_n_4374 ( .a(n_4374), .o(FE_OCPN3571_n_4374) );
in01s02 FE_OCPC3572_n_4374 ( .a(FE_OCPN3571_n_4374), .o(FE_OCPN3572_n_4374) );
in01s01 FE_OCPC3573_n_30345 ( .a(n_30345), .o(FE_OCPN3573_n_30345) );
in01s01 FE_OCPC3574_n_30345 ( .a(FE_OCPN3573_n_30345), .o(FE_OCPN3574_n_30345) );
in01s01 FE_OCPC3575_n_3625 ( .a(FE_OCP_RBN5852_n_3625), .o(FE_OCPN3575_n_3625) );
in01s01 FE_OCPC3576_n_3625 ( .a(FE_OCPN3575_n_3625), .o(FE_OCPN3576_n_3625) );
in01s01 FE_OCPC3577_n_23354 ( .a(FE_RN_1793_0), .o(FE_OCPN3577_n_23354) );
in01s02 FE_OCPC3578_n_23354 ( .a(FE_OCPN3577_n_23354), .o(FE_OCPN3578_n_23354) );
in01s01 FE_OCPC3579_n_25370 ( .a(n_25370), .o(FE_OCPN3579_n_25370) );
in01s01 FE_OCPC3580_n_25370 ( .a(FE_OCPN3579_n_25370), .o(FE_OCPN3580_n_25370) );
in01s01 FE_OCPC3581_n_39747 ( .a(n_39747), .o(FE_OCPN3581_n_39747) );
in01s01 FE_OCPC3582_n_39747 ( .a(FE_OCPN3581_n_39747), .o(FE_OCPN3582_n_39747) );
in01s01 FE_OCPC3583_n_4556 ( .a(FE_OCPN1663_n_4556), .o(FE_OCPN3583_n_4556) );
in01s02 FE_OCPC3584_n_4556 ( .a(FE_OCPN3583_n_4556), .o(FE_OCPN3584_n_4556) );
in01s01 FE_OCPC3585_n_31704 ( .a(n_31704), .o(FE_OCPN3585_n_31704) );
in01s02 FE_OCPC3586_n_31704 ( .a(FE_OCPN3585_n_31704), .o(FE_OCPN3586_n_31704) );
in01s01 FE_OCPC3589_n_21419 ( .a(n_21419), .o(FE_OCPN3589_n_21419) );
in01s01 FE_OCPC3592_n_45301 ( .a(n_45300), .o(FE_OCPN3592_n_45301) );
in01s01 FE_OCPC4514_n_21343 ( .a(n_21343), .o(FE_OCPN4514_n_21343) );
in01s01 FE_OCPC4515_n_21343 ( .a(FE_OCPN4514_n_21343), .o(FE_OCPN4515_n_21343) );
in01s20 FE_OCPC4519_n_32820 ( .a(n_32820), .o(FE_OCPN4519_n_32820) );
in01s20 FE_OCPC4520_n_32820 ( .a(FE_OCPN4519_n_32820), .o(FE_OCPN4520_n_32820) );
in01m02 FE_OCPC4521_n_13015 ( .a(n_13015), .o(FE_OCPN4521_n_13015) );
in01s04 FE_OCPC4522_n_13015 ( .a(FE_OCPN4521_n_13015), .o(FE_OCPN4522_n_13015) );
in01s01 FE_OCPC4523_n_7360 ( .a(n_7360), .o(FE_OCPN4523_n_7360) );
in01s02 FE_OCPC4524_n_7360 ( .a(FE_OCPN4523_n_7360), .o(FE_OCPN4524_n_7360) );
in01s01 FE_OCPC4525_n_8099 ( .a(n_8099), .o(FE_OCPN4525_n_8099) );
in01s01 FE_OCPC4526_n_8099 ( .a(FE_OCPN4525_n_8099), .o(FE_OCPN4526_n_8099) );
in01s01 FE_OCPC4527_n_18117 ( .a(n_18117), .o(FE_OCPN4527_n_18117) );
in01s02 FE_OCPC4528_n_18117 ( .a(FE_OCPN4527_n_18117), .o(FE_OCPN4528_n_18117) );
in01s01 FE_OCPC4529_FE_OCP_RBN2748_n_8474 ( .a(FE_OCP_RBN2748_n_8474), .o(FE_OCPN4529_FE_OCP_RBN2748_n_8474) );
in01s01 FE_OCPC4532_n_3319 ( .a(n_3319), .o(FE_OCPN4532_n_3319) );
in01s01 FE_OCPC4533_n_3319 ( .a(FE_OCPN4532_n_3319), .o(FE_OCPN4533_n_3319) );
in01s01 FE_OCPC4534_n_9012 ( .a(n_9012), .o(FE_OCPN4534_n_9012) );
in01s01 FE_OCPC4535_n_9012 ( .a(FE_OCPN4534_n_9012), .o(FE_OCPN4535_n_9012) );
in01s01 FE_OCPC4536_n_14543 ( .a(n_14543), .o(FE_OCPN4536_n_14543) );
in01s01 FE_OCPC4538_n_20332 ( .a(n_20332), .o(FE_OCPN4538_n_20332) );
in01s01 FE_OCPC4539_n_20332 ( .a(FE_OCPN4538_n_20332), .o(FE_OCPN4539_n_20332) );
in01s01 FE_OCPC4542_FE_OCP_RBN2812_n_8835 ( .a(FE_OCP_RBN2812_n_8835), .o(FE_OCPN4542_FE_OCP_RBN2812_n_8835) );
in01s01 FE_OCPC4544_FE_OCP_RBN2850_n_3645 ( .a(FE_OCP_RBN2850_n_3645), .o(FE_OCPN4544_FE_OCP_RBN2850_n_3645) );
in01s01 FE_OCPC4545_FE_OCP_RBN2850_n_3645 ( .a(FE_OCPN4544_FE_OCP_RBN2850_n_3645), .o(FE_OCPN4545_FE_OCP_RBN2850_n_3645) );
in01s02 FE_OCPC4546_n_4727 ( .a(n_4727), .o(FE_OCPN4546_n_4727) );
in01s02 FE_OCPC4547_n_4727 ( .a(FE_OCPN4546_n_4727), .o(FE_OCPN4547_n_4727) );
in01s01 FE_OCPC4548_FE_OCP_RBN3086_n_10015 ( .a(FE_OCP_RBN3086_n_10015), .o(FE_OCPN4548_FE_OCP_RBN3086_n_10015) );
in01s01 FE_OCPC4549_FE_OCP_RBN3086_n_10015 ( .a(FE_OCPN4548_FE_OCP_RBN3086_n_10015), .o(FE_OCPN4549_FE_OCP_RBN3086_n_10015) );
in01s01 FE_OCPC4550_n_10545 ( .a(n_10545), .o(FE_OCPN4550_n_10545) );
in01s01 FE_OCPC4551_n_10545 ( .a(FE_OCPN4550_n_10545), .o(FE_OCPN4551_n_10545) );
in01s02 FE_OCPC4827_FE_OCP_RBN4275_n_3700 ( .a(FE_OCP_RBN5872_n_3700), .o(FE_OCPN4827_FE_OCP_RBN4275_n_3700) );
in01s04 FE_OCPC4828_FE_OCP_RBN4275_n_3700 ( .a(FE_OCPN4827_FE_OCP_RBN4275_n_3700), .o(FE_OCPN4828_FE_OCP_RBN4275_n_3700) );
in01s01 FE_OCPC4829_n_5603 ( .a(n_5603), .o(FE_OCPN4829_n_5603) );
in01s01 FE_OCPC4830_n_5603 ( .a(FE_OCPN4829_n_5603), .o(FE_OCPN4830_n_5603) );
in01s01 FE_OCPC4831_n_22294 ( .a(n_22294), .o(FE_OCPN4831_n_22294) );
in01s01 FE_OCPC4832_n_22294 ( .a(FE_OCPN4831_n_22294), .o(FE_OCPN4832_n_22294) );
in01s02 FE_OCPC4833_n_32863 ( .a(n_32863), .o(FE_OCPN4833_n_32863) );
in01s01 FE_OCPC4835_n_36034 ( .a(n_36034), .o(FE_OCPN4835_n_36034) );
in01s01 FE_OCPC4836_n_36034 ( .a(FE_OCPN4835_n_36034), .o(FE_OCPN4836_n_36034) );
in01s01 FE_OCPC4843_FE_OFN4779_n_44490 ( .a(FE_OFN4779_n_44490), .o(FE_OCPN4843_FE_OFN4779_n_44490) );
in01s01 FE_OCPC4844_FE_OFN4779_n_44490 ( .a(FE_OCPN4843_FE_OFN4779_n_44490), .o(FE_OCPN4844_FE_OFN4779_n_44490) );
in01m03 FE_OCPC4845_FE_OFN4779_n_44490 ( .a(FE_OCPN4843_FE_OFN4779_n_44490), .o(FE_OCPN4845_FE_OFN4779_n_44490) );
in01s01 FE_OCPC4846_FE_OFN4778_n_44490 ( .a(FE_OFN4778_n_44490), .o(FE_OCPN4846_FE_OFN4778_n_44490) );
in01s02 FE_OCPC4847_FE_OFN4778_n_44490 ( .a(FE_OCPN4846_FE_OFN4778_n_44490), .o(FE_OCPN4847_FE_OFN4778_n_44490) );
in01s01 FE_OCPC4848_n_28460 ( .a(n_28460), .o(FE_OCPN4848_n_28460) );
in01s01 FE_OCPC4849_n_28460 ( .a(FE_OCPN4848_n_28460), .o(FE_OCPN4849_n_28460) );
in01s01 FE_OCPC4850_n_47235 ( .a(n_47235), .o(FE_OCPN4850_n_47235) );
in01s01 FE_OCPC4851_n_47235 ( .a(FE_OCPN4850_n_47235), .o(FE_OCPN4851_n_47235) );
in01s01 FE_OCPC4852_n_29502 ( .a(n_29502), .o(FE_OCPN4852_n_29502) );
in01s01 FE_OCPC4853_n_29502 ( .a(FE_OCPN4852_n_29502), .o(FE_OCPN4853_n_29502) );
in01s01 FE_OCPC4854_n_34369 ( .a(n_34297), .o(FE_OCPN4854_n_34369) );
in01s01 FE_OCPC4855_n_34369 ( .a(FE_OCPN4854_n_34369), .o(FE_OCPN4855_n_34369) );
in01s01 FE_OCPC4856_n_14317 ( .a(n_14317), .o(FE_OCPN4856_n_14317) );
in01s01 FE_OCPC4857_n_14317 ( .a(FE_OCPN4856_n_14317), .o(FE_OCPN4857_n_14317) );
in01s01 FE_OCPC4858_n_10369 ( .a(n_10369), .o(FE_OCPN4858_n_10369) );
in01s01 FE_OCPC4859_n_10369 ( .a(FE_OCPN4858_n_10369), .o(FE_OCPN4859_n_10369) );
in01s01 FE_OCPC4926_n_1452 ( .a(n_1452), .o(FE_OCPN4926_n_1452) );
in01s01 FE_OCPC4927_n_1452 ( .a(FE_OCPN4926_n_1452), .o(FE_OCPN4927_n_1452) );
in01s01 FE_OCPC4928_n_16143 ( .a(n_16143), .o(FE_OCPN4928_n_16143) );
in01s01 FE_OCPC4929_n_16143 ( .a(FE_OCPN4928_n_16143), .o(FE_OCPN4929_n_16143) );
in01s01 FE_OCPC4930_n_20275 ( .a(n_20275), .o(FE_OCPN4930_n_20275) );
in01s02 FE_OCPC4931_n_20275 ( .a(FE_OCPN4930_n_20275), .o(FE_OCPN4931_n_20275) );
in01s01 FE_OCPC4932_n_47023 ( .a(n_47023), .o(FE_OCPN4932_n_47023) );
in01s01 FE_OCPC4933_n_47023 ( .a(FE_OCPN4932_n_47023), .o(FE_OCPN4933_n_47023) );
in01s06 FE_OCPC4934_n_11993 ( .a(n_11993), .o(FE_OCPN4934_n_11993) );
in01s10 FE_OCPC4935_n_11993 ( .a(FE_OCPN4934_n_11993), .o(FE_OCPN4935_n_11993) );
in01s01 FE_OCPC4936_n_13570 ( .a(n_13570), .o(FE_OCPN4936_n_13570) );
in01s01 FE_OCPC4937_n_13570 ( .a(FE_OCPN4936_n_13570), .o(FE_OCPN4937_n_13570) );
in01s01 FE_OCPC5094_n_679 ( .a(n_679), .o(FE_OCPN5094_n_679) );
in01s01 FE_OCPC5095_n_679 ( .a(FE_OCPN5094_n_679), .o(FE_OCPN5095_n_679) );
in01s01 FE_OCPC5096_n_694 ( .a(n_694), .o(FE_OCPN5096_n_694) );
in01s01 FE_OCPC5097_n_694 ( .a(FE_OCPN5096_n_694), .o(FE_OCPN5097_n_694) );
in01s01 FE_OCPC5098_n_1282 ( .a(n_1282), .o(FE_OCPN5098_n_1282) );
in01s01 FE_OCPC5099_n_1282 ( .a(FE_OCPN5098_n_1282), .o(FE_OCPN5099_n_1282) );
in01s01 FE_OCPC5100_n_18918 ( .a(n_18918), .o(FE_OCPN5100_n_18918) );
in01s01 FE_OCPC5101_n_18918 ( .a(FE_OCPN5100_n_18918), .o(FE_OCPN5101_n_18918) );
in01s01 FE_OCPC5102_FE_OCP_RBN5029_n_18678 ( .a(FE_OCP_RBN5029_n_18678), .o(FE_OCPN5102_FE_OCP_RBN5029_n_18678) );
in01s01 FE_OCPC5104_n_30371 ( .a(n_30371), .o(FE_OCPN5104_n_30371) );
in01s01 FE_OCPC5105_n_30371 ( .a(FE_OCPN5104_n_30371), .o(FE_OCPN5105_n_30371) );
in01s01 FE_OCPC5106_n_31804 ( .a(n_31804), .o(FE_OCPN5106_n_31804) );
in01s01 FE_OCPC5107_n_31804 ( .a(FE_OCPN5106_n_31804), .o(FE_OCPN5107_n_31804) );
in01s01 FE_OCPC5108_n_29715 ( .a(n_29715), .o(FE_OCPN5108_n_29715) );
in01s01 FE_OCPC5109_n_29715 ( .a(FE_OCPN5108_n_29715), .o(FE_OCPN5109_n_29715) );
in01s01 FE_OCPC5110_n_25973 ( .a(n_25973), .o(FE_OCPN5110_n_25973) );
in01s01 FE_OCPC5111_n_25973 ( .a(FE_OCPN5110_n_25973), .o(FE_OCPN5111_n_25973) );
in01m10 FE_OCPC5112_n_22249 ( .a(n_22249), .o(FE_OCPN5112_n_22249) );
in01s06 FE_OCPC5113_n_22249 ( .a(FE_OCPN5112_n_22249), .o(FE_OCPN5113_n_22249) );
in01s10 FE_OCPC5114_n_22249 ( .a(FE_OCPN5112_n_22249), .o(FE_OCPN5114_n_22249) );
in01s01 FE_OCPC5119_n_25595 ( .a(n_25595), .o(FE_OCPN5119_n_25595) );
in01s01 FE_OCPC5120_n_25595 ( .a(FE_OCPN5119_n_25595), .o(FE_OCPN5120_n_25595) );
in01s01 FE_OCPC5121_n_44438 ( .a(n_44438), .o(FE_OCPN5121_n_44438) );
in01s01 FE_OCPC5122_n_44438 ( .a(FE_OCPN5121_n_44438), .o(FE_OCPN5122_n_44438) );
in01s01 FE_OCPC5123_n_31197 ( .a(n_31197), .o(FE_OCPN5123_n_31197) );
in01s01 FE_OCPC5124_n_31197 ( .a(FE_OCPN5123_n_31197), .o(FE_OCPN5124_n_31197) );
in01s01 FE_OCPC5125_n_16111 ( .a(n_16111), .o(FE_OCPN5125_n_16111) );
in01s01 FE_OCPC5126_n_16111 ( .a(FE_OCPN5125_n_16111), .o(FE_OCPN5126_n_16111) );
in01s02 FE_OCPC5127_n_22280 ( .a(n_22280), .o(FE_OCPN5127_n_22280) );
in01s02 FE_OCPC5128_n_22280 ( .a(FE_OCPN5127_n_22280), .o(FE_OCPN5128_n_22280) );
in01s01 FE_OCPC5129_FE_OFN1198_n_27014 ( .a(FE_OFN1198_n_27014), .o(FE_OCPN5129_FE_OFN1198_n_27014) );
in01s02 FE_OCPC5130_FE_OFN1198_n_27014 ( .a(FE_OCPN5129_FE_OFN1198_n_27014), .o(FE_OCPN5130_FE_OFN1198_n_27014) );
in01s01 FE_OCPC5131_n_29081 ( .a(n_29081), .o(FE_OCPN5131_n_29081) );
in01s01 FE_OCPC5132_n_29081 ( .a(FE_OCPN5131_n_29081), .o(FE_OCPN5132_n_29081) );
in01s01 FE_OCPC5133_n_27667 ( .a(n_27667), .o(FE_OCPN5133_n_27667) );
in01s01 FE_OCPC5134_n_27667 ( .a(FE_OCPN5133_n_27667), .o(FE_OCPN5134_n_27667) );
in01s01 FE_OCPC5135_n_12795 ( .a(n_12795), .o(FE_OCPN5135_n_12795) );
in01s01 FE_OCPC5136_n_12795 ( .a(FE_OCPN5135_n_12795), .o(FE_OCPN5136_n_12795) );
in01s01 FE_OCPC5219_n_10300 ( .a(n_10300), .o(FE_OCPN5219_n_10300) );
in01s01 FE_OCPC5221_FE_OFN753_n_13889 ( .a(FE_OFN753_n_13889), .o(FE_OCPN5221_FE_OFN753_n_13889) );
in01s01 FE_OCPC5222_FE_OFN753_n_13889 ( .a(FE_OCPN5221_FE_OFN753_n_13889), .o(FE_OCPN5222_FE_OFN753_n_13889) );
in01s01 FE_OCPC5223_n_10357 ( .a(n_10357), .o(FE_OCPN5223_n_10357) );
in01s01 FE_OCPC5225_n_25509 ( .a(n_25509), .o(FE_OCPN5225_n_25509) );
in01s01 FE_OCPC5226_n_25509 ( .a(FE_OCPN5225_n_25509), .o(FE_OCPN5226_n_25509) );
in01s01 FE_OCPC5227_n_33917 ( .a(n_33917), .o(FE_OCPN5227_n_33917) );
in01s01 FE_OCPC5228_n_33917 ( .a(FE_OCPN5227_n_33917), .o(FE_OCPN5228_n_33917) );
in01s01 FE_OCPC5229_n_30587 ( .a(n_30587), .o(FE_OCPN5229_n_30587) );
in01s01 FE_OCPC5230_n_30587 ( .a(FE_OCPN5229_n_30587), .o(FE_OCPN5230_n_30587) );
in01s01 FE_OCPC5231_n_35594 ( .a(n_35594), .o(FE_OCPN5231_n_35594) );
in01s01 FE_OCPC5233_n_27018 ( .a(n_27018), .o(FE_OCPN5233_n_27018) );
in01s01 FE_OCPC5234_n_27018 ( .a(FE_OCPN5233_n_27018), .o(FE_OCPN5234_n_27018) );
in01s01 FE_OCPC5235_n_44162 ( .a(n_44162), .o(FE_OCPN5235_n_44162) );
in01s01 FE_OCPC5237_n_22383 ( .a(n_22383), .o(FE_OCPN5237_n_22383) );
in01s02 FE_OCPC5238_n_22383 ( .a(FE_OCPN5237_n_22383), .o(FE_OCPN5238_n_22383) );
in01s01 FE_OCPC5239_n_26428 ( .a(n_26428), .o(FE_OCPN5239_n_26428) );
in01s01 FE_OCPC5240_n_26428 ( .a(FE_OCPN5239_n_26428), .o(FE_OCPN5240_n_26428) );
in01s01 FE_OCPC5241_n_30859 ( .a(n_30859), .o(FE_OCPN5241_n_30859) );
in01s01 FE_OCPC5242_n_30859 ( .a(FE_OCPN5241_n_30859), .o(FE_OCPN5242_n_30859) );
in01s01 FE_OCPC5243_n_21790 ( .a(n_21790), .o(FE_OCPN5243_n_21790) );
in01s01 FE_OCPC5244_n_21790 ( .a(FE_OCPN5243_n_21790), .o(FE_OCPN5244_n_21790) );
in01s01 FE_OCPC5245_n_18974 ( .a(n_18974), .o(FE_OCPN5245_n_18974) );
in01s01 FE_OCPC5246_n_18974 ( .a(FE_OCPN5245_n_18974), .o(FE_OCPN5246_n_18974) );
in01s01 FE_OCPC5247_FE_OFN4715_n_18642 ( .a(FE_OFN4715_n_18642), .o(FE_OCPN5247_FE_OFN4715_n_18642) );
in01s01 FE_OCPC5248_FE_OFN4715_n_18642 ( .a(FE_OCPN5247_FE_OFN4715_n_18642), .o(FE_OCPN5248_FE_OFN4715_n_18642) );
in01s01 FE_OCPC5249_n_20852 ( .a(n_20852), .o(FE_OCPN5249_n_20852) );
in01s01 FE_OCPC5250_n_20852 ( .a(FE_OCPN5249_n_20852), .o(FE_OCPN5250_n_20852) );
in01s01 FE_OCPC5251_n_30859 ( .a(n_30859), .o(FE_OCPN5251_n_30859) );
in01s01 FE_OCPC5252_n_30859 ( .a(FE_OCPN5251_n_30859), .o(FE_OCPN5252_n_30859) );
in01s01 FE_OCPC5253_n_31871 ( .a(n_31871), .o(FE_OCPN5253_n_31871) );
in01s02 FE_OCPC5254_n_31871 ( .a(FE_OCPN5253_n_31871), .o(FE_OCPN5254_n_31871) );
in01s01 FE_OCPC5257_n_13590 ( .a(n_13590), .o(FE_OCPN5257_n_13590) );
in01s01 FE_OCPC5258_n_13590 ( .a(FE_OCPN5257_n_13590), .o(FE_OCPN5258_n_13590) );
in01s01 FE_OCPC5259_n_30614 ( .a(n_30614), .o(FE_OCPN5259_n_30614) );
in01s01 FE_OCPC5260_n_30614 ( .a(FE_OCPN5259_n_30614), .o(FE_OCPN5260_n_30614) );
in01s01 FE_OCPC5261_n_27536 ( .a(n_27536), .o(FE_OCPN5261_n_27536) );
in01s01 FE_OCPC5262_n_27536 ( .a(FE_OCPN5261_n_27536), .o(FE_OCPN5262_n_27536) );
in01s01 FE_OCPC5263_n_14977 ( .a(n_14977), .o(FE_OCPN5263_n_14977) );
in01s01 FE_OCPC5264_n_14977 ( .a(FE_OCPN5263_n_14977), .o(FE_OCPN5264_n_14977) );
in01s01 FE_OCPC5265_n_20852 ( .a(n_20852), .o(FE_OCPN5265_n_20852) );
in01s01 FE_OCPC5267_n_34852 ( .a(n_34852), .o(FE_OCPN5267_n_34852) );
in01s01 FE_OCPC5268_n_34852 ( .a(FE_OCPN5267_n_34852), .o(FE_OCPN5268_n_34852) );
in01s01 FE_OCPC5269_n_18557 ( .a(n_18557), .o(FE_OCPN5269_n_18557) );
in01s01 FE_OCPC5270_n_18557 ( .a(FE_OCPN5269_n_18557), .o(FE_OCPN5270_n_18557) );
in01s01 FE_OCPC5271_n_21434 ( .a(n_21434), .o(FE_OCPN5271_n_21434) );
in01s01 FE_OCPC5272_n_21434 ( .a(FE_OCPN5271_n_21434), .o(FE_OCPN5272_n_21434) );
in01s02 FE_OCPC5273_FE_RN_366_0 ( .a(FE_RN_366_0), .o(FE_OCPN5273_FE_RN_366_0) );
in01s02 FE_OCPC5274_FE_RN_366_0 ( .a(FE_OCPN5273_FE_RN_366_0), .o(FE_OCPN5274_FE_RN_366_0) );
in01s01 FE_OCPC5275_n_23590 ( .a(n_23590), .o(FE_OCPN5275_n_23590) );
in01s01 FE_OCPC5276_n_23590 ( .a(FE_OCPN5275_n_23590), .o(FE_OCPN5276_n_23590) );
in01s01 FE_OCPC5277_n_13329 ( .a(n_13329), .o(FE_OCPN5277_n_13329) );
in01s01 FE_OCPC5279_n_30614 ( .a(FE_OCPN5260_n_30614), .o(FE_OCPN5279_n_30614) );
in01s01 FE_OCPC5280_n_30614 ( .a(FE_OCPN5279_n_30614), .o(FE_OCPN5280_n_30614) );
in01s01 FE_OCPC5281_n_24425 ( .a(n_24425), .o(FE_OCPN5281_n_24425) );
in01s01 FE_OCPC5283_n_24425 ( .a(n_24425), .o(FE_OCPN5283_n_24425) );
in01s01 FE_OCPC5284_n_24425 ( .a(FE_OCPN5283_n_24425), .o(FE_OCPN5284_n_24425) );
in01s01 FE_OCPC5285_n_30708 ( .a(FE_OCPN1763_n_30708), .o(FE_OCPN5285_n_30708) );
in01s01 FE_OCPC5286_n_30708 ( .a(FE_OCPN5285_n_30708), .o(FE_OCPN5286_n_30708) );
in01s01 FE_OCPC5287_n_27315 ( .a(n_27315), .o(FE_OCPN5287_n_27315) );
in01s01 FE_OCPC5288_n_27315 ( .a(FE_OCPN5287_n_27315), .o(FE_OCPN5288_n_27315) );
in01s01 FE_OCPC5289_n_26125 ( .a(n_26125), .o(FE_OCPN5289_n_26125) );
in01s01 FE_OCPC5290_n_26125 ( .a(FE_OCPN5289_n_26125), .o(FE_OCPN5290_n_26125) );
in01s01 FE_OCPC5291_n_21790 ( .a(n_21790), .o(FE_OCPN5291_n_21790) );
in01s01 FE_OCPC5292_n_21790 ( .a(FE_OCPN5291_n_21790), .o(FE_OCPN5292_n_21790) );
in01s01 FE_OCPC5293_n_30584 ( .a(n_30584), .o(FE_OCPN5293_n_30584) );
in01s01 FE_OCPC5294_n_30584 ( .a(FE_OCPN5293_n_30584), .o(FE_OCPN5294_n_30584) );
in01s01 FE_OCPC5295_FE_OCP_RBN1105_n_18746 ( .a(FE_OCP_RBN1105_n_18746), .o(FE_OCPN5295_FE_OCP_RBN1105_n_18746) );
in01s01 FE_OCPC5296_FE_OCP_RBN1105_n_18746 ( .a(FE_OCPN5295_FE_OCP_RBN1105_n_18746), .o(FE_OCPN5296_FE_OCP_RBN1105_n_18746) );
in01s01 FE_OCPC5297_n_29866 ( .a(n_29866), .o(FE_OCPN5297_n_29866) );
in01s01 FE_OCPC5298_n_29866 ( .a(FE_OCPN5297_n_29866), .o(FE_OCPN5298_n_29866) );
in01s01 FE_OCPC5299_n_27130 ( .a(n_27130), .o(FE_OCPN5299_n_27130) );
in01s02 FE_OCPC5300_n_27130 ( .a(FE_OCPN5299_n_27130), .o(FE_OCPN5300_n_27130) );
in01s01 FE_OCPC5305_n_22338 ( .a(n_22338), .o(FE_OCPN5305_n_22338) );
in01s02 FE_OCPC5306_n_22338 ( .a(FE_OCPN5305_n_22338), .o(FE_OCPN5306_n_22338) );
in01s01 FE_OCPC5363_n_24221 ( .a(n_24221), .o(FE_OCPN5363_n_24221) );
in01s01 FE_OCPC5364_n_24221 ( .a(FE_OCPN5363_n_24221), .o(FE_OCPN5364_n_24221) );
in01s01 FE_OCPC6268_n_30599 ( .a(n_30599), .o(FE_OCPN6268_n_30599) );
in01s01 FE_OCPC6269_n_30599 ( .a(FE_OCPN6268_n_30599), .o(FE_OCPN6269_n_30599) );
in01m06 FE_OCPC6276_n_45450 ( .a(FE_OCPN867_n_45450), .o(FE_OCPN6276_n_45450) );
in01s40 FE_OCPC6277_n_45450 ( .a(FE_OCPN6276_n_45450), .o(FE_OCPN6277_n_45450) );
in01s01 FE_OCPC6278_FE_OCP_RBN1594_n_13557 ( .a(FE_OCP_RBN1594_n_13557), .o(FE_OCPN6278_FE_OCP_RBN1594_n_13557) );
in01s01 FE_OCPC6279_FE_OCP_RBN1594_n_13557 ( .a(FE_OCPN6278_FE_OCP_RBN1594_n_13557), .o(FE_OCPN6279_FE_OCP_RBN1594_n_13557) );
in01s01 FE_OCPC6280_n_30612 ( .a(FE_OCPN1376_n_30612), .o(FE_OCPN6280_n_30612) );
in01s01 FE_OCPC6281_n_30612 ( .a(FE_OCPN6280_n_30612), .o(FE_OCPN6281_n_30612) );
in01s01 FE_OCPC6282_FE_OCP_RBN2783_n_8664 ( .a(FE_OCP_RBN2783_n_8664), .o(FE_OCPN6282_FE_OCP_RBN2783_n_8664) );
in01s01 FE_OCPC6283_FE_OCP_RBN2783_n_8664 ( .a(FE_OCPN6282_FE_OCP_RBN2783_n_8664), .o(FE_OCPN6283_FE_OCP_RBN2783_n_8664) );
in01s01 FE_OCPC6284_FE_OCP_RBN1602_n_14638 ( .a(FE_OCP_RBN1602_n_14638), .o(FE_OCPN6284_FE_OCP_RBN1602_n_14638) );
in01s01 FE_OCPC6285_FE_OCP_RBN1602_n_14638 ( .a(FE_OCPN6284_FE_OCP_RBN1602_n_14638), .o(FE_OCPN6285_FE_OCP_RBN1602_n_14638) );
in01s01 FE_OCPC6286_FE_OCP_RBN6082_n_5454 ( .a(FE_OCP_RBN6082_n_5454), .o(FE_OCPN6286_FE_OCP_RBN6082_n_5454) );
in01s01 FE_OCPC6287_FE_OCP_RBN6082_n_5454 ( .a(FE_OCPN6286_FE_OCP_RBN6082_n_5454), .o(FE_OCPN6287_FE_OCP_RBN6082_n_5454) );
in01s01 FE_OCPC6288_FE_OCP_RBN3263_n_5531 ( .a(FE_OCP_RBN3263_n_5531), .o(FE_OCPN6288_FE_OCP_RBN3263_n_5531) );
in01s01 FE_OCPC6289_FE_OCP_RBN3263_n_5531 ( .a(FE_OCPN6288_FE_OCP_RBN3263_n_5531), .o(FE_OCPN6289_FE_OCP_RBN3263_n_5531) );
in01s02 FE_OCPC6900_FE_OCP_RBN4472_n_31819 ( .a(FE_OCP_RBN4472_n_31819), .o(FE_OCPN6900_FE_OCP_RBN4472_n_31819) );
in01s02 FE_OCPC6901_FE_OCP_RBN4472_n_31819 ( .a(FE_OCPN6900_FE_OCP_RBN4472_n_31819), .o(FE_OCPN6901_FE_OCP_RBN4472_n_31819) );
in01s01 FE_OCPC6908_n_32525 ( .a(n_32525), .o(FE_OCPN6908_n_32525) );
in01s01 FE_OCPC6909_n_32525 ( .a(FE_OCPN6908_n_32525), .o(FE_OCPN6909_n_32525) );
in01s01 FE_OCPC6910_n_1444 ( .a(n_1444), .o(FE_OCPN6910_n_1444) );
in01s01 FE_OCPC6911_n_1444 ( .a(FE_OCPN6910_n_1444), .o(FE_OCPN6911_n_1444) );
in01s01 FE_OCPC6912_n_1715 ( .a(n_1715), .o(FE_OCPN6912_n_1715) );
in01s01 FE_OCPC6913_n_1715 ( .a(FE_OCPN6912_n_1715), .o(FE_OCPN6913_n_1715) );
in01s10 FE_OCPC6914_n_23112 ( .a(n_23112), .o(FE_OCPN6914_n_23112) );
in01s10 FE_OCPC6915_n_23112 ( .a(FE_OCPN6914_n_23112), .o(FE_OCPN6915_n_23112) );
in01s01 FE_OCPC6916_n_28460 ( .a(n_28460), .o(FE_OCPN6916_n_28460) );
in01s01 FE_OCPC6917_n_28460 ( .a(FE_OCPN6916_n_28460), .o(FE_OCPN6917_n_28460) );
in01s01 FE_OCPC6918_n_7726 ( .a(n_7726), .o(FE_OCPN6918_n_7726) );
in01s01 FE_OCPC6919_n_7726 ( .a(FE_OCPN6918_n_7726), .o(FE_OCPN6919_n_7726) );
in01s01 FE_OCPC6920_n_3580 ( .a(n_3580), .o(FE_OCPN6920_n_3580) );
in01s01 FE_OCPC6921_n_3580 ( .a(FE_OCPN6920_n_3580), .o(FE_OCPN6921_n_3580) );
in01m02 FE_OCPC6922_n_39185 ( .a(n_39185), .o(FE_OCPN6922_n_39185) );
in01m04 FE_OCPC6923_n_39185 ( .a(FE_OCPN6922_n_39185), .o(FE_OCPN6923_n_39185) );
in01s01 FE_OCPC6924_n_45081 ( .a(n_45081), .o(FE_OCPN6924_n_45081) );
in01s01 FE_OCPC6925_n_45081 ( .a(FE_OCPN6924_n_45081), .o(FE_OCPN6925_n_45081) );
in01s01 FE_OCPC6926_n_26464 ( .a(n_26464), .o(FE_OCPN6926_n_26464) );
in01s01 FE_OCPC6927_n_26464 ( .a(FE_OCPN6926_n_26464), .o(FE_OCPN6927_n_26464) );
in01s01 FE_OCPC6928_FE_OCP_RBN1152_n_20910 ( .a(FE_OCP_RBN1152_n_20910), .o(FE_OCPN6928_FE_OCP_RBN1152_n_20910) );
in01s01 FE_OCPC6929_FE_OCP_RBN1152_n_20910 ( .a(FE_OCPN6928_FE_OCP_RBN1152_n_20910), .o(FE_OCPN6929_FE_OCP_RBN1152_n_20910) );
in01s01 FE_OCPC6930_n_22156 ( .a(n_22156), .o(FE_OCPN6930_n_22156) );
in01s01 FE_OCPC6931_n_22156 ( .a(FE_OCPN6930_n_22156), .o(FE_OCPN6931_n_22156) );
in01s01 FE_OCPC6932_FE_OCP_RBN6087_n_10852 ( .a(FE_OCP_RBN6087_n_10852), .o(FE_OCPN6932_FE_OCP_RBN6087_n_10852) );
in01s01 FE_OCPC6933_FE_OCP_RBN6087_n_10852 ( .a(FE_OCPN6932_FE_OCP_RBN6087_n_10852), .o(FE_OCPN6933_FE_OCP_RBN6087_n_10852) );
in01s01 FE_OCPC6934_FE_OCP_RBN6066_n_26081 ( .a(FE_OCP_RBN6066_n_26081), .o(FE_OCPN6934_FE_OCP_RBN6066_n_26081) );
in01s01 FE_OCPC6935_FE_OCP_RBN6066_n_26081 ( .a(FE_OCPN6934_FE_OCP_RBN6066_n_26081), .o(FE_OCPN6935_FE_OCP_RBN6066_n_26081) );
in01s01 FE_OCPC7082_n_28891 ( .a(n_28891), .o(FE_OCPN7082_n_28891) );
in01s01 FE_OCPC7083_n_28891 ( .a(FE_OCPN7082_n_28891), .o(FE_OCPN7083_n_28891) );
in01s02 FE_OCPC7084_n_45697 ( .a(n_45697), .o(FE_OCPN7084_n_45697) );
in01m01 FE_OCPC7085_n_45697 ( .a(FE_OCPN7084_n_45697), .o(FE_OCPN7085_n_45697) );
in01s01 FE_OCPC7086_n_6263 ( .a(n_6263), .o(FE_OCPN7086_n_6263) );
in01s01 FE_OCPC7087_n_6263 ( .a(FE_OCPN7086_n_6263), .o(FE_OCPN7087_n_6263) );
in01s01 FE_OCPC7088_n_20979 ( .a(n_20979), .o(FE_OCPN7088_n_20979) );
in01s01 FE_OCPC7089_n_20979 ( .a(FE_OCPN7088_n_20979), .o(FE_OCPN7089_n_20979) );
in01s40 FE_OCPC833_n_45450 ( .a(FE_OCPN1202_n_45450), .o(FE_OCPN833_n_45450) );
in01s03 FE_OCPC835_n_45450 ( .a(FE_OCPN6277_n_45450), .o(FE_OCPN835_n_45450) );
in01s10 FE_OCPC836_n_45450 ( .a(FE_OCPN835_n_45450), .o(FE_OCPN836_n_45450) );
in01s02 FE_OCPC837_n_44672 ( .a(n_44672), .o(FE_OCPN837_n_44672) );
in01s01 FE_OCPC838_n_44672 ( .a(FE_OCPN837_n_44672), .o(FE_OCPN838_n_44672) );
in01s02 FE_OCPC839_n_44672 ( .a(FE_OCPN837_n_44672), .o(FE_OCPN839_n_44672) );
in01s01 FE_OCPC846_n_12799 ( .a(n_12799), .o(FE_OCPN846_n_12799) );
in01s01 FE_OCPC847_n_12799 ( .a(FE_OCPN846_n_12799), .o(FE_OCPN847_n_12799) );
in01s01 FE_OCPC848_n_7712 ( .a(n_7712), .o(FE_OCPN848_n_7712) );
in01s02 FE_OCPC849_n_7712 ( .a(FE_OCPN848_n_7712), .o(FE_OCPN849_n_7712) );
in01s01 FE_OCPC850_n_7712 ( .a(FE_OCPN848_n_7712), .o(FE_OCPN850_n_7712) );
in01s01 FE_OCPC858_n_7802 ( .a(FE_OCP_RBN5612_n_7730), .o(FE_OCPN858_n_7802) );
in01s01 FE_OCPC861_n_7743 ( .a(FE_OCP_RBN6600_n_7708), .o(FE_OCPN861_n_7743) );
in01s01 FE_OCPC865_n_32892 ( .a(FE_OCP_RBN2454_n_32860), .o(FE_OCPN865_n_32892) );
in01s10 FE_OCPC866_n_45450 ( .a(FE_OCP_RBN5513_n_44365), .o(FE_OCPN866_n_45450) );
in01s40 FE_OCPC867_n_45450 ( .a(FE_OCPN866_n_45450), .o(FE_OCPN867_n_45450) );
in01s06 FE_OCPC868_n_45003 ( .a(n_45003), .o(FE_OCPN868_n_45003) );
in01s06 FE_OCPC869_n_45003 ( .a(FE_OCPN868_n_45003), .o(FE_OCPN869_n_45003) );
in01s01 FE_OCPC870_n_24098 ( .a(FE_OCP_RBN5615_n_24070), .o(FE_OCPN870_n_24098) );
in01s01 FE_OCPC871_n_24098 ( .a(FE_OCPN870_n_24098), .o(FE_OCPN871_n_24098) );
in01m02 FE_OCPC872_n_42202 ( .a(n_42202), .o(FE_OCPN872_n_42202) );
in01s04 FE_OCPC873_n_42202 ( .a(FE_OCPN872_n_42202), .o(FE_OCPN873_n_42202) );
in01s01 FE_OCPC877_n_43022 ( .a(n_43022), .o(FE_OCPN877_n_43022) );
in01s04 FE_OCPC878_n_43022 ( .a(FE_OCPN877_n_43022), .o(FE_OCPN878_n_43022) );
in01s01 FE_OCPC880_n_44593 ( .a(FE_OCP_RBN4243_n_44594), .o(FE_OCPN880_n_44593) );
in01s01 FE_OCPC881_n_44776 ( .a(n_44776), .o(FE_OCPN881_n_44776) );
in01s02 FE_OCPC882_n_44776 ( .a(FE_OCPN881_n_44776), .o(FE_OCPN882_n_44776) );
in01s01 FE_OCPC883_n_41540 ( .a(n_41540), .o(FE_OCPN883_n_41540) );
in01s02 FE_OCPC884_n_41540 ( .a(FE_OCPN883_n_41540), .o(FE_OCPN884_n_41540) );
in01s01 FE_OCPC889_n_44223 ( .a(FE_OCP_RBN4904_n_44256), .o(FE_OCPN889_n_44223) );
in01s03 FE_OCPC890_n_44223 ( .a(FE_OCPN889_n_44223), .o(FE_OCPN890_n_44223) );
in01f06 FE_OCPC894_n_28471 ( .a(FE_OCPN893_n_28471), .o(FE_OCPN894_n_28471) );
in01f06 FE_OCPC896_n_28506 ( .a(FE_OCPN895_n_28506), .o(FE_OCPN896_n_28506) );
in01s03 FE_OCPC899_n_16923 ( .a(n_16923), .o(FE_OCPN899_n_16923) );
in01s06 FE_OCPC900_n_16923 ( .a(FE_OCPN899_n_16923), .o(FE_OCPN900_n_16923) );
in01s01 FE_OCPC901_n_47020 ( .a(n_47020), .o(FE_OCPN901_n_47020) );
in01s01 FE_OCPC902_n_47020 ( .a(FE_OCPN901_n_47020), .o(FE_OCPN902_n_47020) );
in01s03 FE_OCPC904_n_21955 ( .a(FE_OCPN903_n_21955), .o(FE_OCPN904_n_21955) );
in01s02 FE_OCPC905_n_21956 ( .a(n_21956), .o(FE_OCPN905_n_21956) );
in01s03 FE_OCPC906_n_21956 ( .a(FE_OCPN905_n_21956), .o(FE_OCPN906_n_21956) );
in01s01 FE_OCPC907_n_46956 ( .a(n_46956), .o(FE_OCPN907_n_46956) );
in01s01 FE_OCPC908_n_46956 ( .a(FE_OCPN907_n_46956), .o(FE_OCPN908_n_46956) );
in01m02 FE_OCPC914_n_8091 ( .a(n_8091), .o(FE_OCPN914_n_8091) );
in01f02 FE_OCPC916_n_8753 ( .a(n_8753), .o(FE_OCPN916_n_8753) );
in01f04 FE_OCPC917_n_8753 ( .a(FE_OCPN916_n_8753), .o(FE_OCPN917_n_8753) );
in01s01 FE_OCPC918_n_17042 ( .a(n_17042), .o(FE_OCPN918_n_17042) );
in01s01 FE_OCPC919_n_17042 ( .a(FE_OCPN918_n_17042), .o(FE_OCPN919_n_17042) );
in01s01 FE_OCPC924_n_13962 ( .a(FE_OCP_RBN2819_n_13962), .o(FE_OCPN924_n_13962) );
in01s06 FE_OCPC926_n_12914 ( .a(FE_OCP_RBN2541_n_12880), .o(FE_OCPN926_n_12914) );
in01s01 FE_OCPC928_n_12880 ( .a(FE_OCP_RBN2539_n_12880), .o(FE_OCPN928_n_12880) );
in01s01 FE_OCPC929_n_12880 ( .a(FE_OCPN928_n_12880), .o(FE_OCPN929_n_12880) );
in01s01 FE_OCPC930_n_7817 ( .a(FE_OCP_RBN5609_n_7730), .o(FE_OCPN930_n_7817) );
in01s02 FE_OCPC931_n_7817 ( .a(FE_OCPN930_n_7817), .o(FE_OCPN931_n_7817) );
in01s02 FE_OCPC935_n_7802 ( .a(FE_OCP_RBN2614_FE_OCPN857_n_7802), .o(FE_OCPN935_n_7802) );
in01s01 FE_OCPC936_n_17684 ( .a(n_17684), .o(FE_OCPN936_n_17684) );
in01s06 FE_OCPC937_n_17684 ( .a(FE_OCPN936_n_17684), .o(FE_OCPN937_n_17684) );
in01f02 FE_OCPC938_n_23577 ( .a(n_23577), .o(FE_OCPN938_n_23577) );
in01f04 FE_OCPC939_n_23577 ( .a(FE_OCPN938_n_23577), .o(FE_OCPN939_n_23577) );
in01s01 FE_OCPC940_n_39096 ( .a(FE_OCP_RBN4329_n_38878), .o(FE_OCPN940_n_39096) );
in01s01 FE_OCPC941_n_39096 ( .a(FE_OCPN940_n_39096), .o(FE_OCPN941_n_39096) );
in01s06 FE_OCPC942_n_31466 ( .a(n_31466), .o(FE_OCPN942_n_31466) );
in01m03 FE_OCPC943_n_31466 ( .a(FE_OCPN942_n_31466), .o(FE_OCPN943_n_31466) );
in01f10 FE_OCPC945_n_27287 ( .a(FE_OCP_RBN6219_n_27110), .o(FE_OCPN945_n_27287) );
in01s06 FE_OCPC950_n_44180 ( .a(FE_OCP_RBN3171_n_44211), .o(FE_OCPN950_n_44180) );
in01s01 FE_OCPUNCOC1742_n_29375 ( .a(FE_OCP_DRV_N5141_n_29375), .o(FE_OCPUNCON1742_n_29375) );
in01s01 FE_OCPUNCOC1743_n_29375 ( .a(FE_OCPUNCON1742_n_29375), .o(FE_OCPUNCON1743_n_29375) );
in01s01 FE_OCPUNCOC1744_n_29420 ( .a(n_29420), .o(FE_OCPUNCON1744_n_29420) );
in01s01 FE_OCPUNCOC1745_n_29420 ( .a(FE_OCPUNCON1744_n_29420), .o(FE_OCPUNCON1745_n_29420) );
in01s01 FE_OCPUNCOC1746_n_34137 ( .a(n_34137), .o(FE_OCPUNCON1746_n_34137) );
in01s01 FE_OCPUNCOC1747_n_34137 ( .a(FE_OCPUNCON1746_n_34137), .o(FE_OCPUNCON1747_n_34137) );
in01s01 FE_OCPUNCOC1748_n_19807 ( .a(n_19807), .o(FE_OCPUNCON1748_n_19807) );
in01s01 FE_OCPUNCOC1749_n_19807 ( .a(FE_OCPUNCON1748_n_19807), .o(FE_OCPUNCON1749_n_19807) );
in01s01 FE_OCPUNCOC1750_n_33904 ( .a(FE_OCPUNCON7063_n_33904), .o(FE_OCPUNCON1750_n_33904) );
in01s01 FE_OCPUNCOC1752_n_35382 ( .a(n_35382), .o(FE_OCPUNCON1752_n_35382) );
in01s01 FE_OCPUNCOC1753_n_35382 ( .a(FE_OCPUNCON1752_n_35382), .o(FE_OCPUNCON1753_n_35382) );
in01s01 FE_OCPUNCOC1754_n_35420 ( .a(n_35420), .o(FE_OCPUNCON1754_n_35420) );
in01s01 FE_OCPUNCOC1755_n_35420 ( .a(FE_OCPUNCON1754_n_35420), .o(FE_OCPUNCON1755_n_35420) );
in01s01 FE_OCPUNCOC1756_n_35482 ( .a(n_35482), .o(FE_OCPUNCON1756_n_35482) );
in01s01 FE_OCPUNCOC1757_n_35482 ( .a(FE_OCPUNCON1756_n_35482), .o(FE_OCPUNCON1757_n_35482) );
in01s01 FE_OCPUNCOC1758_n_35644 ( .a(n_35644), .o(FE_OCPUNCON1758_n_35644) );
in01s01 FE_OCPUNCOC1759_n_35644 ( .a(FE_OCPUNCON1758_n_35644), .o(FE_OCPUNCON1759_n_35644) );
in01s01 FE_OCPUNCOC3465_n_29391 ( .a(n_29391), .o(FE_OCPUNCON3465_n_29391) );
in01s01 FE_OCPUNCOC3466_n_29391 ( .a(FE_OCPUNCON3465_n_29391), .o(FE_OCPUNCON3466_n_29391) );
in01s01 FE_OCPUNCOC3467_n_29644 ( .a(n_29644), .o(FE_OCPUNCON3467_n_29644) );
in01s01 FE_OCPUNCOC3468_n_29644 ( .a(FE_OCPUNCON3467_n_29644), .o(FE_OCPUNCON3468_n_29644) );
in01s01 FE_OCPUNCOC3469_n_28654 ( .a(n_28654), .o(FE_OCPUNCON3469_n_28654) );
in01s01 FE_OCPUNCOC3470_n_28654 ( .a(FE_OCPUNCON3469_n_28654), .o(FE_OCPUNCON3470_n_28654) );
in01s01 FE_OCPUNCOC3471_n_24962 ( .a(n_24962), .o(FE_OCPUNCON3471_n_24962) );
in01s01 FE_OCPUNCOC3472_n_24962 ( .a(FE_OCPUNCON3471_n_24962), .o(FE_OCPUNCON3472_n_24962) );
in01s01 FE_OCPUNCOC3473_n_28656 ( .a(n_28656), .o(FE_OCPUNCON3473_n_28656) );
in01s01 FE_OCPUNCOC3475_n_29812 ( .a(n_29812), .o(FE_OCPUNCON3475_n_29812) );
in01s01 FE_OCPUNCOC3476_n_29812 ( .a(FE_OCPUNCON3475_n_29812), .o(FE_OCPUNCON3476_n_29812) );
in01s01 FE_OCPUNCOC3477_n_29844 ( .a(n_29844), .o(FE_OCPUNCON3477_n_29844) );
in01s01 FE_OCPUNCOC3478_n_29844 ( .a(FE_OCPUNCON3477_n_29844), .o(FE_OCPUNCON3478_n_29844) );
in01s01 FE_OCPUNCOC3479_n_28872 ( .a(n_28872), .o(FE_OCPUNCON3479_n_28872) );
in01s01 FE_OCPUNCOC3480_n_28872 ( .a(FE_OCPUNCON3479_n_28872), .o(FE_OCPUNCON3480_n_28872) );
in01s01 FE_OCPUNCOC3481_n_21058 ( .a(n_21058), .o(FE_OCPUNCON3481_n_21058) );
in01s01 FE_OCPUNCOC3483_n_35500 ( .a(FE_OCPUNCON7065_n_35500), .o(FE_OCPUNCON3483_n_35500) );
in01s01 FE_OCPUNCOC3484_n_35500 ( .a(FE_OCPUNCON3483_n_35500), .o(FE_OCPUNCON3484_n_35500) );
in01s01 FE_OCPUNCOC3485_n_31012 ( .a(n_31012), .o(FE_OCPUNCON3485_n_31012) );
in01s01 FE_OCPUNCOC3487_n_21458 ( .a(n_21458), .o(FE_OCPUNCON3487_n_21458) );
in01s01 FE_OCPUNCOC3488_n_21458 ( .a(FE_OCPUNCON3487_n_21458), .o(FE_OCPUNCON3488_n_21458) );
in01s01 FE_OCPUNCOC3489_n_34327 ( .a(n_34327), .o(FE_OCPUNCON3489_n_34327) );
in01s01 FE_OCPUNCOC3490_n_34327 ( .a(FE_OCPUNCON3489_n_34327), .o(FE_OCPUNCON3490_n_34327) );
in01s01 FE_OCPUNCOC3491_n_30322 ( .a(FE_OCP_DRV_N5161_n_30322), .o(FE_OCPUNCON3491_n_30322) );
in01s01 FE_OCPUNCOC4497_n_34182 ( .a(n_34182), .o(FE_OCPUNCON4497_n_34182) );
in01s01 FE_OCPUNCOC4498_n_34182 ( .a(FE_OCPUNCON4497_n_34182), .o(FE_OCPUNCON4498_n_34182) );
in01s01 FE_OCPUNCOC5301_n_17836 ( .a(n_17836), .o(FE_OCPUNCON5301_n_17836) );
in01s01 FE_OCPUNCOC5302_n_17836 ( .a(FE_OCPUNCON5301_n_17836), .o(FE_OCPUNCON5302_n_17836) );
in01s01 FE_OCPUNCOC6886_n_19961 ( .a(n_19961), .o(FE_OCPUNCON6886_n_19961) );
in01s01 FE_OCPUNCOC6887_n_19961 ( .a(FE_OCPUNCON6886_n_19961), .o(FE_OCPUNCON6887_n_19961) );
in01s01 FE_OCPUNCOC7058_n_34058 ( .a(n_34058), .o(FE_OCPUNCON7058_n_34058) );
in01s01 FE_OCPUNCOC7059_n_34058 ( .a(FE_OCPUNCON7058_n_34058), .o(FE_OCPUNCON7059_n_34058) );
in01s01 FE_OCPUNCOC7060_n_34222 ( .a(n_34222), .o(FE_OCPUNCON7060_n_34222) );
in01s01 FE_OCPUNCOC7061_n_34222 ( .a(FE_OCPUNCON7060_n_34222), .o(FE_OCPUNCON7061_n_34222) );
in01s01 FE_OCPUNCOC7062_n_33904 ( .a(n_33904), .o(FE_OCPUNCON7062_n_33904) );
in01s01 FE_OCPUNCOC7063_n_33904 ( .a(FE_OCPUNCON7062_n_33904), .o(FE_OCPUNCON7063_n_33904) );
in01s01 FE_OCPUNCOC7064_n_35500 ( .a(n_35500), .o(FE_OCPUNCON7064_n_35500) );
in01s01 FE_OCPUNCOC7065_n_35500 ( .a(FE_OCPUNCON7064_n_35500), .o(FE_OCPUNCON7065_n_35500) );
in01s01 FE_OCPUNCOC7066_n_34151 ( .a(n_34151), .o(FE_OCPUNCON7066_n_34151) );
in01s01 FE_OCPUNCOC7067_n_34151 ( .a(FE_OCPUNCON7066_n_34151), .o(FE_OCPUNCON7067_n_34151) );
in01s01 FE_OCPUNCOC7068_n_21493 ( .a(n_21493), .o(FE_OCPUNCON7068_n_21493) );
in01s01 FE_OCPUNCOC7069_n_21493 ( .a(FE_OCPUNCON7068_n_21493), .o(FE_OCPUNCON7069_n_21493) );
in01s01 FE_OCPUNCOC7070_n_21788 ( .a(n_21788), .o(FE_OCPUNCON7070_n_21788) );
in01s01 FE_OCPUNCOC7071_n_21788 ( .a(FE_OCPUNCON7070_n_21788), .o(FE_OCPUNCON7071_n_21788) );
in01s01 FE_OCPUNCOC7072_n_31583 ( .a(n_31583), .o(FE_OCPUNCON7072_n_31583) );
in01s01 FE_OCPUNCOC7073_n_31583 ( .a(FE_OCPUNCON7072_n_31583), .o(FE_OCPUNCON7073_n_31583) );
in01s01 FE_OCP_DRV_C1405_n_43514 ( .a(n_43514), .o(FE_OCP_DRV_N1405_n_43514) );
in01s01 FE_OCP_DRV_C1406_n_43514 ( .a(FE_OCP_DRV_N1405_n_43514), .o(FE_OCP_DRV_N1406_n_43514) );
in01s01 FE_OCP_DRV_C1407_n_28550 ( .a(n_28550), .o(FE_OCP_DRV_N1407_n_28550) );
in01s02 FE_OCP_DRV_C1409_n_12416 ( .a(n_12416), .o(FE_OCP_DRV_N1409_n_12416) );
in01s02 FE_OCP_DRV_C1410_n_12416 ( .a(FE_OCP_DRV_N1409_n_12416), .o(FE_OCP_DRV_N1410_n_12416) );
in01s01 FE_OCP_DRV_C1411_n_12570 ( .a(n_12570), .o(FE_OCP_DRV_N1411_n_12570) );
in01s02 FE_OCP_DRV_C1412_n_12570 ( .a(FE_OCP_DRV_N1411_n_12570), .o(FE_OCP_DRV_N1412_n_12570) );
in01s01 FE_OCP_DRV_C1413_n_33673 ( .a(n_33673), .o(FE_OCP_DRV_N1413_n_33673) );
in01s01 FE_OCP_DRV_C1414_n_33673 ( .a(FE_OCP_DRV_N1413_n_33673), .o(FE_OCP_DRV_N1414_n_33673) );
in01s01 FE_OCP_DRV_C1416_n_34051 ( .a(FE_OCPN1373_n_34051), .o(FE_OCP_DRV_N1416_n_34051) );
in01s01 FE_OCP_DRV_C1417_n_32985 ( .a(n_32985), .o(FE_OCP_DRV_N1417_n_32985) );
in01s01 FE_OCP_DRV_C1419_n_24747 ( .a(n_24747), .o(FE_OCP_DRV_N1419_n_24747) );
in01s01 FE_OCP_DRV_C1420_n_24747 ( .a(FE_OCP_DRV_N1419_n_24747), .o(FE_OCP_DRV_N1420_n_24747) );
in01s01 FE_OCP_DRV_C1421_n_35367 ( .a(n_35367), .o(FE_OCP_DRV_N1421_n_35367) );
in01s01 FE_OCP_DRV_C1423_n_35292 ( .a(n_35292), .o(FE_OCP_DRV_N1423_n_35292) );
in01s01 FE_OCP_DRV_C1424_n_35292 ( .a(FE_OCP_DRV_N1423_n_35292), .o(FE_OCP_DRV_N1424_n_35292) );
in01s01 FE_OCP_DRV_C1425_n_24158 ( .a(n_24158), .o(FE_OCP_DRV_N1425_n_24158) );
in01s01 FE_OCP_DRV_C1426_n_24158 ( .a(FE_OCP_DRV_N1425_n_24158), .o(FE_OCP_DRV_N1426_n_24158) );
in01s01 FE_OCP_DRV_C1427_n_35312 ( .a(n_35312), .o(FE_OCP_DRV_N1427_n_35312) );
in01s01 FE_OCP_DRV_C1428_n_35312 ( .a(FE_OCP_DRV_N1427_n_35312), .o(FE_OCP_DRV_N1428_n_35312) );
in01s01 FE_OCP_DRV_C1429_n_22126 ( .a(n_22126), .o(FE_OCP_DRV_N1429_n_22126) );
in01s01 FE_OCP_DRV_C1430_n_22126 ( .a(FE_OCP_DRV_N1429_n_22126), .o(FE_OCP_DRV_N1430_n_22126) );
in01s01 FE_OCP_DRV_C1431_n_26850 ( .a(n_26850), .o(FE_OCP_DRV_N1431_n_26850) );
in01s01 FE_OCP_DRV_C1432_n_26850 ( .a(FE_OCP_DRV_N1431_n_26850), .o(FE_OCP_DRV_N1432_n_26850) );
in01s01 FE_OCP_DRV_C1433_n_21283 ( .a(n_21283), .o(FE_OCP_DRV_N1433_n_21283) );
in01s01 FE_OCP_DRV_C1434_n_21283 ( .a(FE_OCP_DRV_N1433_n_21283), .o(FE_OCP_DRV_N1434_n_21283) );
in01s01 FE_OCP_DRV_C1437_n_17643 ( .a(n_17643), .o(FE_OCP_DRV_N1437_n_17643) );
in01s01 FE_OCP_DRV_C1438_n_17643 ( .a(FE_OCP_DRV_N1437_n_17643), .o(FE_OCP_DRV_N1438_n_17643) );
in01s01 FE_OCP_DRV_C1439_n_19010 ( .a(FE_OCP_DRV_N5356_n_19010), .o(FE_OCP_DRV_N1439_n_19010) );
in01s01 FE_OCP_DRV_C1440_n_19010 ( .a(FE_OCP_DRV_N1439_n_19010), .o(FE_OCP_DRV_N1440_n_19010) );
in01s01 FE_OCP_DRV_C1441_n_17836 ( .a(FE_OCPUNCON5302_n_17836), .o(FE_OCP_DRV_N1441_n_17836) );
in01s01 FE_OCP_DRV_C1443_n_19138 ( .a(n_19138), .o(FE_OCP_DRV_N1443_n_19138) );
in01s01 FE_OCP_DRV_C1444_n_19138 ( .a(FE_OCP_DRV_N1443_n_19138), .o(FE_OCP_DRV_N1444_n_19138) );
in01s01 FE_OCP_DRV_C1445_n_19314 ( .a(n_19314), .o(FE_OCP_DRV_N1445_n_19314) );
in01s01 FE_OCP_DRV_C1446_n_19314 ( .a(FE_OCP_DRV_N1445_n_19314), .o(FE_OCP_DRV_N1446_n_19314) );
in01s01 FE_OCP_DRV_C1447_n_19354 ( .a(FE_OCP_DRV_N6903_n_19354), .o(FE_OCP_DRV_N1447_n_19354) );
in01s01 FE_OCP_DRV_C1448_n_19354 ( .a(FE_OCP_DRV_N1447_n_19354), .o(FE_OCP_DRV_N1448_n_19354) );
in01s01 FE_OCP_DRV_C1449_n_19384 ( .a(FE_OFN4804_n_19384), .o(FE_OCP_DRV_N1449_n_19384) );
in01s01 FE_OCP_DRV_C1450_n_19384 ( .a(FE_OCP_DRV_N1449_n_19384), .o(FE_OCP_DRV_N1450_n_19384) );
in01s01 FE_OCP_DRV_C1451_n_12585 ( .a(n_12585), .o(FE_OCP_DRV_N1451_n_12585) );
in01s01 FE_OCP_DRV_C1452_n_12585 ( .a(FE_OCP_DRV_N1451_n_12585), .o(FE_OCP_DRV_N1452_n_12585) );
in01s01 FE_OCP_DRV_C1453_n_19590 ( .a(n_19590), .o(FE_OCP_DRV_N1453_n_19590) );
in01s01 FE_OCP_DRV_C1454_n_19590 ( .a(FE_OCP_DRV_N1453_n_19590), .o(FE_OCP_DRV_N1454_n_19590) );
in01s01 FE_OCP_DRV_C1455_n_19562 ( .a(n_19562), .o(FE_OCP_DRV_N1455_n_19562) );
in01s01 FE_OCP_DRV_C1456_n_19562 ( .a(FE_OCP_DRV_N1455_n_19562), .o(FE_OCP_DRV_N1456_n_19562) );
in01s01 FE_OCP_DRV_C1457_n_19665 ( .a(n_19665), .o(FE_OCP_DRV_N1457_n_19665) );
in01s01 FE_OCP_DRV_C1458_n_19665 ( .a(FE_OCP_DRV_N1457_n_19665), .o(FE_OCP_DRV_N1458_n_19665) );
in01s01 FE_OCP_DRV_C1459_n_18111 ( .a(n_18111), .o(FE_OCP_DRV_N1459_n_18111) );
in01s01 FE_OCP_DRV_C1460_n_18111 ( .a(FE_OCP_DRV_N1459_n_18111), .o(FE_OCP_DRV_N1460_n_18111) );
in01s01 FE_OCP_DRV_C1461_n_29777 ( .a(n_29777), .o(FE_OCP_DRV_N1461_n_29777) );
in01s01 FE_OCP_DRV_C1462_n_29777 ( .a(FE_OCP_DRV_N1461_n_29777), .o(FE_OCP_DRV_N1462_n_29777) );
in01s01 FE_OCP_DRV_C1463_n_19751 ( .a(n_19751), .o(FE_OCP_DRV_N1463_n_19751) );
in01s01 FE_OCP_DRV_C1464_n_19751 ( .a(FE_OCP_DRV_N1463_n_19751), .o(FE_OCP_DRV_N1464_n_19751) );
in01s01 FE_OCP_DRV_C1465_n_29860 ( .a(n_29860), .o(FE_OCP_DRV_N1465_n_29860) );
in01s01 FE_OCP_DRV_C1466_n_29860 ( .a(FE_OCP_DRV_N1465_n_29860), .o(FE_OCP_DRV_N1466_n_29860) );
in01s01 FE_OCP_DRV_C1467_n_28775 ( .a(n_28775), .o(FE_OCP_DRV_N1467_n_28775) );
in01s01 FE_OCP_DRV_C1468_n_28775 ( .a(FE_OCP_DRV_N1467_n_28775), .o(FE_OCP_DRV_N1468_n_28775) );
in01s01 FE_OCP_DRV_C1469_n_25022 ( .a(n_25022), .o(FE_OCP_DRV_N1469_n_25022) );
in01s01 FE_OCP_DRV_C1470_n_25022 ( .a(FE_OCP_DRV_N1469_n_25022), .o(FE_OCP_DRV_N1470_n_25022) );
in01s01 FE_OCP_DRV_C1471_n_25044 ( .a(n_25044), .o(FE_OCP_DRV_N1471_n_25044) );
in01s01 FE_OCP_DRV_C1472_n_25044 ( .a(FE_OCP_DRV_N1471_n_25044), .o(FE_OCP_DRV_N1472_n_25044) );
in01s01 FE_OCP_DRV_C1473_n_23792 ( .a(n_23792), .o(FE_OCP_DRV_N1473_n_23792) );
in01s01 FE_OCP_DRV_C1474_n_23792 ( .a(FE_OCP_DRV_N1473_n_23792), .o(FE_OCP_DRV_N1474_n_23792) );
in01s01 FE_OCP_DRV_C1475_n_23887 ( .a(n_23887), .o(FE_OCP_DRV_N1475_n_23887) );
in01s01 FE_OCP_DRV_C1476_n_23887 ( .a(FE_OCP_DRV_N1475_n_23887), .o(FE_OCP_DRV_N1476_n_23887) );
in01s01 FE_OCP_DRV_C1477_n_35106 ( .a(n_35106), .o(FE_OCP_DRV_N1477_n_35106) );
in01s01 FE_OCP_DRV_C1478_n_35106 ( .a(FE_OCP_DRV_N1477_n_35106), .o(FE_OCP_DRV_N1478_n_35106) );
in01s01 FE_OCP_DRV_C1479_n_30917 ( .a(n_30917), .o(FE_OCP_DRV_N1479_n_30917) );
in01s01 FE_OCP_DRV_C1480_n_30917 ( .a(FE_OCP_DRV_N1479_n_30917), .o(FE_OCP_DRV_N1480_n_30917) );
in01s01 FE_OCP_DRV_C1481_n_26296 ( .a(n_26296), .o(FE_OCP_DRV_N1481_n_26296) );
in01s01 FE_OCP_DRV_C1482_n_26296 ( .a(FE_OCP_DRV_N1481_n_26296), .o(FE_OCP_DRV_N1482_n_26296) );
in01s01 FE_OCP_DRV_C1483_n_35427 ( .a(n_35427), .o(FE_OCP_DRV_N1483_n_35427) );
in01s01 FE_OCP_DRV_C1484_n_35427 ( .a(FE_OCP_DRV_N1483_n_35427), .o(FE_OCP_DRV_N1484_n_35427) );
in01s01 FE_OCP_DRV_C1485_n_21639 ( .a(n_21639), .o(FE_OCP_DRV_N1485_n_21639) );
in01s01 FE_OCP_DRV_C1486_n_21639 ( .a(FE_OCP_DRV_N1485_n_21639), .o(FE_OCP_DRV_N1486_n_21639) );
in01s01 FE_OCP_DRV_C1487_n_24848 ( .a(n_24848), .o(FE_OCP_DRV_N1487_n_24848) );
in01s01 FE_OCP_DRV_C1488_n_24848 ( .a(FE_OCP_DRV_N1487_n_24848), .o(FE_OCP_DRV_N1488_n_24848) );
in01s01 FE_OCP_DRV_C1489_n_26656 ( .a(n_26656), .o(FE_OCP_DRV_N1489_n_26656) );
in01s01 FE_OCP_DRV_C1490_n_26656 ( .a(FE_OCP_DRV_N1489_n_26656), .o(FE_OCP_DRV_N1490_n_26656) );
in01s01 FE_OCP_DRV_C1491_n_31445 ( .a(n_31445), .o(FE_OCP_DRV_N1491_n_31445) );
in01s01 FE_OCP_DRV_C1492_n_31445 ( .a(FE_OCP_DRV_N1491_n_31445), .o(FE_OCP_DRV_N1492_n_31445) );
in01s01 FE_OCP_DRV_C1493_n_20059 ( .a(n_20059), .o(FE_OCP_DRV_N1493_n_20059) );
in01s01 FE_OCP_DRV_C1494_n_20059 ( .a(FE_OCP_DRV_N1493_n_20059), .o(FE_OCP_DRV_N1494_n_20059) );
in01s01 FE_OCP_DRV_C1495_n_31473 ( .a(n_31473), .o(FE_OCP_DRV_N1495_n_31473) );
in01s01 FE_OCP_DRV_C1496_n_31473 ( .a(FE_OCP_DRV_N1495_n_31473), .o(FE_OCP_DRV_N1496_n_31473) );
in01s01 FE_OCP_DRV_C1497_n_34924 ( .a(n_34924), .o(FE_OCP_DRV_N1497_n_34924) );
in01s01 FE_OCP_DRV_C1498_n_34924 ( .a(FE_OCP_DRV_N1497_n_34924), .o(FE_OCP_DRV_N1498_n_34924) );
in01s01 FE_OCP_DRV_C1499_n_15605 ( .a(n_15605), .o(FE_OCP_DRV_N1499_n_15605) );
in01s01 FE_OCP_DRV_C1500_n_15605 ( .a(FE_OCP_DRV_N1499_n_15605), .o(FE_OCP_DRV_N1500_n_15605) );
in01s01 FE_OCP_DRV_C1501_n_15979 ( .a(n_15979), .o(FE_OCP_DRV_N1501_n_15979) );
in01s01 FE_OCP_DRV_C1502_n_15979 ( .a(FE_OCP_DRV_N1501_n_15979), .o(FE_OCP_DRV_N1502_n_15979) );
in01s01 FE_OCP_DRV_C1503_n_16106 ( .a(n_16106), .o(FE_OCP_DRV_N1503_n_16106) );
in01s01 FE_OCP_DRV_C1504_n_16106 ( .a(FE_OCP_DRV_N1503_n_16106), .o(FE_OCP_DRV_N1504_n_16106) );
in01s01 FE_OCP_DRV_C1505_n_16183 ( .a(n_16183), .o(FE_OCP_DRV_N1505_n_16183) );
in01s01 FE_OCP_DRV_C1506_n_16183 ( .a(FE_OCP_DRV_N1505_n_16183), .o(FE_OCP_DRV_N1506_n_16183) );
in01s01 FE_OCP_DRV_C1507_n_26491 ( .a(n_26491), .o(FE_OCP_DRV_N1507_n_26491) );
in01s01 FE_OCP_DRV_C1508_n_26491 ( .a(FE_OCP_DRV_N1507_n_26491), .o(FE_OCP_DRV_N1508_n_26491) );
in01s02 FE_OCP_DRV_C1509_n_36387 ( .a(n_36387), .o(FE_OCP_DRV_N1509_n_36387) );
in01s01 FE_OCP_DRV_C1510_n_36387 ( .a(FE_OCP_DRV_N1509_n_36387), .o(FE_OCP_DRV_N1510_n_36387) );
in01s01 FE_OCP_DRV_C1511_n_26582 ( .a(n_26582), .o(FE_OCP_DRV_N1511_n_26582) );
in01s01 FE_OCP_DRV_C1512_n_26582 ( .a(FE_OCP_DRV_N1511_n_26582), .o(FE_OCP_DRV_N1512_n_26582) );
in01s01 FE_OCP_DRV_C1513_n_26786 ( .a(n_26786), .o(FE_OCP_DRV_N1513_n_26786) );
in01s01 FE_OCP_DRV_C1514_n_26786 ( .a(FE_OCP_DRV_N1513_n_26786), .o(FE_OCP_DRV_N1514_n_26786) );
in01s01 FE_OCP_DRV_C1515_n_21706 ( .a(n_21706), .o(FE_OCP_DRV_N1515_n_21706) );
in01s01 FE_OCP_DRV_C1516_n_21706 ( .a(FE_OCP_DRV_N1515_n_21706), .o(FE_OCP_DRV_N1516_n_21706) );
in01s01 FE_OCP_DRV_C1517_n_21851 ( .a(n_21851), .o(FE_OCP_DRV_N1517_n_21851) );
in01s01 FE_OCP_DRV_C1518_n_21851 ( .a(FE_OCP_DRV_N1517_n_21851), .o(FE_OCP_DRV_N1518_n_21851) );
in01s01 FE_OCP_DRV_C1519_n_26761 ( .a(n_26761), .o(FE_OCP_DRV_N1519_n_26761) );
in01s01 FE_OCP_DRV_C1520_n_26761 ( .a(FE_OCP_DRV_N1519_n_26761), .o(FE_OCP_DRV_N1520_n_26761) );
in01s01 FE_OCP_DRV_C1521_n_26807 ( .a(n_26807), .o(FE_OCP_DRV_N1521_n_26807) );
in01s01 FE_OCP_DRV_C1522_n_26807 ( .a(FE_OCP_DRV_N1521_n_26807), .o(FE_OCP_DRV_N1522_n_26807) );
in01s01 FE_OCP_DRV_C1523_n_31435 ( .a(FE_OFN5077_n_31435), .o(FE_OCP_DRV_N1523_n_31435) );
in01s01 FE_OCP_DRV_C1524_n_31435 ( .a(FE_OCP_DRV_N1523_n_31435), .o(FE_OCP_DRV_N1524_n_31435) );
in01s01 FE_OCP_DRV_C1760_n_20145 ( .a(n_20145), .o(FE_OCP_DRV_N1760_n_20145) );
in01s01 FE_OCP_DRV_C1761_n_20145 ( .a(FE_OCP_DRV_N1760_n_20145), .o(FE_OCP_DRV_N1761_n_20145) );
in01s01 FE_OCP_DRV_C1879_n_28164 ( .a(n_28164), .o(FE_OCP_DRV_N1879_n_28164) );
in01s01 FE_OCP_DRV_C1880_n_28164 ( .a(FE_OCP_DRV_N1879_n_28164), .o(FE_OCP_DRV_N1880_n_28164) );
in01s01 FE_OCP_DRV_C1881_n_32758 ( .a(n_32758), .o(FE_OCP_DRV_N1881_n_32758) );
in01s01 FE_OCP_DRV_C1882_n_32758 ( .a(FE_OCP_DRV_N1881_n_32758), .o(FE_OCP_DRV_N1882_n_32758) );
in01s01 FE_OCP_DRV_C1883_n_24361 ( .a(n_24361), .o(FE_OCP_DRV_N1883_n_24361) );
in01s01 FE_OCP_DRV_C1884_n_24361 ( .a(FE_OCP_DRV_N1883_n_24361), .o(FE_OCP_DRV_N1884_n_24361) );
in01s01 FE_OCP_DRV_C1885_n_34009 ( .a(n_34009), .o(FE_OCP_DRV_N1885_n_34009) );
in01s01 FE_OCP_DRV_C1886_n_34009 ( .a(FE_OCP_DRV_N1885_n_34009), .o(FE_OCP_DRV_N1886_n_34009) );
in01s01 FE_OCP_DRV_C1887_n_33756 ( .a(n_33756), .o(FE_OCP_DRV_N1887_n_33756) );
in01s01 FE_OCP_DRV_C1888_n_33756 ( .a(FE_OCP_DRV_N1887_n_33756), .o(FE_OCP_DRV_N1888_n_33756) );
in01s01 FE_OCP_DRV_C1889_n_29317 ( .a(n_29317), .o(FE_OCP_DRV_N1889_n_29317) );
in01s01 FE_OCP_DRV_C1891_n_29573 ( .a(n_29573), .o(FE_OCP_DRV_N1891_n_29573) );
in01s01 FE_OCP_DRV_C1892_n_29573 ( .a(FE_OCP_DRV_N1891_n_29573), .o(FE_OCP_DRV_N1892_n_29573) );
in01s01 FE_OCP_DRV_C1893_n_33221 ( .a(n_33221), .o(FE_OCP_DRV_N1893_n_33221) );
in01s01 FE_OCP_DRV_C1894_n_33221 ( .a(FE_OCP_DRV_N1893_n_33221), .o(FE_OCP_DRV_N1894_n_33221) );
in01s01 FE_OCP_DRV_C1895_n_19855 ( .a(n_19855), .o(FE_OCP_DRV_N1895_n_19855) );
in01s01 FE_OCP_DRV_C1896_n_19855 ( .a(FE_OCP_DRV_N1895_n_19855), .o(FE_OCP_DRV_N1896_n_19855) );
in01s01 FE_OCP_DRV_C1897_n_18287 ( .a(FE_OFN5072_n_18287), .o(FE_OCP_DRV_N1897_n_18287) );
in01s01 FE_OCP_DRV_C1898_n_18287 ( .a(FE_OCP_DRV_N1897_n_18287), .o(FE_OCP_DRV_N1898_n_18287) );
in01s01 FE_OCP_DRV_C1899_n_23668 ( .a(n_23668), .o(FE_OCP_DRV_N1899_n_23668) );
in01s01 FE_OCP_DRV_C1900_n_23668 ( .a(FE_OCP_DRV_N1899_n_23668), .o(FE_OCP_DRV_N1900_n_23668) );
in01s06 FE_OCP_DRV_C3493_n_40837 ( .a(n_40837), .o(FE_OCP_DRV_N3493_n_40837) );
in01s06 FE_OCP_DRV_C3494_n_40837 ( .a(FE_OCP_DRV_N3493_n_40837), .o(FE_OCP_DRV_N3494_n_40837) );
in01s01 FE_OCP_DRV_C3495_n_33156 ( .a(n_33156), .o(FE_OCP_DRV_N3495_n_33156) );
in01s01 FE_OCP_DRV_C3496_n_33156 ( .a(FE_OCP_DRV_N3495_n_33156), .o(FE_OCP_DRV_N3496_n_33156) );
in01s01 FE_OCP_DRV_C3497_n_7233 ( .a(n_7233), .o(FE_OCP_DRV_N3497_n_7233) );
in01s01 FE_OCP_DRV_C3498_n_7233 ( .a(FE_OCP_DRV_N3497_n_7233), .o(FE_OCP_DRV_N3498_n_7233) );
in01s01 FE_OCP_DRV_C3499_n_7204 ( .a(n_7204), .o(FE_OCP_DRV_N3499_n_7204) );
in01s01 FE_OCP_DRV_C3500_n_7204 ( .a(FE_OCP_DRV_N3499_n_7204), .o(FE_OCP_DRV_N3500_n_7204) );
in01s01 FE_OCP_DRV_C3501_n_29140 ( .a(n_29140), .o(FE_OCP_DRV_N3501_n_29140) );
in01s01 FE_OCP_DRV_C3502_n_29140 ( .a(FE_OCP_DRV_N3501_n_29140), .o(FE_OCP_DRV_N3502_n_29140) );
in01s01 FE_OCP_DRV_C3504_FE_OCP_RBN1807_n_13010 ( .a(FE_OCP_DRV_N4501_FE_OCP_RBN1807_n_13010), .o(FE_OCP_DRV_N3504_FE_OCP_RBN1807_n_13010) );
in01s01 FE_OCP_DRV_C3505_n_8189 ( .a(n_8189), .o(FE_OCP_DRV_N3505_n_8189) );
in01s02 FE_OCP_DRV_C3506_n_8189 ( .a(FE_OCP_DRV_N3505_n_8189), .o(FE_OCP_DRV_N3506_n_8189) );
in01s01 FE_OCP_DRV_C3507_n_13329 ( .a(n_13329), .o(FE_OCP_DRV_N3507_n_13329) );
in01s01 FE_OCP_DRV_C3508_n_13329 ( .a(FE_OCP_DRV_N3507_n_13329), .o(FE_OCP_DRV_N3508_n_13329) );
in01s01 FE_OCP_DRV_C3509_n_35315 ( .a(n_35315), .o(FE_OCP_DRV_N3509_n_35315) );
in01s01 FE_OCP_DRV_C3510_n_35315 ( .a(FE_OCP_DRV_N3509_n_35315), .o(FE_OCP_DRV_N3510_n_35315) );
in01s01 FE_OCP_DRV_C3511_n_30318 ( .a(n_30318), .o(FE_OCP_DRV_N3511_n_30318) );
in01s01 FE_OCP_DRV_C3512_n_30318 ( .a(FE_OCP_DRV_N3511_n_30318), .o(FE_OCP_DRV_N3512_n_30318) );
in01s01 FE_OCP_DRV_C3513_n_14650 ( .a(n_14650), .o(FE_OCP_DRV_N3513_n_14650) );
in01s02 FE_OCP_DRV_C3514_n_14650 ( .a(FE_OCP_DRV_N3513_n_14650), .o(FE_OCP_DRV_N3514_n_14650) );
in01s01 FE_OCP_DRV_C3515_n_31504 ( .a(n_31504), .o(FE_OCP_DRV_N3515_n_31504) );
in01s01 FE_OCP_DRV_C3516_n_31504 ( .a(FE_OCP_DRV_N3515_n_31504), .o(FE_OCP_DRV_N3516_n_31504) );
in01s01 FE_OCP_DRV_C3517_n_39785 ( .a(n_39785), .o(FE_OCP_DRV_N3517_n_39785) );
in01s01 FE_OCP_DRV_C3518_n_39785 ( .a(FE_OCP_DRV_N3517_n_39785), .o(FE_OCP_DRV_N3518_n_39785) );
in01s02 FE_OCP_DRV_C3519_n_43153 ( .a(n_43153), .o(FE_OCP_DRV_N3519_n_43153) );
in01m04 FE_OCP_DRV_C3520_n_43153 ( .a(FE_OCP_DRV_N3519_n_43153), .o(FE_OCP_DRV_N3520_n_43153) );
in01s02 FE_OCP_DRV_C3521_n_43538 ( .a(n_43538), .o(FE_OCP_DRV_N3521_n_43538) );
in01s04 FE_OCP_DRV_C3522_n_43538 ( .a(FE_OCP_DRV_N3521_n_43538), .o(FE_OCP_DRV_N3522_n_43538) );
in01s01 FE_OCP_DRV_C3523_FE_OCP_RBN3021_n_15319 ( .a(FE_OCP_RBN3021_n_15319), .o(FE_OCP_DRV_N3523_FE_OCP_RBN3021_n_15319) );
in01s01 FE_OCP_DRV_C3524_FE_OCP_RBN3021_n_15319 ( .a(FE_OCP_DRV_N3523_FE_OCP_RBN3021_n_15319), .o(FE_OCP_DRV_N3524_FE_OCP_RBN3021_n_15319) );
in01s01 FE_OCP_DRV_C3525_n_17031 ( .a(n_17031), .o(FE_OCP_DRV_N3525_n_17031) );
in01s01 FE_OCP_DRV_C3526_n_17031 ( .a(FE_OCP_DRV_N3525_n_17031), .o(FE_OCP_DRV_N3526_n_17031) );
in01s01 FE_OCP_DRV_C3527_n_17071 ( .a(n_17071), .o(FE_OCP_DRV_N3527_n_17071) );
in01s01 FE_OCP_DRV_C3528_n_17071 ( .a(FE_OCP_DRV_N3527_n_17071), .o(FE_OCP_DRV_N3528_n_17071) );
in01s01 FE_OCP_DRV_C3533_n_18559 ( .a(n_18559), .o(FE_OCP_DRV_N3533_n_18559) );
in01s01 FE_OCP_DRV_C3534_n_18559 ( .a(FE_OCP_DRV_N3533_n_18559), .o(FE_OCP_DRV_N3534_n_18559) );
in01s01 FE_OCP_DRV_C3535_n_19053 ( .a(n_19053), .o(FE_OCP_DRV_N3535_n_19053) );
in01s01 FE_OCP_DRV_C3536_n_19053 ( .a(FE_OCP_DRV_N3535_n_19053), .o(FE_OCP_DRV_N3536_n_19053) );
in01s01 FE_OCP_DRV_C3537_n_21763 ( .a(n_21763), .o(FE_OCP_DRV_N3537_n_21763) );
in01s01 FE_OCP_DRV_C3538_n_21763 ( .a(FE_OCP_DRV_N3537_n_21763), .o(FE_OCP_DRV_N3538_n_21763) );
in01s01 FE_OCP_DRV_C3539_n_20146 ( .a(n_20146), .o(FE_OCP_DRV_N3539_n_20146) );
in01s01 FE_OCP_DRV_C3540_n_20146 ( .a(FE_OCP_DRV_N3539_n_20146), .o(FE_OCP_DRV_N3540_n_20146) );
in01s01 FE_OCP_DRV_C4499_n_13785 ( .a(n_13785), .o(FE_OCP_DRV_N4499_n_13785) );
in01s02 FE_OCP_DRV_C4500_n_13785 ( .a(FE_OCP_DRV_N4499_n_13785), .o(FE_OCP_DRV_N4500_n_13785) );
in01s01 FE_OCP_DRV_C4501_FE_OCP_RBN1807_n_13010 ( .a(FE_OCP_RBN1807_n_13010), .o(FE_OCP_DRV_N4501_FE_OCP_RBN1807_n_13010) );
in01s01 FE_OCP_DRV_C4502_FE_OCP_RBN1807_n_13010 ( .a(FE_OCP_DRV_N4501_FE_OCP_RBN1807_n_13010), .o(FE_OCP_DRV_N4502_FE_OCP_RBN1807_n_13010) );
in01s01 FE_OCP_DRV_C4503_n_28888 ( .a(n_28888), .o(FE_OCP_DRV_N4503_n_28888) );
in01s01 FE_OCP_DRV_C4505_n_13476 ( .a(n_13476), .o(FE_OCP_DRV_N4505_n_13476) );
in01s02 FE_OCP_DRV_C4507_n_15099 ( .a(n_15099), .o(FE_OCP_DRV_N4507_n_15099) );
in01s04 FE_OCP_DRV_C4508_n_15099 ( .a(FE_OCP_DRV_N4507_n_15099), .o(FE_OCP_DRV_N4508_n_15099) );
in01s01 FE_OCP_DRV_C4510_n_21343 ( .a(FE_OCPN4514_n_21343), .o(FE_OCP_DRV_N4510_n_21343) );
in01s01 FE_OCP_DRV_C5140_n_29375 ( .a(n_29375), .o(FE_OCP_DRV_N5140_n_29375) );
in01s01 FE_OCP_DRV_C5141_n_29375 ( .a(FE_OCP_DRV_N5140_n_29375), .o(FE_OCP_DRV_N5141_n_29375) );
in01s01 FE_OCP_DRV_C5142_n_28426 ( .a(n_28426), .o(FE_OCP_DRV_N5142_n_28426) );
in01s01 FE_OCP_DRV_C5143_n_28426 ( .a(FE_OCP_DRV_N5142_n_28426), .o(FE_OCP_DRV_N5143_n_28426) );
in01s01 FE_OCP_DRV_C5144_n_28349 ( .a(n_28349), .o(FE_OCP_DRV_N5144_n_28349) );
in01s01 FE_OCP_DRV_C5145_n_28349 ( .a(FE_OCP_DRV_N5144_n_28349), .o(FE_OCP_DRV_N5145_n_28349) );
in01s01 FE_OCP_DRV_C5146_n_29765 ( .a(n_29765), .o(FE_OCP_DRV_N5146_n_29765) );
in01s01 FE_OCP_DRV_C5147_n_29765 ( .a(FE_OCP_DRV_N5146_n_29765), .o(FE_OCP_DRV_N5147_n_29765) );
in01s01 FE_OCP_DRV_C5148_n_31125 ( .a(n_31125), .o(FE_OCP_DRV_N5148_n_31125) );
in01s01 FE_OCP_DRV_C5149_n_31125 ( .a(FE_OCP_DRV_N5148_n_31125), .o(FE_OCP_DRV_N5149_n_31125) );
in01s01 FE_OCP_DRV_C5150_n_31264 ( .a(n_31264), .o(FE_OCP_DRV_N5150_n_31264) );
in01s01 FE_OCP_DRV_C5151_n_31264 ( .a(FE_OCP_DRV_N5150_n_31264), .o(FE_OCP_DRV_N5151_n_31264) );
in01s01 FE_OCP_DRV_C5152_n_31164 ( .a(n_31164), .o(FE_OCP_DRV_N5152_n_31164) );
in01s01 FE_OCP_DRV_C5153_n_31164 ( .a(FE_OCP_DRV_N5152_n_31164), .o(FE_OCP_DRV_N5153_n_31164) );
in01s01 FE_OCP_DRV_C5154_n_31206 ( .a(n_31206), .o(FE_OCP_DRV_N5154_n_31206) );
in01s01 FE_OCP_DRV_C5155_n_31206 ( .a(FE_OCP_DRV_N5154_n_31206), .o(FE_OCP_DRV_N5155_n_31206) );
in01s01 FE_OCP_DRV_C5156_n_25100 ( .a(n_25100), .o(FE_OCP_DRV_N5156_n_25100) );
in01s01 FE_OCP_DRV_C5157_n_25100 ( .a(FE_OCP_DRV_N5156_n_25100), .o(FE_OCP_DRV_N5157_n_25100) );
in01s01 FE_OCP_DRV_C5158_n_26801 ( .a(n_26801), .o(FE_OCP_DRV_N5158_n_26801) );
in01s01 FE_OCP_DRV_C5159_n_26801 ( .a(FE_OCP_DRV_N5158_n_26801), .o(FE_OCP_DRV_N5159_n_26801) );
in01s01 FE_OCP_DRV_C5160_n_30322 ( .a(n_30322), .o(FE_OCP_DRV_N5160_n_30322) );
in01s01 FE_OCP_DRV_C5161_n_30322 ( .a(FE_OCP_DRV_N5160_n_30322), .o(FE_OCP_DRV_N5161_n_30322) );
in01s01 FE_OCP_DRV_C5303_n_29892 ( .a(n_29892), .o(FE_OCP_DRV_N5303_n_29892) );
in01s01 FE_OCP_DRV_C5304_n_29892 ( .a(FE_OCP_DRV_N5303_n_29892), .o(FE_OCP_DRV_N5304_n_29892) );
in01s01 FE_OCP_DRV_C5353_n_18860 ( .a(n_18860), .o(FE_OCP_DRV_N5353_n_18860) );
in01s01 FE_OCP_DRV_C5354_n_18860 ( .a(FE_OCP_DRV_N5353_n_18860), .o(FE_OCP_DRV_N5354_n_18860) );
in01s01 FE_OCP_DRV_C5355_n_19010 ( .a(n_19010), .o(FE_OCP_DRV_N5355_n_19010) );
in01s01 FE_OCP_DRV_C5356_n_19010 ( .a(FE_OCP_DRV_N5355_n_19010), .o(FE_OCP_DRV_N5356_n_19010) );
in01s01 FE_OCP_DRV_C5357_n_12436 ( .a(n_12436), .o(FE_OCP_DRV_N5357_n_12436) );
in01s01 FE_OCP_DRV_C5358_n_12436 ( .a(FE_OCP_DRV_N5357_n_12436), .o(FE_OCP_DRV_N5358_n_12436) );
in01s01 FE_OCP_DRV_C5359_n_13495 ( .a(n_13495), .o(FE_OCP_DRV_N5359_n_13495) );
in01s01 FE_OCP_DRV_C5360_n_13495 ( .a(FE_OCP_DRV_N5359_n_13495), .o(FE_OCP_DRV_N5360_n_13495) );
in01s01 FE_OCP_DRV_C5361_n_21732 ( .a(n_21732), .o(FE_OCP_DRV_N5361_n_21732) );
in01s01 FE_OCP_DRV_C5362_n_21732 ( .a(FE_OCP_DRV_N5361_n_21732), .o(FE_OCP_DRV_N5362_n_21732) );
in01s01 FE_OCP_DRV_C6260_n_37471 ( .a(n_37471), .o(FE_OCP_DRV_N6260_n_37471) );
in01s01 FE_OCP_DRV_C6261_n_37471 ( .a(FE_OCP_DRV_N6260_n_37471), .o(FE_OCP_DRV_N6261_n_37471) );
in01s01 FE_OCP_DRV_C6262_FE_OCP_RBN5603_n_29056 ( .a(FE_OCP_RBN5603_n_29056), .o(FE_OCP_DRV_N6262_FE_OCP_RBN5603_n_29056) );
in01s01 FE_OCP_DRV_C6263_FE_OCP_RBN5603_n_29056 ( .a(FE_OCP_DRV_N6262_FE_OCP_RBN5603_n_29056), .o(FE_OCP_DRV_N6263_FE_OCP_RBN5603_n_29056) );
in01s01 FE_OCP_DRV_C6264_n_9014 ( .a(n_9014), .o(FE_OCP_DRV_N6264_n_9014) );
in01s01 FE_OCP_DRV_C6266_FE_OCP_RBN1823_n_19434 ( .a(FE_OCP_RBN1823_n_19434), .o(FE_OCP_DRV_N6266_FE_OCP_RBN1823_n_19434) );
in01s01 FE_OCP_DRV_C6270_n_13264 ( .a(n_13264), .o(FE_OCP_DRV_N6270_n_13264) );
in01s01 FE_OCP_DRV_C6271_n_13264 ( .a(FE_OCP_DRV_N6270_n_13264), .o(FE_OCP_DRV_N6271_n_13264) );
in01s01 FE_OCP_DRV_C6272_n_13330 ( .a(n_13330), .o(FE_OCP_DRV_N6272_n_13330) );
in01s01 FE_OCP_DRV_C6273_n_13330 ( .a(FE_OCP_DRV_N6272_n_13330), .o(FE_OCP_DRV_N6273_n_13330) );
in01s01 FE_OCP_DRV_C6274_n_28582 ( .a(n_28582), .o(FE_OCP_DRV_N6274_n_28582) );
in01s01 FE_OCP_DRV_C6275_n_28582 ( .a(FE_OCP_DRV_N6274_n_28582), .o(FE_OCP_DRV_N6275_n_28582) );
in01s01 FE_OCP_DRV_C6884_n_28829 ( .a(FE_OCP_DRV_N6885_n_28829), .o(FE_OCP_DRV_N6884_n_28829) );
in01s01 FE_OCP_DRV_C6885_n_28829 ( .a(n_28829), .o(FE_OCP_DRV_N6885_n_28829) );
in01s01 FE_OCP_DRV_C6888_n_33945 ( .a(n_33945), .o(FE_OCP_DRV_N6888_n_33945) );
in01s01 FE_OCP_DRV_C6889_n_33945 ( .a(FE_OCP_DRV_N6888_n_33945), .o(FE_OCP_DRV_N6889_n_33945) );
in01s01 FE_OCP_DRV_C6890_n_34296 ( .a(n_34296), .o(FE_OCP_DRV_N6890_n_34296) );
in01s01 FE_OCP_DRV_C6891_n_34296 ( .a(FE_OCP_DRV_N6890_n_34296), .o(FE_OCP_DRV_N6891_n_34296) );
in01s01 FE_OCP_DRV_C6892_FE_OCPN6281_n_30612 ( .a(FE_OCPN6281_n_30612), .o(FE_OCP_DRV_N6892_FE_OCPN6281_n_30612) );
in01s01 FE_OCP_DRV_C6893_FE_OCPN6281_n_30612 ( .a(FE_OCP_DRV_N6892_FE_OCPN6281_n_30612), .o(FE_OCP_DRV_N6893_FE_OCPN6281_n_30612) );
in01m04 FE_OCP_DRV_C6894_n_15391 ( .a(n_15391), .o(FE_OCP_DRV_N6894_n_15391) );
in01f04 FE_OCP_DRV_C6895_n_15391 ( .a(FE_OCP_DRV_N6894_n_15391), .o(FE_OCP_DRV_N6895_n_15391) );
in01s01 FE_OCP_DRV_C6896_FE_OCPN1679_n_27315 ( .a(FE_OCPN1679_n_27315), .o(FE_OCP_DRV_N6896_FE_OCPN1679_n_27315) );
in01s01 FE_OCP_DRV_C6897_FE_OCPN1679_n_27315 ( .a(FE_OCP_DRV_N6896_FE_OCPN1679_n_27315), .o(FE_OCP_DRV_N6897_FE_OCPN1679_n_27315) );
in01s01 FE_OCP_DRV_C6898_FE_OCPN5276_n_23590 ( .a(FE_OCPN5276_n_23590), .o(FE_OCP_DRV_N6898_FE_OCPN5276_n_23590) );
in01s01 FE_OCP_DRV_C6899_FE_OCPN5276_n_23590 ( .a(FE_OCP_DRV_N6898_FE_OCPN5276_n_23590), .o(FE_OCP_DRV_N6899_FE_OCPN5276_n_23590) );
in01s01 FE_OCP_DRV_C6902_n_19354 ( .a(n_19354), .o(FE_OCP_DRV_N6902_n_19354) );
in01s01 FE_OCP_DRV_C6903_n_19354 ( .a(FE_OCP_DRV_N6902_n_19354), .o(FE_OCP_DRV_N6903_n_19354) );
in01s01 FE_OCP_DRV_C6904_n_33945 ( .a(n_33945), .o(FE_OCP_DRV_N6904_n_33945) );
in01s01 FE_OCP_DRV_C6906_n_34096 ( .a(n_34096), .o(FE_OCP_DRV_N6906_n_34096) );
in01s01 FE_OCP_DRV_C6907_n_34096 ( .a(FE_OCP_DRV_N6906_n_34096), .o(FE_OCP_DRV_N6907_n_34096) );
in01s01 FE_OCP_DRV_C7074_n_7116 ( .a(n_7116), .o(FE_OCP_DRV_N7074_n_7116) );
in01s01 FE_OCP_DRV_C7076_n_10105 ( .a(n_10105), .o(FE_OCP_DRV_N7076_n_10105) );
in01s01 FE_OCP_DRV_C7077_n_10105 ( .a(FE_OCP_DRV_N7076_n_10105), .o(FE_OCP_DRV_N7077_n_10105) );
in01s01 FE_OCP_DRV_C7078_n_8992 ( .a(n_8992), .o(FE_OCP_DRV_N7078_n_8992) );
in01s01 FE_OCP_DRV_C7079_n_8992 ( .a(FE_OCP_DRV_N7078_n_8992), .o(FE_OCP_DRV_N7079_n_8992) );
in01s01 FE_OCP_DRV_C7080_n_27130 ( .a(n_27130), .o(FE_OCP_DRV_N7080_n_27130) );
in01s01 FE_OCP_DRV_C7081_n_27130 ( .a(FE_OCP_DRV_N7080_n_27130), .o(FE_OCP_DRV_N7081_n_27130) );
in01s02 FE_OCP_RBC1001_n_24079 ( .a(n_24079), .o(FE_OCP_RBN1001_n_24079) );
in01s01 FE_OCP_RBC1002_n_24079 ( .a(FE_OCP_RBN1001_n_24079), .o(FE_OCP_RBN1002_n_24079) );
in01s01 FE_OCP_RBC1003_n_24079 ( .a(FE_OCP_RBN1002_n_24079), .o(FE_OCP_RBN1003_n_24079) );
in01m04 FE_OCP_RBC1004_n_25545 ( .a(n_25545), .o(FE_OCP_RBN1004_n_25545) );
in01m06 FE_OCP_RBC1005_n_25545 ( .a(FE_OCP_RBN1004_n_25545), .o(FE_OCP_RBN1005_n_25545) );
in01m02 FE_OCP_RBC1006_n_24094 ( .a(n_24094), .o(FE_OCP_RBN1006_n_24094) );
in01m02 FE_OCP_RBC1007_n_24175 ( .a(n_24175), .o(FE_OCP_RBN1007_n_24175) );
in01s01 FE_OCP_RBC1009_n_24175 ( .a(FE_OCP_RBN2622_n_24175), .o(FE_OCP_RBN1009_n_24175) );
in01s01 FE_OCP_RBC1010_n_24175 ( .a(FE_OCP_RBN2622_n_24175), .o(FE_OCP_RBN1010_n_24175) );
in01f02 FE_OCP_RBC1011_n_24246 ( .a(n_24246), .o(FE_OCP_RBN1011_n_24246) );
in01m02 FE_OCP_RBC1012_n_25826 ( .a(n_25826), .o(FE_OCP_RBN1012_n_25826) );
in01s01 FE_OCP_RBC1013_n_25826 ( .a(n_25826), .o(FE_OCP_RBN1013_n_25826) );
in01s01 FE_OCP_RBC1014_n_25826 ( .a(FE_OCP_RBN1013_n_25826), .o(FE_OCP_RBN1014_n_25826) );
in01s01 FE_OCP_RBC1015_n_25826 ( .a(FE_OCP_RBN1014_n_25826), .o(FE_OCP_RBN1015_n_25826) );
in01s02 FE_OCP_RBC1016_n_13601 ( .a(n_13601), .o(FE_OCP_RBN1016_n_13601) );
in01s01 FE_OCP_RBC1017_n_24165 ( .a(n_24165), .o(FE_OCP_RBN1017_n_24165) );
in01f02 FE_OCP_RBC1018_n_24165 ( .a(n_24165), .o(FE_OCP_RBN1018_n_24165) );
in01s02 FE_OCP_RBC1019_n_24165 ( .a(FE_OCP_RBN1017_n_24165), .o(FE_OCP_RBN1019_n_24165) );
in01s02 FE_OCP_RBC1020_n_24181 ( .a(n_24181), .o(FE_OCP_RBN1020_n_24181) );
in01s01 FE_OCP_RBC1021_n_24181 ( .a(FE_OCP_RBN1020_n_24181), .o(FE_OCP_RBN1021_n_24181) );
in01s01 FE_OCP_RBC1022_n_24181 ( .a(FE_OCP_RBN1021_n_24181), .o(FE_OCP_RBN1022_n_24181) );
in01s01 FE_OCP_RBC1023_n_24125 ( .a(n_24125), .o(FE_OCP_RBN1023_n_24125) );
in01s01 FE_OCP_RBC1024_n_24125 ( .a(n_24125), .o(FE_OCP_RBN1024_n_24125) );
in01s03 FE_OCP_RBC1025_n_17417 ( .a(n_17417), .o(FE_OCP_RBN1025_n_17417) );
in01s03 FE_OCP_RBC1026_n_17417 ( .a(FE_OCP_RBN1025_n_17417), .o(FE_OCP_RBN1026_n_17417) );
in01s01 FE_OCP_RBC1027_n_17417 ( .a(FE_OCP_RBN1025_n_17417), .o(FE_OCP_RBN1027_n_17417) );
in01s01 FE_OCP_RBC1028_n_17417 ( .a(FE_OCP_RBN1027_n_17417), .o(FE_OCP_RBN1028_n_17417) );
in01s01 FE_OCP_RBC1032_n_25844 ( .a(FE_OCP_RBN1172_n_25817), .o(FE_OCP_RBN1032_n_25844) );
in01s01 FE_OCP_RBC1034_n_25844 ( .a(FE_OCP_RBN1032_n_25844), .o(FE_OCP_RBN1034_n_25844) );
in01s02 FE_OCP_RBC1035_FE_RN_557_0 ( .a(FE_RN_557_0), .o(FE_OCP_RBN1035_FE_RN_557_0) );
in01f02 FE_OCP_RBC1036_FE_RN_557_0 ( .a(FE_RN_557_0), .o(FE_OCP_RBN1036_FE_RN_557_0) );
in01s01 FE_OCP_RBC1037_n_45533 ( .a(n_45533), .o(FE_OCP_RBN1037_n_45533) );
in01s01 FE_OCP_RBC1038_n_45533 ( .a(FE_OCP_RBN1037_n_45533), .o(FE_OCP_RBN1038_n_45533) );
in01s01 FE_OCP_RBC1039_n_45533 ( .a(FE_OCP_RBN1038_n_45533), .o(FE_OCP_RBN1039_n_45533) );
in01s02 FE_OCP_RBC1040_n_26158 ( .a(n_26158), .o(FE_OCP_RBN1040_n_26158) );
in01s01 FE_OCP_RBC1105_n_18746 ( .a(n_18746), .o(FE_OCP_RBN1105_n_18746) );
in01s06 FE_OCP_RBC1109_n_44061 ( .a(FE_OCP_RBN5179_n_44061), .o(FE_OCP_RBN1109_n_44061) );
in01s02 FE_OCP_RBC1118_delay_xor_ln22_unr15_stage6_stallmux_q_0_ ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_0_), .o(FE_OCP_RBN1118_delay_xor_ln22_unr15_stage6_stallmux_q_0_) );
in01s40 FE_OCP_RBC1120_delay_xor_ln22_unr12_stage5_stallmux_q_2_ ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_2_), .o(FE_OCP_RBN1120_delay_xor_ln22_unr12_stage5_stallmux_q_2_) );
in01s10 FE_OCP_RBC1121_delay_xor_ln22_unr12_stage5_stallmux_q_2_ ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_2_), .o(FE_OCP_RBN1121_delay_xor_ln22_unr12_stage5_stallmux_q_2_) );
in01s01 FE_OCP_RBC1130_n_18918 ( .a(n_18918), .o(FE_OCP_RBN1130_n_18918) );
in01s04 FE_OCP_RBC1131_n_19077 ( .a(n_19077), .o(FE_OCP_RBN1131_n_19077) );
in01s01 FE_OCP_RBC1132_n_19077 ( .a(n_19077), .o(FE_OCP_RBN1132_n_19077) );
in01s01 FE_OCP_RBC1133_n_19077 ( .a(FE_OCP_RBN1132_n_19077), .o(FE_OCP_RBN1133_n_19077) );
in01s02 FE_OCP_RBC1134_n_19077 ( .a(FE_OCP_RBN1132_n_19077), .o(FE_OCP_RBN1134_n_19077) );
in01m02 FE_OCP_RBC1137_n_19270 ( .a(n_19270), .o(FE_OCP_RBN1137_n_19270) );
in01s01 FE_OCP_RBC1138_n_19270 ( .a(n_19270), .o(FE_OCP_RBN1138_n_19270) );
in01s01 FE_OCP_RBC1139_n_19270 ( .a(FE_OCPN1665_FE_OCP_RBN1138_n_19270), .o(FE_OCP_RBN1139_n_19270) );
in01s01 FE_OCP_RBC1140_n_19270 ( .a(FE_OCP_RBN1139_n_19270), .o(FE_OCP_RBN1140_n_19270) );
in01s01 FE_OCP_RBC1146_n_19353 ( .a(FE_OCP_RBN2064_n_19353), .o(FE_OCP_RBN1146_n_19353) );
in01s01 FE_OCP_RBC1150_n_18981 ( .a(FE_OCP_RBN7033_n_18981), .o(FE_OCP_RBN1150_n_18981) );
in01m02 FE_OCP_RBC1151_FE_RN_533_0 ( .a(FE_RN_533_0), .o(FE_OCP_RBN1151_FE_RN_533_0) );
in01s01 FE_OCP_RBC1152_n_20910 ( .a(n_20910), .o(FE_OCP_RBN1152_n_20910) );
in01s04 FE_OCP_RBC1153_n_20910 ( .a(n_20910), .o(FE_OCP_RBN1153_n_20910) );
in01s01 FE_OCP_RBC1157_n_20336 ( .a(FE_OCP_RBN7043_n_20336), .o(FE_OCP_RBN1157_n_20336) );
in01m04 FE_OCP_RBC1159_n_20763 ( .a(n_20763), .o(FE_OCP_RBN1159_n_20763) );
in01s01 FE_OCP_RBC1160_n_20763 ( .a(n_20763), .o(FE_OCP_RBN1160_n_20763) );
in01s01 FE_OCP_RBC1161_n_20763 ( .a(FE_OCP_RBN1160_n_20763), .o(FE_OCP_RBN1161_n_20763) );
in01s01 FE_OCP_RBC1162_n_20763 ( .a(FE_OCP_RBN1161_n_20763), .o(FE_OCP_RBN1162_n_20763) );
in01s01 FE_OCP_RBC1163_n_24471 ( .a(n_24471), .o(FE_OCP_RBN1163_n_24471) );
in01f02 FE_OCP_RBC1164_n_24471 ( .a(n_24471), .o(FE_OCP_RBN1164_n_24471) );
in01s01 FE_OCP_RBC1166_n_25889 ( .a(FE_OCP_RBN4367_n_25889), .o(FE_OCP_RBN1166_n_25889) );
in01s02 FE_OCP_RBC1170_n_21318 ( .a(n_21318), .o(FE_OCP_RBN1170_n_21318) );
in01s02 FE_OCP_RBC1171_n_25817 ( .a(n_25817), .o(FE_OCP_RBN1171_n_25817) );
in01s01 FE_OCP_RBC1172_n_25817 ( .a(FE_OCP_RBN1171_n_25817), .o(FE_OCP_RBN1172_n_25817) );
in01f04 FE_OCP_RBC1173_n_22476 ( .a(n_22476), .o(FE_OCP_RBN1173_n_22476) );
in01s02 FE_OCP_RBC1175_n_27593 ( .a(n_27593), .o(FE_OCP_RBN1175_n_27593) );
in01s06 FE_OCP_RBC1176_n_27593 ( .a(n_27593), .o(FE_OCP_RBN1176_n_27593) );
in01m02 FE_OCP_RBC1589_n_13460 ( .a(n_13460), .o(FE_OCP_RBN1589_n_13460) );
in01s01 FE_OCP_RBC1590_n_13557 ( .a(n_13557), .o(FE_OCP_RBN1590_n_13557) );
in01f02 FE_OCP_RBC1591_n_13557 ( .a(n_13557), .o(FE_OCP_RBN1591_n_13557) );
in01s02 FE_OCP_RBC1592_n_13557 ( .a(FE_OCP_RBN1590_n_13557), .o(FE_OCP_RBN1592_n_13557) );
in01s01 FE_OCP_RBC1593_n_13557 ( .a(FE_OCP_RBN1592_n_13557), .o(FE_OCP_RBN1593_n_13557) );
in01s01 FE_OCP_RBC1594_n_13557 ( .a(FE_OCP_RBN1592_n_13557), .o(FE_OCP_RBN1594_n_13557) );
in01f02 FE_OCP_RBC1595_n_14823 ( .a(n_14823), .o(FE_OCP_RBN1595_n_14823) );
in01s01 FE_OCP_RBC1596_n_14823 ( .a(n_14823), .o(FE_OCP_RBN1596_n_14823) );
in01f02 FE_OCP_RBC1597_n_14763 ( .a(n_14763), .o(FE_OCP_RBN1597_n_14763) );
in01s01 FE_OCP_RBC1598_n_14763 ( .a(n_14763), .o(FE_OCP_RBN1598_n_14763) );
in01s01 FE_OCP_RBC1599_n_14763 ( .a(FE_OCP_RBN1598_n_14763), .o(FE_OCP_RBN1599_n_14763) );
in01s01 FE_OCP_RBC1600_n_14763 ( .a(FE_OCP_RBN1599_n_14763), .o(FE_OCP_RBN1600_n_14763) );
in01f02 FE_OCP_RBC1601_n_14638 ( .a(n_14638), .o(FE_OCP_RBN1601_n_14638) );
in01s01 FE_OCP_RBC1602_n_14638 ( .a(n_14638), .o(FE_OCP_RBN1602_n_14638) );
in01s01 FE_OCP_RBC1603_n_20995 ( .a(n_20995), .o(FE_OCP_RBN1603_n_20995) );
in01s01 FE_OCP_RBC1604_n_20995 ( .a(n_20995), .o(FE_OCP_RBN1604_n_20995) );
in01m06 FE_OCP_RBC1803_n_32647 ( .a(n_32647), .o(FE_OCP_RBN1803_n_32647) );
in01s06 FE_OCP_RBC1804_n_27825 ( .a(n_27825), .o(FE_OCP_RBN1804_n_27825) );
in01f08 FE_OCP_RBC1805_n_27934 ( .a(n_27934), .o(FE_OCP_RBN1805_n_27934) );
in01s01 FE_OCP_RBC1807_n_13010 ( .a(n_13010), .o(FE_OCP_RBN1807_n_13010) );
in01f02 FE_OCP_RBC1808_n_28968 ( .a(n_28968), .o(FE_OCP_RBN1808_n_28968) );
in01m01 FE_OCP_RBC1809_n_18754 ( .a(n_18754), .o(FE_OCP_RBN1809_n_18754) );
in01f04 FE_OCP_RBC1810_n_18754 ( .a(n_18754), .o(FE_OCP_RBN1810_n_18754) );
in01m02 FE_OCP_RBC1811_n_33750 ( .a(n_33750), .o(FE_OCP_RBN1811_n_33750) );
in01s01 FE_OCP_RBC1812_n_33750 ( .a(n_33750), .o(FE_OCP_RBN1812_n_33750) );
in01s01 FE_OCP_RBC1813_n_33846 ( .a(n_33846), .o(FE_OCP_RBN1813_n_33846) );
in01s02 FE_OCP_RBC1814_n_33846 ( .a(n_33846), .o(FE_OCP_RBN1814_n_33846) );
in01s04 FE_OCP_RBC1815_n_33873 ( .a(n_33873), .o(FE_OCP_RBN1815_n_33873) );
in01s01 FE_OCP_RBC1816_n_33873 ( .a(n_33873), .o(FE_OCP_RBN1816_n_33873) );
in01m06 FE_OCP_RBC1817_n_19178 ( .a(n_19178), .o(FE_OCP_RBN1817_n_19178) );
in01s01 FE_OCP_RBC1818_n_13858 ( .a(n_13858), .o(FE_OCP_RBN1818_n_13858) );
in01s01 FE_OCP_RBC1819_n_13858 ( .a(n_13858), .o(FE_OCP_RBN1819_n_13858) );
in01s01 FE_OCP_RBC1820_n_13858 ( .a(FE_OCP_RBN1818_n_13858), .o(FE_OCP_RBN1820_n_13858) );
in01s01 FE_OCP_RBC1821_n_13858 ( .a(FE_OCP_RBN1818_n_13858), .o(FE_OCP_RBN1821_n_13858) );
in01f04 FE_OCP_RBC1822_n_24473 ( .a(n_24473), .o(FE_OCP_RBN1822_n_24473) );
in01s01 FE_OCP_RBC1823_n_19434 ( .a(n_19434), .o(FE_OCP_RBN1823_n_19434) );
in01m02 FE_OCP_RBC1824_n_19434 ( .a(n_19434), .o(FE_OCP_RBN1824_n_19434) );
in01s01 FE_OCP_RBC1825_n_19513 ( .a(n_19513), .o(FE_OCP_RBN1825_n_19513) );
in01m02 FE_OCP_RBC1826_n_19513 ( .a(n_19513), .o(FE_OCP_RBN1826_n_19513) );
in01m02 FE_OCP_RBC1827_n_19538 ( .a(n_19538), .o(FE_OCP_RBN1827_n_19538) );
in01f06 FE_OCP_RBC1829_n_19528 ( .a(n_19528), .o(FE_OCP_RBN1829_n_19528) );
in01s01 FE_OCP_RBC1831_n_19663 ( .a(FE_OCP_RBN5705_n_19663), .o(FE_OCP_RBN1831_n_19663) );
in01f01 FE_OCP_RBC1832_n_14197 ( .a(n_14197), .o(FE_OCP_RBN1832_n_14197) );
in01s02 FE_OCP_RBC1833_n_14197 ( .a(n_14197), .o(FE_OCP_RBN1833_n_14197) );
in01f01 FE_OCP_RBC1834_n_14664 ( .a(n_14664), .o(FE_OCP_RBN1834_n_14664) );
in01f02 FE_OCP_RBC1836_n_20209 ( .a(n_20209), .o(FE_OCP_RBN1836_n_20209) );
in01f02 FE_OCP_RBC1837_n_20215 ( .a(n_20215), .o(FE_OCP_RBN1837_n_20215) );
in01s01 FE_OCP_RBC1838_n_20273 ( .a(n_20273), .o(FE_OCP_RBN1838_n_20273) );
in01s02 FE_OCP_RBC1839_n_20273 ( .a(n_20273), .o(FE_OCP_RBN1839_n_20273) );
in01f02 FE_OCP_RBC1840_n_20439 ( .a(n_20439), .o(FE_OCP_RBN1840_n_20439) );
in01m02 FE_OCP_RBC1841_FE_RN_442_0 ( .a(FE_RN_442_0), .o(FE_OCP_RBN1841_FE_RN_442_0) );
in01s01 FE_OCP_RBC1842_FE_RN_442_0 ( .a(FE_RN_442_0), .o(FE_OCP_RBN1842_FE_RN_442_0) );
in01f02 FE_OCP_RBC1843_n_20640 ( .a(n_20640), .o(FE_OCP_RBN1843_n_20640) );
in01m02 FE_OCP_RBC1844_n_20616 ( .a(n_20616), .o(FE_OCP_RBN1844_n_20616) );
in01s01 FE_OCP_RBC1845_n_30492 ( .a(n_30492), .o(FE_OCP_RBN1845_n_30492) );
in01m02 FE_OCP_RBC1846_n_30492 ( .a(n_30492), .o(FE_OCP_RBN1846_n_30492) );
in01m04 FE_OCP_RBC1847_n_30428 ( .a(n_30428), .o(FE_OCP_RBN1847_n_30428) );
in01m02 FE_OCP_RBC1848_FE_RN_578_0 ( .a(FE_RN_578_0), .o(FE_OCP_RBN1848_FE_RN_578_0) );
in01f02 FE_OCP_RBC1849_FE_RN_578_0 ( .a(FE_RN_578_0), .o(FE_OCP_RBN1849_FE_RN_578_0) );
in01f01 FE_OCP_RBC1850_n_25898 ( .a(n_25898), .o(FE_OCP_RBN1850_n_25898) );
in01f02 FE_OCP_RBC1851_n_25898 ( .a(n_25898), .o(FE_OCP_RBN1851_n_25898) );
in01f02 FE_OCP_RBC1855_n_20879 ( .a(n_20879), .o(FE_OCP_RBN1855_n_20879) );
in01m04 FE_OCP_RBC1856_n_30731 ( .a(n_30731), .o(FE_OCP_RBN1856_n_30731) );
in01s01 FE_OCP_RBC1857_n_30731 ( .a(FE_OCP_RBN1856_n_30731), .o(FE_OCP_RBN1857_n_30731) );
in01s01 FE_OCP_RBC1859_n_30731 ( .a(FE_OCP_RBN1857_n_30731), .o(FE_OCP_RBN1859_n_30731) );
in01f02 FE_OCP_RBC1862_n_26049 ( .a(n_26049), .o(FE_OCP_RBN1862_n_26049) );
in01m02 FE_OCP_RBC1864_n_21163 ( .a(n_21163), .o(FE_OCP_RBN1864_n_21163) );
in01s01 FE_OCP_RBC1865_n_21163 ( .a(n_21163), .o(FE_OCP_RBN1865_n_21163) );
in01s01 FE_OCP_RBC1866_n_26407 ( .a(n_26407), .o(FE_OCP_RBN1866_n_26407) );
in01s02 FE_OCP_RBC1867_n_26407 ( .a(n_26407), .o(FE_OCP_RBN1867_n_26407) );
in01m04 FE_OCP_RBC1868_n_21358 ( .a(n_21358), .o(FE_OCP_RBN1868_n_21358) );
in01s01 FE_OCP_RBC1869_n_21358 ( .a(n_21358), .o(FE_OCP_RBN1869_n_21358) );
in01s02 FE_OCP_RBC1871_n_36489 ( .a(n_36489), .o(FE_OCP_RBN1871_n_36489) );
in01s01 FE_OCP_RBC1872_n_36489 ( .a(n_36489), .o(FE_OCP_RBN1872_n_36489) );
in01m01 FE_OCP_RBC1875_n_17689 ( .a(n_17689), .o(FE_OCP_RBN1875_n_17689) );
in01m02 FE_OCP_RBC1876_n_27723 ( .a(n_27723), .o(FE_OCP_RBN1876_n_27723) );
in01m02 FE_OCP_RBC1877_n_32382 ( .a(n_32382), .o(FE_OCP_RBN1877_n_32382) );
in01s01 FE_OCP_RBC1878_n_27804 ( .a(n_27804), .o(FE_OCP_RBN1878_n_27804) );
in01s03 FE_OCP_RBC2028_n_44722 ( .a(FE_OCP_RBN7128_n_44722), .o(FE_OCP_RBN2028_n_44722) );
in01s40 FE_OCP_RBC2029_n_44722 ( .a(FE_OCP_RBN7128_n_44722), .o(FE_OCP_RBN2029_n_44722) );
in01s06 FE_OCP_RBC2030_n_44722 ( .a(FE_OCP_RBN7128_n_44722), .o(FE_OCP_RBN2030_n_44722) );
in01s06 FE_OCP_RBC2034_n_44722 ( .a(FE_OCP_RBN2029_n_44722), .o(FE_OCP_RBN2034_n_44722) );
in01s06 FE_OCP_RBC2037_n_44722 ( .a(FE_OCP_RBN2034_n_44722), .o(FE_OCP_RBN2037_n_44722) );
in01s06 FE_OCP_RBC2038_n_44722 ( .a(FE_OCP_RBN2034_n_44722), .o(FE_OCP_RBN2038_n_44722) );
in01s40 FE_OCP_RBC2039_n_44722 ( .a(FE_OCP_RBN2417_n_44722), .o(FE_OCP_RBN2039_n_44722) );
in01s01 FE_OCP_RBC2040_n_28268 ( .a(n_28268), .o(FE_OCP_RBN2040_n_28268) );
in01s01 FE_OCP_RBC2041_n_18269 ( .a(n_18269), .o(FE_OCP_RBN2041_n_18269) );
in01s02 FE_OCP_RBC2042_n_18269 ( .a(FE_OCP_RBN2041_n_18269), .o(FE_OCP_RBN2042_n_18269) );
in01s02 FE_OCP_RBC2043_n_18269 ( .a(FE_OCP_RBN2042_n_18269), .o(FE_OCP_RBN2043_n_18269) );
in01s01 FE_OCP_RBC2044_n_12907 ( .a(n_12907), .o(FE_OCP_RBN2044_n_12907) );
in01s01 FE_OCP_RBC2045_n_12907 ( .a(n_12907), .o(FE_OCP_RBN2045_n_12907) );
in01s04 FE_OCP_RBC2046_n_12907 ( .a(n_12907), .o(FE_OCP_RBN2046_n_12907) );
in01s01 FE_OCP_RBC2049_n_29056 ( .a(FE_OCP_DRV_N6263_FE_OCP_RBN5603_n_29056), .o(FE_OCP_RBN2049_n_29056) );
in01f02 FE_OCP_RBC2050_n_13694 ( .a(n_13694), .o(FE_OCP_RBN2050_n_13694) );
in01s01 FE_OCP_RBC2055_n_13784 ( .a(n_13784), .o(FE_OCP_RBN2055_n_13784) );
in01s02 FE_OCP_RBC2056_n_13784 ( .a(FE_OCP_RBN2055_n_13784), .o(FE_OCP_RBN2056_n_13784) );
in01s01 FE_OCP_RBC2057_n_13784 ( .a(FE_OCP_RBN2056_n_13784), .o(FE_OCP_RBN2057_n_13784) );
in01s01 FE_OCP_RBC2058_n_13784 ( .a(FE_OCP_RBN2056_n_13784), .o(FE_OCP_RBN2058_n_13784) );
in01f02 FE_OCP_RBC2059_n_29380 ( .a(n_29380), .o(FE_OCP_RBN2059_n_29380) );
in01s02 FE_OCP_RBC2060_n_29380 ( .a(n_29380), .o(FE_OCP_RBN2060_n_29380) );
in01f02 FE_OCP_RBC2061_n_13813 ( .a(n_13813), .o(FE_OCP_RBN2061_n_13813) );
in01s01 FE_OCP_RBC2062_n_19353 ( .a(n_19353), .o(FE_OCP_RBN2062_n_19353) );
in01m04 FE_OCP_RBC2063_n_19353 ( .a(n_19353), .o(FE_OCP_RBN2063_n_19353) );
in01s01 FE_OCP_RBC2064_n_19353 ( .a(FE_OCP_RBN2062_n_19353), .o(FE_OCP_RBN2064_n_19353) );
in01f02 FE_OCP_RBC2065_n_13913 ( .a(n_13913), .o(FE_OCP_RBN2065_n_13913) );
in01m02 FE_OCP_RBC2066_n_14069 ( .a(n_14069), .o(FE_OCP_RBN2066_n_14069) );
in01s01 FE_OCP_RBC2067_n_14069 ( .a(n_14069), .o(FE_OCP_RBN2067_n_14069) );
in01s02 FE_OCP_RBC2068_n_14069 ( .a(FE_OCP_RBN2067_n_14069), .o(FE_OCP_RBN2068_n_14069) );
in01s01 FE_OCP_RBC2069_n_14069 ( .a(FE_OCP_RBN2068_n_14069), .o(FE_OCP_RBN2069_n_14069) );
in01s02 FE_OCP_RBC2070_n_14069 ( .a(FE_OCP_RBN2068_n_14069), .o(FE_OCP_RBN2070_n_14069) );
in01f01 FE_OCP_RBC2071_n_14120 ( .a(n_14120), .o(FE_OCP_RBN2071_n_14120) );
in01s01 FE_OCP_RBC2073_n_14120 ( .a(FE_OCP_RBN5727_n_14120), .o(FE_OCP_RBN2073_n_14120) );
in01f04 FE_OCP_RBC2074_n_29603 ( .a(n_29603), .o(FE_OCP_RBN2074_n_29603) );
in01m04 FE_OCP_RBC2075_n_14093 ( .a(n_14093), .o(FE_OCP_RBN2075_n_14093) );
in01m02 FE_OCP_RBC2076_n_14149 ( .a(n_14149), .o(FE_OCP_RBN2076_n_14149) );
in01s01 FE_OCP_RBC2077_n_14149 ( .a(n_14149), .o(FE_OCP_RBN2077_n_14149) );
in01s02 FE_OCP_RBC2078_n_14149 ( .a(FE_OCP_RBN2077_n_14149), .o(FE_OCP_RBN2078_n_14149) );
in01s01 FE_OCP_RBC2079_n_14149 ( .a(FE_OCP_RBN2078_n_14149), .o(FE_OCP_RBN2079_n_14149) );
in01s01 FE_OCP_RBC2080_n_14554 ( .a(n_14554), .o(FE_OCP_RBN2080_n_14554) );
in01s01 FE_OCP_RBC2081_n_14554 ( .a(FE_OCP_RBN2080_n_14554), .o(FE_OCP_RBN2081_n_14554) );
in01s01 FE_OCP_RBC2082_n_14554 ( .a(FE_OCP_RBN2081_n_14554), .o(FE_OCP_RBN2082_n_14554) );
in01f01 FE_OCP_RBC2083_n_14611 ( .a(n_14611), .o(FE_OCP_RBN2083_n_14611) );
in01s02 FE_OCP_RBC2084_n_19970 ( .a(n_19970), .o(FE_OCP_RBN2084_n_19970) );
in01f03 FE_OCP_RBC2085_n_14911 ( .a(n_14911), .o(FE_OCP_RBN2085_n_14911) );
in01s01 FE_OCP_RBC2086_n_14911 ( .a(n_14911), .o(FE_OCP_RBN2086_n_14911) );
in01s01 FE_OCP_RBC2087_n_14911 ( .a(FE_OCP_RBN2085_n_14911), .o(FE_OCP_RBN2087_n_14911) );
in01f02 FE_OCP_RBC2089_n_14964 ( .a(n_14964), .o(FE_OCP_RBN2089_n_14964) );
in01f01 FE_OCP_RBC2090_n_14908 ( .a(n_14908), .o(FE_OCP_RBN2090_n_14908) );
in01f01 FE_OCP_RBC2091_n_14909 ( .a(n_14909), .o(FE_OCP_RBN2091_n_14909) );
in01s01 FE_OCP_RBC2092_n_14991 ( .a(n_14991), .o(FE_OCP_RBN2092_n_14991) );
in01m02 FE_OCP_RBC2093_n_14991 ( .a(n_14991), .o(FE_OCP_RBN2093_n_14991) );
in01s01 FE_OCP_RBC2094_n_47175 ( .a(n_47175), .o(FE_OCP_RBN2094_n_47175) );
in01m02 FE_OCP_RBC2095_n_20325 ( .a(n_20325), .o(FE_OCP_RBN2095_n_20325) );
in01s01 FE_OCP_RBC2096_n_20325 ( .a(n_20325), .o(FE_OCP_RBN2096_n_20325) );
in01s01 FE_OCP_RBC2097_n_20325 ( .a(FE_OCP_RBN2096_n_20325), .o(FE_OCP_RBN2097_n_20325) );
in01s01 FE_OCP_RBC2098_n_20325 ( .a(FE_OCP_RBN2097_n_20325), .o(FE_OCP_RBN2098_n_20325) );
in01s02 FE_OCP_RBC2101_n_15083 ( .a(n_15083), .o(FE_OCP_RBN2101_n_15083) );
in01s01 FE_OCP_RBC2102_n_15083 ( .a(n_15083), .o(FE_OCP_RBN2102_n_15083) );
in01s02 FE_OCP_RBC2103_n_15286 ( .a(n_15286), .o(FE_OCP_RBN2103_n_15286) );
in01f02 FE_OCP_RBC2104_n_30465 ( .a(n_30465), .o(FE_OCP_RBN2104_n_30465) );
in01s01 FE_OCP_RBC2105_n_30465 ( .a(n_30465), .o(FE_OCP_RBN2105_n_30465) );
in01s01 FE_OCP_RBC2106_n_30619 ( .a(n_30619), .o(FE_OCP_RBN2106_n_30619) );
in01f02 FE_OCP_RBC2107_n_30747 ( .a(n_30747), .o(FE_OCP_RBN2107_n_30747) );
in01f04 FE_OCP_RBC2108_n_15911 ( .a(n_15911), .o(FE_OCP_RBN2108_n_15911) );
in01s01 FE_OCP_RBC2109_n_15911 ( .a(n_15911), .o(FE_OCP_RBN2109_n_15911) );
in01s01 FE_OCP_RBC2110_n_15911 ( .a(FE_OCP_RBN2109_n_15911), .o(FE_OCP_RBN2110_n_15911) );
in01s01 FE_OCP_RBC2111_n_15911 ( .a(FE_OCP_RBN2110_n_15911), .o(FE_OCP_RBN2111_n_15911) );
in01s02 FE_OCP_RBC2112_n_20935 ( .a(n_20935), .o(FE_OCP_RBN2112_n_20935) );
in01s01 FE_OCP_RBC2113_n_20935 ( .a(FE_OCP_RBN2112_n_20935), .o(FE_OCP_RBN2113_n_20935) );
in01s01 FE_OCP_RBC2114_n_20935 ( .a(FE_OCP_RBN2113_n_20935), .o(FE_OCP_RBN2114_n_20935) );
in01s01 FE_OCP_RBC2115_n_20935 ( .a(FE_OCP_RBN2113_n_20935), .o(FE_OCP_RBN2115_n_20935) );
in01s01 FE_OCP_RBC2118_n_22351 ( .a(n_22351), .o(FE_OCP_RBN2118_n_22351) );
in01s40 FE_OCP_RBC2250_n_44061 ( .a(FE_OCP_RBN5179_n_44061), .o(FE_OCP_RBN2250_n_44061) );
in01s01 FE_OCP_RBC2258_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2258_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s01 FE_OCP_RBC2259_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2259_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s01 FE_OCP_RBC2260_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2260_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s01 FE_OCP_RBC2261_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(FE_OCP_RBN5465_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2261_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s01 FE_OCP_RBC2262_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(FE_OCP_RBN2261_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2262_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s01 FE_OCP_RBC2263_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(FE_OCP_RBN2261_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2263_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s01 FE_OCP_RBC2264_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(FE_OCP_RBN2261_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2264_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s01 FE_OCP_RBC2265_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(FE_OCP_RBN2261_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2265_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s01 FE_OCP_RBC2266_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(FE_OCP_RBN2261_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2266_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s01 FE_OCP_RBC2267_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(FE_OCP_RBN2261_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2267_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s01 FE_OCP_RBC2268_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(FE_OCP_RBN2261_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2268_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01m10 FE_OCP_RBC2270_delay_xor_ln22_unr15_stage6_stallmux_q_2_ ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_2_), .o(FE_OCP_RBN2270_delay_xor_ln22_unr15_stage6_stallmux_q_2_) );
in01s40 FE_OCP_RBC2271_delay_xor_ln22_unr15_stage6_stallmux_q_5_ ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_5_), .o(FE_OCP_RBN2271_delay_xor_ln22_unr15_stage6_stallmux_q_5_) );
in01s10 FE_OCP_RBC2272_delay_xor_ln22_unr15_stage6_stallmux_q_5_ ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_5_), .o(FE_OCP_RBN2272_delay_xor_ln22_unr15_stage6_stallmux_q_5_) );
in01m03 FE_OCP_RBC2282_delay_sub_ln23_unr21_stage7_stallmux_q_1_ ( .a(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(FE_OCP_RBN2282_delay_sub_ln23_unr21_stage7_stallmux_q_1_) );
in01s10 FE_OCP_RBC2311_delay_sub_ln23_unr25_stage8_stallmux_q_1_ ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .o(FE_OCP_RBN2311_delay_sub_ln23_unr25_stage8_stallmux_q_1_) );
in01s10 FE_OCP_RBC2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_ ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_) );
in01s01 FE_OCP_RBC2337_delay_sub_ln21_0_unr23_stage9_stallmux_q_20_ ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_20_), .o(FE_OCP_RBN2337_delay_sub_ln21_0_unr23_stage9_stallmux_q_20_) );
in01s01 FE_OCP_RBC2338_delay_sub_ln21_0_unr23_stage9_stallmux_q_20_ ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_20_), .o(FE_OCP_RBN2338_delay_sub_ln21_0_unr23_stage9_stallmux_q_20_) );
in01s06 FE_OCP_RBC2369_n_44061 ( .a(FE_OCP_RBN3871_n_44061), .o(FE_OCP_RBN2369_n_44061) );
in01s01 FE_OCP_RBC2377_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN5412_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN2377_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s01 FE_OCP_RBC2378_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN5412_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN2378_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s01 FE_OCP_RBC2382_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN6509_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN2382_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01m06 FE_OCP_RBC2385_n_22820 ( .a(n_22820), .o(FE_OCP_RBN2385_n_22820) );
in01s02 FE_OCP_RBC2386_n_22650 ( .a(n_22650), .o(FE_OCP_RBN2386_n_22650) );
in01m20 FE_OCP_RBC2387_n_23227 ( .a(n_23227), .o(FE_OCP_RBN2387_n_23227) );
in01m20 FE_OCP_RBC2388_n_23227 ( .a(FE_OCP_RBN2387_n_23227), .o(FE_OCP_RBN2388_n_23227) );
in01s01 FE_OCP_RBC2389_n_23227 ( .a(FE_OCP_RBN2387_n_23227), .o(FE_OCP_RBN2389_n_23227) );
in01m08 FE_OCP_RBC2390_FE_RN_1364_0 ( .a(FE_RN_1364_0), .o(FE_OCP_RBN2390_FE_RN_1364_0) );
in01s06 FE_OCP_RBC2392_n_16970 ( .a(n_16970), .o(FE_OCP_RBN2392_n_16970) );
in01m03 FE_OCP_RBC2393_n_45697 ( .a(n_45697), .o(FE_OCP_RBN2393_n_45697) );
in01s10 FE_OCP_RBC2394_n_45697 ( .a(FE_OCP_RBN2393_n_45697), .o(FE_OCP_RBN2394_n_45697) );
in01s01 FE_OCP_RBC2395_n_45697 ( .a(FE_OCP_RBN2393_n_45697), .o(FE_OCP_RBN2395_n_45697) );
in01s01 FE_OCP_RBC2396_n_45697 ( .a(FE_OCP_RBN2394_n_45697), .o(FE_OCP_RBN2396_n_45697) );
in01s01 FE_OCP_RBC2397_n_45697 ( .a(FE_OCP_RBN2394_n_45697), .o(FE_OCP_RBN2397_n_45697) );
in01s01 FE_OCP_RBC2398_n_45697 ( .a(FE_OCP_RBN2395_n_45697), .o(FE_OCP_RBN2398_n_45697) );
in01s06 FE_OCP_RBC2399_n_45697 ( .a(FE_OCP_RBN2396_n_45697), .o(FE_OCP_RBN2399_n_45697) );
in01s01 FE_OCP_RBC2400_n_45697 ( .a(FE_OCP_RBN2397_n_45697), .o(FE_OCP_RBN2400_n_45697) );
in01s01 FE_OCP_RBC2401_n_45697 ( .a(FE_OCP_RBN2399_n_45697), .o(FE_OCP_RBN2401_n_45697) );
in01s02 FE_OCP_RBC2402_n_45697 ( .a(FE_OCP_RBN2400_n_45697), .o(FE_OCP_RBN2402_n_45697) );
in01s02 FE_OCP_RBC2404_n_45697 ( .a(FE_OCP_RBN2401_n_45697), .o(FE_OCP_RBN2404_n_45697) );
in01s01 FE_OCP_RBC2405_n_45697 ( .a(FE_OCP_RBN2402_n_45697), .o(FE_OCP_RBN2405_n_45697) );
in01s01 FE_OCP_RBC2406_n_45697 ( .a(FE_OCP_RBN2405_n_45697), .o(FE_OCP_RBN2406_n_45697) );
in01s02 FE_OCP_RBC2407_n_6635 ( .a(n_6635), .o(FE_OCP_RBN2407_n_6635) );
in01m06 FE_OCP_RBC2410_n_40631 ( .a(n_40631), .o(FE_OCP_RBN2410_n_40631) );
in01s06 FE_OCP_RBC2411_n_44722 ( .a(FE_OCP_RBN2029_n_44722), .o(FE_OCP_RBN2411_n_44722) );
in01s06 FE_OCP_RBC2412_n_44722 ( .a(FE_OCP_RBN2029_n_44722), .o(FE_OCP_RBN2412_n_44722) );
in01s40 FE_OCP_RBC2413_n_44722 ( .a(FE_OCP_RBN2029_n_44722), .o(FE_OCP_RBN2413_n_44722) );
in01s20 FE_OCP_RBC2414_n_44722 ( .a(FE_OCP_RBN2411_n_44722), .o(FE_OCP_RBN2414_n_44722) );
in01s10 FE_OCP_RBC2415_n_44722 ( .a(FE_OCP_RBN2412_n_44722), .o(FE_OCP_RBN2415_n_44722) );
in01s80 FE_OCP_RBC2416_n_44722 ( .a(FE_OCP_RBN2413_n_44722), .o(FE_OCP_RBN2416_n_44722) );
in01s06 FE_OCP_RBC2417_n_44722 ( .a(FE_OCP_RBN2413_n_44722), .o(FE_OCP_RBN2417_n_44722) );
in01s06 FE_OCP_RBC2418_n_44083 ( .a(n_44083), .o(FE_OCP_RBN2418_n_44083) );
in01s40 FE_OCP_RBC2422_n_23023 ( .a(n_23023), .o(FE_OCP_RBN2422_n_23023) );
in01s01 FE_OCP_RBC2423_n_32554 ( .a(n_32554), .o(FE_OCP_RBN2423_n_32554) );
in01s02 FE_OCP_RBC2426_n_11907 ( .a(n_11907), .o(FE_OCP_RBN2426_n_11907) );
in01s06 FE_OCP_RBC2427_n_11907 ( .a(n_11907), .o(FE_OCP_RBN2427_n_11907) );
in01m06 FE_OCP_RBC2428_n_37207 ( .a(n_37207), .o(FE_OCP_RBN2428_n_37207) );
in01m02 FE_OCP_RBC2429_FE_RN_107_0 ( .a(FE_RN_107_0), .o(FE_OCP_RBN2429_FE_RN_107_0) );
in01s08 FE_OCP_RBC2430_FE_RN_107_0 ( .a(FE_RN_107_0), .o(FE_OCP_RBN2430_FE_RN_107_0) );
in01m06 FE_OCP_RBC2431_FE_RN_107_0 ( .a(FE_RN_107_0), .o(FE_OCP_RBN2431_FE_RN_107_0) );
in01f10 FE_OCP_RBC2432_FE_RN_107_0 ( .a(FE_RN_107_0), .o(FE_OCP_RBN2432_FE_RN_107_0) );
in01f20 FE_OCP_RBC2433_FE_RN_107_0 ( .a(FE_OCP_RBN2432_FE_RN_107_0), .o(FE_OCP_RBN2433_FE_RN_107_0) );
in01m04 FE_OCP_RBC2434_n_32702 ( .a(n_32702), .o(FE_OCP_RBN2434_n_32702) );
in01s80 FE_OCP_RBC2435_FE_OCPN833_n_45450 ( .a(FE_OCPN833_n_45450), .o(FE_OCP_RBN2435_FE_OCPN833_n_45450) );
in01s80 FE_OCP_RBC2436_FE_OCPN833_n_45450 ( .a(FE_OCP_RBN2435_FE_OCPN833_n_45450), .o(FE_OCP_RBN2436_FE_OCPN833_n_45450) );
in01s01 FE_OCP_RBC2437_FE_OCPN833_n_45450 ( .a(FE_OCP_RBN2436_FE_OCPN833_n_45450), .o(FE_OCP_RBN2437_FE_OCPN833_n_45450) );
in01m03 FE_OCP_RBC2438_FE_OCPN833_n_45450 ( .a(FE_OCP_RBN2436_FE_OCPN833_n_45450), .o(FE_OCP_RBN2438_FE_OCPN833_n_45450) );
in01s01 FE_OCP_RBC2439_n_6937 ( .a(n_6937), .o(FE_OCP_RBN2439_n_6937) );
in01f20 FE_OCP_RBC2440_n_44798 ( .a(n_44798), .o(FE_OCP_RBN2440_n_44798) );
in01s04 FE_OCP_RBC2441_n_44798 ( .a(n_44798), .o(FE_OCP_RBN2441_n_44798) );
in01s06 FE_OCP_RBC2442_n_44798 ( .a(FE_OCP_RBN2440_n_44798), .o(FE_OCP_RBN2442_n_44798) );
in01f20 FE_OCP_RBC2443_n_44798 ( .a(FE_OCP_RBN2440_n_44798), .o(FE_OCP_RBN2443_n_44798) );
in01m02 FE_OCP_RBC2444_n_1675 ( .a(n_1675), .o(FE_OCP_RBN2444_n_1675) );
in01s01 FE_OCP_RBC2445_n_1675 ( .a(n_1675), .o(FE_OCP_RBN2445_n_1675) );
in01s10 FE_OCP_RBC2446_n_23079 ( .a(n_23079), .o(FE_OCP_RBN2446_n_23079) );
in01s06 FE_OCP_RBC2447_n_12312 ( .a(n_12312), .o(FE_OCP_RBN2447_n_12312) );
in01s01 FE_OCP_RBC2448_n_23246 ( .a(n_23246), .o(FE_OCP_RBN2448_n_23246) );
in01m08 FE_OCP_RBC2449_n_23246 ( .a(n_23246), .o(FE_OCP_RBN2449_n_23246) );
in01f02 FE_OCP_RBC2450_n_23246 ( .a(n_23246), .o(FE_OCP_RBN2450_n_23246) );
in01s08 FE_OCP_RBC2451_n_32860 ( .a(n_32860), .o(FE_OCP_RBN2451_n_32860) );
in01m08 FE_OCP_RBC2452_n_32860 ( .a(n_32860), .o(FE_OCP_RBN2452_n_32860) );
in01s02 FE_OCP_RBC2453_n_32860 ( .a(n_32860), .o(FE_OCP_RBN2453_n_32860) );
in01s01 FE_OCP_RBC2454_n_32860 ( .a(FE_OCP_RBN2451_n_32860), .o(FE_OCP_RBN2454_n_32860) );
in01s01 FE_OCP_RBC2460_n_12365 ( .a(n_12365), .o(FE_OCP_RBN2460_n_12365) );
in01s06 FE_OCP_RBC2461_n_12365 ( .a(n_12365), .o(FE_OCP_RBN2461_n_12365) );
in01m08 FE_OCP_RBC2462_n_23345 ( .a(n_23345), .o(FE_OCP_RBN2462_n_23345) );
in01f03 FE_OCP_RBC2463_n_37449 ( .a(n_37449), .o(FE_OCP_RBN2463_n_37449) );
in01s01 FE_OCP_RBC2464_n_7129 ( .a(n_7129), .o(FE_OCP_RBN2464_n_7129) );
in01s08 FE_OCP_RBC2467_n_33034 ( .a(FE_OCP_RBN4005_n_33015), .o(FE_OCP_RBN2467_n_33034) );
in01m04 FE_OCP_RBC2468_n_33034 ( .a(FE_OCP_RBN4005_n_33015), .o(FE_OCP_RBN2468_n_33034) );
in01s08 FE_OCP_RBC2469_n_33034 ( .a(FE_OCP_RBN4005_n_33015), .o(FE_OCP_RBN2469_n_33034) );
in01s01 FE_OCP_RBC2476_n_33034 ( .a(FE_OCP_RBN4018_n_33034), .o(FE_OCP_RBN2476_n_33034) );
in01s01 FE_OCP_RBC2477_n_33034 ( .a(FE_OCP_RBN2476_n_33034), .o(FE_OCP_RBN2477_n_33034) );
in01s01 FE_OCP_RBC2478_n_1862 ( .a(n_1862), .o(FE_OCP_RBN2478_n_1862) );
in01m06 FE_OCP_RBC2479_n_47245 ( .a(n_47245), .o(FE_OCP_RBN2479_n_47245) );
in01m04 FE_OCP_RBC2480_FE_RN_734_0 ( .a(FE_RN_734_0), .o(FE_OCP_RBN2480_FE_RN_734_0) );
in01s01 FE_OCP_RBC2481_FE_RN_734_0 ( .a(FE_RN_734_0), .o(FE_OCP_RBN2481_FE_RN_734_0) );
in01f04 FE_OCP_RBC2482_n_37509 ( .a(n_37509), .o(FE_OCP_RBN2482_n_37509) );
in01s06 FE_OCP_RBC2483_FE_RN_657_0 ( .a(FE_RN_657_0), .o(FE_OCP_RBN2483_FE_RN_657_0) );
in01s02 FE_OCP_RBC2484_FE_RN_657_0 ( .a(FE_RN_657_0), .o(FE_OCP_RBN2484_FE_RN_657_0) );
in01f03 FE_OCP_RBC2485_n_41213 ( .a(n_41213), .o(FE_OCP_RBN2485_n_41213) );
in01m06 FE_OCP_RBC2490_FE_RN_1367_0 ( .a(FE_OCP_RBN6554_n_28458), .o(FE_OCP_RBN2490_FE_RN_1367_0) );
in01s01 FE_OCP_RBC2491_FE_RN_1367_0 ( .a(FE_OCP_RBN6554_n_28458), .o(FE_OCP_RBN2491_FE_RN_1367_0) );
in01s02 FE_OCP_RBC2492_FE_RN_1367_0 ( .a(FE_OCP_RBN6554_n_28458), .o(FE_OCP_RBN2492_FE_RN_1367_0) );
in01s01 FE_OCP_RBC2494_n_7349 ( .a(n_7349), .o(FE_OCP_RBN2494_n_7349) );
in01m08 FE_OCP_RBC2495_n_18242 ( .a(n_18242), .o(FE_OCP_RBN2495_n_18242) );
in01m08 FE_OCP_RBC2496_n_18242 ( .a(FE_OCP_RBN2495_n_18242), .o(FE_OCP_RBN2496_n_18242) );
in01s06 FE_OCP_RBC2497_n_18242 ( .a(FE_OCP_RBN2496_n_18242), .o(FE_OCP_RBN2497_n_18242) );
in01f02 FE_OCP_RBC2498_n_37624 ( .a(n_37624), .o(FE_OCP_RBN2498_n_37624) );
in01s01 FE_OCP_RBC2499_FE_RN_1553_0 ( .a(FE_RN_1553_0), .o(FE_OCP_RBN2499_FE_RN_1553_0) );
in01s01 FE_OCP_RBC2500_n_28773 ( .a(n_28773), .o(FE_OCP_RBN2500_n_28773) );
in01s01 FE_OCP_RBC2502_n_33226 ( .a(FE_OCP_RBN6561_n_33208), .o(FE_OCP_RBN2502_n_33226) );
in01s01 FE_OCP_RBC2503_n_33226 ( .a(FE_OCP_RBN6561_n_33208), .o(FE_OCP_RBN2503_n_33226) );
in01s06 FE_OCP_RBC2505_n_33226 ( .a(FE_OCP_RBN6562_n_33208), .o(FE_OCP_RBN2505_n_33226) );
in01s01 FE_OCP_RBC2506_n_33226 ( .a(FE_OCP_RBN2505_n_33226), .o(FE_OCP_RBN2506_n_33226) );
in01s01 FE_OCP_RBC2507_n_37720 ( .a(n_37720), .o(FE_OCP_RBN2507_n_37720) );
in01m06 FE_OCP_RBC2508_n_37720 ( .a(n_37720), .o(FE_OCP_RBN2508_n_37720) );
in01m08 FE_OCP_RBC2509_n_41215 ( .a(n_41215), .o(FE_OCP_RBN2509_n_41215) );
in01s01 FE_OCP_RBC2510_n_12800 ( .a(n_12800), .o(FE_OCP_RBN2510_n_12800) );
in01s01 FE_OCP_RBC2511_n_12800 ( .a(FE_OCP_RBN2510_n_12800), .o(FE_OCP_RBN2511_n_12800) );
in01s01 FE_OCP_RBC2512_n_12800 ( .a(FE_OCP_RBN2511_n_12800), .o(FE_OCP_RBN2512_n_12800) );
in01s01 FE_OCP_RBC2513_n_28699 ( .a(n_28699), .o(FE_OCP_RBN2513_n_28699) );
in01s01 FE_OCP_RBC2514_n_28699 ( .a(n_28699), .o(FE_OCP_RBN2514_n_28699) );
in01f01 FE_OCP_RBC2515_n_45120 ( .a(n_45120), .o(FE_OCP_RBN2515_n_45120) );
in01m06 FE_OCP_RBC2517_n_45120 ( .a(n_45120), .o(FE_OCP_RBN2517_n_45120) );
in01s01 FE_OCP_RBC2519_n_12721 ( .a(FE_OCP_RBN4047_n_12721), .o(FE_OCP_RBN2519_n_12721) );
in01s01 FE_OCP_RBC2521_n_12721 ( .a(FE_OCP_RBN4047_n_12721), .o(FE_OCP_RBN2521_n_12721) );
in01s02 FE_OCP_RBC2522_n_12721 ( .a(FE_OCP_RBN2521_n_12721), .o(FE_OCP_RBN2522_n_12721) );
in01s01 FE_OCP_RBC2523_n_29017 ( .a(n_29017), .o(FE_OCP_RBN2523_n_29017) );
in01m06 FE_OCP_RBC2524_n_28749 ( .a(n_28749), .o(FE_OCP_RBN2524_n_28749) );
in01s02 FE_OCP_RBC2526_n_2086 ( .a(n_2086), .o(FE_OCP_RBN2526_n_2086) );
in01s01 FE_OCP_RBC2528_n_2097 ( .a(n_2097), .o(FE_OCP_RBN2528_n_2097) );
in01m01 FE_OCP_RBC2529_n_12731 ( .a(n_12731), .o(FE_OCP_RBN2529_n_12731) );
in01m02 FE_OCP_RBC2530_n_13151 ( .a(n_13151), .o(FE_OCP_RBN2530_n_13151) );
in01s01 FE_OCP_RBC2531_n_33372 ( .a(n_33372), .o(FE_OCP_RBN2531_n_33372) );
in01s06 FE_OCP_RBC2532_n_33372 ( .a(n_33372), .o(FE_OCP_RBN2532_n_33372) );
in01s01 FE_OCP_RBC2533_n_33372 ( .a(n_33372), .o(FE_OCP_RBN2533_n_33372) );
in01s01 FE_OCP_RBC2534_n_33372 ( .a(FE_OCP_RBN2533_n_33372), .o(FE_OCP_RBN2534_n_33372) );
in01m04 FE_OCP_RBC2535_n_33568 ( .a(n_33568), .o(FE_OCP_RBN2535_n_33568) );
in01s04 FE_OCP_RBC2536_n_12880 ( .a(n_12880), .o(FE_OCP_RBN2536_n_12880) );
in01s20 FE_OCP_RBC2537_n_12880 ( .a(n_12880), .o(FE_OCP_RBN2537_n_12880) );
in01s01 FE_OCP_RBC2538_n_12880 ( .a(n_12880), .o(FE_OCP_RBN2538_n_12880) );
in01s10 FE_OCP_RBC2539_n_12880 ( .a(FE_OCP_RBN2536_n_12880), .o(FE_OCP_RBN2539_n_12880) );
in01s20 FE_OCP_RBC2540_n_12880 ( .a(FE_OCP_RBN2537_n_12880), .o(FE_OCP_RBN2540_n_12880) );
in01m02 FE_OCP_RBC2541_n_12880 ( .a(FE_OCP_RBN2537_n_12880), .o(FE_OCP_RBN2541_n_12880) );
in01m06 FE_OCP_RBC2542_n_12921 ( .a(n_12921), .o(FE_OCP_RBN2542_n_12921) );
in01f04 FE_OCP_RBC2543_n_33584 ( .a(n_33584), .o(FE_OCP_RBN2543_n_33584) );
in01s01 FE_OCP_RBC2544_n_33584 ( .a(n_33584), .o(FE_OCP_RBN2544_n_33584) );
in01s06 FE_OCP_RBC2548_n_44881 ( .a(FE_OCP_RBN6574_n_44875), .o(FE_OCP_RBN2548_n_44881) );
in01s10 FE_OCP_RBC2549_n_44881 ( .a(FE_OCP_RBN2548_n_44881), .o(FE_OCP_RBN2549_n_44881) );
in01s02 FE_OCP_RBC2550_n_33664 ( .a(n_33664), .o(FE_OCP_RBN2550_n_33664) );
in01s01 FE_OCP_RBC2551_n_33664 ( .a(n_33664), .o(FE_OCP_RBN2551_n_33664) );
in01s01 FE_OCP_RBC2552_n_33697 ( .a(n_33697), .o(FE_OCP_RBN2552_n_33697) );
in01s01 FE_OCP_RBC2553_n_33697 ( .a(n_33697), .o(FE_OCP_RBN2553_n_33697) );
in01s02 FE_OCP_RBC2554_n_13141 ( .a(n_13141), .o(FE_OCP_RBN2554_n_13141) );
in01m04 FE_OCP_RBC2555_n_13141 ( .a(n_13141), .o(FE_OCP_RBN2555_n_13141) );
in01f02 FE_OCP_RBC2556_n_13141 ( .a(n_13141), .o(FE_OCP_RBN2556_n_13141) );
in01s01 FE_OCP_RBC2557_n_13141 ( .a(n_13141), .o(FE_OCP_RBN2557_n_13141) );
in01m04 FE_OCP_RBC2558_n_7665 ( .a(n_7665), .o(FE_OCP_RBN2558_n_7665) );
in01m08 FE_OCP_RBC2559_n_13084 ( .a(n_13084), .o(FE_OCP_RBN2559_n_13084) );
in01s01 FE_OCP_RBC2560_n_13084 ( .a(FE_OCP_RBN2559_n_13084), .o(FE_OCP_RBN2560_n_13084) );
in01s01 FE_OCP_RBC2561_n_13084 ( .a(FE_OCP_RBN2559_n_13084), .o(FE_OCP_RBN2561_n_13084) );
in01s06 FE_OCP_RBC2562_n_13084 ( .a(FE_OCP_RBN2559_n_13084), .o(FE_OCP_RBN2562_n_13084) );
in01s01 FE_OCP_RBC2563_n_13084 ( .a(FE_OCP_RBN2561_n_13084), .o(FE_OCP_RBN2563_n_13084) );
in01m01 FE_OCP_RBC2564_n_29110 ( .a(n_29110), .o(FE_OCP_RBN2564_n_29110) );
in01f01 FE_OCP_RBC2565_n_29110 ( .a(n_29110), .o(FE_OCP_RBN2565_n_29110) );
in01m02 FE_OCP_RBC2566_n_29163 ( .a(n_29163), .o(FE_OCP_RBN2566_n_29163) );
in01s01 FE_OCP_RBC2567_n_29163 ( .a(n_29163), .o(FE_OCP_RBN2567_n_29163) );
in01m02 FE_OCP_RBC2570_n_33735 ( .a(n_33735), .o(FE_OCP_RBN2570_n_33735) );
in01s01 FE_OCP_RBC2571_n_2430 ( .a(n_2430), .o(FE_OCP_RBN2571_n_2430) );
in01s01 FE_OCP_RBC2573_n_2558 ( .a(n_2558), .o(FE_OCP_RBN2573_n_2558) );
in01s01 FE_OCP_RBC2574_n_2558 ( .a(n_2558), .o(FE_OCP_RBN2574_n_2558) );
in01s02 FE_OCP_RBC2579_n_13154 ( .a(n_13154), .o(FE_OCP_RBN2579_n_13154) );
in01f06 FE_OCP_RBC2580_n_13154 ( .a(n_13154), .o(FE_OCP_RBN2580_n_13154) );
in01s02 FE_OCP_RBC2581_n_37913 ( .a(n_37913), .o(FE_OCP_RBN2581_n_37913) );
in01f02 FE_OCP_RBC2582_n_29091 ( .a(n_29091), .o(FE_OCP_RBN2582_n_29091) );
in01f04 FE_OCP_RBC2583_n_29091 ( .a(FE_OCP_RBN2582_n_29091), .o(FE_OCP_RBN2583_n_29091) );
in01s01 FE_OCP_RBC2584_n_29091 ( .a(FE_OCP_RBN2583_n_29091), .o(FE_OCP_RBN2584_n_29091) );
in01s01 FE_OCP_RBC2587_n_7743 ( .a(FE_OCP_RBN6600_n_7708), .o(FE_OCP_RBN2587_n_7743) );
in01s01 FE_OCP_RBC2588_n_7743 ( .a(FE_OCP_RBN6600_n_7708), .o(FE_OCP_RBN2588_n_7743) );
in01s01 FE_OCP_RBC2592_n_7743 ( .a(FE_OCP_RBN4143_n_7743), .o(FE_OCP_RBN2592_n_7743) );
in01s01 FE_OCP_RBC2593_n_7743 ( .a(FE_OCP_RBN2588_n_7743), .o(FE_OCP_RBN2593_n_7743) );
in01s01 FE_OCP_RBC2595_n_7743 ( .a(FE_OCP_RBN2588_n_7743), .o(FE_OCP_RBN2595_n_7743) );
in01s01 FE_OCP_RBC2597_n_7743 ( .a(FE_OCP_RBN4145_n_7743), .o(FE_OCP_RBN2597_n_7743) );
in01s01 FE_OCP_RBC2598_n_7743 ( .a(FE_OCP_RBN2592_n_7743), .o(FE_OCP_RBN2598_n_7743) );
in01s01 FE_OCP_RBC2599_n_7743 ( .a(FE_OCP_RBN2592_n_7743), .o(FE_OCP_RBN2599_n_7743) );
in01s01 FE_OCP_RBC2601_n_13483 ( .a(FE_OCP_RBN4120_n_13483), .o(FE_OCP_RBN2601_n_13483) );
in01s01 FE_OCP_RBC2602_n_13483 ( .a(FE_OCP_RBN2601_n_13483), .o(FE_OCP_RBN2602_n_13483) );
in01s01 FE_OCP_RBC2604_FE_OCPN855_n_7721 ( .a(FE_OCP_RBN6601_n_7708), .o(FE_OCP_RBN2604_FE_OCPN855_n_7721) );
in01s01 FE_OCP_RBC2605_FE_OCPN855_n_7721 ( .a(FE_OCP_RBN2604_FE_OCPN855_n_7721), .o(FE_OCP_RBN2605_FE_OCPN855_n_7721) );
in01s01 FE_OCP_RBC2607_FE_OCPN855_n_7721 ( .a(FE_OCP_RBN5647_FE_OCPN855_n_7721), .o(FE_OCP_RBN2607_FE_OCPN855_n_7721) );
in01s01 FE_OCP_RBC2608_FE_OCPN855_n_7721 ( .a(FE_OCP_RBN2607_FE_OCPN855_n_7721), .o(FE_OCP_RBN2608_FE_OCPN855_n_7721) );
in01s01 FE_OCP_RBC2609_n_47235 ( .a(n_47235), .o(FE_OCP_RBN2609_n_47235) );
in01f02 FE_OCP_RBC2610_n_29298 ( .a(n_29298), .o(FE_OCP_RBN2610_n_29298) );
in01s01 FE_OCP_RBC2611_n_29298 ( .a(n_29298), .o(FE_OCP_RBN2611_n_29298) );
in01s06 FE_OCP_RBC2612_FE_OCPN857_n_7802 ( .a(FE_OCP_RBN5612_n_7730), .o(FE_OCP_RBN2612_FE_OCPN857_n_7802) );
in01s02 FE_OCP_RBC2613_FE_OCPN857_n_7802 ( .a(FE_OCP_RBN2612_FE_OCPN857_n_7802), .o(FE_OCP_RBN2613_FE_OCPN857_n_7802) );
in01s01 FE_OCP_RBC2614_FE_OCPN857_n_7802 ( .a(FE_OCP_RBN2612_FE_OCPN857_n_7802), .o(FE_OCP_RBN2614_FE_OCPN857_n_7802) );
in01s01 FE_OCP_RBC2616_FE_OCPN857_n_7802 ( .a(FE_OCP_RBN2613_FE_OCPN857_n_7802), .o(FE_OCP_RBN2616_FE_OCPN857_n_7802) );
in01s01 FE_OCP_RBC2620_n_24175 ( .a(FE_OCP_RBN6624_n_24175), .o(FE_OCP_RBN2620_n_24175) );
in01s01 FE_OCP_RBC2621_n_24175 ( .a(FE_OCP_RBN2620_n_24175), .o(FE_OCP_RBN2621_n_24175) );
in01s01 FE_OCP_RBC2622_n_24175 ( .a(FE_OCP_RBN2620_n_24175), .o(FE_OCP_RBN2622_n_24175) );
in01s02 FE_OCP_RBC2627_n_2737 ( .a(FE_OCP_RBN5661_n_2438), .o(FE_OCP_RBN2627_n_2737) );
in01s02 FE_OCP_RBC2629_n_2737 ( .a(FE_OCP_RBN5659_n_2438), .o(FE_OCP_RBN2629_n_2737) );
in01m03 FE_OCP_RBC2630_n_2737 ( .a(FE_OCP_RBN5659_n_2438), .o(FE_OCP_RBN2630_n_2737) );
in01s02 FE_OCP_RBC2631_n_9003 ( .a(n_9003), .o(FE_OCP_RBN2631_n_9003) );
in01s01 FE_OCP_RBC2632_n_9003 ( .a(FE_OCP_RBN2631_n_9003), .o(FE_OCP_RBN2632_n_9003) );
in01s01 FE_OCP_RBC2633_n_9003 ( .a(FE_OCP_RBN2631_n_9003), .o(FE_OCP_RBN2633_n_9003) );
in01s01 FE_OCP_RBC2634_n_9003 ( .a(FE_OCP_RBN2632_n_9003), .o(FE_OCP_RBN2634_n_9003) );
in01s01 FE_OCP_RBC2635_n_29371 ( .a(n_29371), .o(FE_OCP_RBN2635_n_29371) );
in01s03 FE_OCP_RBC2636_n_29371 ( .a(n_29371), .o(FE_OCP_RBN2636_n_29371) );
in01s01 FE_OCP_RBC2637_n_33954 ( .a(n_33954), .o(FE_OCP_RBN2637_n_33954) );
in01m02 FE_OCP_RBC2638_n_33954 ( .a(n_33954), .o(FE_OCP_RBN2638_n_33954) );
in01m01 FE_OCP_RBC2639_n_13667 ( .a(n_13667), .o(FE_OCP_RBN2639_n_13667) );
in01s01 FE_OCP_RBC2640_n_13667 ( .a(n_13667), .o(FE_OCP_RBN2640_n_13667) );
in01s01 FE_OCP_RBC2641_n_13667 ( .a(FE_OCP_RBN2640_n_13667), .o(FE_OCP_RBN2641_n_13667) );
in01s01 FE_OCP_RBC2642_n_13667 ( .a(FE_OCP_RBN2640_n_13667), .o(FE_OCP_RBN2642_n_13667) );
in01s01 FE_OCP_RBC2644_n_13667 ( .a(FE_OCP_RBN2641_n_13667), .o(FE_OCP_RBN2644_n_13667) );
in01s04 FE_OCP_RBC2645_n_2747 ( .a(n_2747), .o(FE_OCP_RBN2645_n_2747) );
in01s01 FE_OCP_RBC2646_n_2747 ( .a(n_2747), .o(FE_OCP_RBN2646_n_2747) );
in01m01 FE_OCP_RBC2649_n_8073 ( .a(n_8073), .o(FE_OCP_RBN2649_n_8073) );
in01s01 FE_OCP_RBC2650_n_29470 ( .a(n_29470), .o(FE_OCP_RBN2650_n_29470) );
in01m04 FE_OCP_RBC2651_n_29470 ( .a(n_29470), .o(FE_OCP_RBN2651_n_29470) );
in01s01 FE_OCP_RBC2652_n_29448 ( .a(n_29448), .o(FE_OCP_RBN2652_n_29448) );
in01m06 FE_OCP_RBC2653_n_29448 ( .a(n_29448), .o(FE_OCP_RBN2653_n_29448) );
in01s06 FE_OCP_RBC2654_FE_OCPN914_n_8091 ( .a(FE_OCPN914_n_8091), .o(FE_OCP_RBN2654_FE_OCPN914_n_8091) );
in01s01 FE_OCP_RBC2655_FE_OCPN914_n_8091 ( .a(FE_OCP_RBN2654_FE_OCPN914_n_8091), .o(FE_OCP_RBN2655_FE_OCPN914_n_8091) );
in01s01 FE_OCP_RBC2656_FE_OCPN914_n_8091 ( .a(FE_OCP_RBN2655_FE_OCPN914_n_8091), .o(FE_OCP_RBN2656_FE_OCPN914_n_8091) );
in01s01 FE_OCP_RBC2659_n_2832 ( .a(n_2832), .o(FE_OCP_RBN2659_n_2832) );
in01s01 FE_OCP_RBC2661_n_9304 ( .a(FE_OCP_RBN6635_n_9304), .o(FE_OCP_RBN2661_n_9304) );
in01s04 FE_OCP_RBC2662_n_19393 ( .a(n_19393), .o(FE_OCP_RBN2662_n_19393) );
in01m02 FE_OCP_RBC2663_n_19393 ( .a(n_19393), .o(FE_OCP_RBN2663_n_19393) );
in01s02 FE_OCP_RBC2664_n_24372 ( .a(n_24372), .o(FE_OCP_RBN2664_n_24372) );
in01s01 FE_OCP_RBC2665_n_24372 ( .a(n_24372), .o(FE_OCP_RBN2665_n_24372) );
in01s01 FE_OCP_RBC2666_n_24372 ( .a(n_24372), .o(FE_OCP_RBN2666_n_24372) );
in01s04 FE_OCP_RBC2667_n_24408 ( .a(n_24408), .o(FE_OCP_RBN2667_n_24408) );
in01s04 FE_OCP_RBC2668_n_29500 ( .a(n_29500), .o(FE_OCP_RBN2668_n_29500) );
in01f02 FE_OCP_RBC2669_n_29500 ( .a(n_29500), .o(FE_OCP_RBN2669_n_29500) );
in01s01 FE_OCP_RBC2670_n_46991 ( .a(n_46991), .o(FE_OCP_RBN2670_n_46991) );
in01s01 FE_OCP_RBC2672_n_38534 ( .a(n_38534), .o(FE_OCP_RBN2672_n_38534) );
in01m02 FE_OCP_RBC2673_n_38534 ( .a(n_38534), .o(FE_OCP_RBN2673_n_38534) );
in01s01 FE_OCP_RBC2674_n_8163 ( .a(n_8163), .o(FE_OCP_RBN2674_n_8163) );
in01s01 FE_OCP_RBC2675_n_8163 ( .a(n_8163), .o(FE_OCP_RBN2675_n_8163) );
in01s01 FE_OCP_RBC2676_n_8163 ( .a(FE_OCP_RBN2675_n_8163), .o(FE_OCP_RBN2676_n_8163) );
in01s01 FE_OCP_RBC2677_n_8163 ( .a(FE_OCP_RBN2676_n_8163), .o(FE_OCP_RBN2677_n_8163) );
in01s01 FE_OCP_RBC2678_n_8163 ( .a(FE_OCP_RBN2676_n_8163), .o(FE_OCP_RBN2678_n_8163) );
in01s01 FE_OCP_RBC2680_n_38515 ( .a(FE_OCP_RBN5690_n_38515), .o(FE_OCP_RBN2680_n_38515) );
in01s01 FE_OCP_RBC2681_n_38515 ( .a(FE_OCP_RBN2680_n_38515), .o(FE_OCP_RBN2681_n_38515) );
in01s01 FE_OCP_RBC2682_n_38515 ( .a(FE_OCP_RBN2680_n_38515), .o(FE_OCP_RBN2682_n_38515) );
in01f02 FE_OCP_RBC2683_n_13818 ( .a(n_13818), .o(FE_OCP_RBN2683_n_13818) );
in01s01 FE_OCP_RBC2684_n_13818 ( .a(n_13818), .o(FE_OCP_RBN2684_n_13818) );
in01m08 FE_OCP_RBC2687_n_44100 ( .a(n_44100), .o(FE_OCP_RBN2687_n_44100) );
in01s02 FE_OCP_RBC2688_n_44100 ( .a(FE_OCP_RBN2687_n_44100), .o(FE_OCP_RBN2688_n_44100) );
in01m10 FE_OCP_RBC2689_n_44100 ( .a(FE_OCP_RBN2687_n_44100), .o(FE_OCP_RBN2689_n_44100) );
in01s04 FE_OCP_RBC2690_n_8221 ( .a(n_8221), .o(FE_OCP_RBN2690_n_8221) );
in01s01 FE_OCP_RBC2691_n_8221 ( .a(FE_OCP_RBN2690_n_8221), .o(FE_OCP_RBN2691_n_8221) );
in01s01 FE_OCP_RBC2692_n_8221 ( .a(FE_OCP_RBN2691_n_8221), .o(FE_OCP_RBN2692_n_8221) );
in01s01 FE_OCP_RBC2693_n_24436 ( .a(n_24436), .o(FE_OCP_RBN2693_n_24436) );
in01s04 FE_OCP_RBC2694_n_24436 ( .a(n_24436), .o(FE_OCP_RBN2694_n_24436) );
in01s01 FE_OCP_RBC2695_n_24436 ( .a(n_24436), .o(FE_OCP_RBN2695_n_24436) );
in01f02 FE_OCP_RBC2696_n_13703 ( .a(n_13703), .o(FE_OCP_RBN2696_n_13703) );
in01s02 FE_OCP_RBC2697_n_13703 ( .a(n_13703), .o(FE_OCP_RBN2697_n_13703) );
in01s02 FE_OCP_RBC2701_n_8187 ( .a(FE_OCP_RBN6656_n_8187), .o(FE_OCP_RBN2701_n_8187) );
in01s02 FE_OCP_RBC2702_FE_RN_299_0 ( .a(FE_RN_299_0), .o(FE_OCP_RBN2702_FE_RN_299_0) );
in01f02 FE_OCP_RBC2703_FE_RN_984_0 ( .a(FE_RN_984_0), .o(FE_OCP_RBN2703_FE_RN_984_0) );
in01s04 FE_OCP_RBC2704_n_24510 ( .a(n_24510), .o(FE_OCP_RBN2704_n_24510) );
in01s01 FE_OCP_RBC2705_n_47023 ( .a(n_47023), .o(FE_OCP_RBN2705_n_47023) );
in01s01 FE_OCP_RBC2706_n_47023 ( .a(n_47023), .o(FE_OCP_RBN2706_n_47023) );
in01s02 FE_OCP_RBC2708_n_24505 ( .a(n_24505), .o(FE_OCP_RBN2708_n_24505) );
in01s01 FE_OCP_RBC2709_n_24505 ( .a(n_24505), .o(FE_OCP_RBN2709_n_24505) );
in01s01 FE_OCP_RBC2711_n_19599 ( .a(FE_OCP_RBN4182_n_19599), .o(FE_OCP_RBN2711_n_19599) );
in01m02 FE_OCP_RBC2712_n_24501 ( .a(n_24501), .o(FE_OCP_RBN2712_n_24501) );
in01s01 FE_OCP_RBC2713_n_24501 ( .a(FE_OCP_RBN2712_n_24501), .o(FE_OCP_RBN2713_n_24501) );
in01s01 FE_OCP_RBC2714_n_24501 ( .a(FE_OCP_RBN2713_n_24501), .o(FE_OCP_RBN2714_n_24501) );
in01s01 FE_OCP_RBC2715_n_24501 ( .a(FE_OCP_RBN2713_n_24501), .o(FE_OCP_RBN2715_n_24501) );
in01m02 FE_OCP_RBC2716_n_8242 ( .a(n_8242), .o(FE_OCP_RBN2716_n_8242) );
in01s01 FE_OCP_RBC2717_n_8242 ( .a(FE_OCP_RBN2716_n_8242), .o(FE_OCP_RBN2717_n_8242) );
in01s01 FE_OCP_RBC2719_n_8242 ( .a(FE_OCP_RBN2717_n_8242), .o(FE_OCP_RBN2719_n_8242) );
in01s02 FE_OCP_RBC2720_n_19601 ( .a(n_19601), .o(FE_OCP_RBN2720_n_19601) );
in01s01 FE_OCP_RBC2721_n_19601 ( .a(n_19601), .o(FE_OCP_RBN2721_n_19601) );
in01m04 FE_OCP_RBC2722_n_8243 ( .a(n_8243), .o(FE_OCP_RBN2722_n_8243) );
in01s02 FE_OCP_RBC2723_FE_RN_522_0 ( .a(FE_RN_522_0), .o(FE_OCP_RBN2723_FE_RN_522_0) );
in01s04 FE_OCP_RBC2724_n_14018 ( .a(n_14018), .o(FE_OCP_RBN2724_n_14018) );
in01s01 FE_OCP_RBC2725_n_14018 ( .a(n_14018), .o(FE_OCP_RBN2725_n_14018) );
in01s02 FE_OCP_RBC2726_n_14018 ( .a(FE_OCP_RBN2725_n_14018), .o(FE_OCP_RBN2726_n_14018) );
in01s02 FE_OCP_RBC2727_n_14018 ( .a(FE_OCP_RBN2726_n_14018), .o(FE_OCP_RBN2727_n_14018) );
in01m04 FE_OCP_RBC2728_n_14072 ( .a(n_14072), .o(FE_OCP_RBN2728_n_14072) );
in01s01 FE_OCP_RBC2729_n_14072 ( .a(FE_OCP_RBN2728_n_14072), .o(FE_OCP_RBN2729_n_14072) );
in01s01 FE_OCP_RBC2730_n_14072 ( .a(FE_OCP_RBN2729_n_14072), .o(FE_OCP_RBN2730_n_14072) );
in01s01 FE_OCP_RBC2731_n_14072 ( .a(FE_OCP_RBN2729_n_14072), .o(FE_OCP_RBN2731_n_14072) );
in01m01 FE_OCP_RBC2732_n_29657 ( .a(n_29657), .o(FE_OCP_RBN2732_n_29657) );
in01m04 FE_OCP_RBC2733_n_29657 ( .a(n_29657), .o(FE_OCP_RBN2733_n_29657) );
in01s02 FE_OCP_RBC2734_n_8402 ( .a(n_8402), .o(FE_OCP_RBN2734_n_8402) );
in01s01 FE_OCP_RBC2735_n_8402 ( .a(FE_OCP_RBN2734_n_8402), .o(FE_OCP_RBN2735_n_8402) );
in01s01 FE_OCP_RBC2737_n_8402 ( .a(FE_OCP_RBN5738_n_8402), .o(FE_OCP_RBN2737_n_8402) );
in01m02 FE_OCP_RBC2739_n_8300 ( .a(n_8300), .o(FE_OCP_RBN2739_n_8300) );
in01s02 FE_OCP_RBC2740_n_8398 ( .a(n_8398), .o(FE_OCP_RBN2740_n_8398) );
in01m02 FE_OCP_RBC2741_n_14114 ( .a(n_14114), .o(FE_OCP_RBN2741_n_14114) );
in01s01 FE_OCP_RBC2742_n_14114 ( .a(FE_OCP_RBN2741_n_14114), .o(FE_OCP_RBN2742_n_14114) );
in01s02 FE_OCP_RBC2743_n_14114 ( .a(FE_OCP_RBN2742_n_14114), .o(FE_OCP_RBN2743_n_14114) );
in01s01 FE_OCP_RBC2744_n_14114 ( .a(FE_OCP_RBN2743_n_14114), .o(FE_OCP_RBN2744_n_14114) );
in01s02 FE_OCP_RBC2745_n_19747 ( .a(n_19747), .o(FE_OCP_RBN2745_n_19747) );
in01m01 FE_OCP_RBC2746_n_19747 ( .a(n_19747), .o(FE_OCP_RBN2746_n_19747) );
in01s02 FE_OCP_RBC2747_n_8474 ( .a(n_8474), .o(FE_OCP_RBN2747_n_8474) );
in01s01 FE_OCP_RBC2748_n_8474 ( .a(FE_OCP_RBN2747_n_8474), .o(FE_OCP_RBN2748_n_8474) );
in01s04 FE_OCP_RBC2749_n_14157 ( .a(n_14157), .o(FE_OCP_RBN2749_n_14157) );
in01s01 FE_OCP_RBC2750_n_14157 ( .a(n_14157), .o(FE_OCP_RBN2750_n_14157) );
in01s01 FE_OCP_RBC2751_FE_RN_1223_0 ( .a(FE_RN_1223_0), .o(FE_OCP_RBN2751_FE_RN_1223_0) );
in01s01 FE_OCP_RBC2752_FE_RN_1223_0 ( .a(FE_RN_1223_0), .o(FE_OCP_RBN2752_FE_RN_1223_0) );
in01s01 FE_OCP_RBC2753_n_3016 ( .a(n_3016), .o(FE_OCP_RBN2753_n_3016) );
in01s02 FE_OCP_RBC2754_n_3016 ( .a(n_3016), .o(FE_OCP_RBN2754_n_3016) );
in01s01 FE_OCP_RBC2756_n_13796 ( .a(FE_OCP_RBN4188_n_13765), .o(FE_OCP_RBN2756_n_13796) );
in01s01 FE_OCP_RBC2757_n_13796 ( .a(FE_OCP_RBN4189_n_13765), .o(FE_OCP_RBN2757_n_13796) );
in01s10 FE_OCP_RBC2758_n_13796 ( .a(FE_OCP_RBN4189_n_13765), .o(FE_OCP_RBN2758_n_13796) );
in01s01 FE_OCP_RBC2759_n_13796 ( .a(FE_OCP_RBN4189_n_13765), .o(FE_OCP_RBN2759_n_13796) );
in01s01 FE_OCP_RBC2760_n_13796 ( .a(FE_OCP_RBN4189_n_13765), .o(FE_OCP_RBN2760_n_13796) );
in01s01 FE_OCP_RBC2762_n_13796 ( .a(FE_OCP_RBN2760_n_13796), .o(FE_OCP_RBN2762_n_13796) );
in01s02 FE_OCP_RBC2765_n_38530 ( .a(n_38530), .o(FE_OCP_RBN2765_n_38530) );
in01s01 FE_OCP_RBC2766_n_38530 ( .a(n_38530), .o(FE_OCP_RBN2766_n_38530) );
in01s01 FE_OCP_RBC2767_n_3035 ( .a(n_3035), .o(FE_OCP_RBN2767_n_3035) );
in01s02 FE_OCP_RBC2768_n_3167 ( .a(n_3167), .o(FE_OCP_RBN2768_n_3167) );
in01s02 FE_OCP_RBC2769_n_3238 ( .a(n_3238), .o(FE_OCP_RBN2769_n_3238) );
in01s01 FE_OCP_RBC2771_n_4336 ( .a(FE_OCP_RBN5741_n_4336), .o(FE_OCP_RBN2771_n_4336) );
in01s04 FE_OCP_RBC2772_n_45521 ( .a(n_45521), .o(FE_OCP_RBN2772_n_45521) );
in01s01 FE_OCP_RBC2775_n_8637 ( .a(FE_OCP_RBN5748_n_8637), .o(FE_OCP_RBN2775_n_8637) );
in01s01 FE_OCP_RBC2776_n_8637 ( .a(FE_OCP_RBN2775_n_8637), .o(FE_OCP_RBN2776_n_8637) );
in01s01 FE_OCP_RBC2778_n_8599 ( .a(FE_OCP_RBN5750_n_8599), .o(FE_OCP_RBN2778_n_8599) );
in01s01 FE_OCP_RBC2779_n_8599 ( .a(FE_OCP_RBN2778_n_8599), .o(FE_OCP_RBN2779_n_8599) );
in01s02 FE_OCP_RBC2780_n_8664 ( .a(n_8664), .o(FE_OCP_RBN2780_n_8664) );
in01s02 FE_OCP_RBC2781_n_8664 ( .a(n_8664), .o(FE_OCP_RBN2781_n_8664) );
in01s01 FE_OCP_RBC2782_n_8664 ( .a(FE_OCP_RBN2780_n_8664), .o(FE_OCP_RBN2782_n_8664) );
in01s01 FE_OCP_RBC2783_n_8664 ( .a(FE_OCP_RBN2782_n_8664), .o(FE_OCP_RBN2783_n_8664) );
in01s02 FE_OCP_RBC2785_n_8767 ( .a(n_8767), .o(FE_OCP_RBN2785_n_8767) );
in01s01 FE_OCP_RBC2786_n_8767 ( .a(n_8767), .o(FE_OCP_RBN2786_n_8767) );
in01s01 FE_OCP_RBC2789_n_8767 ( .a(FE_OCP_RBN2786_n_8767), .o(FE_OCP_RBN2789_n_8767) );
in01s01 FE_OCP_RBC2790_n_8767 ( .a(FE_OCP_RBN2789_n_8767), .o(FE_OCP_RBN2790_n_8767) );
in01f02 FE_OCP_RBC2791_FE_RN_368_0 ( .a(FE_RN_368_0), .o(FE_OCP_RBN2791_FE_RN_368_0) );
in01s01 FE_OCP_RBC2796_n_3250 ( .a(n_3250), .o(FE_OCP_RBN2796_n_3250) );
in01s02 FE_OCP_RBC2797_n_8530 ( .a(n_8530), .o(FE_OCP_RBN2797_n_8530) );
in01s04 FE_OCP_RBC2798_n_8817 ( .a(n_8817), .o(FE_OCP_RBN2798_n_8817) );
in01m04 FE_OCP_RBC2799_n_8817 ( .a(n_8817), .o(FE_OCP_RBN2799_n_8817) );
in01s01 FE_OCP_RBC2800_n_8817 ( .a(n_8817), .o(FE_OCP_RBN2800_n_8817) );
in01s02 FE_OCP_RBC2803_n_3220 ( .a(n_3220), .o(FE_OCP_RBN2803_n_3220) );
in01s02 FE_OCP_RBC2804_n_3261 ( .a(n_3261), .o(FE_OCP_RBN2804_n_3261) );
in01s01 FE_OCP_RBC2808_n_3338 ( .a(FE_OCP_RBN5770_n_3338), .o(FE_OCP_RBN2808_n_3338) );
in01s02 FE_OCP_RBC2810_n_8542 ( .a(n_8542), .o(FE_OCP_RBN2810_n_8542) );
in01s02 FE_OCP_RBC2811_n_8542 ( .a(FE_OCP_RBN2810_n_8542), .o(FE_OCP_RBN2811_n_8542) );
in01s01 FE_OCP_RBC2812_n_8835 ( .a(n_8835), .o(FE_OCP_RBN2812_n_8835) );
in01m02 FE_OCP_RBC2813_n_8835 ( .a(n_8835), .o(FE_OCP_RBN2813_n_8835) );
in01s01 FE_OCP_RBC2814_n_14441 ( .a(n_14441), .o(FE_OCP_RBN2814_n_14441) );
in01m02 FE_OCP_RBC2815_n_14441 ( .a(n_14441), .o(FE_OCP_RBN2815_n_14441) );
in01s01 FE_OCP_RBC2816_n_34509 ( .a(n_34509), .o(FE_OCP_RBN2816_n_34509) );
in01s02 FE_OCP_RBC2817_n_8939 ( .a(n_8939), .o(FE_OCP_RBN2817_n_8939) );
in01s01 FE_OCP_RBC2819_n_13962 ( .a(FE_OCP_RBN5776_n_13796), .o(FE_OCP_RBN2819_n_13962) );
in01s01 FE_OCP_RBC2820_n_13962 ( .a(FE_OCP_RBN4205_n_13796), .o(FE_OCP_RBN2820_n_13962) );
in01s01 FE_OCP_RBC2825_n_13962 ( .a(FE_OCP_RBN6695_n_13796), .o(FE_OCP_RBN2825_n_13962) );
in01s03 FE_OCP_RBC2828_n_13962 ( .a(FE_OCP_RBN6696_n_13796), .o(FE_OCP_RBN2828_n_13962) );
in01s01 FE_OCP_RBC2829_n_13962 ( .a(FE_OCP_RBN5797_n_13962), .o(FE_OCP_RBN2829_n_13962) );
in01s01 FE_OCP_RBC2830_n_13962 ( .a(FE_OCP_RBN2825_n_13962), .o(FE_OCP_RBN2830_n_13962) );
in01s40 FE_OCP_RBC2832_n_13962 ( .a(FE_OCP_RBN4232_n_13962), .o(FE_OCP_RBN2832_n_13962) );
in01s03 FE_OCP_RBC2833_n_13962 ( .a(FE_OCP_RBN4232_n_13962), .o(FE_OCP_RBN2833_n_13962) );
in01s03 FE_OCP_RBC2834_n_13962 ( .a(FE_OCP_RBN2828_n_13962), .o(FE_OCP_RBN2834_n_13962) );
in01s02 FE_OCP_RBC2835_n_13962 ( .a(FE_OCP_RBN2829_n_13962), .o(FE_OCP_RBN2835_n_13962) );
in01s40 FE_OCP_RBC2836_n_13962 ( .a(FE_OCP_RBN2832_n_13962), .o(FE_OCP_RBN2836_n_13962) );
in01s40 FE_OCP_RBC2837_n_13962 ( .a(FE_OCP_RBN2836_n_13962), .o(FE_OCP_RBN2837_n_13962) );
in01s02 FE_OCP_RBC2838_n_13962 ( .a(FE_OCP_RBN2836_n_13962), .o(FE_OCP_RBN2838_n_13962) );
in01f02 FE_OCP_RBC2839_n_8974 ( .a(n_8974), .o(FE_OCP_RBN2839_n_8974) );
in01s01 FE_OCP_RBC2841_n_9044 ( .a(n_9044), .o(FE_OCP_RBN2841_n_9044) );
in01m02 FE_OCP_RBC2842_n_9044 ( .a(n_9044), .o(FE_OCP_RBN2842_n_9044) );
in01s01 FE_OCP_RBC2845_n_47018 ( .a(FE_OCP_RBN5808_n_47018), .o(FE_OCP_RBN2845_n_47018) );
in01s01 FE_OCP_RBC2846_n_47018 ( .a(FE_OCP_RBN2845_n_47018), .o(FE_OCP_RBN2846_n_47018) );
in01s01 FE_OCP_RBC2847_n_47018 ( .a(FE_OCP_RBN2845_n_47018), .o(FE_OCP_RBN2847_n_47018) );
in01s01 FE_OCP_RBC2850_n_3645 ( .a(FE_OCP_RBN5811_n_3645), .o(FE_OCP_RBN2850_n_3645) );
in01s02 FE_OCP_RBC2851_n_4905 ( .a(n_4905), .o(FE_OCP_RBN2851_n_4905) );
in01s01 FE_OCP_RBC2852_n_4905 ( .a(n_4905), .o(FE_OCP_RBN2852_n_4905) );
in01s01 FE_OCP_RBC2853_n_4905 ( .a(FE_OCP_RBN2852_n_4905), .o(FE_OCP_RBN2853_n_4905) );
in01f01 FE_OCP_RBC2854_n_8692 ( .a(n_8692), .o(FE_OCP_RBN2854_n_8692) );
in01m02 FE_OCP_RBC2856_n_8755 ( .a(n_8755), .o(FE_OCP_RBN2856_n_8755) );
in01m02 FE_OCP_RBC2857_n_9082 ( .a(n_9082), .o(FE_OCP_RBN2857_n_9082) );
in01s01 FE_OCP_RBC2858_n_9082 ( .a(FE_OCP_RBN2857_n_9082), .o(FE_OCP_RBN2858_n_9082) );
in01s01 FE_OCP_RBC2859_n_9082 ( .a(FE_OCP_RBN2858_n_9082), .o(FE_OCP_RBN2859_n_9082) );
in01s04 FE_OCP_RBC2860_n_29800 ( .a(n_29800), .o(FE_OCP_RBN2860_n_29800) );
in01m06 FE_OCP_RBC2861_n_44921 ( .a(n_44921), .o(FE_OCP_RBN2861_n_44921) );
in01m02 FE_OCP_RBC2863_n_3468 ( .a(n_3468), .o(FE_OCP_RBN2863_n_3468) );
in01s01 FE_OCP_RBC2864_n_8714 ( .a(n_8714), .o(FE_OCP_RBN2864_n_8714) );
in01f02 FE_OCP_RBC2865_n_8850 ( .a(n_8850), .o(FE_OCP_RBN2865_n_8850) );
in01s01 FE_OCP_RBC2866_n_9347 ( .a(n_9347), .o(FE_OCP_RBN2866_n_9347) );
in01s02 FE_OCP_RBC2867_n_9347 ( .a(n_9347), .o(FE_OCP_RBN2867_n_9347) );
in01s02 FE_OCP_RBC2868_n_9188 ( .a(n_9188), .o(FE_OCP_RBN2868_n_9188) );
in01s01 FE_OCP_RBC2869_n_9188 ( .a(n_9188), .o(FE_OCP_RBN2869_n_9188) );
in01s01 FE_OCP_RBC2880_n_3539 ( .a(n_3539), .o(FE_OCP_RBN2880_n_3539) );
in01f01 FE_OCP_RBC2881_n_8872 ( .a(n_8872), .o(FE_OCP_RBN2881_n_8872) );
in01f06 FE_OCP_RBC2884_n_20127 ( .a(n_20127), .o(FE_OCP_RBN2884_n_20127) );
in01s02 FE_OCP_RBC2885_n_8806 ( .a(n_8806), .o(FE_OCP_RBN2885_n_8806) );
in01m02 FE_OCP_RBC2886_n_9017 ( .a(n_9017), .o(FE_OCP_RBN2886_n_9017) );
in01s02 FE_OCP_RBC2887_n_9492 ( .a(n_9492), .o(FE_OCP_RBN2887_n_9492) );
in01s01 FE_OCP_RBC2888_n_9492 ( .a(n_9492), .o(FE_OCP_RBN2888_n_9492) );
in01s01 FE_OCP_RBC2889_n_9492 ( .a(n_9492), .o(FE_OCP_RBN2889_n_9492) );
in01f02 FE_OCP_RBC2890_n_14460 ( .a(n_14460), .o(FE_OCP_RBN2890_n_14460) );
in01s01 FE_OCP_RBC2891_n_14460 ( .a(n_14460), .o(FE_OCP_RBN2891_n_14460) );
in01s01 FE_OCP_RBC2892_n_14460 ( .a(FE_OCP_RBN2891_n_14460), .o(FE_OCP_RBN2892_n_14460) );
in01s04 FE_OCP_RBC2895_n_35003 ( .a(n_35003), .o(FE_OCP_RBN2895_n_35003) );
in01s01 FE_OCP_RBC2896_n_35003 ( .a(n_35003), .o(FE_OCP_RBN2896_n_35003) );
in01f02 FE_OCP_RBC2897_n_38750 ( .a(n_38750), .o(FE_OCP_RBN2897_n_38750) );
in01s01 FE_OCP_RBC2899_n_3807 ( .a(FE_OCP_RBN5856_n_3807), .o(FE_OCP_RBN2899_n_3807) );
in01s01 FE_OCP_RBC2900_n_3807 ( .a(FE_OCP_RBN2899_n_3807), .o(FE_OCP_RBN2900_n_3807) );
in01s02 FE_OCP_RBC2901_n_3643 ( .a(n_3643), .o(FE_OCP_RBN2901_n_3643) );
in01s01 FE_OCP_RBC2902_n_8902 ( .a(n_8902), .o(FE_OCP_RBN2902_n_8902) );
in01s01 FE_OCP_RBC2903_n_8902 ( .a(n_8902), .o(FE_OCP_RBN2903_n_8902) );
in01f02 FE_OCP_RBC2904_n_14590 ( .a(n_14590), .o(FE_OCP_RBN2904_n_14590) );
in01s01 FE_OCP_RBC2905_n_14590 ( .a(n_14590), .o(FE_OCP_RBN2905_n_14590) );
in01s02 FE_OCP_RBC2907_n_25238 ( .a(FE_OCP_RBN5925_n_25211), .o(FE_OCP_RBN2907_n_25238) );
in01m10 FE_OCP_RBC2910_n_25178 ( .a(n_25178), .o(FE_OCP_RBN2910_n_25178) );
in01f01 FE_OCP_RBC2911_n_25178 ( .a(n_25178), .o(FE_OCP_RBN2911_n_25178) );
in01s01 FE_OCP_RBC2915_n_3878 ( .a(FE_OCP_RBN5868_n_3704), .o(FE_OCP_RBN2915_n_3878) );
in01s01 FE_OCP_RBC2920_n_3878 ( .a(FE_OCP_RBN6766_n_3704), .o(FE_OCP_RBN2920_n_3878) );
in01s01 FE_OCP_RBC2921_n_3878 ( .a(FE_OCP_RBN6766_n_3704), .o(FE_OCP_RBN2921_n_3878) );
in01s02 FE_OCP_RBC2922_n_9030 ( .a(n_9030), .o(FE_OCP_RBN2922_n_9030) );
in01s01 FE_OCP_RBC2923_n_9070 ( .a(n_9070), .o(FE_OCP_RBN2923_n_9070) );
in01s01 FE_OCP_RBC2924_n_9198 ( .a(FE_OCP_RBN6750_n_9198), .o(FE_OCP_RBN2924_n_9198) );
in01f02 FE_OCP_RBC2926_n_14684 ( .a(n_14684), .o(FE_OCP_RBN2926_n_14684) );
in01s01 FE_OCP_RBC2927_n_14684 ( .a(n_14684), .o(FE_OCP_RBN2927_n_14684) );
in01s02 FE_OCP_RBC2928_n_14923 ( .a(n_14923), .o(FE_OCP_RBN2928_n_14923) );
in01s01 FE_OCP_RBC2929_n_34971 ( .a(n_34971), .o(FE_OCP_RBN2929_n_34971) );
in01m08 FE_OCP_RBC2930_n_34971 ( .a(n_34971), .o(FE_OCP_RBN2930_n_34971) );
in01s01 FE_OCP_RBC2932_n_9075 ( .a(FE_OCP_RBN6759_n_9075), .o(FE_OCP_RBN2932_n_9075) );
in01s01 FE_OCP_RBC2933_n_9075 ( .a(FE_OCP_RBN2932_n_9075), .o(FE_OCP_RBN2933_n_9075) );
in01s01 FE_OCP_RBC2934_n_9075 ( .a(FE_OCP_RBN2932_n_9075), .o(FE_OCP_RBN2934_n_9075) );
in01m04 FE_OCP_RBC2935_n_25401 ( .a(n_25401), .o(FE_OCP_RBN2935_n_25401) );
in01s01 FE_OCP_RBC2936_n_8981 ( .a(n_8981), .o(FE_OCP_RBN2936_n_8981) );
in01m02 FE_OCP_RBC2937_n_8981 ( .a(n_8981), .o(FE_OCP_RBN2937_n_8981) );
in01s02 FE_OCP_RBC2938_n_47013 ( .a(n_47013), .o(FE_OCP_RBN2938_n_47013) );
in01s01 FE_OCP_RBC2939_n_47013 ( .a(n_47013), .o(FE_OCP_RBN2939_n_47013) );
in01s01 FE_OCP_RBC2941_n_4101 ( .a(FE_OCP_RBN5918_n_4101), .o(FE_OCP_RBN2941_n_4101) );
in01s01 FE_OCP_RBC2942_n_4101 ( .a(FE_OCP_RBN2941_n_4101), .o(FE_OCP_RBN2942_n_4101) );
in01m01 FE_OCP_RBC2943_n_20242 ( .a(n_20242), .o(FE_OCP_RBN2943_n_20242) );
in01s02 FE_OCP_RBC2944_n_20242 ( .a(n_20242), .o(FE_OCP_RBN2944_n_20242) );
in01s01 FE_OCP_RBC2950_n_4158 ( .a(n_4158), .o(FE_OCP_RBN2950_n_4158) );
in01s01 FE_OCP_RBC2951_n_3867 ( .a(n_3867), .o(FE_OCP_RBN2951_n_3867) );
in01s01 FE_OCP_RBC2952_n_3867 ( .a(n_3867), .o(FE_OCP_RBN2952_n_3867) );
in01s01 FE_OCP_RBC2953_n_3841 ( .a(n_3841), .o(FE_OCP_RBN2953_n_3841) );
in01s01 FE_OCP_RBC2960_n_4046 ( .a(FE_OCP_RBN6777_n_4046), .o(FE_OCP_RBN2960_n_4046) );
in01s01 FE_OCP_RBC2961_n_4046 ( .a(FE_OCP_RBN6777_n_4046), .o(FE_OCP_RBN2961_n_4046) );
in01s10 FE_OCP_RBC2962_n_4046 ( .a(FE_OCP_RBN6784_n_4046), .o(FE_OCP_RBN2962_n_4046) );
in01s01 FE_OCP_RBC2963_n_4046 ( .a(FE_OCP_RBN6783_n_4046), .o(FE_OCP_RBN2963_n_4046) );
in01s01 FE_OCP_RBC2964_n_4046 ( .a(FE_OCP_RBN2960_n_4046), .o(FE_OCP_RBN2964_n_4046) );
in01s01 FE_OCP_RBC2965_n_4046 ( .a(FE_OCP_RBN2962_n_4046), .o(FE_OCP_RBN2965_n_4046) );
in01s01 FE_OCP_RBC2966_n_4046 ( .a(FE_OCP_RBN2963_n_4046), .o(FE_OCP_RBN2966_n_4046) );
in01s01 FE_OCP_RBC2967_n_4046 ( .a(FE_OCP_RBN2965_n_4046), .o(FE_OCP_RBN2967_n_4046) );
in01s01 FE_OCP_RBC2968_n_4046 ( .a(FE_OCP_RBN2967_n_4046), .o(FE_OCP_RBN2968_n_4046) );
in01s01 FE_OCP_RBC2969_n_4046 ( .a(FE_OCP_RBN2968_n_4046), .o(FE_OCP_RBN2969_n_4046) );
in01s01 FE_OCP_RBC2970_n_9676 ( .a(n_9676), .o(FE_OCP_RBN2970_n_9676) );
in01s01 FE_OCP_RBC2971_n_9676 ( .a(n_9676), .o(FE_OCP_RBN2971_n_9676) );
in01s01 FE_OCP_RBC2973_n_14768 ( .a(FE_OCP_RBN4319_n_14768), .o(FE_OCP_RBN2973_n_14768) );
in01s01 FE_OCP_RBC2976_n_25295 ( .a(n_25295), .o(FE_OCP_RBN2976_n_25295) );
in01s01 FE_OCP_RBC2977_n_25509 ( .a(n_25509), .o(FE_OCP_RBN2977_n_25509) );
in01s01 FE_OCP_RBC2978_n_25562 ( .a(n_25562), .o(FE_OCP_RBN2978_n_25562) );
in01m01 FE_OCP_RBC2979_n_35213 ( .a(n_35213), .o(FE_OCP_RBN2979_n_35213) );
in01s01 FE_OCP_RBC2980_n_35213 ( .a(n_35213), .o(FE_OCP_RBN2980_n_35213) );
in01f02 FE_OCP_RBC2981_n_14814 ( .a(n_14814), .o(FE_OCP_RBN2981_n_14814) );
in01s01 FE_OCP_RBC2982_n_14814 ( .a(FE_OCP_RBN2981_n_14814), .o(FE_OCP_RBN2982_n_14814) );
in01s01 FE_OCP_RBC2983_n_14814 ( .a(FE_OCP_RBN2982_n_14814), .o(FE_OCP_RBN2983_n_14814) );
in01s01 FE_OCP_RBC2984_n_9247 ( .a(n_9247), .o(FE_OCP_RBN2984_n_9247) );
in01f02 FE_OCP_RBC2985_n_9247 ( .a(n_9247), .o(FE_OCP_RBN2985_n_9247) );
in01s01 FE_OCP_RBC2987_n_4238 ( .a(n_4238), .o(FE_OCP_RBN2987_n_4238) );
in01s02 FE_OCP_RBC2988_n_9182 ( .a(n_9182), .o(FE_OCP_RBN2988_n_9182) );
in01s01 FE_OCP_RBC2989_n_9182 ( .a(n_9182), .o(FE_OCP_RBN2989_n_9182) );
in01s01 FE_OCP_RBC2990_n_4041 ( .a(n_4041), .o(FE_OCP_RBN2990_n_4041) );
in01s01 FE_OCP_RBC2991_n_4041 ( .a(n_4041), .o(FE_OCP_RBN2991_n_4041) );
in01s02 FE_OCP_RBC2992_n_9413 ( .a(n_9413), .o(FE_OCP_RBN2992_n_9413) );
in01s01 FE_OCP_RBC2999_n_20374 ( .a(n_20374), .o(FE_OCP_RBN2999_n_20374) );
in01s01 FE_OCP_RBC3000_n_20374 ( .a(n_20374), .o(FE_OCP_RBN3000_n_20374) );
in01s02 FE_OCP_RBC3001_n_20400 ( .a(n_20400), .o(FE_OCP_RBN3001_n_20400) );
in01s02 FE_OCP_RBC3002_n_20400 ( .a(n_20400), .o(FE_OCP_RBN3002_n_20400) );
in01s02 FE_OCP_RBC3003_n_20432 ( .a(n_20432), .o(FE_OCP_RBN3003_n_20432) );
in01s01 FE_OCP_RBC3005_n_14905 ( .a(FE_OCP_RBN5968_n_14905), .o(FE_OCP_RBN3005_n_14905) );
in01s01 FE_OCP_RBC3006_n_14905 ( .a(FE_OCP_RBN3005_n_14905), .o(FE_OCP_RBN3006_n_14905) );
in01s01 FE_OCP_RBC3007_n_15206 ( .a(n_15206), .o(FE_OCP_RBN3007_n_15206) );
in01f02 FE_OCP_RBC3008_n_15206 ( .a(n_15206), .o(FE_OCP_RBN3008_n_15206) );
in01s02 FE_OCP_RBC3011_n_9565 ( .a(n_9565), .o(FE_OCP_RBN3011_n_9565) );
in01s01 FE_OCP_RBC3012_n_14985 ( .a(n_14985), .o(FE_OCP_RBN3012_n_14985) );
in01m02 FE_OCP_RBC3013_n_14985 ( .a(n_14985), .o(FE_OCP_RBN3013_n_14985) );
in01s01 FE_OCP_RBC3014_n_15055 ( .a(n_15055), .o(FE_OCP_RBN3014_n_15055) );
in01s02 FE_OCP_RBC3015_n_15300 ( .a(n_15300), .o(FE_OCP_RBN3015_n_15300) );
in01s01 FE_OCP_RBC3016_n_15300 ( .a(n_15300), .o(FE_OCP_RBN3016_n_15300) );
in01s10 FE_OCP_RBC3017_n_20404 ( .a(n_20404), .o(FE_OCP_RBN3017_n_20404) );
in01s10 FE_OCP_RBC3018_n_20404 ( .a(FE_OCP_RBN3017_n_20404), .o(FE_OCP_RBN3018_n_20404) );
in01s01 FE_OCP_RBC3021_n_15319 ( .a(n_15319), .o(FE_OCP_RBN3021_n_15319) );
in01s01 FE_OCP_RBC3022_n_15319 ( .a(n_15319), .o(FE_OCP_RBN3022_n_15319) );
in01s02 FE_OCP_RBC3023_n_47011 ( .a(n_47011), .o(FE_OCP_RBN3023_n_47011) );
in01s01 FE_OCP_RBC3024_n_47011 ( .a(n_47011), .o(FE_OCP_RBN3024_n_47011) );
in01s01 FE_OCP_RBC3025_n_4065 ( .a(n_4065), .o(FE_OCP_RBN3025_n_4065) );
in01s01 FE_OCP_RBC3026_n_4699 ( .a(FE_OCP_RBN4340_n_4403), .o(FE_OCP_RBN3026_n_4699) );
in01m02 FE_OCP_RBC3028_n_9584 ( .a(n_9584), .o(FE_OCP_RBN3028_n_9584) );
in01s01 FE_OCP_RBC3029_n_9584 ( .a(n_9584), .o(FE_OCP_RBN3029_n_9584) );
in01s01 FE_OCP_RBC3030_n_9624 ( .a(n_9624), .o(FE_OCP_RBN3030_n_9624) );
in01m02 FE_OCP_RBC3031_n_9624 ( .a(n_9624), .o(FE_OCP_RBN3031_n_9624) );
in01s06 FE_OCP_RBC3032_n_15150 ( .a(FE_OCP_RBN5948_n_14982), .o(FE_OCP_RBN3032_n_15150) );
in01m02 FE_OCP_RBC3033_n_9629 ( .a(n_9629), .o(FE_OCP_RBN3033_n_9629) );
in01s01 FE_OCP_RBC3034_n_9629 ( .a(n_9629), .o(FE_OCP_RBN3034_n_9629) );
in01s01 FE_OCP_RBC3036_n_15079 ( .a(FE_OCP_RBN5985_n_15079), .o(FE_OCP_RBN3036_n_15079) );
in01s01 FE_OCP_RBC3037_n_15079 ( .a(FE_OCP_RBN3036_n_15079), .o(FE_OCP_RBN3037_n_15079) );
in01s01 FE_OCP_RBC3039_n_9494 ( .a(n_9494), .o(FE_OCP_RBN3039_n_9494) );
in01f08 FE_OCP_RBC3040_n_45139 ( .a(n_45139), .o(FE_OCP_RBN3040_n_45139) );
in01s06 FE_OCP_RBC3041_n_45139 ( .a(FE_OCP_RBN3040_n_45139), .o(FE_OCP_RBN3041_n_45139) );
in01s01 FE_OCP_RBC3042_n_4296 ( .a(n_4296), .o(FE_OCP_RBN3042_n_4296) );
in01s01 FE_OCP_RBC3043_n_4296 ( .a(n_4296), .o(FE_OCP_RBN3043_n_4296) );
in01s02 FE_OCP_RBC3044_n_4449 ( .a(n_4449), .o(FE_OCP_RBN3044_n_4449) );
in01m02 FE_OCP_RBC3045_n_9621 ( .a(n_9621), .o(FE_OCP_RBN3045_n_9621) );
in01s01 FE_OCP_RBC3048_n_15200 ( .a(n_15200), .o(FE_OCP_RBN3048_n_15200) );
in01f02 FE_OCP_RBC3049_n_15200 ( .a(n_15200), .o(FE_OCP_RBN3049_n_15200) );
in01s01 FE_OCP_RBC3050_n_4376 ( .a(n_4376), .o(FE_OCP_RBN3050_n_4376) );
in01s10 FE_OCP_RBC3052_n_10100 ( .a(n_10100), .o(FE_OCP_RBN3052_n_10100) );
in01s01 FE_OCP_RBC3057_n_10100 ( .a(FE_OCP_RBN4355_n_10100), .o(FE_OCP_RBN3057_n_10100) );
in01f02 FE_OCP_RBC3058_n_15595 ( .a(n_15595), .o(FE_OCP_RBN3058_n_15595) );
in01s01 FE_OCP_RBC3059_n_15595 ( .a(FE_OCP_RBN3058_n_15595), .o(FE_OCP_RBN3059_n_15595) );
in01s01 FE_OCP_RBC3060_n_15595 ( .a(FE_OCP_RBN3059_n_15595), .o(FE_OCP_RBN3060_n_15595) );
in01m01 FE_OCP_RBC3061_n_30575 ( .a(n_30575), .o(FE_OCP_RBN3061_n_30575) );
in01f02 FE_OCP_RBC3062_n_9859 ( .a(n_9859), .o(FE_OCP_RBN3062_n_9859) );
in01s01 FE_OCP_RBC3063_n_9859 ( .a(n_9859), .o(FE_OCP_RBN3063_n_9859) );
in01s01 FE_OCP_RBC3064_n_9892 ( .a(n_9892), .o(FE_OCP_RBN3064_n_9892) );
in01m02 FE_OCP_RBC3065_n_9892 ( .a(n_9892), .o(FE_OCP_RBN3065_n_9892) );
in01s01 FE_OCP_RBC3066_n_4294 ( .a(n_4294), .o(FE_OCP_RBN3066_n_4294) );
in01s02 FE_OCP_RBC3067_n_4294 ( .a(n_4294), .o(FE_OCP_RBN3067_n_4294) );
in01m02 FE_OCP_RBC3068_n_9910 ( .a(n_9910), .o(FE_OCP_RBN3068_n_9910) );
in01s01 FE_OCP_RBC3069_n_9910 ( .a(n_9910), .o(FE_OCP_RBN3069_n_9910) );
in01f02 FE_OCP_RBC3070_n_15275 ( .a(n_15275), .o(FE_OCP_RBN3070_n_15275) );
in01f02 FE_OCP_RBC3071_n_15433 ( .a(n_15433), .o(FE_OCP_RBN3071_n_15433) );
in01s01 FE_OCP_RBC3072_n_15433 ( .a(n_15433), .o(FE_OCP_RBN3072_n_15433) );
in01f02 FE_OCP_RBC3073_n_15706 ( .a(n_15706), .o(FE_OCP_RBN3073_n_15706) );
in01s01 FE_OCP_RBC3074_n_15706 ( .a(FE_OCP_RBN3073_n_15706), .o(FE_OCP_RBN3074_n_15706) );
in01s01 FE_OCP_RBC3075_n_15706 ( .a(FE_OCP_RBN3074_n_15706), .o(FE_OCP_RBN3075_n_15706) );
in01f04 FE_OCP_RBC3076_n_25816 ( .a(n_25816), .o(FE_OCP_RBN3076_n_25816) );
in01s01 FE_OCP_RBC3077_n_25816 ( .a(FE_OCP_RBN3076_n_25816), .o(FE_OCP_RBN3077_n_25816) );
in01s02 FE_OCP_RBC3078_n_25816 ( .a(FE_OCP_RBN3077_n_25816), .o(FE_OCP_RBN3078_n_25816) );
in01m04 FE_OCP_RBC3079_n_30643 ( .a(n_30643), .o(FE_OCP_RBN3079_n_30643) );
in01s01 FE_OCP_RBC3080_n_30643 ( .a(n_30643), .o(FE_OCP_RBN3080_n_30643) );
in01m06 FE_OCP_RBC3081_n_39514 ( .a(n_39514), .o(FE_OCP_RBN3081_n_39514) );
in01f02 FE_OCP_RBC3082_n_15314 ( .a(n_15314), .o(FE_OCP_RBN3082_n_15314) );
in01s01 FE_OCP_RBC3083_n_15314 ( .a(FE_OCP_RBN3082_n_15314), .o(FE_OCP_RBN3083_n_15314) );
in01s01 FE_OCP_RBC3084_n_15314 ( .a(FE_OCP_RBN3083_n_15314), .o(FE_OCP_RBN3084_n_15314) );
in01s01 FE_OCP_RBC3086_n_10015 ( .a(n_10015), .o(FE_OCP_RBN3086_n_10015) );
in01s01 FE_OCP_RBC3087_n_4458 ( .a(n_4458), .o(FE_OCP_RBN3087_n_4458) );
in01s02 FE_OCP_RBC3088_n_4458 ( .a(n_4458), .o(FE_OCP_RBN3088_n_4458) );
in01s01 FE_OCP_RBC3089_n_4872 ( .a(n_4872), .o(FE_OCP_RBN3089_n_4872) );
in01s01 FE_OCP_RBC3090_n_4872 ( .a(n_4872), .o(FE_OCP_RBN3090_n_4872) );
in01f02 FE_OCP_RBC3091_n_10023 ( .a(n_10023), .o(FE_OCP_RBN3091_n_10023) );
in01s01 FE_OCP_RBC3092_n_10023 ( .a(n_10023), .o(FE_OCP_RBN3092_n_10023) );
in01s01 FE_OCP_RBC3093_n_10023 ( .a(FE_OCP_RBN3092_n_10023), .o(FE_OCP_RBN3093_n_10023) );
in01s01 FE_OCP_RBC3094_n_10023 ( .a(FE_OCP_RBN3093_n_10023), .o(FE_OCP_RBN3094_n_10023) );
in01s01 FE_OCP_RBC3095_n_10023 ( .a(FE_OCP_RBN3093_n_10023), .o(FE_OCP_RBN3095_n_10023) );
in01f04 FE_OCP_RBC3098_n_15561 ( .a(n_15561), .o(FE_OCP_RBN3098_n_15561) );
in01f04 FE_OCP_RBC3099_n_15561 ( .a(FE_OCP_RBN3098_n_15561), .o(FE_OCP_RBN3099_n_15561) );
in01s06 FE_OCP_RBC3102_n_15768 ( .a(n_15768), .o(FE_OCP_RBN3102_n_15768) );
in01s03 FE_OCP_RBC3103_n_20710 ( .a(n_20710), .o(FE_OCP_RBN3103_n_20710) );
in01f02 FE_OCP_RBC3105_n_25819 ( .a(n_25819), .o(FE_OCP_RBN3105_n_25819) );
in01f04 FE_OCP_RBC3106_n_25849 ( .a(n_25849), .o(FE_OCP_RBN3106_n_25849) );
in01f06 FE_OCP_RBC3107_n_39531 ( .a(n_39531), .o(FE_OCP_RBN3107_n_39531) );
in01s01 FE_OCP_RBC3108_n_39531 ( .a(n_39531), .o(FE_OCP_RBN3108_n_39531) );
in01m02 FE_OCP_RBC3109_n_15817 ( .a(n_15817), .o(FE_OCP_RBN3109_n_15817) );
in01s01 FE_OCP_RBC3110_n_15817 ( .a(FE_OCP_RBN3109_n_15817), .o(FE_OCP_RBN3110_n_15817) );
in01s01 FE_OCP_RBC3111_n_15817 ( .a(FE_OCP_RBN3110_n_15817), .o(FE_OCP_RBN3111_n_15817) );
in01s02 FE_OCP_RBC3112_n_10025 ( .a(n_10025), .o(FE_OCP_RBN3112_n_10025) );
in01f02 FE_OCP_RBC3113_n_10195 ( .a(n_10195), .o(FE_OCP_RBN3113_n_10195) );
in01f02 FE_OCP_RBC3114_n_10198 ( .a(n_10198), .o(FE_OCP_RBN3114_n_10198) );
in01s01 FE_OCP_RBC3115_n_10198 ( .a(FE_OCP_RBN3114_n_10198), .o(FE_OCP_RBN3115_n_10198) );
in01s01 FE_OCP_RBC3116_n_10198 ( .a(FE_OCP_RBN3115_n_10198), .o(FE_OCP_RBN3116_n_10198) );
in01s01 FE_OCP_RBC3118_n_20812 ( .a(n_20812), .o(FE_OCP_RBN3118_n_20812) );
in01s02 FE_OCP_RBC3120_n_4751 ( .a(n_4751), .o(FE_OCP_RBN3120_n_4751) );
in01s01 FE_OCP_RBC3121_n_4751 ( .a(n_4751), .o(FE_OCP_RBN3121_n_4751) );
in01s01 FE_OCP_RBC3122_n_4784 ( .a(n_4784), .o(FE_OCP_RBN3122_n_4784) );
in01s02 FE_OCP_RBC3123_n_4784 ( .a(n_4784), .o(FE_OCP_RBN3123_n_4784) );
in01m02 FE_OCP_RBC3124_n_5121 ( .a(n_5121), .o(FE_OCP_RBN3124_n_5121) );
in01m02 FE_OCP_RBC3125_n_15856 ( .a(n_15856), .o(FE_OCP_RBN3125_n_15856) );
in01s01 FE_OCP_RBC3126_n_21051 ( .a(n_21051), .o(FE_OCP_RBN3126_n_21051) );
in01s02 FE_OCP_RBC3127_n_21051 ( .a(n_21051), .o(FE_OCP_RBN3127_n_21051) );
in01s01 FE_OCP_RBC3128_n_21051 ( .a(n_21051), .o(FE_OCP_RBN3128_n_21051) );
in01s01 FE_OCP_RBC3129_n_21051 ( .a(FE_OCP_RBN3127_n_21051), .o(FE_OCP_RBN3129_n_21051) );
in01s02 FE_OCP_RBC3130_n_21051 ( .a(FE_OCP_RBN3128_n_21051), .o(FE_OCP_RBN3130_n_21051) );
in01s02 FE_OCP_RBC3131_n_21051 ( .a(FE_OCP_RBN3129_n_21051), .o(FE_OCP_RBN3131_n_21051) );
in01s01 FE_OCP_RBC3134_n_46982 ( .a(n_46982), .o(FE_OCP_RBN3134_n_46982) );
in01s01 FE_OCP_RBC3135_n_10274 ( .a(n_10274), .o(FE_OCP_RBN3135_n_10274) );
in01m01 FE_OCP_RBC3136_n_10274 ( .a(n_10274), .o(FE_OCP_RBN3136_n_10274) );
in01s01 FE_OCP_RBC3137_n_10326 ( .a(n_10326), .o(FE_OCP_RBN3137_n_10326) );
in01f02 FE_OCP_RBC3138_n_10326 ( .a(n_10326), .o(FE_OCP_RBN3138_n_10326) );
in01m02 FE_OCP_RBC3140_n_30849 ( .a(n_30849), .o(FE_OCP_RBN3140_n_30849) );
in01s01 FE_OCP_RBC3141_n_30849 ( .a(n_30849), .o(FE_OCP_RBN3141_n_30849) );
in01s01 FE_OCP_RBC3143_n_4858 ( .a(FE_OCP_RBN6026_n_4858), .o(FE_OCP_RBN3143_n_4858) );
in01s01 FE_OCP_RBC3144_n_4858 ( .a(FE_OCP_RBN3143_n_4858), .o(FE_OCP_RBN3144_n_4858) );
in01s02 FE_OCP_RBC3145_n_5085 ( .a(n_5085), .o(FE_OCP_RBN3145_n_5085) );
in01s02 FE_OCP_RBC3146_n_10369 ( .a(n_10369), .o(FE_OCP_RBN3146_n_10369) );
in01s01 FE_OCP_RBC3147_n_10369 ( .a(FE_OCPN4859_n_10369), .o(FE_OCP_RBN3147_n_10369) );
in01s02 FE_OCP_RBC3148_n_15584 ( .a(n_15584), .o(FE_OCP_RBN3148_n_15584) );
in01f02 FE_OCP_RBC3149_n_15553 ( .a(n_15553), .o(FE_OCP_RBN3149_n_15553) );
in01s04 FE_OCP_RBC3150_n_25925 ( .a(n_25925), .o(FE_OCP_RBN3150_n_25925) );
in01s01 FE_OCP_RBC3152_n_46962 ( .a(FE_OCP_RBN6034_n_46962), .o(FE_OCP_RBN3152_n_46962) );
in01m04 FE_OCP_RBC3153_n_15804 ( .a(n_15804), .o(FE_OCP_RBN3153_n_15804) );
in01s02 FE_OCP_RBC3154_n_15804 ( .a(n_15804), .o(FE_OCP_RBN3154_n_15804) );
in01s01 FE_OCP_RBC3155_n_4925 ( .a(n_4925), .o(FE_OCP_RBN3155_n_4925) );
in01s01 FE_OCP_RBC3156_n_4925 ( .a(n_4925), .o(FE_OCP_RBN3156_n_4925) );
in01s01 FE_OCP_RBC3160_n_10399 ( .a(FE_OCP_RBN6037_n_10399), .o(FE_OCP_RBN3160_n_10399) );
in01s01 FE_OCP_RBC3161_n_10399 ( .a(FE_OCP_RBN3160_n_10399), .o(FE_OCP_RBN3161_n_10399) );
in01s02 FE_OCP_RBC3167_n_44211 ( .a(FE_OCP_RBN6044_n_35487), .o(FE_OCP_RBN3167_n_44211) );
in01s10 FE_OCP_RBC3168_n_44211 ( .a(FE_OCP_RBN6045_n_35487), .o(FE_OCP_RBN3168_n_44211) );
in01s01 FE_OCP_RBC3169_n_44211 ( .a(FE_OCP_RBN6045_n_35487), .o(FE_OCP_RBN3169_n_44211) );
in01s06 FE_OCP_RBC3170_n_44211 ( .a(FE_OCP_RBN6045_n_35487), .o(FE_OCP_RBN3170_n_44211) );
in01m08 FE_OCP_RBC3171_n_44211 ( .a(FE_OCP_RBN6045_n_35487), .o(FE_OCP_RBN3171_n_44211) );
in01s04 FE_OCP_RBC3172_n_10134 ( .a(n_10134), .o(FE_OCP_RBN3172_n_10134) );
in01s02 FE_OCP_RBC3173_n_26178 ( .a(n_26178), .o(FE_OCP_RBN3173_n_26178) );
in01s02 FE_OCP_RBC3174_n_26158 ( .a(n_26158), .o(FE_OCP_RBN3174_n_26158) );
in01m02 FE_OCP_RBC3175_n_31001 ( .a(n_31001), .o(FE_OCP_RBN3175_n_31001) );
in01s02 FE_OCP_RBC3176_n_39640 ( .a(n_39640), .o(FE_OCP_RBN3176_n_39640) );
in01s01 FE_OCP_RBC3177_n_39640 ( .a(n_39640), .o(FE_OCP_RBN3177_n_39640) );
in01s04 FE_OCP_RBC3178_n_16088 ( .a(n_16088), .o(FE_OCP_RBN3178_n_16088) );
in01s01 FE_OCP_RBC3179_n_16088 ( .a(n_16088), .o(FE_OCP_RBN3179_n_16088) );
in01s02 FE_OCP_RBC3180_n_4959 ( .a(n_4959), .o(FE_OCP_RBN3180_n_4959) );
in01s01 FE_OCP_RBC3181_n_10477 ( .a(n_10477), .o(FE_OCP_RBN3181_n_10477) );
in01m02 FE_OCP_RBC3182_n_10477 ( .a(n_10477), .o(FE_OCP_RBN3182_n_10477) );
in01s02 FE_OCP_RBC3185_n_15599 ( .a(FE_OCP_RBN6828_n_15514), .o(FE_OCP_RBN3185_n_15599) );
in01s02 FE_OCP_RBC3186_n_15599 ( .a(FE_OCP_RBN3185_n_15599), .o(FE_OCP_RBN3186_n_15599) );
in01s02 FE_OCP_RBC3190_n_15599 ( .a(FE_OCP_RBN6844_n_15599), .o(FE_OCP_RBN3190_n_15599) );
in01s01 FE_OCP_RBC3192_n_15599 ( .a(FE_OCP_RBN6847_n_15599), .o(FE_OCP_RBN3192_n_15599) );
in01s03 FE_OCP_RBC3193_n_15599 ( .a(FE_OCP_RBN6848_n_15599), .o(FE_OCP_RBN3193_n_15599) );
in01s01 FE_OCP_RBC3194_n_15599 ( .a(FE_OCP_RBN6848_n_15599), .o(FE_OCP_RBN3194_n_15599) );
in01s01 FE_OCP_RBC3195_n_15599 ( .a(FE_OCP_RBN3192_n_15599), .o(FE_OCP_RBN3195_n_15599) );
in01s02 FE_OCP_RBC3196_n_15599 ( .a(FE_OCP_RBN3193_n_15599), .o(FE_OCP_RBN3196_n_15599) );
in01s01 FE_OCP_RBC3197_n_15599 ( .a(FE_OCP_RBN3193_n_15599), .o(FE_OCP_RBN3197_n_15599) );
in01s01 FE_OCP_RBC3198_n_15599 ( .a(FE_OCP_RBN3193_n_15599), .o(FE_OCP_RBN3198_n_15599) );
in01s01 FE_OCP_RBC3199_n_15599 ( .a(FE_OCP_RBN3198_n_15599), .o(FE_OCP_RBN3199_n_15599) );
in01s04 FE_OCP_RBC3202_n_15900 ( .a(n_15900), .o(FE_OCP_RBN3202_n_15900) );
in01s01 FE_OCP_RBC3203_n_15900 ( .a(n_15900), .o(FE_OCP_RBN3203_n_15900) );
in01s01 FE_OCP_RBC3204_n_15900 ( .a(FE_OCP_RBN3203_n_15900), .o(FE_OCP_RBN3204_n_15900) );
in01s03 FE_OCP_RBC3205_n_26042 ( .a(n_26042), .o(FE_OCP_RBN3205_n_26042) );
in01s01 FE_OCP_RBC3206_n_35517 ( .a(n_35517), .o(FE_OCP_RBN3206_n_35517) );
in01s02 FE_OCP_RBC3207_n_39662 ( .a(n_39662), .o(FE_OCP_RBN3207_n_39662) );
in01s01 FE_OCP_RBC3209_n_5221 ( .a(n_5221), .o(FE_OCP_RBN3209_n_5221) );
in01s01 FE_OCP_RBC3210_n_21203 ( .a(n_21203), .o(FE_OCP_RBN3210_n_21203) );
in01s02 FE_OCP_RBC3211_n_21203 ( .a(n_21203), .o(FE_OCP_RBN3211_n_21203) );
in01m02 FE_OCP_RBC3212_n_10568 ( .a(n_10568), .o(FE_OCP_RBN3212_n_10568) );
in01s01 FE_OCP_RBC3213_n_10568 ( .a(FE_OCP_RBN3212_n_10568), .o(FE_OCP_RBN3213_n_10568) );
in01s01 FE_OCP_RBC3214_n_10568 ( .a(FE_OCP_RBN3213_n_10568), .o(FE_OCP_RBN3214_n_10568) );
in01s02 FE_OCP_RBC3215_n_5003 ( .a(n_5003), .o(FE_OCP_RBN3215_n_5003) );
in01s01 FE_OCP_RBC3216_n_5003 ( .a(n_5003), .o(FE_OCP_RBN3216_n_5003) );
in01m02 FE_OCP_RBC3217_n_15758 ( .a(n_15758), .o(FE_OCP_RBN3217_n_15758) );
in01m02 FE_OCP_RBC3218_n_15992 ( .a(n_15992), .o(FE_OCP_RBN3218_n_15992) );
in01s01 FE_OCP_RBC3219_n_15992 ( .a(FE_OCP_RBN3218_n_15992), .o(FE_OCP_RBN3219_n_15992) );
in01s01 FE_OCP_RBC3220_n_15992 ( .a(FE_OCP_RBN3219_n_15992), .o(FE_OCP_RBN3220_n_15992) );
in01s03 FE_OCP_RBC3221_n_21242 ( .a(n_21242), .o(FE_OCP_RBN3221_n_21242) );
in01s01 FE_OCP_RBC3222_n_21242 ( .a(n_21242), .o(FE_OCP_RBN3222_n_21242) );
in01s04 FE_OCP_RBC3224_n_39575 ( .a(n_39575), .o(FE_OCP_RBN3224_n_39575) );
in01s01 FE_OCP_RBC3225_n_39575 ( .a(FE_OCP_RBN3224_n_39575), .o(FE_OCP_RBN3225_n_39575) );
in01s01 FE_OCP_RBC3226_n_39575 ( .a(FE_OCP_RBN3225_n_39575), .o(FE_OCP_RBN3226_n_39575) );
in01s02 FE_OCP_RBC3227_n_10644 ( .a(n_10644), .o(FE_OCP_RBN3227_n_10644) );
in01s01 FE_OCP_RBC3228_n_10644 ( .a(FE_OCP_RBN3227_n_10644), .o(FE_OCP_RBN3228_n_10644) );
in01s01 FE_OCP_RBC3229_n_10644 ( .a(FE_OCP_RBN3228_n_10644), .o(FE_OCP_RBN3229_n_10644) );
in01m02 FE_OCP_RBC3230_n_31107 ( .a(n_31107), .o(FE_OCP_RBN3230_n_31107) );
in01s01 FE_OCP_RBC3231_n_31107 ( .a(n_31107), .o(FE_OCP_RBN3231_n_31107) );
in01s01 FE_OCP_RBC3233_n_16041 ( .a(FE_OCP_RBN6071_n_16041), .o(FE_OCP_RBN3233_n_16041) );
in01s01 FE_OCP_RBC3234_n_16041 ( .a(FE_OCP_RBN3233_n_16041), .o(FE_OCP_RBN3234_n_16041) );
in01s01 FE_OCP_RBC3235_n_16041 ( .a(FE_OCP_RBN3233_n_16041), .o(FE_OCP_RBN3235_n_16041) );
in01s01 FE_OCP_RBC3236_n_5130 ( .a(n_5130), .o(FE_OCP_RBN3236_n_5130) );
in01s01 FE_OCP_RBC3237_n_5130 ( .a(n_5130), .o(FE_OCP_RBN3237_n_5130) );
in01s01 FE_OCP_RBC3238_n_5307 ( .a(n_5307), .o(FE_OCP_RBN3238_n_5307) );
in01s01 FE_OCP_RBC3239_n_5307 ( .a(n_5307), .o(FE_OCP_RBN3239_n_5307) );
in01m02 FE_OCP_RBC3240_n_10612 ( .a(n_10612), .o(FE_OCP_RBN3240_n_10612) );
in01s01 FE_OCP_RBC3241_n_10612 ( .a(n_10612), .o(FE_OCP_RBN3241_n_10612) );
in01s02 FE_OCP_RBC3242_n_10676 ( .a(n_10676), .o(FE_OCP_RBN3242_n_10676) );
in01s01 FE_OCP_RBC3243_n_10676 ( .a(n_10676), .o(FE_OCP_RBN3243_n_10676) );
in01s02 FE_OCP_RBC3244_n_21269 ( .a(n_21269), .o(FE_OCP_RBN3244_n_21269) );
in01s02 FE_OCP_RBC3245_n_21351 ( .a(n_21351), .o(FE_OCP_RBN3245_n_21351) );
in01m02 FE_OCP_RBC3246_n_26169 ( .a(n_26169), .o(FE_OCP_RBN3246_n_26169) );
in01s01 FE_OCP_RBC3247_n_26169 ( .a(n_26169), .o(FE_OCP_RBN3247_n_26169) );
in01f02 FE_OCP_RBC3248_n_39697 ( .a(n_39697), .o(FE_OCP_RBN3248_n_39697) );
in01m08 FE_OCP_RBC3249_n_39697 ( .a(n_39697), .o(FE_OCP_RBN3249_n_39697) );
in01s04 FE_OCP_RBC3250_n_21312 ( .a(n_21312), .o(FE_OCP_RBN3250_n_21312) );
in01s01 FE_OCP_RBC3251_n_21312 ( .a(n_21312), .o(FE_OCP_RBN3251_n_21312) );
in01s02 FE_OCP_RBC3252_n_26276 ( .a(n_26276), .o(FE_OCP_RBN3252_n_26276) );
in01s01 FE_OCP_RBC3253_n_26276 ( .a(n_26276), .o(FE_OCP_RBN3253_n_26276) );
in01s02 FE_OCP_RBC3254_n_5478 ( .a(n_5478), .o(FE_OCP_RBN3254_n_5478) );
in01s01 FE_OCP_RBC3255_n_10454 ( .a(n_10454), .o(FE_OCP_RBN3255_n_10454) );
in01m01 FE_OCP_RBC3256_n_16113 ( .a(n_16113), .o(FE_OCP_RBN3256_n_16113) );
in01m02 FE_OCP_RBC3257_n_42998 ( .a(n_42998), .o(FE_OCP_RBN3257_n_42998) );
in01f02 FE_OCP_RBC3258_n_42998 ( .a(n_42998), .o(FE_OCP_RBN3258_n_42998) );
in01s01 FE_OCP_RBC3259_n_21360 ( .a(n_21360), .o(FE_OCP_RBN3259_n_21360) );
in01s01 FE_OCP_RBC3260_n_21360 ( .a(n_21360), .o(FE_OCP_RBN3260_n_21360) );
in01s02 FE_OCP_RBC3261_n_21360 ( .a(n_21360), .o(FE_OCP_RBN3261_n_21360) );
in01s01 FE_OCP_RBC3263_n_5531 ( .a(n_5531), .o(FE_OCP_RBN3263_n_5531) );
in01s01 FE_OCP_RBC3265_n_10852 ( .a(FE_OCP_RBN6087_n_10852), .o(FE_OCP_RBN3265_n_10852) );
in01s06 FE_OCP_RBC3266_n_26160 ( .a(n_26160), .o(FE_OCP_RBN3266_n_26160) );
in01s01 FE_OCP_RBC3269_n_26160 ( .a(FE_OCP_RBN4405_n_26160), .o(FE_OCP_RBN3269_n_26160) );
in01m02 FE_OCP_RBC3272_n_31239 ( .a(n_31239), .o(FE_OCP_RBN3272_n_31239) );
in01s01 FE_OCP_RBC3273_n_31239 ( .a(n_31239), .o(FE_OCP_RBN3273_n_31239) );
in01f02 FE_OCP_RBC3274_n_26464 ( .a(n_26464), .o(FE_OCP_RBN3274_n_26464) );
in01s01 FE_OCP_RBC3275_n_26464 ( .a(FE_OCPN6927_n_26464), .o(FE_OCP_RBN3275_n_26464) );
in01s01 FE_OCP_RBC3276_n_5284 ( .a(n_5284), .o(FE_OCP_RBN3276_n_5284) );
in01s02 FE_OCP_RBC3277_n_5284 ( .a(n_5284), .o(FE_OCP_RBN3277_n_5284) );
in01m02 FE_OCP_RBC3279_FE_RN_1496_0 ( .a(FE_RN_1496_0), .o(FE_OCP_RBN3279_FE_RN_1496_0) );
in01s01 FE_OCP_RBC3281_n_5614 ( .a(n_5614), .o(FE_OCP_RBN3281_n_5614) );
in01f02 FE_OCP_RBC3283_n_26316 ( .a(n_26316), .o(FE_OCP_RBN3283_n_26316) );
in01s04 FE_OCP_RBC3284_n_39674 ( .a(n_39674), .o(FE_OCP_RBN3284_n_39674) );
in01s01 FE_OCP_RBC3285_n_39674 ( .a(n_39674), .o(FE_OCP_RBN3285_n_39674) );
in01s01 FE_OCP_RBC3286_n_5656 ( .a(n_5656), .o(FE_OCP_RBN3286_n_5656) );
in01m02 FE_OCP_RBC3287_n_5656 ( .a(n_5656), .o(FE_OCP_RBN3287_n_5656) );
in01s04 FE_OCP_RBC3288_n_10915 ( .a(n_10915), .o(FE_OCP_RBN3288_n_10915) );
in01s01 FE_OCP_RBC3289_n_10915 ( .a(n_10915), .o(FE_OCP_RBN3289_n_10915) );
in01s06 FE_OCP_RBC3290_n_35539 ( .a(n_35539), .o(FE_OCP_RBN3290_n_35539) );
in01s02 FE_OCP_RBC3291_n_35539 ( .a(FE_OCP_RBN3290_n_35539), .o(FE_OCP_RBN3291_n_35539) );
in01s03 FE_OCP_RBC3292_n_35539 ( .a(FE_OCP_RBN3290_n_35539), .o(FE_OCP_RBN3292_n_35539) );
in01s01 FE_OCP_RBC3293_n_35539 ( .a(FE_OCP_RBN3290_n_35539), .o(FE_OCP_RBN3293_n_35539) );
in01s01 FE_OCP_RBC3294_n_35539 ( .a(FE_OCP_RBN3290_n_35539), .o(FE_OCP_RBN3294_n_35539) );
in01s02 FE_OCP_RBC3295_n_35539 ( .a(FE_OCP_RBN3291_n_35539), .o(FE_OCP_RBN3295_n_35539) );
in01s01 FE_OCP_RBC3297_n_35539 ( .a(FE_OCP_RBN3292_n_35539), .o(FE_OCP_RBN3297_n_35539) );
in01s01 FE_OCP_RBC3298_n_35539 ( .a(FE_OCP_RBN3293_n_35539), .o(FE_OCP_RBN3298_n_35539) );
in01s02 FE_OCP_RBC3299_n_35539 ( .a(FE_OCP_RBN3294_n_35539), .o(FE_OCP_RBN3299_n_35539) );
in01s02 FE_OCP_RBC3300_n_35539 ( .a(FE_OCP_RBN3297_n_35539), .o(FE_OCP_RBN3300_n_35539) );
in01s01 FE_OCP_RBC3301_n_35539 ( .a(FE_OCP_RBN3298_n_35539), .o(FE_OCP_RBN3301_n_35539) );
in01s01 FE_OCP_RBC3302_n_35539 ( .a(FE_OCP_RBN3301_n_35539), .o(FE_OCP_RBN3302_n_35539) );
in01s01 FE_OCP_RBC3303_n_35539 ( .a(FE_OCP_RBN3302_n_35539), .o(FE_OCP_RBN3303_n_35539) );
in01s10 FE_OCP_RBC3306_n_43022 ( .a(FE_OCP_RBN6109_n_43022), .o(FE_OCP_RBN3306_n_43022) );
in01s04 FE_OCP_RBC3307_n_43022 ( .a(FE_OCP_RBN6110_n_43022), .o(FE_OCP_RBN3307_n_43022) );
in01s01 FE_OCP_RBC3308_n_43022 ( .a(FE_OCP_RBN6110_n_43022), .o(FE_OCP_RBN3308_n_43022) );
in01s01 FE_OCP_RBC3309_n_43022 ( .a(FE_OCP_RBN3306_n_43022), .o(FE_OCP_RBN3309_n_43022) );
in01s10 FE_OCP_RBC3310_n_43022 ( .a(FE_OCP_RBN3306_n_43022), .o(FE_OCP_RBN3310_n_43022) );
in01s06 FE_OCP_RBC3311_n_43022 ( .a(FE_OCP_RBN3306_n_43022), .o(FE_OCP_RBN3311_n_43022) );
in01s03 FE_OCP_RBC3312_n_43022 ( .a(FE_OCP_RBN3307_n_43022), .o(FE_OCP_RBN3312_n_43022) );
in01s01 FE_OCP_RBC3313_n_43022 ( .a(FE_OCP_RBN3308_n_43022), .o(FE_OCP_RBN3313_n_43022) );
in01s01 FE_OCP_RBC3315_n_43022 ( .a(FE_OCP_RBN3313_n_43022), .o(FE_OCP_RBN3315_n_43022) );
in01s01 FE_OCP_RBC3318_n_5555 ( .a(FE_OCP_RBN6119_n_5555), .o(FE_OCP_RBN3318_n_5555) );
in01s01 FE_OCP_RBC3319_n_5555 ( .a(FE_OCP_RBN3318_n_5555), .o(FE_OCP_RBN3319_n_5555) );
in01f03 FE_OCP_RBC3320_n_42959 ( .a(n_42959), .o(FE_OCP_RBN3320_n_42959) );
in01s01 FE_OCP_RBC3321_n_42959 ( .a(n_42959), .o(FE_OCP_RBN3321_n_42959) );
in01s02 FE_OCP_RBC3322_n_5586 ( .a(n_5586), .o(FE_OCP_RBN3322_n_5586) );
in01s02 FE_OCP_RBC3324_n_5813 ( .a(n_5813), .o(FE_OCP_RBN3324_n_5813) );
in01s01 FE_OCP_RBC3325_n_5813 ( .a(FE_OCP_RBN3324_n_5813), .o(FE_OCP_RBN3325_n_5813) );
in01s01 FE_OCP_RBC3326_n_5813 ( .a(FE_OCP_RBN3325_n_5813), .o(FE_OCP_RBN3326_n_5813) );
in01m02 FE_OCP_RBC3327_n_21616 ( .a(n_21616), .o(FE_OCP_RBN3327_n_21616) );
in01m04 FE_OCP_RBC3328_n_21616 ( .a(FE_OCP_RBN3327_n_21616), .o(FE_OCP_RBN3328_n_21616) );
in01f02 FE_OCP_RBC3329_n_39685 ( .a(n_39685), .o(FE_OCP_RBN3329_n_39685) );
in01s01 FE_OCP_RBC3330_n_11087 ( .a(n_11087), .o(FE_OCP_RBN3330_n_11087) );
in01s02 FE_OCP_RBC3331_n_11087 ( .a(n_11087), .o(FE_OCP_RBN3331_n_11087) );
in01s10 FE_OCP_RBC3333_n_39942 ( .a(FE_OCP_RBN4431_n_39942), .o(FE_OCP_RBN3333_n_39942) );
in01s02 FE_OCP_RBC3336_n_39942 ( .a(FE_OCP_RBN3333_n_39942), .o(FE_OCP_RBN3336_n_39942) );
in01s01 FE_OCP_RBC3337_n_39942 ( .a(FE_OCP_RBN6853_n_39793), .o(FE_OCP_RBN3337_n_39942) );
in01s01 FE_OCP_RBC3339_n_39942 ( .a(FE_OCP_RBN4429_n_39942), .o(FE_OCP_RBN3339_n_39942) );
in01s01 FE_OCP_RBC3340_n_39942 ( .a(FE_OCP_RBN4429_n_39942), .o(FE_OCP_RBN3340_n_39942) );
in01s03 FE_OCP_RBC3341_n_39942 ( .a(FE_OCP_RBN3336_n_39942), .o(FE_OCP_RBN3341_n_39942) );
in01s02 FE_OCP_RBC3342_n_39942 ( .a(FE_OCP_RBN3336_n_39942), .o(FE_OCP_RBN3342_n_39942) );
in01m01 FE_OCP_RBC3343_n_39942 ( .a(FE_OCP_RBN4429_n_39942), .o(FE_OCP_RBN3343_n_39942) );
in01s02 FE_OCP_RBC3344_n_39942 ( .a(FE_OCP_RBN3343_n_39942), .o(FE_OCP_RBN3344_n_39942) );
in01s02 FE_OCP_RBC3345_n_39942 ( .a(FE_OCP_RBN3343_n_39942), .o(FE_OCP_RBN3345_n_39942) );
in01s02 FE_OCP_RBC3346_n_47269 ( .a(n_47269), .o(FE_OCP_RBN3346_n_47269) );
in01s02 FE_OCP_RBC3347_n_47269 ( .a(n_47269), .o(FE_OCP_RBN3347_n_47269) );
in01s01 FE_OCP_RBC3348_n_47269 ( .a(n_47269), .o(FE_OCP_RBN3348_n_47269) );
in01s01 FE_OCP_RBC3351_n_21812 ( .a(n_21812), .o(FE_OCP_RBN3351_n_21812) );
in01s02 FE_OCP_RBC3352_FE_OFN760_n_46337 ( .a(FE_OCP_RBN6163_n_46337), .o(FE_OCP_RBN3352_FE_OFN760_n_46337) );
in01f06 FE_OCP_RBC3355_FE_RN_1058_0 ( .a(FE_RN_1058_0), .o(FE_OCP_RBN3355_FE_RN_1058_0) );
in01m08 FE_OCP_RBC3356_FE_RN_1058_0 ( .a(FE_OCP_RBN3355_FE_RN_1058_0), .o(FE_OCP_RBN3356_FE_RN_1058_0) );
in01m04 FE_OCP_RBC3357_n_6013 ( .a(n_6013), .o(FE_OCP_RBN3357_n_6013) );
in01s03 FE_OCP_RBC3358_n_11275 ( .a(n_11275), .o(FE_OCP_RBN3358_n_11275) );
in01m02 FE_OCP_RBC3359_n_11275 ( .a(n_11275), .o(FE_OCP_RBN3359_n_11275) );
in01f04 FE_OCP_RBC3360_n_16596 ( .a(n_16596), .o(FE_OCP_RBN3360_n_16596) );
in01f02 FE_OCP_RBC3361_n_21847 ( .a(n_21847), .o(FE_OCP_RBN3361_n_21847) );
in01s01 FE_OCP_RBC3362_n_21951 ( .a(n_21951), .o(FE_OCP_RBN3362_n_21951) );
in01m04 FE_OCP_RBC3365_n_31520 ( .a(FE_OCP_RBN6139_n_31520), .o(FE_OCP_RBN3365_n_31520) );
in01m02 FE_OCP_RBC3368_n_31520 ( .a(FE_OCP_RBN3365_n_31520), .o(FE_OCP_RBN3368_n_31520) );
in01s01 FE_OCP_RBC3369_n_31520 ( .a(FE_OCP_RBN3365_n_31520), .o(FE_OCP_RBN3369_n_31520) );
in01s01 FE_OCP_RBC3370_n_31520 ( .a(FE_OCP_RBN3365_n_31520), .o(FE_OCP_RBN3370_n_31520) );
in01s01 FE_OCP_RBC3371_n_36490 ( .a(n_36490), .o(FE_OCP_RBN3371_n_36490) );
in01s06 FE_OCP_RBC3372_n_43046 ( .a(n_43046), .o(FE_OCP_RBN3372_n_43046) );
in01s06 FE_OCP_RBC3373_n_43046 ( .a(n_43046), .o(FE_OCP_RBN3373_n_43046) );
in01s02 FE_OCP_RBC3374_n_43046 ( .a(n_43046), .o(FE_OCP_RBN3374_n_43046) );
in01s01 FE_OCP_RBC3375_n_43046 ( .a(n_43046), .o(FE_OCP_RBN3375_n_43046) );
in01s06 FE_OCP_RBC3377_n_44342 ( .a(FE_OCP_RBN6162_FE_RN_1136_0), .o(FE_OCP_RBN3377_n_44342) );
in01m02 FE_OCP_RBC3380_n_6034 ( .a(n_6034), .o(FE_OCP_RBN3380_n_6034) );
in01s04 FE_OCP_RBC3381_n_36547 ( .a(n_36547), .o(FE_OCP_RBN3381_n_36547) );
in01s04 FE_OCP_RBC3382_n_11405 ( .a(n_11405), .o(FE_OCP_RBN3382_n_11405) );
in01s01 FE_OCP_RBC3383_n_11405 ( .a(n_11405), .o(FE_OCP_RBN3383_n_11405) );
in01m08 FE_OCP_RBC3384_n_11439 ( .a(n_11439), .o(FE_OCP_RBN3384_n_11439) );
in01s02 FE_OCP_RBC3386_n_11439 ( .a(FE_OCP_RBN3384_n_11439), .o(FE_OCP_RBN3386_n_11439) );
in01s01 FE_OCP_RBC3387_n_17130 ( .a(n_17130), .o(FE_OCP_RBN3387_n_17130) );
in01m10 FE_OCP_RBC3388_n_31819 ( .a(n_31819), .o(FE_OCP_RBN3388_n_31819) );
in01s04 FE_OCP_RBC3390_n_31819 ( .a(n_31819), .o(FE_OCP_RBN3390_n_31819) );
in01s06 FE_OCP_RBC3391_n_31819 ( .a(n_31819), .o(FE_OCP_RBN3391_n_31819) );
in01s01 FE_OCP_RBC3394_FE_RN_1094_0 ( .a(FE_RN_1094_0), .o(FE_OCP_RBN3394_FE_RN_1094_0) );
in01f04 FE_OCP_RBC3395_FE_RN_1094_0 ( .a(FE_RN_1094_0), .o(FE_OCP_RBN3395_FE_RN_1094_0) );
in01s02 FE_OCP_RBC3396_n_11486 ( .a(n_11486), .o(FE_OCP_RBN3396_n_11486) );
in01s06 FE_OCP_RBC3398_n_11486 ( .a(n_11486), .o(FE_OCP_RBN3398_n_11486) );
in01s01 FE_OCP_RBC3401_n_17233 ( .a(n_17233), .o(FE_OCP_RBN3401_n_17233) );
in01s01 FE_OCP_RBC3402_n_43775 ( .a(n_43775), .o(FE_OCP_RBN3402_n_43775) );
in01m04 FE_OCP_RBC3403_n_6205 ( .a(n_6205), .o(FE_OCP_RBN3403_n_6205) );
in01m06 FE_OCP_RBC3404_n_6205 ( .a(FE_OCP_RBN3403_n_6205), .o(FE_OCP_RBN3404_n_6205) );
in01s01 FE_OCP_RBC3405_n_6205 ( .a(FE_OCP_RBN3404_n_6205), .o(FE_OCP_RBN3405_n_6205) );
in01f04 FE_OCP_RBC3406_n_32143 ( .a(n_32143), .o(FE_OCP_RBN3406_n_32143) );
in01s01 FE_OCP_RBC3407_n_11560 ( .a(n_11560), .o(FE_OCP_RBN3407_n_11560) );
in01s01 FE_OCP_RBC3408_n_22604 ( .a(n_22604), .o(FE_OCP_RBN3408_n_22604) );
in01s01 FE_OCP_RBC3409_n_32072 ( .a(n_32072), .o(FE_OCP_RBN3409_n_32072) );
in01s02 FE_OCP_RBC3410_n_36706 ( .a(n_36706), .o(FE_OCP_RBN3410_n_36706) );
in01s01 FE_OCP_RBC3411_n_43811 ( .a(n_43811), .o(FE_OCP_RBN3411_n_43811) );
in01s01 FE_OCP_RBC3412_n_43829 ( .a(n_43829), .o(FE_OCP_RBN3412_n_43829) );
in01s01 FE_OCP_RBC3413_FE_OCPN891_n_31944 ( .a(FE_OCP_RBN6879_n_31819), .o(FE_OCP_RBN3413_FE_OCPN891_n_31944) );
in01s01 FE_OCP_RBC3414_FE_OCPN891_n_31944 ( .a(FE_OCP_RBN6879_n_31819), .o(FE_OCP_RBN3414_FE_OCPN891_n_31944) );
in01s02 FE_OCP_RBC3416_n_22564 ( .a(n_22564), .o(FE_OCP_RBN3416_n_22564) );
in01f03 FE_OCP_RBC3417_n_22564 ( .a(n_22564), .o(FE_OCP_RBN3417_n_22564) );
in01m02 FE_OCP_RBC3418_n_27590 ( .a(n_27590), .o(FE_OCP_RBN3418_n_27590) );
in01s02 FE_OCP_RBC3419_n_32130 ( .a(n_32130), .o(FE_OCP_RBN3419_n_32130) );
in01s01 FE_OCP_RBC3420_n_40300 ( .a(n_40300), .o(FE_OCP_RBN3420_n_40300) );
in01f02 FE_OCP_RBC3421_n_32254 ( .a(n_32254), .o(FE_OCP_RBN3421_n_32254) );
in01s02 FE_OCP_RBC3424_FE_RN_1622_0 ( .a(FE_RN_1622_0), .o(FE_OCP_RBN3424_FE_RN_1622_0) );
in01s01 FE_OCP_RBC3425_n_11754 ( .a(n_11754), .o(FE_OCP_RBN3425_n_11754) );
in01s02 FE_OCP_RBC3426_n_11810 ( .a(n_11810), .o(FE_OCP_RBN3426_n_11810) );
in01s01 FE_OCP_RBC3427_n_17510 ( .a(n_17510), .o(FE_OCP_RBN3427_n_17510) );
in01s01 FE_OCP_RBC3428_n_32180 ( .a(n_32180), .o(FE_OCP_RBN3428_n_32180) );
in01s01 FE_OCP_RBC3429_n_36664 ( .a(n_36664), .o(FE_OCP_RBN3429_n_36664) );
in01f02 FE_OCP_RBC3430_n_40563 ( .a(n_40563), .o(FE_OCP_RBN3430_n_40563) );
in01f02 FE_OCP_RBC3431_n_43880 ( .a(n_43880), .o(FE_OCP_RBN3431_n_43880) );
in01m02 FE_OCP_RBC3432_n_32239 ( .a(n_32239), .o(FE_OCP_RBN3432_n_32239) );
in01s01 FE_OCP_RBC3434_n_6379 ( .a(n_6379), .o(FE_OCP_RBN3434_n_6379) );
in01s01 FE_OCP_RBC3435_n_6379 ( .a(n_6379), .o(FE_OCP_RBN3435_n_6379) );
in01s01 FE_OCP_RBC3436_n_6485 ( .a(n_6485), .o(FE_OCP_RBN3436_n_6485) );
in01m02 FE_OCP_RBC3437_n_11980 ( .a(n_11980), .o(FE_OCP_RBN3437_n_11980) );
in01s01 FE_OCP_RBC3438_n_32232 ( .a(n_32232), .o(FE_OCP_RBN3438_n_32232) );
in01m02 FE_OCP_RBC3441_n_32266 ( .a(n_32266), .o(FE_OCP_RBN3441_n_32266) );
in01s01 FE_OCP_RBC3442_n_32266 ( .a(n_32266), .o(FE_OCP_RBN3442_n_32266) );
in01s01 FE_OCP_RBC3443_n_6471 ( .a(n_6471), .o(FE_OCP_RBN3443_n_6471) );
in01s04 FE_OCP_RBC3444_n_6513 ( .a(n_6513), .o(FE_OCP_RBN3444_n_6513) );
in01s01 FE_OCP_RBC3445_n_6513 ( .a(n_6513), .o(FE_OCP_RBN3445_n_6513) );
in01s02 FE_OCP_RBC3446_n_6513 ( .a(n_6513), .o(FE_OCP_RBN3446_n_6513) );
in01s02 FE_OCP_RBC3449_n_43777 ( .a(n_43777), .o(FE_OCP_RBN3449_n_43777) );
in01m02 FE_OCP_RBC3450_n_17697 ( .a(n_17697), .o(FE_OCP_RBN3450_n_17697) );
in01m02 FE_OCP_RBC3451_n_22710 ( .a(n_22710), .o(FE_OCP_RBN3451_n_22710) );
in01m04 FE_OCP_RBC3453_n_27632 ( .a(n_27632), .o(FE_OCP_RBN3453_n_27632) );
in01s01 FE_OCP_RBC3454_n_6557 ( .a(n_6557), .o(FE_OCP_RBN3454_n_6557) );
in01s01 FE_OCP_RBC3455_n_6557 ( .a(n_6557), .o(FE_OCP_RBN3455_n_6557) );
in01m02 FE_OCP_RBC3456_n_22709 ( .a(n_22709), .o(FE_OCP_RBN3456_n_22709) );
in01s02 FE_OCP_RBC3458_n_12196 ( .a(n_12196), .o(FE_OCP_RBN3458_n_12196) );
in01s01 FE_OCP_RBC3463_n_32316 ( .a(n_32316), .o(FE_OCP_RBN3463_n_32316) );
in01f02 FE_OCP_RBC3464_n_43836 ( .a(n_43836), .o(FE_OCP_RBN3464_n_43836) );
in01s06 FE_OCP_RBC3702_n_11788 ( .a(n_11788), .o(FE_OCP_RBN3702_n_11788) );
in01s01 FE_OCP_RBC3703_n_12904 ( .a(n_12904), .o(FE_OCP_RBN3703_n_12904) );
in01s01 FE_OCP_RBC3706_n_18716 ( .a(n_18716), .o(FE_OCP_RBN3706_n_18716) );
in01s01 FE_OCP_RBC3707_n_18716 ( .a(FE_OCP_RBN3706_n_18716), .o(FE_OCP_RBN3707_n_18716) );
in01f01 FE_OCP_RBC3709_n_29055 ( .a(n_29055), .o(FE_OCP_RBN3709_n_29055) );
in01s01 FE_OCP_RBC3710_n_29055 ( .a(n_29055), .o(FE_OCP_RBN3710_n_29055) );
in01s02 FE_OCP_RBC3711_n_19116 ( .a(n_19116), .o(FE_OCP_RBN3711_n_19116) );
in01f02 FE_OCP_RBC3713_n_19241 ( .a(n_19241), .o(FE_OCP_RBN3713_n_19241) );
in01s01 FE_OCP_RBC3714_n_19241 ( .a(FE_OCP_RBN3713_n_19241), .o(FE_OCP_RBN3714_n_19241) );
in01s01 FE_OCP_RBC3715_n_19241 ( .a(FE_OCP_RBN3714_n_19241), .o(FE_OCP_RBN3715_n_19241) );
in01s01 FE_OCP_RBC3716_n_19241 ( .a(FE_OCP_RBN3714_n_19241), .o(FE_OCP_RBN3716_n_19241) );
in01s02 FE_OCP_RBC3717_n_19535 ( .a(n_19535), .o(FE_OCP_RBN3717_n_19535) );
in01f02 FE_OCP_RBC3718_n_20621 ( .a(n_20621), .o(FE_OCP_RBN3718_n_20621) );
in01s01 FE_OCP_RBC3719_n_20621 ( .a(n_20621), .o(FE_OCP_RBN3719_n_20621) );
in01s02 FE_OCP_RBC3720_n_20621 ( .a(FE_OCP_RBN3719_n_20621), .o(FE_OCP_RBN3720_n_20621) );
in01s02 FE_OCP_RBC3721_n_20621 ( .a(FE_OCP_RBN3720_n_20621), .o(FE_OCP_RBN3721_n_20621) );
in01f02 FE_OCP_RBC3722_n_30776 ( .a(n_30776), .o(FE_OCP_RBN3722_n_30776) );
in01m02 FE_OCP_RBC3723_n_21442 ( .a(n_21442), .o(FE_OCP_RBN3723_n_21442) );
in01s01 FE_OCP_RBC3762_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN3762_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s03 FE_OCP_RBC3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s06 FE_OCP_RBC3815_n_45209 ( .a(n_45209), .o(FE_OCP_RBN3815_n_45209) );
in01s40 FE_OCP_RBC3818_n_45622 ( .a(n_45622), .o(FE_OCP_RBN3818_n_45622) );
in01f20 FE_OCP_RBC3844_delay_sub_ln23_unr13_stage5_stallmux_q_1_ ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(FE_OCP_RBN3844_delay_sub_ln23_unr13_stage5_stallmux_q_1_) );
in01f20 FE_OCP_RBC3845_delay_sub_ln23_unr13_stage5_stallmux_q_1_ ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(FE_OCP_RBN3845_delay_sub_ln23_unr13_stage5_stallmux_q_1_) );
in01s80 FE_OCP_RBC3871_n_44061 ( .a(FE_OCP_RBN6467_n_44061), .o(FE_OCP_RBN3871_n_44061) );
in01s01 FE_OCP_RBC3879_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN3879_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s01 FE_OCP_RBC3881_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN3881_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s40 FE_OCP_RBC3938_n_46254 ( .a(FE_OCP_RBN3939_n_46254), .o(FE_OCP_RBN3938_n_46254) );
in01s40 FE_OCP_RBC3939_n_46254 ( .a(n_46254), .o(FE_OCP_RBN3939_n_46254) );
in01s10 FE_OCP_RBC3963_delay_sub_ln21_unr24_stage9_stallmux_q_8_ ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(FE_OCP_RBN3963_delay_sub_ln21_unr24_stage9_stallmux_q_8_) );
in01s80 FE_OCP_RBC3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_ ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_) );
in01s20 FE_OCP_RBC3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_ ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_) );
in01s80 FE_OCP_RBC3966_n_44061 ( .a(FE_OCP_RBN3871_n_44061), .o(FE_OCP_RBN3966_n_44061) );
in01s20 FE_OCP_RBC3967_n_44061 ( .a(FE_OCP_RBN3871_n_44061), .o(FE_OCP_RBN3967_n_44061) );
in01s80 FE_OCP_RBC3968_n_44061 ( .a(FE_OCP_RBN3966_n_44061), .o(FE_OCP_RBN3968_n_44061) );
in01s10 FE_OCP_RBC3975_n_45224 ( .a(FE_OCP_RBN6523_n_45224), .o(FE_OCP_RBN3975_n_45224) );
in01s01 FE_OCP_RBC3976_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN6513_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN3976_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s40 FE_OCP_RBC3979_n_22972 ( .a(n_22972), .o(FE_OCP_RBN3979_n_22972) );
in01s20 FE_OCP_RBC3980_n_32436 ( .a(n_32436), .o(FE_OCP_RBN3980_n_32436) );
in01s06 FE_OCP_RBC3982_n_27911 ( .a(n_27911), .o(FE_OCP_RBN3982_n_27911) );
in01s10 FE_OCP_RBC3984_n_32791 ( .a(FE_OCP_RBN6532_n_32791), .o(FE_OCP_RBN3984_n_32791) );
in01s01 FE_OCP_RBC3985_FE_RN_158_0 ( .a(FE_RN_158_0), .o(FE_OCP_RBN3985_FE_RN_158_0) );
in01s10 FE_OCP_RBC3986_FE_RN_158_0 ( .a(FE_RN_158_0), .o(FE_OCP_RBN3986_FE_RN_158_0) );
in01s06 FE_OCP_RBC3988_n_32772 ( .a(n_32772), .o(FE_OCP_RBN3988_n_32772) );
in01s06 FE_OCP_RBC3989_n_32772 ( .a(n_32772), .o(FE_OCP_RBN3989_n_32772) );
in01s10 FE_OCP_RBC3990_n_32772 ( .a(n_32772), .o(FE_OCP_RBN3990_n_32772) );
in01s06 FE_OCP_RBC3991_FE_RN_1579_0 ( .a(FE_RN_1579_0), .o(FE_OCP_RBN3991_FE_RN_1579_0) );
in01s01 FE_OCP_RBC3997_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN6512_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN3997_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01m03 FE_OCP_RBC3998_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN6512_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN3998_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01s04 FE_OCP_RBC4002_n_33015 ( .a(n_33015), .o(FE_OCP_RBN4002_n_33015) );
in01s04 FE_OCP_RBC4003_n_33015 ( .a(n_33015), .o(FE_OCP_RBN4003_n_33015) );
in01s06 FE_OCP_RBC4004_n_33015 ( .a(n_33015), .o(FE_OCP_RBN4004_n_33015) );
in01s08 FE_OCP_RBC4005_n_33015 ( .a(FE_OCP_RBN4004_n_33015), .o(FE_OCP_RBN4005_n_33015) );
in01s01 FE_OCP_RBC4006_n_32860 ( .a(FE_OCP_RBN2452_n_32860), .o(FE_OCP_RBN4006_n_32860) );
in01s02 FE_OCP_RBC4007_n_32860 ( .a(FE_OCP_RBN2452_n_32860), .o(FE_OCP_RBN4007_n_32860) );
in01s01 FE_OCP_RBC4008_n_32860 ( .a(FE_OCP_RBN2452_n_32860), .o(FE_OCP_RBN4008_n_32860) );
in01s02 FE_OCP_RBC4009_n_32860 ( .a(FE_OCP_RBN4006_n_32860), .o(FE_OCP_RBN4009_n_32860) );
in01s01 FE_OCP_RBC4011_n_1864 ( .a(n_1864), .o(FE_OCP_RBN4011_n_1864) );
in01s04 FE_OCP_RBC4012_n_1864 ( .a(n_1864), .o(FE_OCP_RBN4012_n_1864) );
in01s06 FE_OCP_RBC4013_n_33034 ( .a(FE_OCP_RBN2467_n_33034), .o(FE_OCP_RBN4013_n_33034) );
in01s08 FE_OCP_RBC4014_n_33034 ( .a(FE_OCP_RBN2467_n_33034), .o(FE_OCP_RBN4014_n_33034) );
in01s04 FE_OCP_RBC4015_n_33034 ( .a(FE_OCP_RBN2467_n_33034), .o(FE_OCP_RBN4015_n_33034) );
in01s01 FE_OCP_RBC4016_n_33034 ( .a(FE_OCP_RBN2467_n_33034), .o(FE_OCP_RBN4016_n_33034) );
in01m04 FE_OCP_RBC4017_n_33034 ( .a(FE_OCP_RBN4014_n_33034), .o(FE_OCP_RBN4017_n_33034) );
in01m01 FE_OCP_RBC4018_n_33034 ( .a(FE_OCP_RBN4014_n_33034), .o(FE_OCP_RBN4018_n_33034) );
in01s10 FE_OCP_RBC4019_n_33034 ( .a(FE_OCP_RBN4014_n_33034), .o(FE_OCP_RBN4019_n_33034) );
in01s01 FE_OCP_RBC4020_n_33034 ( .a(FE_OCP_RBN4016_n_33034), .o(FE_OCP_RBN4020_n_33034) );
in01s01 FE_OCP_RBC4021_n_33034 ( .a(FE_OCP_RBN4020_n_33034), .o(FE_OCP_RBN4021_n_33034) );
in01s01 FE_OCP_RBC4022_n_33034 ( .a(FE_OCP_RBN4020_n_33034), .o(FE_OCP_RBN4022_n_33034) );
in01s02 FE_OCP_RBC4023_n_37577 ( .a(n_37577), .o(FE_OCP_RBN4023_n_37577) );
in01s01 FE_OCP_RBC4024_n_37577 ( .a(FE_OCP_RBN4023_n_37577), .o(FE_OCP_RBN4024_n_37577) );
in01s01 FE_OCP_RBC4025_n_37577 ( .a(FE_OCP_RBN4024_n_37577), .o(FE_OCP_RBN4025_n_37577) );
in01s01 FE_OCP_RBC4026_n_37577 ( .a(FE_OCP_RBN4025_n_37577), .o(FE_OCP_RBN4026_n_37577) );
in01s01 FE_OCP_RBC4027_n_37577 ( .a(FE_OCP_RBN4026_n_37577), .o(FE_OCP_RBN4027_n_37577) );
in01m10 FE_OCP_RBC4028_n_28458 ( .a(n_28458), .o(FE_OCP_RBN4028_n_28458) );
in01s01 FE_OCP_RBC4030_n_28458 ( .a(FE_OCP_RBN4028_n_28458), .o(FE_OCP_RBN4030_n_28458) );
in01s01 FE_OCP_RBC4031_n_28458 ( .a(FE_OCP_RBN6552_n_28458), .o(FE_OCP_RBN4031_n_28458) );
in01f06 FE_OCP_RBC4032_n_37690 ( .a(n_37690), .o(FE_OCP_RBN4032_n_37690) );
in01m02 FE_OCP_RBC4033_n_37690 ( .a(n_37690), .o(FE_OCP_RBN4033_n_37690) );
in01m02 FE_OCP_RBC4034_n_37690 ( .a(n_37690), .o(FE_OCP_RBN4034_n_37690) );
in01s02 FE_OCP_RBC4035_n_28651 ( .a(n_28651), .o(FE_OCP_RBN4035_n_28651) );
in01s04 FE_OCP_RBC4036_n_28651 ( .a(n_28651), .o(FE_OCP_RBN4036_n_28651) );
in01s02 FE_OCP_RBC4037_n_12904 ( .a(FE_OCP_RBN3703_n_12904), .o(FE_OCP_RBN4037_n_12904) );
in01s02 FE_OCP_RBC4038_n_2059 ( .a(n_2059), .o(FE_OCP_RBN4038_n_2059) );
in01s02 FE_OCP_RBC4040_n_37707 ( .a(n_37707), .o(FE_OCP_RBN4040_n_37707) );
in01s01 FE_OCP_RBC4041_n_37707 ( .a(FE_OCP_RBN4040_n_37707), .o(FE_OCP_RBN4041_n_37707) );
in01s01 FE_OCP_RBC4042_n_37707 ( .a(FE_OCP_RBN4041_n_37707), .o(FE_OCP_RBN4042_n_37707) );
in01f06 FE_OCP_RBC4043_n_41258 ( .a(n_41258), .o(FE_OCP_RBN4043_n_41258) );
in01m06 FE_OCP_RBC4044_n_41298 ( .a(n_41298), .o(FE_OCP_RBN4044_n_41298) );
in01f02 FE_OCP_RBC4045_n_41298 ( .a(n_41298), .o(FE_OCP_RBN4045_n_41298) );
in01s01 FE_OCP_RBC4046_n_41298 ( .a(n_41298), .o(FE_OCP_RBN4046_n_41298) );
in01s10 FE_OCP_RBC4047_n_12721 ( .a(FE_OCP_RBN5578_n_12753), .o(FE_OCP_RBN4047_n_12721) );
in01s20 FE_OCP_RBC4048_n_12721 ( .a(FE_OCP_RBN4047_n_12721), .o(FE_OCP_RBN4048_n_12721) );
in01s02 FE_OCP_RBC4049_n_33491 ( .a(n_33491), .o(FE_OCP_RBN4049_n_33491) );
in01s01 FE_OCP_RBC4052_n_2086 ( .a(FE_OCP_RBN2526_n_2086), .o(FE_OCP_RBN4052_n_2086) );
in01s02 FE_OCP_RBC4053_n_2086 ( .a(FE_OCP_RBN2526_n_2086), .o(FE_OCP_RBN4053_n_2086) );
in01s01 FE_OCP_RBC4054_n_41325 ( .a(n_41325), .o(FE_OCP_RBN4054_n_41325) );
in01m02 FE_OCP_RBC4055_n_41325 ( .a(n_41325), .o(FE_OCP_RBN4055_n_41325) );
in01s01 FE_OCP_RBC4058_n_44875 ( .a(FE_OCP_RBN5600_n_44875), .o(FE_OCP_RBN4058_n_44875) );
in01s01 FE_OCP_RBC4059_n_44875 ( .a(FE_OCP_RBN6575_n_44875), .o(FE_OCP_RBN4059_n_44875) );
in01s01 FE_OCP_RBC4060_n_44875 ( .a(FE_OCP_RBN6571_n_44875), .o(FE_OCP_RBN4060_n_44875) );
in01s02 FE_OCP_RBC4061_n_44030 ( .a(n_44030), .o(FE_OCP_RBN4061_n_44030) );
in01s01 FE_OCP_RBC4062_n_44030 ( .a(n_44030), .o(FE_OCP_RBN4062_n_44030) );
in01s01 FE_OCP_RBC4063_n_7558 ( .a(n_7558), .o(FE_OCP_RBN4063_n_7558) );
in01s01 FE_OCP_RBC4064_n_7558 ( .a(n_7558), .o(FE_OCP_RBN4064_n_7558) );
in01s01 FE_OCP_RBC4065_n_7558 ( .a(n_7558), .o(FE_OCP_RBN4065_n_7558) );
in01s02 FE_OCP_RBC4066_n_7558 ( .a(FE_OCP_RBN4063_n_7558), .o(FE_OCP_RBN4066_n_7558) );
in01f04 FE_OCP_RBC4067_n_18829 ( .a(n_18829), .o(FE_OCP_RBN4067_n_18829) );
in01m02 FE_OCP_RBC4068_n_18829 ( .a(n_18829), .o(FE_OCP_RBN4068_n_18829) );
in01s01 FE_OCP_RBC4070_n_29292 ( .a(n_29292), .o(FE_OCP_RBN4070_n_29292) );
in01s06 FE_OCP_RBC4071_n_2289 ( .a(n_2289), .o(FE_OCP_RBN4071_n_2289) );
in01s10 FE_OCP_RBC4072_n_2289 ( .a(n_2289), .o(FE_OCP_RBN4072_n_2289) );
in01s10 FE_OCP_RBC4073_n_2289 ( .a(FE_OCP_RBN4072_n_2289), .o(FE_OCP_RBN4073_n_2289) );
in01s01 FE_OCP_RBC4074_n_2289 ( .a(FE_OCP_RBN6610_n_2289), .o(FE_OCP_RBN4074_n_2289) );
in01s08 FE_OCP_RBC4075_n_7708 ( .a(n_7708), .o(FE_OCP_RBN4075_n_7708) );
in01s01 FE_OCP_RBC4080_n_7708 ( .a(FE_OCP_RBN6596_n_7708), .o(FE_OCP_RBN4080_n_7708) );
in01s01 FE_OCP_RBC4081_n_18899 ( .a(n_18899), .o(FE_OCP_RBN4081_n_18899) );
in01f02 FE_OCP_RBC4082_n_18899 ( .a(n_18899), .o(FE_OCP_RBN4082_n_18899) );
in01f01 FE_OCP_RBC4083_n_13453 ( .a(n_13453), .o(FE_OCP_RBN4083_n_13453) );
in01s01 FE_OCP_RBC4084_n_13453 ( .a(FE_OCP_RBN4083_n_13453), .o(FE_OCP_RBN4084_n_13453) );
in01s10 FE_OCP_RBC4087_n_12880 ( .a(FE_OCP_RBN2540_n_12880), .o(FE_OCP_RBN4087_n_12880) );
in01s01 FE_OCP_RBC4088_n_12880 ( .a(FE_OCP_RBN4087_n_12880), .o(FE_OCP_RBN4088_n_12880) );
in01s03 FE_OCP_RBC4089_n_12880 ( .a(FE_OCP_RBN4087_n_12880), .o(FE_OCP_RBN4089_n_12880) );
in01s01 FE_OCP_RBC4090_n_12880 ( .a(FE_OCP_RBN4087_n_12880), .o(FE_OCP_RBN4090_n_12880) );
in01s01 FE_OCP_RBC4091_n_12880 ( .a(FE_OCP_RBN4088_n_12880), .o(FE_OCP_RBN4091_n_12880) );
in01s03 FE_OCP_RBC4092_n_12880 ( .a(FE_OCP_RBN4089_n_12880), .o(FE_OCP_RBN4092_n_12880) );
in01s01 FE_OCP_RBC4093_n_12880 ( .a(FE_OCP_RBN4090_n_12880), .o(FE_OCP_RBN4093_n_12880) );
in01s01 FE_OCP_RBC4094_n_12880 ( .a(FE_OCP_RBN4090_n_12880), .o(FE_OCP_RBN4094_n_12880) );
in01s01 FE_OCP_RBC4095_n_12880 ( .a(FE_OCP_RBN4090_n_12880), .o(FE_OCP_RBN4095_n_12880) );
in01s01 FE_OCP_RBC4096_n_12880 ( .a(FE_OCP_RBN4091_n_12880), .o(FE_OCP_RBN4096_n_12880) );
in01s03 FE_OCP_RBC4097_n_12880 ( .a(FE_OCP_RBN4092_n_12880), .o(FE_OCP_RBN4097_n_12880) );
in01s01 FE_OCP_RBC4098_n_12880 ( .a(FE_OCP_RBN4097_n_12880), .o(FE_OCP_RBN4098_n_12880) );
in01s03 FE_OCP_RBC4099_n_12880 ( .a(FE_OCP_RBN4097_n_12880), .o(FE_OCP_RBN4099_n_12880) );
in01m01 FE_OCP_RBC4100_n_12880 ( .a(FE_OCP_RBN4098_n_12880), .o(FE_OCP_RBN4100_n_12880) );
in01s03 FE_OCP_RBC4101_n_12880 ( .a(FE_OCP_RBN4099_n_12880), .o(FE_OCP_RBN4101_n_12880) );
in01s03 FE_OCP_RBC4102_n_12880 ( .a(FE_OCP_RBN4101_n_12880), .o(FE_OCP_RBN4102_n_12880) );
in01s01 FE_OCP_RBC4103_n_12880 ( .a(FE_OCP_RBN4101_n_12880), .o(FE_OCP_RBN4103_n_12880) );
in01s01 FE_OCP_RBC4104_n_12880 ( .a(FE_OCP_RBN4101_n_12880), .o(FE_OCP_RBN4104_n_12880) );
in01s01 FE_OCP_RBC4105_n_12880 ( .a(FE_OCP_RBN4102_n_12880), .o(FE_OCP_RBN4105_n_12880) );
in01s01 FE_OCP_RBC4106_n_12880 ( .a(FE_OCP_RBN4105_n_12880), .o(FE_OCP_RBN4106_n_12880) );
in01s01 FE_OCP_RBC4107_n_12880 ( .a(FE_OCP_RBN4106_n_12880), .o(FE_OCP_RBN4107_n_12880) );
in01s01 FE_OCP_RBC4108_n_12880 ( .a(FE_OCP_RBN4107_n_12880), .o(FE_OCP_RBN4108_n_12880) );
in01s01 FE_OCP_RBC4109_n_12880 ( .a(FE_OCP_RBN4107_n_12880), .o(FE_OCP_RBN4109_n_12880) );
in01s01 FE_OCP_RBC4110_n_12880 ( .a(FE_OCP_RBN2541_n_12880), .o(FE_OCP_RBN4110_n_12880) );
in01s01 FE_OCP_RBC4111_n_12880 ( .a(FE_OCP_RBN4110_n_12880), .o(FE_OCP_RBN4111_n_12880) );
in01s06 FE_OCP_RBC4112_n_12880 ( .a(FE_OCP_RBN4111_n_12880), .o(FE_OCP_RBN4112_n_12880) );
in01m02 FE_OCP_RBC4113_n_33533 ( .a(n_33533), .o(FE_OCP_RBN4113_n_33533) );
in01m02 FE_OCP_RBC4114_n_33533 ( .a(n_33533), .o(FE_OCP_RBN4114_n_33533) );
in01s08 FE_OCP_RBC4115_n_41381 ( .a(n_41381), .o(FE_OCP_RBN4115_n_41381) );
in01s02 FE_OCP_RBC4118_n_45487 ( .a(n_45487), .o(FE_OCP_RBN4118_n_45487) );
in01s01 FE_OCP_RBC4120_n_13483 ( .a(n_13483), .o(FE_OCP_RBN4120_n_13483) );
in01m02 FE_OCP_RBC4130_n_24077 ( .a(n_24077), .o(FE_OCP_RBN4130_n_24077) );
in01s02 FE_OCP_RBC4131_n_24077 ( .a(n_24077), .o(FE_OCP_RBN4131_n_24077) );
in01s01 FE_OCP_RBC4132_n_38028 ( .a(n_38028), .o(FE_OCP_RBN4132_n_38028) );
in01s02 FE_OCP_RBC4133_n_38028 ( .a(FE_OCP_RBN4132_n_38028), .o(FE_OCP_RBN4133_n_38028) );
in01s01 FE_OCP_RBC4135_n_7743 ( .a(FE_OCP_RBN6600_n_7708), .o(FE_OCP_RBN4135_n_7743) );
in01s01 FE_OCP_RBC4136_n_7743 ( .a(FE_OCP_RBN6600_n_7708), .o(FE_OCP_RBN4136_n_7743) );
in01s01 FE_OCP_RBC4137_n_7743 ( .a(FE_OCP_RBN6600_n_7708), .o(FE_OCP_RBN4137_n_7743) );
in01s06 FE_OCP_RBC4138_n_7743 ( .a(FE_OCP_RBN5634_n_7708), .o(FE_OCP_RBN4138_n_7743) );
in01s02 FE_OCP_RBC4139_n_7743 ( .a(FE_OCP_RBN5636_n_7708), .o(FE_OCP_RBN4139_n_7743) );
in01s01 FE_OCP_RBC4140_n_7743 ( .a(FE_OCP_RBN5634_n_7708), .o(FE_OCP_RBN4140_n_7743) );
in01s02 FE_OCP_RBC4141_n_7743 ( .a(FE_OCP_RBN4135_n_7743), .o(FE_OCP_RBN4141_n_7743) );
in01s06 FE_OCP_RBC4142_n_7743 ( .a(FE_OCP_RBN4138_n_7743), .o(FE_OCP_RBN4142_n_7743) );
in01s01 FE_OCP_RBC4143_n_7743 ( .a(FE_OCP_RBN4140_n_7743), .o(FE_OCP_RBN4143_n_7743) );
in01s01 FE_OCP_RBC4144_n_7743 ( .a(FE_OCP_RBN4140_n_7743), .o(FE_OCP_RBN4144_n_7743) );
in01s01 FE_OCP_RBC4145_n_7743 ( .a(FE_OCP_RBN4141_n_7743), .o(FE_OCP_RBN4145_n_7743) );
in01s10 FE_OCP_RBC4146_n_7743 ( .a(FE_OCP_RBN4142_n_7743), .o(FE_OCP_RBN4146_n_7743) );
in01s02 FE_OCP_RBC4147_n_3217 ( .a(n_3217), .o(FE_OCP_RBN4147_n_3217) );
in01s04 FE_OCP_RBC4148_n_24173 ( .a(n_24173), .o(FE_OCP_RBN4148_n_24173) );
in01s01 FE_OCP_RBC4149_n_24173 ( .a(n_24173), .o(FE_OCP_RBN4149_n_24173) );
in01s01 FE_OCP_RBC4150_n_13616 ( .a(n_13616), .o(FE_OCP_RBN4150_n_13616) );
in01f02 FE_OCP_RBC4151_n_13616 ( .a(n_13616), .o(FE_OCP_RBN4151_n_13616) );
in01s01 FE_OCP_RBC4152_n_13616 ( .a(FE_OCP_RBN4150_n_13616), .o(FE_OCP_RBN4152_n_13616) );
in01m04 FE_OCP_RBC4153_n_29378 ( .a(n_29378), .o(FE_OCP_RBN4153_n_29378) );
in01s01 FE_OCP_RBC4154_n_29378 ( .a(FE_OCP_RBN4153_n_29378), .o(FE_OCP_RBN4154_n_29378) );
in01s01 FE_OCP_RBC4156_n_29378 ( .a(FE_OCP_RBN4154_n_29378), .o(FE_OCP_RBN4156_n_29378) );
in01s01 FE_OCP_RBC4157_n_24222 ( .a(n_24222), .o(FE_OCP_RBN4157_n_24222) );
in01s02 FE_OCP_RBC4158_n_24222 ( .a(n_24222), .o(FE_OCP_RBN4158_n_24222) );
in01s01 FE_OCP_RBC4159_FE_OCPN857_n_7802 ( .a(FE_OCP_RBN2613_FE_OCPN857_n_7802), .o(FE_OCP_RBN4159_FE_OCPN857_n_7802) );
in01s01 FE_OCP_RBC4160_FE_OCPN857_n_7802 ( .a(FE_OCP_RBN2613_FE_OCPN857_n_7802), .o(FE_OCP_RBN4160_FE_OCPN857_n_7802) );
in01s01 FE_OCP_RBC4161_FE_OCPN857_n_7802 ( .a(FE_OCP_RBN2613_FE_OCPN857_n_7802), .o(FE_OCP_RBN4161_FE_OCPN857_n_7802) );
in01s02 FE_OCP_RBC4162_FE_OCPN857_n_7802 ( .a(FE_OCP_RBN2613_FE_OCPN857_n_7802), .o(FE_OCP_RBN4162_FE_OCPN857_n_7802) );
in01s02 FE_OCP_RBC4163_n_3390 ( .a(n_3390), .o(FE_OCP_RBN4163_n_3390) );
in01s02 FE_OCP_RBC4164_n_3390 ( .a(FE_OCP_RBN4163_n_3390), .o(FE_OCP_RBN4164_n_3390) );
in01s02 FE_OCP_RBC4165_n_3494 ( .a(n_3494), .o(FE_OCP_RBN4165_n_3494) );
in01s01 FE_OCP_RBC4166_n_3494 ( .a(FE_OCP_RBN4165_n_3494), .o(FE_OCP_RBN4166_n_3494) );
in01s01 FE_OCP_RBC4167_n_3494 ( .a(FE_OCP_RBN4165_n_3494), .o(FE_OCP_RBN4167_n_3494) );
in01s01 FE_OCP_RBC4168_n_29553 ( .a(n_29553), .o(FE_OCP_RBN4168_n_29553) );
in01m02 FE_OCP_RBC4169_n_29553 ( .a(n_29553), .o(FE_OCP_RBN4169_n_29553) );
in01s01 FE_OCP_RBC4170_n_19390 ( .a(n_19390), .o(FE_OCP_RBN4170_n_19390) );
in01s02 FE_OCP_RBC4171_n_19390 ( .a(n_19390), .o(FE_OCP_RBN4171_n_19390) );
in01m02 FE_OCP_RBC4172_n_38545 ( .a(n_38545), .o(FE_OCP_RBN4172_n_38545) );
in01s01 FE_OCP_RBC4173_n_38545 ( .a(n_38545), .o(FE_OCP_RBN4173_n_38545) );
in01m02 FE_OCP_RBC4174_FE_OCPN1913_n_2669 ( .a(FE_OCPN1913_n_2669), .o(FE_OCP_RBN4174_FE_OCPN1913_n_2669) );
in01s01 FE_OCP_RBC4175_n_3626 ( .a(n_3626), .o(FE_OCP_RBN4175_n_3626) );
in01s02 FE_OCP_RBC4176_n_3626 ( .a(n_3626), .o(FE_OCP_RBN4176_n_3626) );
in01f02 FE_OCP_RBC4177_n_38586 ( .a(n_38586), .o(FE_OCP_RBN4177_n_38586) );
in01s01 FE_OCP_RBC4178_n_38586 ( .a(n_38586), .o(FE_OCP_RBN4178_n_38586) );
in01s02 FE_OCP_RBC4179_n_38592 ( .a(n_38592), .o(FE_OCP_RBN4179_n_38592) );
in01s01 FE_OCP_RBC4180_n_38592 ( .a(n_38592), .o(FE_OCP_RBN4180_n_38592) );
in01s02 FE_OCP_RBC4181_n_19599 ( .a(n_19599), .o(FE_OCP_RBN4181_n_19599) );
in01s01 FE_OCP_RBC4182_n_19599 ( .a(n_19599), .o(FE_OCP_RBN4182_n_19599) );
in01s02 FE_OCP_RBC4184_n_24467 ( .a(n_24467), .o(FE_OCP_RBN4184_n_24467) );
in01f02 FE_OCP_RBC4185_n_8288 ( .a(n_8288), .o(FE_OCP_RBN4185_n_8288) );
in01s01 FE_OCP_RBC4186_n_8288 ( .a(n_8288), .o(FE_OCP_RBN4186_n_8288) );
in01s02 FE_OCP_RBC4187_n_8621 ( .a(n_8621), .o(FE_OCP_RBN4187_n_8621) );
in01f08 FE_OCP_RBC4188_n_13765 ( .a(n_13765), .o(FE_OCP_RBN4188_n_13765) );
in01s10 FE_OCP_RBC4189_n_13765 ( .a(FE_OCP_RBN4188_n_13765), .o(FE_OCP_RBN4189_n_13765) );
in01m02 FE_OCP_RBC4190_n_14279 ( .a(n_14279), .o(FE_OCP_RBN4190_n_14279) );
in01s06 FE_OCP_RBC4191_n_34285 ( .a(n_34285), .o(FE_OCP_RBN4191_n_34285) );
in01m02 FE_OCP_RBC4192_n_38537 ( .a(n_38537), .o(FE_OCP_RBN4192_n_38537) );
in01s01 FE_OCP_RBC4193_n_38537 ( .a(n_38537), .o(FE_OCP_RBN4193_n_38537) );
in01s03 FE_OCP_RBC4194_n_38683 ( .a(n_38683), .o(FE_OCP_RBN4194_n_38683) );
in01s02 FE_OCP_RBC4195_n_38683 ( .a(n_38683), .o(FE_OCP_RBN4195_n_38683) );
in01s01 FE_OCP_RBC4198_n_13796 ( .a(FE_OCP_RBN2758_n_13796), .o(FE_OCP_RBN4198_n_13796) );
in01m10 FE_OCP_RBC4199_n_13796 ( .a(FE_OCP_RBN2758_n_13796), .o(FE_OCP_RBN4199_n_13796) );
in01s02 FE_OCP_RBC4200_n_13796 ( .a(FE_OCP_RBN2758_n_13796), .o(FE_OCP_RBN4200_n_13796) );
in01s02 FE_OCP_RBC4201_n_13796 ( .a(FE_OCP_RBN4198_n_13796), .o(FE_OCP_RBN4201_n_13796) );
in01s01 FE_OCP_RBC4202_n_13796 ( .a(FE_OCP_RBN4199_n_13796), .o(FE_OCP_RBN4202_n_13796) );
in01s10 FE_OCP_RBC4203_n_13796 ( .a(FE_OCP_RBN4199_n_13796), .o(FE_OCP_RBN4203_n_13796) );
in01s01 FE_OCP_RBC4204_n_13796 ( .a(FE_OCP_RBN4199_n_13796), .o(FE_OCP_RBN4204_n_13796) );
in01m08 FE_OCP_RBC4205_n_13796 ( .a(FE_OCP_RBN4199_n_13796), .o(FE_OCP_RBN4205_n_13796) );
in01s01 FE_OCP_RBC4206_n_13796 ( .a(FE_OCP_RBN4201_n_13796), .o(FE_OCP_RBN4206_n_13796) );
in01s01 FE_OCP_RBC4208_n_13796 ( .a(FE_OCP_RBN4206_n_13796), .o(FE_OCP_RBN4208_n_13796) );
in01s01 FE_OCP_RBC4209_n_13796 ( .a(FE_OCP_RBN4208_n_13796), .o(FE_OCP_RBN4209_n_13796) );
in01s01 FE_OCP_RBC4210_n_13796 ( .a(FE_OCP_RBN4208_n_13796), .o(FE_OCP_RBN4210_n_13796) );
in01s01 FE_OCP_RBC4211_n_8767 ( .a(FE_OCP_RBN2786_n_8767), .o(FE_OCP_RBN4211_n_8767) );
in01m02 FE_OCP_RBC4212_n_3343 ( .a(n_3343), .o(FE_OCP_RBN4212_n_3343) );
in01s02 FE_OCP_RBC4213_n_3386 ( .a(n_3386), .o(FE_OCP_RBN4213_n_3386) );
in01s02 FE_OCP_RBC4214_FE_OCPN3565_n_10214 ( .a(FE_OCPN3565_n_10214), .o(FE_OCP_RBN4214_FE_OCPN3565_n_10214) );
in01s01 FE_OCP_RBC4215_FE_OCPN3565_n_10214 ( .a(FE_OCP_RBN4214_FE_OCPN3565_n_10214), .o(FE_OCP_RBN4215_FE_OCPN3565_n_10214) );
in01s01 FE_OCP_RBC4216_FE_OCPN3565_n_10214 ( .a(FE_OCP_RBN4215_FE_OCPN3565_n_10214), .o(FE_OCP_RBN4216_FE_OCPN3565_n_10214) );
in01s02 FE_OCP_RBC4217_n_8597 ( .a(n_8597), .o(FE_OCP_RBN4217_n_8597) );
in01s01 FE_OCP_RBC4218_n_8597 ( .a(n_8597), .o(FE_OCP_RBN4218_n_8597) );
in01s01 FE_OCP_RBC4219_n_8594 ( .a(n_8594), .o(FE_OCP_RBN4219_n_8594) );
in01s01 FE_OCP_RBC4220_n_8594 ( .a(n_8594), .o(FE_OCP_RBN4220_n_8594) );
in01m02 FE_OCP_RBC4221_n_8732 ( .a(n_8732), .o(FE_OCP_RBN4221_n_8732) );
in01s01 FE_OCP_RBC4222_n_8732 ( .a(n_8732), .o(FE_OCP_RBN4222_n_8732) );
in01m02 FE_OCP_RBC4223_n_8784 ( .a(n_8784), .o(FE_OCP_RBN4223_n_8784) );
in01m02 FE_OCP_RBC4224_n_8799 ( .a(n_8799), .o(FE_OCP_RBN4224_n_8799) );
in01s01 FE_OCP_RBC4226_n_13962 ( .a(FE_OCP_RBN5774_n_13796), .o(FE_OCP_RBN4226_n_13962) );
in01s01 FE_OCP_RBC4228_n_13962 ( .a(FE_OCP_RBN5774_n_13796), .o(FE_OCP_RBN4228_n_13962) );
in01s06 FE_OCP_RBC4229_n_13962 ( .a(FE_OCP_RBN5774_n_13796), .o(FE_OCP_RBN4229_n_13962) );
in01s01 FE_OCP_RBC4231_n_13962 ( .a(FE_OCP_RBN4229_n_13962), .o(FE_OCP_RBN4231_n_13962) );
in01s40 FE_OCP_RBC4232_n_13962 ( .a(FE_OCP_RBN6693_n_13796), .o(FE_OCP_RBN4232_n_13962) );
in01s01 FE_OCP_RBC4234_n_13962 ( .a(FE_OCP_RBN4231_n_13962), .o(FE_OCP_RBN4234_n_13962) );
in01m02 FE_OCP_RBC4235_n_9089 ( .a(n_9089), .o(FE_OCP_RBN4235_n_9089) );
in01s02 FE_OCP_RBC4236_n_9089 ( .a(n_9089), .o(FE_OCP_RBN4236_n_9089) );
in01s02 FE_OCP_RBC4237_n_8781 ( .a(n_8781), .o(FE_OCP_RBN4237_n_8781) );
in01s01 FE_OCP_RBC4238_n_8781 ( .a(n_8781), .o(FE_OCP_RBN4238_n_8781) );
in01s01 FE_OCP_RBC4239_n_44594 ( .a(n_44594), .o(FE_OCP_RBN4239_n_44594) );
in01s06 FE_OCP_RBC4240_n_44594 ( .a(n_44594), .o(FE_OCP_RBN4240_n_44594) );
in01s01 FE_OCP_RBC4241_n_44594 ( .a(n_44594), .o(FE_OCP_RBN4241_n_44594) );
in01s01 FE_OCP_RBC4242_n_44594 ( .a(n_44594), .o(FE_OCP_RBN4242_n_44594) );
in01s01 FE_OCP_RBC4243_n_44594 ( .a(FE_OCP_RBN4241_n_44594), .o(FE_OCP_RBN4243_n_44594) );
in01s01 FE_OCP_RBC4244_n_44594 ( .a(FE_OCP_RBN4242_n_44594), .o(FE_OCP_RBN4244_n_44594) );
in01m04 FE_OCP_RBC4246_n_8904 ( .a(FE_OFN5066_n_8904), .o(FE_OCP_RBN4246_n_8904) );
in01s01 FE_OCP_RBC4247_n_8904 ( .a(FE_OFN5066_n_8904), .o(FE_OCP_RBN4247_n_8904) );
in01f01 FE_OCP_RBC4248_n_14573 ( .a(n_14573), .o(FE_OCP_RBN4248_n_14573) );
in01f01 FE_OCP_RBC4249_n_14697 ( .a(n_14697), .o(FE_OCP_RBN4249_n_14697) );
in01s01 FE_OCP_RBC4251_n_8687 ( .a(FE_OCP_RBN5818_n_8687), .o(FE_OCP_RBN4251_n_8687) );
in01s01 FE_OCP_RBC4252_n_8687 ( .a(FE_OCP_RBN5818_n_8687), .o(FE_OCP_RBN4252_n_8687) );
in01s01 FE_OCP_RBC4253_n_8687 ( .a(FE_OCP_RBN4251_n_8687), .o(FE_OCP_RBN4253_n_8687) );
in01s01 FE_OCP_RBC4254_n_3705 ( .a(n_3705), .o(FE_OCP_RBN4254_n_3705) );
in01m08 FE_OCP_RBC4255_n_3705 ( .a(n_3705), .o(FE_OCP_RBN4255_n_3705) );
in01s01 FE_OCP_RBC4256_n_3705 ( .a(n_3705), .o(FE_OCP_RBN4256_n_3705) );
in01f02 FE_OCP_RBC4258_n_34921 ( .a(n_34921), .o(FE_OCP_RBN4258_n_34921) );
in01s01 FE_OCP_RBC4259_n_34921 ( .a(FE_OCP_RBN4258_n_34921), .o(FE_OCP_RBN4259_n_34921) );
in01s01 FE_OCP_RBC4260_n_34921 ( .a(FE_OCP_RBN4259_n_34921), .o(FE_OCP_RBN4260_n_34921) );
in01s02 FE_OCP_RBC4261_n_34878 ( .a(n_34878), .o(FE_OCP_RBN4261_n_34878) );
in01s01 FE_OCP_RBC4262_n_9009 ( .a(n_9009), .o(FE_OCP_RBN4262_n_9009) );
in01f02 FE_OCP_RBC4263_n_9009 ( .a(n_9009), .o(FE_OCP_RBN4263_n_9009) );
in01s01 FE_OCP_RBC4266_FE_RN_998_0 ( .a(FE_OCP_RBN5860_FE_RN_998_0), .o(FE_OCP_RBN4266_FE_RN_998_0) );
in01f02 FE_OCP_RBC4269_n_8872 ( .a(FE_OCP_RBN2881_n_8872), .o(FE_OCP_RBN4269_n_8872) );
in01s02 FE_OCP_RBC4270_n_8872 ( .a(FE_OCP_RBN4269_n_8872), .o(FE_OCP_RBN4270_n_8872) );
in01s01 FE_OCP_RBC4274_n_3700 ( .a(FE_OCP_RBN5871_n_3700), .o(FE_OCP_RBN4274_n_3700) );
in01s01 FE_OCP_RBC4280_n_3848 ( .a(FE_OCP_RBN5877_n_3848), .o(FE_OCP_RBN4280_n_3848) );
in01s01 FE_OCP_RBC4281_n_3848 ( .a(FE_OCP_RBN4280_n_3848), .o(FE_OCP_RBN4281_n_3848) );
in01s01 FE_OCP_RBC4282_n_9243 ( .a(n_9243), .o(FE_OCP_RBN4282_n_9243) );
in01s02 FE_OCP_RBC4283_n_9243 ( .a(n_9243), .o(FE_OCP_RBN4283_n_9243) );
in01s01 FE_OCP_RBC4288_n_44563 ( .a(FE_OCP_RBN6741_n_44563), .o(FE_OCP_RBN4288_n_44563) );
in01s02 FE_OCP_RBC4289_n_47014 ( .a(n_47014), .o(FE_OCP_RBN4289_n_47014) );
in01s01 FE_OCP_RBC4290_n_47014 ( .a(FE_OCP_RBN4289_n_47014), .o(FE_OCP_RBN4290_n_47014) );
in01s01 FE_OCP_RBC4291_n_3909 ( .a(n_3909), .o(FE_OCP_RBN4291_n_3909) );
in01s02 FE_OCP_RBC4292_n_4080 ( .a(n_4080), .o(FE_OCP_RBN4292_n_4080) );
in01s01 FE_OCP_RBC4293_n_4080 ( .a(FE_OCP_RBN4292_n_4080), .o(FE_OCP_RBN4293_n_4080) );
in01s01 FE_OCP_RBC4294_n_4080 ( .a(FE_OCP_RBN4293_n_4080), .o(FE_OCP_RBN4294_n_4080) );
in01s01 FE_OCP_RBC4295_n_4080 ( .a(FE_OCP_RBN4294_n_4080), .o(FE_OCP_RBN4295_n_4080) );
in01s01 FE_OCP_RBC4296_n_4080 ( .a(FE_OCP_RBN4295_n_4080), .o(FE_OCP_RBN4296_n_4080) );
in01s01 FE_OCP_RBC4298_n_25238 ( .a(FE_OCP_RBN5923_n_25211), .o(FE_OCP_RBN4298_n_25238) );
in01s01 FE_OCP_RBC4302_n_44579 ( .a(FE_OCP_RBN6736_n_44579), .o(FE_OCP_RBN4302_n_44579) );
in01s01 FE_OCP_RBC4303_n_44579 ( .a(FE_OCP_RBN6736_n_44579), .o(FE_OCP_RBN4303_n_44579) );
in01s01 FE_OCP_RBC4304_n_44579 ( .a(FE_OCP_RBN4302_n_44579), .o(FE_OCP_RBN4304_n_44579) );
in01s01 FE_OCP_RBC4305_n_44579 ( .a(FE_OCP_RBN4304_n_44579), .o(FE_OCP_RBN4305_n_44579) );
in01s01 FE_OCP_RBC4307_n_25178 ( .a(FE_OCP_RBN2910_n_25178), .o(FE_OCP_RBN4307_n_25178) );
in01m10 FE_OCP_RBC4309_n_25178 ( .a(FE_OCP_RBN2910_n_25178), .o(FE_OCP_RBN4309_n_25178) );
in01s10 FE_OCP_RBC4311_n_25178 ( .a(FE_OCP_RBN5900_n_25178), .o(FE_OCP_RBN4311_n_25178) );
in01m02 FE_OCP_RBC4314_n_9396 ( .a(n_9396), .o(FE_OCP_RBN4314_n_9396) );
in01m02 FE_OCP_RBC4315_n_14881 ( .a(n_14881), .o(FE_OCP_RBN4315_n_14881) );
in01s01 FE_OCP_RBC4316_n_9292 ( .a(n_9292), .o(FE_OCP_RBN4316_n_9292) );
in01m02 FE_OCP_RBC4317_n_9292 ( .a(n_9292), .o(FE_OCP_RBN4317_n_9292) );
in01s01 FE_OCP_RBC4319_n_14768 ( .a(n_14768), .o(FE_OCP_RBN4319_n_14768) );
in01m04 FE_OCP_RBC4322_n_15156 ( .a(n_15156), .o(FE_OCP_RBN4322_n_15156) );
in01m04 FE_OCP_RBC4323_n_15156 ( .a(FE_OCP_RBN4322_n_15156), .o(FE_OCP_RBN4323_n_15156) );
in01s04 FE_OCP_RBC4324_n_15156 ( .a(FE_OCP_RBN4322_n_15156), .o(FE_OCP_RBN4324_n_15156) );
in01s02 FE_OCP_RBC4325_n_20333 ( .a(n_20333), .o(FE_OCP_RBN4325_n_20333) );
in01s01 FE_OCP_RBC4326_n_20333 ( .a(FE_OCP_RBN4325_n_20333), .o(FE_OCP_RBN4326_n_20333) );
in01s04 FE_OCP_RBC4327_n_38878 ( .a(FE_OCP_RBN5896_n_38806), .o(FE_OCP_RBN4327_n_38878) );
in01s10 FE_OCP_RBC4328_n_38878 ( .a(FE_OCP_RBN5895_n_38806), .o(FE_OCP_RBN4328_n_38878) );
in01s06 FE_OCP_RBC4329_n_38878 ( .a(FE_OCP_RBN4328_n_38878), .o(FE_OCP_RBN4329_n_38878) );
in01s02 FE_OCP_RBC4330_n_9102 ( .a(n_9102), .o(FE_OCP_RBN4330_n_9102) );
in01s02 FE_OCP_RBC4334_n_20242 ( .a(FE_OCP_RBN2944_n_20242), .o(FE_OCP_RBN4334_n_20242) );
in01s01 FE_OCP_RBC4335_n_20242 ( .a(FE_OCP_RBN2944_n_20242), .o(FE_OCP_RBN4335_n_20242) );
in01s02 FE_OCP_RBC4337_n_20242 ( .a(FE_OCP_RBN2944_n_20242), .o(FE_OCP_RBN4337_n_20242) );
in01s01 FE_OCP_RBC4338_n_9521 ( .a(n_9521), .o(FE_OCP_RBN4338_n_9521) );
in01s01 FE_OCP_RBC4339_n_4403 ( .a(n_4403), .o(FE_OCP_RBN4339_n_4403) );
in01s01 FE_OCP_RBC4340_n_4403 ( .a(n_4403), .o(FE_OCP_RBN4340_n_4403) );
in01s01 FE_OCP_RBC4341_n_25500 ( .a(n_25500), .o(FE_OCP_RBN4341_n_25500) );
in01s01 FE_OCP_RBC4342_n_4198 ( .a(n_4198), .o(FE_OCP_RBN4342_n_4198) );
in01m02 FE_OCP_RBC4343_n_15071 ( .a(n_15071), .o(FE_OCP_RBN4343_n_15071) );
in01s08 FE_OCP_RBC4344_n_35177 ( .a(n_35177), .o(FE_OCP_RBN4344_n_35177) );
in01s02 FE_OCP_RBC4345_n_4378 ( .a(n_4378), .o(FE_OCP_RBN4345_n_4378) );
in01s02 FE_OCP_RBC4347_n_10017 ( .a(n_10017), .o(FE_OCP_RBN4347_n_10017) );
in01s01 FE_OCP_RBC4348_n_20568 ( .a(n_20568), .o(FE_OCP_RBN4348_n_20568) );
in01s01 FE_OCP_RBC4349_n_9975 ( .a(n_9975), .o(FE_OCP_RBN4349_n_9975) );
in01s01 FE_OCP_RBC4350_n_9975 ( .a(n_9975), .o(FE_OCP_RBN4350_n_9975) );
in01s06 FE_OCP_RBC4351_n_20456 ( .a(n_20456), .o(FE_OCP_RBN4351_n_20456) );
in01s01 FE_OCP_RBC4352_FE_OCPN1263_n_20971 ( .a(FE_OCPN1263_n_20971), .o(FE_OCP_RBN4352_FE_OCPN1263_n_20971) );
in01s01 FE_OCP_RBC4353_FE_OCPN1263_n_20971 ( .a(FE_OCPN1263_n_20971), .o(FE_OCP_RBN4353_FE_OCPN1263_n_20971) );
in01s02 FE_OCP_RBC4354_n_4585 ( .a(n_4585), .o(FE_OCP_RBN4354_n_4585) );
in01s01 FE_OCP_RBC4355_n_10100 ( .a(FE_OCP_RBN3052_n_10100), .o(FE_OCP_RBN4355_n_10100) );
in01s01 FE_OCP_RBC4356_n_10100 ( .a(FE_OCP_RBN3052_n_10100), .o(FE_OCP_RBN4356_n_10100) );
in01s06 FE_OCP_RBC4357_n_10100 ( .a(FE_OCP_RBN3052_n_10100), .o(FE_OCP_RBN4357_n_10100) );
in01s01 FE_OCP_RBC4358_n_10100 ( .a(FE_OCP_RBN4357_n_10100), .o(FE_OCP_RBN4358_n_10100) );
in01s01 FE_OCP_RBC4359_n_10100 ( .a(FE_OCP_RBN4358_n_10100), .o(FE_OCP_RBN4359_n_10100) );
in01s01 FE_OCP_RBC4360_n_20632 ( .a(n_20632), .o(FE_OCP_RBN4360_n_20632) );
in01f01 FE_OCP_RBC4361_FE_RN_1500_0 ( .a(FE_RN_1500_0), .o(FE_OCP_RBN4361_FE_RN_1500_0) );
in01m02 FE_OCP_RBC4362_FE_RN_1500_0 ( .a(FE_RN_1500_0), .o(FE_OCP_RBN4362_FE_RN_1500_0) );
in01s04 FE_OCP_RBC4363_n_39584 ( .a(n_39584), .o(FE_OCP_RBN4363_n_39584) );
in01s03 FE_OCP_RBC4364_n_20710 ( .a(FE_OCP_RBN3103_n_20710), .o(FE_OCP_RBN4364_n_20710) );
in01s01 FE_OCP_RBC4365_n_4692 ( .a(n_4692), .o(FE_OCP_RBN4365_n_4692) );
in01s01 FE_OCP_RBC4366_n_4692 ( .a(n_4692), .o(FE_OCP_RBN4366_n_4692) );
in01s01 FE_OCP_RBC4367_n_25889 ( .a(n_25889), .o(FE_OCP_RBN4367_n_25889) );
in01m04 FE_OCP_RBC4368_n_25889 ( .a(n_25889), .o(FE_OCP_RBN4368_n_25889) );
in01s04 FE_OCP_RBC4369_n_46982 ( .a(n_46982), .o(FE_OCP_RBN4369_n_46982) );
in01s01 FE_OCP_RBC4370_n_46982 ( .a(FE_OCP_RBN4369_n_46982), .o(FE_OCP_RBN4370_n_46982) );
in01s01 FE_OCP_RBC4371_n_5032 ( .a(n_5032), .o(FE_OCP_RBN4371_n_5032) );
in01s01 FE_OCP_RBC4372_n_5048 ( .a(n_5048), .o(FE_OCP_RBN4372_n_5048) );
in01s01 FE_OCP_RBC4373_n_5048 ( .a(FE_OCP_RBN4372_n_5048), .o(FE_OCP_RBN4373_n_5048) );
in01s01 FE_OCP_RBC4374_n_5048 ( .a(FE_OCP_RBN4373_n_5048), .o(FE_OCP_RBN4374_n_5048) );
in01s02 FE_OCP_RBC4375_n_15514 ( .a(n_15514), .o(FE_OCP_RBN4375_n_15514) );
in01f02 FE_OCP_RBC4377_n_15700 ( .a(n_15700), .o(FE_OCP_RBN4377_n_15700) );
in01s01 FE_OCP_RBC4378_n_4956 ( .a(n_4956), .o(FE_OCP_RBN4378_n_4956) );
in01s02 FE_OCP_RBC4379_n_4956 ( .a(n_4956), .o(FE_OCP_RBN4379_n_4956) );
in01s02 FE_OCP_RBC4380_n_5028 ( .a(n_5028), .o(FE_OCP_RBN4380_n_5028) );
in01s02 FE_OCP_RBC4381_n_5041 ( .a(n_5041), .o(FE_OCP_RBN4381_n_5041) );
in01s01 FE_OCP_RBC4382_n_39523 ( .a(n_39523), .o(FE_OCP_RBN4382_n_39523) );
in01s01 FE_OCP_RBC4384_n_5221 ( .a(n_5221), .o(FE_OCP_RBN4384_n_5221) );
in01s01 FE_OCP_RBC4385_n_10570 ( .a(n_10570), .o(FE_OCP_RBN4385_n_10570) );
in01s02 FE_OCP_RBC4387_n_5013 ( .a(n_5013), .o(FE_OCP_RBN4387_n_5013) );
in01s02 FE_OCP_RBC4388_n_26173 ( .a(n_26173), .o(FE_OCP_RBN4388_n_26173) );
in01s01 FE_OCP_RBC4389_n_26173 ( .a(FE_OCP_RBN4388_n_26173), .o(FE_OCP_RBN4389_n_26173) );
in01s01 FE_OCP_RBC4390_n_26173 ( .a(FE_OCP_RBN4389_n_26173), .o(FE_OCP_RBN4390_n_26173) );
in01f06 FE_OCP_RBC4391_n_16230 ( .a(n_16230), .o(FE_OCP_RBN4391_n_16230) );
in01s06 FE_OCP_RBC4392_n_26146 ( .a(n_26146), .o(FE_OCP_RBN4392_n_26146) );
in01s02 FE_OCP_RBC4393_n_10682 ( .a(n_10682), .o(FE_OCP_RBN4393_n_10682) );
in01m04 FE_OCP_RBC4394_n_16146 ( .a(n_16146), .o(FE_OCP_RBN4394_n_16146) );
in01s01 FE_OCP_RBC4395_n_16146 ( .a(FE_OCP_RBN4394_n_16146), .o(FE_OCP_RBN4395_n_16146) );
in01s01 FE_OCP_RBC4396_n_16146 ( .a(FE_OCP_RBN4395_n_16146), .o(FE_OCP_RBN4396_n_16146) );
in01f02 FE_OCP_RBC4398_n_39629 ( .a(n_39629), .o(FE_OCP_RBN4398_n_39629) );
in01s02 FE_OCP_RBC4399_n_5308 ( .a(n_5308), .o(FE_OCP_RBN4399_n_5308) );
in01s02 FE_OCP_RBC4400_n_5532 ( .a(n_5532), .o(FE_OCP_RBN4400_n_5532) );
in01m04 FE_OCP_RBC4401_n_16321 ( .a(n_16321), .o(FE_OCP_RBN4401_n_16321) );
in01s01 FE_OCP_RBC4402_n_43013 ( .a(n_43013), .o(FE_OCP_RBN4402_n_43013) );
in01s06 FE_OCP_RBC4405_n_26160 ( .a(FE_OCP_RBN6097_n_26160), .o(FE_OCP_RBN4405_n_26160) );
in01s04 FE_OCP_RBC4408_n_26394 ( .a(n_26394), .o(FE_OCP_RBN4408_n_26394) );
in01m02 FE_OCP_RBC4409_n_16429 ( .a(n_16429), .o(FE_OCP_RBN4409_n_16429) );
in01s02 FE_OCP_RBC4412_n_26661 ( .a(n_26661), .o(FE_OCP_RBN4412_n_26661) );
in01s01 FE_OCP_RBC4413_n_31117 ( .a(n_31117), .o(FE_OCP_RBN4413_n_31117) );
in01s06 FE_OCP_RBC4414_n_31117 ( .a(n_31117), .o(FE_OCP_RBN4414_n_31117) );
in01s02 FE_OCP_RBC4415_n_31117 ( .a(n_31117), .o(FE_OCP_RBN4415_n_31117) );
in01s01 FE_OCP_RBC4416_n_31117 ( .a(FE_OCP_RBN4413_n_31117), .o(FE_OCP_RBN4416_n_31117) );
in01s01 FE_OCP_RBC4417_n_31117 ( .a(FE_OCP_RBN4413_n_31117), .o(FE_OCP_RBN4417_n_31117) );
in01s02 FE_OCP_RBC4418_n_31117 ( .a(FE_OCP_RBN4414_n_31117), .o(FE_OCP_RBN4418_n_31117) );
in01s06 FE_OCP_RBC4419_n_31117 ( .a(FE_OCP_RBN4414_n_31117), .o(FE_OCP_RBN4419_n_31117) );
in01s01 FE_OCP_RBC4420_n_31117 ( .a(FE_OCP_RBN4415_n_31117), .o(FE_OCP_RBN4420_n_31117) );
in01s01 FE_OCP_RBC4421_n_31117 ( .a(FE_OCP_RBN4415_n_31117), .o(FE_OCP_RBN4421_n_31117) );
in01s01 FE_OCP_RBC4422_n_31117 ( .a(FE_OCP_RBN4420_n_31117), .o(FE_OCP_RBN4422_n_31117) );
in01s01 FE_OCP_RBC4423_n_31117 ( .a(FE_OCP_RBN4420_n_31117), .o(FE_OCP_RBN4423_n_31117) );
in01s01 FE_OCP_RBC4424_n_31117 ( .a(FE_OCP_RBN4420_n_31117), .o(FE_OCP_RBN4424_n_31117) );
in01s01 FE_OCP_RBC4425_n_31117 ( .a(FE_OCP_RBN4421_n_31117), .o(FE_OCP_RBN4425_n_31117) );
in01m04 FE_OCP_RBC4429_n_39942 ( .a(FE_OCP_RBN6852_n_39793), .o(FE_OCP_RBN4429_n_39942) );
in01s10 FE_OCP_RBC4430_n_39942 ( .a(FE_OCP_RBN6852_n_39793), .o(FE_OCP_RBN4430_n_39942) );
in01m10 FE_OCP_RBC4431_n_39942 ( .a(FE_OCP_RBN6852_n_39793), .o(FE_OCP_RBN4431_n_39942) );
in01s02 FE_OCP_RBC4432_n_26160 ( .a(FE_OCP_RBN6858_n_26160), .o(FE_OCP_RBN4432_n_26160) );
in01s01 FE_OCP_RBC4433_n_26160 ( .a(FE_OCP_RBN6858_n_26160), .o(FE_OCP_RBN4433_n_26160) );
in01s03 FE_OCP_RBC4434_n_26160 ( .a(FE_OCP_RBN4432_n_26160), .o(FE_OCP_RBN4434_n_26160) );
in01s01 FE_OCP_RBC4435_n_26160 ( .a(FE_OCP_RBN4433_n_26160), .o(FE_OCP_RBN4435_n_26160) );
in01s01 FE_OCP_RBC4436_n_26160 ( .a(FE_OCP_RBN4433_n_26160), .o(FE_OCP_RBN4436_n_26160) );
in01s01 FE_OCP_RBC4437_n_26160 ( .a(FE_OCP_RBN4436_n_26160), .o(FE_OCP_RBN4437_n_26160) );
in01s01 FE_OCP_RBC4438_n_26160 ( .a(FE_OCP_RBN4436_n_26160), .o(FE_OCP_RBN4438_n_26160) );
in01s01 FE_OCP_RBC4439_n_26160 ( .a(FE_OCP_RBN4436_n_26160), .o(FE_OCP_RBN4439_n_26160) );
in01s02 FE_OCP_RBC4441_n_5891 ( .a(FE_OCP_RBN4440_n_5891), .o(FE_OCP_RBN4441_n_5891) );
in01s02 FE_OCP_RBC4443_n_46424 ( .a(n_46424), .o(FE_OCP_RBN4443_n_46424) );
in01s01 FE_OCP_RBC4445_n_43022 ( .a(FE_OCP_RBN3312_n_43022), .o(FE_OCP_RBN4445_n_43022) );
in01s01 FE_OCP_RBC4446_n_43022 ( .a(FE_OCP_RBN4445_n_43022), .o(FE_OCP_RBN4446_n_43022) );
in01s01 FE_OCP_RBC4447_FE_OFN760_n_46337 ( .a(FE_OCP_RBN6163_n_46337), .o(FE_OCP_RBN4447_FE_OFN760_n_46337) );
in01s01 FE_OCP_RBC4448_FE_OFN760_n_46337 ( .a(FE_OCP_RBN6163_n_46337), .o(FE_OCP_RBN4448_FE_OFN760_n_46337) );
in01s01 FE_OCP_RBC4451_n_5870 ( .a(n_5870), .o(FE_OCP_RBN4451_n_5870) );
in01m04 FE_OCP_RBC4454_n_6102 ( .a(n_6102), .o(FE_OCP_RBN4454_n_6102) );
in01m04 FE_OCP_RBC4455_n_6102 ( .a(n_6102), .o(FE_OCP_RBN4455_n_6102) );
in01s20 FE_OCP_RBC4456_n_43103 ( .a(n_43103), .o(FE_OCP_RBN4456_n_43103) );
in01s10 FE_OCP_RBC4457_n_43103 ( .a(FE_OCP_RBN4456_n_43103), .o(FE_OCP_RBN4457_n_43103) );
in01m02 FE_OCP_RBC4458_FE_RN_1190_0 ( .a(FE_RN_1190_0), .o(FE_OCP_RBN4458_FE_RN_1190_0) );
in01f02 FE_OCP_RBC4459_FE_RN_1190_0 ( .a(FE_RN_1190_0), .o(FE_OCP_RBN4459_FE_RN_1190_0) );
in01s02 FE_OCP_RBC4462_n_44267 ( .a(FE_OCP_RBN6182_n_44267), .o(FE_OCP_RBN4462_n_44267) );
in01s02 FE_OCP_RBC4464_n_44267 ( .a(FE_OCP_RBN6182_n_44267), .o(FE_OCP_RBN4464_n_44267) );
in01s02 FE_OCP_RBC4466_n_44267 ( .a(FE_OCP_RBN6185_n_44267), .o(FE_OCP_RBN4466_n_44267) );
in01s02 FE_OCP_RBC4467_n_44267 ( .a(FE_OCP_RBN6184_n_44267), .o(FE_OCP_RBN4467_n_44267) );
in01s06 FE_OCP_RBC4468_n_44267 ( .a(FE_OCP_RBN4464_n_44267), .o(FE_OCP_RBN4468_n_44267) );
in01s02 FE_OCP_RBC4471_n_31819 ( .a(FE_OCP_RBN3390_n_31819), .o(FE_OCP_RBN4471_n_31819) );
in01s02 FE_OCP_RBC4472_n_31819 ( .a(FE_OCP_RBN3390_n_31819), .o(FE_OCP_RBN4472_n_31819) );
in01s01 FE_OCP_RBC4476_FE_OCPN913_n_43230 ( .a(FE_OCP_RBN6191_n_43103), .o(FE_OCP_RBN4476_FE_OCPN913_n_43230) );
in01s01 FE_OCP_RBC4477_FE_OCPN913_n_43230 ( .a(FE_OCP_RBN6191_n_43103), .o(FE_OCP_RBN4477_FE_OCPN913_n_43230) );
in01s06 FE_OCP_RBC4478_FE_OCPN913_n_43230 ( .a(FE_OCP_RBN6191_n_43103), .o(FE_OCP_RBN4478_FE_OCPN913_n_43230) );
in01s06 FE_OCP_RBC4479_FE_OCPN913_n_43230 ( .a(FE_OCP_RBN6191_n_43103), .o(FE_OCP_RBN4479_FE_OCPN913_n_43230) );
in01s01 FE_OCP_RBC4480_n_11439 ( .a(FE_OCP_RBN3384_n_11439), .o(FE_OCP_RBN4480_n_11439) );
in01s02 FE_OCP_RBC4481_n_11439 ( .a(FE_OCP_RBN3384_n_11439), .o(FE_OCP_RBN4481_n_11439) );
in01s06 FE_OCP_RBC4482_n_11439 ( .a(FE_OCP_RBN3384_n_11439), .o(FE_OCP_RBN4482_n_11439) );
in01s06 FE_OCP_RBC4483_n_11439 ( .a(FE_OCP_RBN4481_n_11439), .o(FE_OCP_RBN4483_n_11439) );
in01s01 FE_OCP_RBC4484_n_22667 ( .a(n_22667), .o(FE_OCP_RBN4484_n_22667) );
in01s01 FE_OCP_RBC4485_n_22667 ( .a(FE_OCP_RBN4484_n_22667), .o(FE_OCP_RBN4485_n_22667) );
in01s02 FE_OCP_RBC4486_n_27145 ( .a(n_27145), .o(FE_OCP_RBN4486_n_27145) );
in01s02 FE_OCP_RBC4487_n_22438 ( .a(n_22438), .o(FE_OCP_RBN4487_n_22438) );
in01m02 FE_OCP_RBC4488_n_6299 ( .a(n_6299), .o(FE_OCP_RBN4488_n_6299) );
in01s02 FE_OCP_RBC4489_n_6299 ( .a(n_6299), .o(FE_OCP_RBN4489_n_6299) );
in01s01 FE_OCP_RBC4490_n_32152 ( .a(n_32152), .o(FE_OCP_RBN4490_n_32152) );
in01m02 FE_OCP_RBC4492_n_22755 ( .a(n_22755), .o(FE_OCP_RBN4492_n_22755) );
in01s01 FE_OCP_RBC4494_n_27555 ( .a(n_27555), .o(FE_OCP_RBN4494_n_27555) );
in01s01 FE_OCP_RBC4495_n_27639 ( .a(n_27639), .o(FE_OCP_RBN4495_n_27639) );
in01s01 FE_OCP_RBC4496_n_27639 ( .a(n_27639), .o(FE_OCP_RBN4496_n_27639) );
in01s40 FE_OCP_RBC4590_n_44847 ( .a(n_44847), .o(FE_OCP_RBN4590_n_44847) );
in01s06 FE_OCP_RBC4593_delay_xor_ln22_unr12_stage5_stallmux_q_1_ ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_1_), .o(FE_OCP_RBN4593_delay_xor_ln22_unr12_stage5_stallmux_q_1_) );
in01s40 FE_OCP_RBC4630_n_44962 ( .a(FE_OCP_RBN7012_n_44962), .o(FE_OCP_RBN4630_n_44962) );
in01s80 FE_OCP_RBC4633_n_44962 ( .a(FE_OCP_RBN7012_n_44962), .o(FE_OCP_RBN4633_n_44962) );
in01s01 FE_OCP_RBC4635_n_33589 ( .a(n_33589), .o(FE_OCP_RBN4635_n_33589) );
in01s01 FE_OCP_RBC4636_n_18600 ( .a(n_18600), .o(FE_OCP_RBN4636_n_18600) );
in01s01 FE_OCP_RBC4637_n_18600 ( .a(FE_OCP_RBN4636_n_18600), .o(FE_OCP_RBN4637_n_18600) );
in01s01 FE_OCP_RBC4639_n_18681 ( .a(n_18681), .o(FE_OCP_RBN4639_n_18681) );
in01s01 FE_OCP_RBC4643_n_35121 ( .a(n_35121), .o(FE_OCP_RBN4643_n_35121) );
in01f02 FE_OCP_RBC4644_n_20420 ( .a(n_20420), .o(FE_OCP_RBN4644_n_20420) );
in01s01 FE_OCP_RBC4645_n_20420 ( .a(n_20420), .o(FE_OCP_RBN4645_n_20420) );
in01m06 FE_OCP_RBC4646_n_22553 ( .a(n_22553), .o(FE_OCP_RBN4646_n_22553) );
in01m06 FE_OCP_RBC4647_n_22553 ( .a(FE_OCP_RBN4646_n_22553), .o(FE_OCP_RBN4647_n_22553) );
in01m02 FE_OCP_RBC4648_n_22625 ( .a(n_22625), .o(FE_OCP_RBN4648_n_22625) );
in01m02 FE_OCP_RBC4649_n_22625 ( .a(n_22625), .o(FE_OCP_RBN4649_n_22625) );
in01f02 FE_OCP_RBC4870_n_35145 ( .a(n_35145), .o(FE_OCP_RBN4870_n_35145) );
in01m01 FE_OCP_RBC4900_n_29056 ( .a(n_29056), .o(FE_OCP_RBN4900_n_29056) );
in01s01 FE_OCP_RBC4902_n_44256 ( .a(n_44256), .o(FE_OCP_RBN4902_n_44256) );
in01m10 FE_OCP_RBC4903_n_44256 ( .a(n_44256), .o(FE_OCP_RBN4903_n_44256) );
in01m10 FE_OCP_RBC4904_n_44256 ( .a(FE_OCP_RBN4903_n_44256), .o(FE_OCP_RBN4904_n_44256) );
in01m08 FE_OCP_RBC4905_n_44256 ( .a(FE_OCP_RBN4903_n_44256), .o(FE_OCP_RBN4905_n_44256) );
in01s03 FE_OCP_RBC4906_n_44256 ( .a(FE_OCP_RBN4904_n_44256), .o(FE_OCP_RBN4906_n_44256) );
in01m10 FE_OCP_RBC4908_n_44222 ( .a(n_44222), .o(FE_OCP_RBN4908_n_44222) );
in01s06 FE_OCP_RBC4909_n_44222 ( .a(FE_OCP_RBN4908_n_44222), .o(FE_OCP_RBN4909_n_44222) );
in01s20 FE_OCP_RBC4910_n_44222 ( .a(FE_OCP_RBN4908_n_44222), .o(FE_OCP_RBN4910_n_44222) );
in01s06 FE_OCP_RBC4912_n_33803 ( .a(FE_OCP_RBN6568_n_33803), .o(FE_OCP_RBN4912_n_33803) );
in01m06 FE_OCP_RBC4913_n_33833 ( .a(n_33833), .o(FE_OCP_RBN4913_n_33833) );
in01f02 FE_OCP_RBC4914_n_33833 ( .a(n_33833), .o(FE_OCP_RBN4914_n_33833) );
in01s02 FE_OCP_RBC4915_n_33503 ( .a(n_33503), .o(FE_OCP_RBN4915_n_33503) );
in01s01 FE_OCP_RBC4916_n_33503 ( .a(FE_OCP_RBN4915_n_33503), .o(FE_OCP_RBN4916_n_33503) );
in01s02 FE_OCP_RBC4917_n_33491 ( .a(FE_OCP_RBN4049_n_33491), .o(FE_OCP_RBN4917_n_33491) );
in01s01 FE_OCP_RBC4918_n_33491 ( .a(FE_OCP_RBN4917_n_33491), .o(FE_OCP_RBN4918_n_33491) );
in01m10 FE_OCP_RBC4919_n_32575 ( .a(n_32575), .o(FE_OCP_RBN4919_n_32575) );
in01s01 FE_OCP_RBC4920_n_33691 ( .a(n_33691), .o(FE_OCP_RBN4920_n_33691) );
in01m02 FE_OCP_RBC4921_n_33691 ( .a(n_33691), .o(FE_OCP_RBN4921_n_33691) );
in01f02 FE_OCP_RBC4923_n_34980 ( .a(n_34980), .o(FE_OCP_RBN4923_n_34980) );
in01s01 FE_OCP_RBC4924_n_34980 ( .a(FE_OCP_RBN4923_n_34980), .o(FE_OCP_RBN4924_n_34980) );
in01s01 FE_OCP_RBC4925_n_34980 ( .a(FE_OCP_RBN4924_n_34980), .o(FE_OCP_RBN4925_n_34980) );
in01s06 FE_OCP_RBC5016_n_12026 ( .a(n_12026), .o(FE_OCP_RBN5016_n_12026) );
in01s06 FE_OCP_RBC5017_n_12026 ( .a(FE_OCP_RBN5016_n_12026), .o(FE_OCP_RBN5017_n_12026) );
in01s10 FE_OCP_RBC5018_n_16972 ( .a(n_16972), .o(FE_OCP_RBN5018_n_16972) );
in01m01 FE_OCP_RBC5019_n_13726 ( .a(n_13726), .o(FE_OCP_RBN5019_n_13726) );
in01s01 FE_OCP_RBC5021_n_13726 ( .a(FE_OCP_RBN6639_n_13726), .o(FE_OCP_RBN5021_n_13726) );
in01s01 FE_OCP_RBC5022_n_29080 ( .a(n_29080), .o(FE_OCP_RBN5022_n_29080) );
in01s02 FE_OCP_RBC5023_n_29080 ( .a(FE_OCP_RBN5022_n_29080), .o(FE_OCP_RBN5023_n_29080) );
in01s01 FE_OCP_RBC5024_n_29080 ( .a(FE_OCP_RBN5023_n_29080), .o(FE_OCP_RBN5024_n_29080) );
in01f02 FE_OCP_RBC5025_n_29053 ( .a(n_29053), .o(FE_OCP_RBN5025_n_29053) );
in01s01 FE_OCP_RBC5026_n_29053 ( .a(n_29053), .o(FE_OCP_RBN5026_n_29053) );
in01f02 FE_OCP_RBC5027_n_18515 ( .a(n_18515), .o(FE_OCP_RBN5027_n_18515) );
in01m01 FE_OCP_RBC5028_n_18515 ( .a(FE_OCP_RBN5027_n_18515), .o(FE_OCP_RBN5028_n_18515) );
in01s01 FE_OCP_RBC5029_n_18678 ( .a(n_18678), .o(FE_OCP_RBN5029_n_18678) );
in01s01 FE_OCP_RBC5030_n_18678 ( .a(n_18678), .o(FE_OCP_RBN5030_n_18678) );
in01s02 FE_OCP_RBC5031_n_18951 ( .a(n_18951), .o(FE_OCP_RBN5031_n_18951) );
in01s06 FE_OCP_RBC5032_n_18951 ( .a(n_18951), .o(FE_OCP_RBN5032_n_18951) );
in01m02 FE_OCP_RBC5033_n_18951 ( .a(n_18951), .o(FE_OCP_RBN5033_n_18951) );
in01m02 FE_OCP_RBC5034_n_19062 ( .a(n_19062), .o(FE_OCP_RBN5034_n_19062) );
in01s01 FE_OCP_RBC5035_n_19055 ( .a(n_19055), .o(FE_OCP_RBN5035_n_19055) );
in01s01 FE_OCP_RBC5037_n_13927 ( .a(n_13927), .o(FE_OCP_RBN5037_n_13927) );
in01f02 FE_OCP_RBC5038_n_13927 ( .a(n_13927), .o(FE_OCP_RBN5038_n_13927) );
in01s01 FE_OCP_RBC5039_n_13927 ( .a(FE_OCP_RBN5037_n_13927), .o(FE_OCP_RBN5039_n_13927) );
in01f08 FE_OCP_RBC5040_n_27827 ( .a(n_27827), .o(FE_OCP_RBN5040_n_27827) );
in01s02 FE_OCP_RBC5041_n_14201 ( .a(n_14201), .o(FE_OCP_RBN5041_n_14201) );
in01f01 FE_OCP_RBC5045_n_14450 ( .a(n_14450), .o(FE_OCP_RBN5045_n_14450) );
in01f01 FE_OCP_RBC5046_n_14450 ( .a(n_14450), .o(FE_OCP_RBN5046_n_14450) );
in01s03 FE_OCP_RBC5047_n_29648 ( .a(n_29648), .o(FE_OCP_RBN5047_n_29648) );
in01s04 FE_OCP_RBC5049_FE_RN_606_0 ( .a(FE_RN_606_0), .o(FE_OCP_RBN5049_FE_RN_606_0) );
in01m02 FE_OCP_RBC5050_FE_RN_606_0 ( .a(FE_RN_606_0), .o(FE_OCP_RBN5050_FE_RN_606_0) );
in01s01 FE_OCP_RBC5051_n_22709 ( .a(FE_OCP_RBN3456_n_22709), .o(FE_OCP_RBN5051_n_22709) );
in01f04 FE_OCP_RBC5053_n_32169 ( .a(n_32169), .o(FE_OCP_RBN5053_n_32169) );
in01m02 FE_OCP_RBC5055_n_32340 ( .a(n_32340), .o(FE_OCP_RBN5055_n_32340) );
in01s02 FE_OCP_RBC5058_n_32427 ( .a(n_32427), .o(FE_OCP_RBN5058_n_32427) );
in01s10 FE_OCP_RBC5175_n_44061 ( .a(FE_OCP_RBN6465_n_44061), .o(FE_OCP_RBN5175_n_44061) );
in01s20 FE_OCP_RBC5179_n_44061 ( .a(FE_OCP_RBN5180_n_44061), .o(FE_OCP_RBN5179_n_44061) );
in01s03 FE_OCP_RBC5180_n_44061 ( .a(n_44061), .o(FE_OCP_RBN5180_n_44061) );
in01s06 FE_OCP_RBC5181_n_44061 ( .a(FE_OCP_RBN5459_n_44061), .o(FE_OCP_RBN5181_n_44061) );
in01m04 FE_OCP_RBC5196_n_25893 ( .a(n_25893), .o(FE_OCP_RBN5196_n_25893) );
in01s01 FE_OCP_RBC5197_n_25893 ( .a(n_25893), .o(FE_OCP_RBN5197_n_25893) );
in01s01 FE_OCP_RBC5198_n_25893 ( .a(FE_OCP_RBN5197_n_25893), .o(FE_OCP_RBN5198_n_25893) );
in01s01 FE_OCP_RBC5199_n_25893 ( .a(FE_OCP_RBN5198_n_25893), .o(FE_OCP_RBN5199_n_25893) );
in01f02 FE_OCP_RBC5200_n_25729 ( .a(n_25729), .o(FE_OCP_RBN5200_n_25729) );
in01s01 FE_OCP_RBC5201_n_25729 ( .a(n_25729), .o(FE_OCP_RBN5201_n_25729) );
in01s01 FE_OCP_RBC5202_n_25729 ( .a(FE_OCP_RBN5201_n_25729), .o(FE_OCP_RBN5202_n_25729) );
in01s01 FE_OCP_RBC5203_n_25729 ( .a(FE_OCP_RBN5202_n_25729), .o(FE_OCP_RBN5203_n_25729) );
in01s01 FE_OCP_RBC5204_n_25729 ( .a(FE_OCP_RBN5203_n_25729), .o(FE_OCP_RBN5204_n_25729) );
in01s01 FE_OCP_RBC5205_n_20504 ( .a(n_20504), .o(FE_OCP_RBN5205_n_20504) );
in01s01 FE_OCP_RBC5206_n_20504 ( .a(FE_OCP_RBN5205_n_20504), .o(FE_OCP_RBN5206_n_20504) );
in01s01 FE_OCP_RBC5207_n_20504 ( .a(FE_OCP_RBN5206_n_20504), .o(FE_OCP_RBN5207_n_20504) );
in01f02 FE_OCP_RBC5208_n_20412 ( .a(n_20412), .o(FE_OCP_RBN5208_n_20412) );
in01s01 FE_OCP_RBC5209_n_20412 ( .a(n_20412), .o(FE_OCP_RBN5209_n_20412) );
in01s01 FE_OCP_RBC5210_n_20412 ( .a(FE_OCP_RBN5209_n_20412), .o(FE_OCP_RBN5210_n_20412) );
in01s01 FE_OCP_RBC5211_n_20412 ( .a(FE_OCP_RBN5210_n_20412), .o(FE_OCP_RBN5211_n_20412) );
in01m02 FE_OCP_RBC5212_n_21987 ( .a(n_21987), .o(FE_OCP_RBN5212_n_21987) );
in01f02 FE_OCP_RBC5213_n_29773 ( .a(n_29773), .o(FE_OCP_RBN5213_n_29773) );
in01m01 FE_OCP_RBC5214_n_22150 ( .a(n_22150), .o(FE_OCP_RBN5214_n_22150) );
in01m02 FE_OCP_RBC5215_n_22150 ( .a(FE_OCP_RBN5214_n_22150), .o(FE_OCP_RBN5215_n_22150) );
in01s02 FE_OCP_RBC5216_n_22212 ( .a(n_22212), .o(FE_OCP_RBN5216_n_22212) );
in01s01 FE_OCP_RBC5217_n_22212 ( .a(FE_OCP_RBN5216_n_22212), .o(FE_OCP_RBN5217_n_22212) );
in01s06 FE_OCP_RBC5322_n_16745 ( .a(n_16745), .o(FE_OCP_RBN5322_n_16745) );
in01m10 FE_OCP_RBC5323_n_27893 ( .a(n_27893), .o(FE_OCP_RBN5323_n_27893) );
in01f10 FE_OCP_RBC5324_n_27885 ( .a(n_27885), .o(FE_OCP_RBN5324_n_27885) );
in01s02 FE_OCP_RBC5325_n_18653 ( .a(n_18653), .o(FE_OCP_RBN5325_n_18653) );
in01m02 FE_OCP_RBC5326_n_29292 ( .a(n_29292), .o(FE_OCP_RBN5326_n_29292) );
in01f02 FE_OCP_RBC5327_FE_RN_2034_0 ( .a(FE_RN_2034_0), .o(FE_OCP_RBN5327_FE_RN_2034_0) );
in01m02 FE_OCP_RBC5328_n_15047 ( .a(n_15047), .o(FE_OCP_RBN5328_n_15047) );
in01s04 FE_OCP_RBC5329_n_15047 ( .a(n_15047), .o(FE_OCP_RBN5329_n_15047) );
in01f02 FE_OCP_RBC5330_n_20678 ( .a(n_20678), .o(FE_OCP_RBN5330_n_20678) );
in01f02 FE_OCP_RBC5331_n_20843 ( .a(n_20843), .o(FE_OCP_RBN5331_n_20843) );
in01s02 FE_OCP_RBC5333_FE_RN_1490_0 ( .a(FE_RN_1490_0), .o(FE_OCP_RBN5333_FE_RN_1490_0) );
in01m02 FE_OCP_RBC5334_FE_RN_1490_0 ( .a(FE_RN_1490_0), .o(FE_OCP_RBN5334_FE_RN_1490_0) );
in01m04 FE_OCP_RBC5335_FE_RN_1144_0 ( .a(FE_RN_1144_0), .o(FE_OCP_RBN5335_FE_RN_1144_0) );
in01f02 FE_OCP_RBC5336_n_30865 ( .a(n_30865), .o(FE_OCP_RBN5336_n_30865) );
in01m02 FE_OCP_RBC5337_FE_RN_2064_0 ( .a(FE_RN_2064_0), .o(FE_OCP_RBN5337_FE_RN_2064_0) );
in01m01 FE_OCP_RBC5338_FE_RN_2064_0 ( .a(FE_RN_2064_0), .o(FE_OCP_RBN5338_FE_RN_2064_0) );
in01m04 FE_OCP_RBC5340_n_21261 ( .a(n_21261), .o(FE_OCP_RBN5340_n_21261) );
in01m06 FE_OCP_RBC5341_n_22068 ( .a(n_22068), .o(FE_OCP_RBN5341_n_22068) );
in01m06 FE_OCP_RBC5342_n_22068 ( .a(FE_OCP_RBN5341_n_22068), .o(FE_OCP_RBN5342_n_22068) );
in01m06 FE_OCP_RBC5343_n_22068 ( .a(FE_OCP_RBN5341_n_22068), .o(FE_OCP_RBN5343_n_22068) );
in01f04 FE_OCP_RBC5344_n_22476 ( .a(FE_OCP_RBN1173_n_22476), .o(FE_OCP_RBN5344_n_22476) );
in01m02 FE_OCP_RBC5345_n_22476 ( .a(FE_OCP_RBN1173_n_22476), .o(FE_OCP_RBN5345_n_22476) );
in01s02 FE_OCP_RBC5346_n_22556 ( .a(n_22556), .o(FE_OCP_RBN5346_n_22556) );
in01m02 FE_OCP_RBC5347_n_22556 ( .a(n_22556), .o(FE_OCP_RBN5347_n_22556) );
in01s01 FE_OCP_RBC5348_FE_RN_627_0 ( .a(FE_RN_627_0), .o(FE_OCP_RBN5348_FE_RN_627_0) );
in01s01 FE_OCP_RBC5349_n_32518 ( .a(n_32518), .o(FE_OCP_RBN5349_n_32518) );
in01m02 FE_OCP_RBC5350_n_22818 ( .a(n_22818), .o(FE_OCP_RBN5350_n_22818) );
in01m02 FE_OCP_RBC5351_n_22903 ( .a(n_22903), .o(FE_OCP_RBN5351_n_22903) );
in01s01 FE_OCP_RBC5352_n_32516 ( .a(n_32516), .o(FE_OCP_RBN5352_n_32516) );
in01s01 FE_OCP_RBC5374_n_28186 ( .a(n_28186), .o(FE_OCP_RBN5374_n_28186) );
in01s03 FE_OCP_RBC5375_n_28123 ( .a(n_28123), .o(FE_OCP_RBN5375_n_28123) );
in01m08 FE_OCP_RBC5376_n_28123 ( .a(n_28123), .o(FE_OCP_RBN5376_n_28123) );
in01s02 FE_OCP_RBC5377_n_19055 ( .a(FE_OCP_RBN5035_n_19055), .o(FE_OCP_RBN5377_n_19055) );
in01s01 FE_OCP_RBC5378_n_19055 ( .a(FE_OCP_RBN5377_n_19055), .o(FE_OCP_RBN5378_n_19055) );
in01s01 FE_OCP_RBC5379_n_19055 ( .a(FE_OCP_RBN5378_n_19055), .o(FE_OCP_RBN5379_n_19055) );
in01f02 FE_OCP_RBC5380_n_19428 ( .a(n_19428), .o(FE_OCP_RBN5380_n_19428) );
in01m01 FE_OCP_RBC5381_n_20123 ( .a(n_20123), .o(FE_OCP_RBN5381_n_20123) );
in01s01 FE_OCP_RBC5382_n_20123 ( .a(n_20123), .o(FE_OCP_RBN5382_n_20123) );
in01s01 FE_OCP_RBC5386_n_20638 ( .a(n_20638), .o(FE_OCP_RBN5386_n_20638) );
in01s01 FE_OCP_RBC5387_n_22149 ( .a(n_22149), .o(FE_OCP_RBN5387_n_22149) );
in01s01 FE_OCP_RBC5388_n_22149 ( .a(FE_OCP_RBN5387_n_22149), .o(FE_OCP_RBN5388_n_22149) );
in01s01 FE_OCP_RBC5391_cordic_combinational_sub_ln23_0_unr12_z_0_ ( .a(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(FE_OCP_RBN5391_cordic_combinational_sub_ln23_0_unr12_z_0_) );
in01s01 FE_OCP_RBC5392_cordic_combinational_sub_ln23_0_unr12_z_0_ ( .a(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(FE_OCP_RBN5392_cordic_combinational_sub_ln23_0_unr12_z_0_) );
in01m06 FE_OCP_RBC5393_cordic_combinational_sub_ln23_0_unr12_z_0_ ( .a(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(FE_OCP_RBN5393_cordic_combinational_sub_ln23_0_unr12_z_0_) );
in01s01 FE_OCP_RBC5394_cordic_combinational_sub_ln23_0_unr12_z_0_ ( .a(FE_OCP_RBN5391_cordic_combinational_sub_ln23_0_unr12_z_0_), .o(FE_OCP_RBN5394_cordic_combinational_sub_ln23_0_unr12_z_0_) );
in01s01 FE_OCP_RBC5395_cordic_combinational_sub_ln23_0_unr12_z_0_ ( .a(FE_OCP_RBN5391_cordic_combinational_sub_ln23_0_unr12_z_0_), .o(FE_OCP_RBN5395_cordic_combinational_sub_ln23_0_unr12_z_0_) );
in01s01 FE_OCP_RBC5412_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN6516_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN5412_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s10 FE_OCP_RBC5434_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN5434_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01m01 FE_OCP_RBC5435_delay_xor_ln22_unr6_stage3_stallmux_q_0_ ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .o(FE_OCP_RBN5435_delay_xor_ln22_unr6_stage3_stallmux_q_0_) );
in01s02 FE_OCP_RBC5436_delay_xor_ln22_unr6_stage3_stallmux_q_0_ ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .o(FE_OCP_RBN5436_delay_xor_ln22_unr6_stage3_stallmux_q_0_) );
in01s01 FE_OCP_RBC5437_delay_xor_ln22_unr6_stage3_stallmux_q_0_ ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .o(FE_OCP_RBN5437_delay_xor_ln22_unr6_stage3_stallmux_q_0_) );
in01s10 FE_OCP_RBC5438_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_ ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .o(FE_OCP_RBN5438_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_) );
in01s10 FE_OCP_RBC5439_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_ ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .o(FE_OCP_RBN5439_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_) );
in01m06 FE_OCP_RBC5441_delay_sub_ln23_0_unr8_stage4_stallmux_q_2_ ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_2_), .o(FE_OCP_RBN5441_delay_sub_ln23_0_unr8_stage4_stallmux_q_2_) );
in01s10 FE_OCP_RBC5442_delay_sub_ln23_unr9_stage4_stallmux_q_3_ ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(FE_OCP_RBN5442_delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
in01s40 FE_OCP_RBC5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_ ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
in01s20 FE_OCP_RBC5445_delay_sub_ln23_unr9_stage4_stallmux_q_3_ ( .a(FE_OCP_RBN5442_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(FE_OCP_RBN5445_delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
in01s06 FE_OCP_RBC5459_n_44061 ( .a(n_44061), .o(FE_OCP_RBN5459_n_44061) );
in01s01 FE_OCP_RBC5465_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN5465_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s02 FE_OCP_RBC5466_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN5466_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s01 FE_OCP_RBC5467_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN5467_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01s06 FE_OCP_RBC5498_n_44610 ( .a(n_44610), .o(FE_OCP_RBN5498_n_44610) );
in01s01 FE_OCP_RBC5503_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN6438_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN5503_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01s01 FE_OCP_RBC5504_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN6438_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN5504_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01s03 FE_OCP_RBC5506_n_44061 ( .a(FE_OCP_RBN6464_n_44061), .o(FE_OCP_RBN5506_n_44061) );
in01s06 FE_OCP_RBC5507_n_44061 ( .a(FE_OCP_RBN5506_n_44061), .o(FE_OCP_RBN5507_n_44061) );
in01m10 FE_OCP_RBC5508_FE_RN_1997_0 ( .a(FE_RN_1997_0), .o(FE_OCP_RBN5508_FE_RN_1997_0) );
in01s02 FE_OCP_RBC5509_FE_RN_1997_0 ( .a(FE_RN_1997_0), .o(FE_OCP_RBN5509_FE_RN_1997_0) );
in01m08 FE_OCP_RBC5510_FE_RN_1997_0 ( .a(FE_OCP_RBN5508_FE_RN_1997_0), .o(FE_OCP_RBN5510_FE_RN_1997_0) );
in01s40 FE_OCP_RBC5511_n_44365 ( .a(FE_OCP_RBN7102_n_44365), .o(FE_OCP_RBN5511_n_44365) );
in01s40 FE_OCP_RBC5512_n_44365 ( .a(FE_OCP_RBN5511_n_44365), .o(FE_OCP_RBN5512_n_44365) );
in01s40 FE_OCP_RBC5513_n_44365 ( .a(FE_OCP_RBN5512_n_44365), .o(FE_OCP_RBN5513_n_44365) );
in01s06 FE_OCP_RBC5514_n_44365 ( .a(FE_OCP_RBN5512_n_44365), .o(FE_OCP_RBN5514_n_44365) );
in01s02 FE_OCP_RBC5515_n_1472 ( .a(n_1472), .o(FE_OCP_RBN5515_n_1472) );
in01s10 FE_OCP_RBC5516_n_32436 ( .a(FE_OCP_RBN3980_n_32436), .o(FE_OCP_RBN5516_n_32436) );
in01s10 FE_OCP_RBC5517_n_32436 ( .a(FE_OCP_RBN5516_n_32436), .o(FE_OCP_RBN5517_n_32436) );
in01s02 FE_OCP_RBC5518_n_32436 ( .a(FE_OCP_RBN5517_n_32436), .o(FE_OCP_RBN5518_n_32436) );
in01m06 FE_OCP_RBC5522_n_23078 ( .a(n_23078), .o(FE_OCP_RBN5522_n_23078) );
in01s10 FE_OCP_RBC5523_n_28058 ( .a(n_28058), .o(FE_OCP_RBN5523_n_28058) );
in01s10 FE_OCP_RBC5524_n_32752 ( .a(n_32752), .o(FE_OCP_RBN5524_n_32752) );
in01s01 FE_OCP_RBC5525_n_36921 ( .a(n_36921), .o(FE_OCP_RBN5525_n_36921) );
in01s10 FE_OCP_RBC5527_n_6760 ( .a(n_6760), .o(FE_OCP_RBN5527_n_6760) );
in01s20 FE_OCP_RBC5528_n_44061 ( .a(FE_OCP_RBN3967_n_44061), .o(FE_OCP_RBN5528_n_44061) );
in01s40 FE_OCP_RBC5529_n_44061 ( .a(FE_OCP_RBN3967_n_44061), .o(FE_OCP_RBN5529_n_44061) );
in01m10 FE_OCP_RBC5530_n_1541 ( .a(n_1541), .o(FE_OCP_RBN5530_n_1541) );
in01f08 FE_OCP_RBC5531_n_27941 ( .a(n_27941), .o(FE_OCP_RBN5531_n_27941) );
in01s10 FE_OCP_RBC5532_n_44083 ( .a(n_44083), .o(FE_OCP_RBN5532_n_44083) );
in01s40 FE_OCP_RBC5533_n_44083 ( .a(n_44083), .o(FE_OCP_RBN5533_n_44083) );
in01s10 FE_OCP_RBC5534_n_44083 ( .a(n_44083), .o(FE_OCP_RBN5534_n_44083) );
in01s10 FE_OCP_RBC5535_n_44083 ( .a(n_44083), .o(FE_OCP_RBN5535_n_44083) );
in01s06 FE_OCP_RBC5536_n_44083 ( .a(n_44083), .o(FE_OCP_RBN5536_n_44083) );
in01s80 FE_OCP_RBC5537_n_44083 ( .a(n_44083), .o(FE_OCP_RBN5537_n_44083) );
in01s06 FE_OCP_RBC5539_n_23307 ( .a(n_23307), .o(FE_OCP_RBN5539_n_23307) );
in01s06 FE_OCP_RBC5540_n_23307 ( .a(n_23307), .o(FE_OCP_RBN5540_n_23307) );
in01f06 FE_OCP_RBC5541_n_23044 ( .a(n_23044), .o(FE_OCP_RBN5541_n_23044) );
in01m03 FE_OCP_RBC5542_n_23044 ( .a(n_23044), .o(FE_OCP_RBN5542_n_23044) );
in01s03 FE_OCP_RBC5543_n_23044 ( .a(n_23044), .o(FE_OCP_RBN5543_n_23044) );
in01s06 FE_OCP_RBC5544_n_45145 ( .a(n_45145), .o(FE_OCP_RBN5544_n_45145) );
in01m10 FE_OCP_RBC5545_n_45145 ( .a(n_45145), .o(FE_OCP_RBN5545_n_45145) );
in01s20 FE_OCP_RBC5546_n_45145 ( .a(n_45145), .o(FE_OCP_RBN5546_n_45145) );
in01s02 FE_OCP_RBC5547_n_1733 ( .a(n_1733), .o(FE_OCP_RBN5547_n_1733) );
in01s02 FE_OCP_RBC5548_FE_OCPN4833_n_32863 ( .a(FE_OCPN4833_n_32863), .o(FE_OCP_RBN5548_FE_OCPN4833_n_32863) );
in01s10 FE_OCP_RBC5549_n_28319 ( .a(n_28319), .o(FE_OCP_RBN5549_n_28319) );
in01s10 FE_OCP_RBC5550_n_17914 ( .a(n_17914), .o(FE_OCP_RBN5550_n_17914) );
in01s01 FE_OCP_RBC5551_n_17914 ( .a(n_17914), .o(FE_OCP_RBN5551_n_17914) );
in01f10 FE_OCP_RBC5552_n_23328 ( .a(n_23328), .o(FE_OCP_RBN5552_n_23328) );
in01s01 FE_OCP_RBC5553_n_1812 ( .a(n_1812), .o(FE_OCP_RBN5553_n_1812) );
in01s01 FE_OCP_RBC5554_n_1822 ( .a(n_1822), .o(FE_OCP_RBN5554_n_1822) );
in01s01 FE_OCP_RBC5555_n_1827 ( .a(n_1827), .o(FE_OCP_RBN5555_n_1827) );
in01s01 FE_OCP_RBC5556_n_37559 ( .a(n_37559), .o(FE_OCP_RBN5556_n_37559) );
in01m02 FE_OCP_RBC5557_n_37559 ( .a(n_37559), .o(FE_OCP_RBN5557_n_37559) );
in01f02 FE_OCP_RBC5558_n_37559 ( .a(n_37559), .o(FE_OCP_RBN5558_n_37559) );
in01s01 FE_OCP_RBC5559_n_1853 ( .a(n_1853), .o(FE_OCP_RBN5559_n_1853) );
in01s01 FE_OCP_RBC5560_n_1889 ( .a(n_1889), .o(FE_OCP_RBN5560_n_1889) );
in01s01 FE_OCP_RBC5561_n_33097 ( .a(n_33097), .o(FE_OCP_RBN5561_n_33097) );
in01s04 FE_OCP_RBC5562_n_33097 ( .a(n_33097), .o(FE_OCP_RBN5562_n_33097) );
in01s01 FE_OCP_RBC5563_n_37551 ( .a(n_37551), .o(FE_OCP_RBN5563_n_37551) );
in01s01 FE_OCP_RBC5564_n_37551 ( .a(n_37551), .o(FE_OCP_RBN5564_n_37551) );
in01s02 FE_OCP_RBC5565_n_2346 ( .a(n_2346), .o(FE_OCP_RBN5565_n_2346) );
in01s02 FE_OCP_RBC5566_n_2346 ( .a(FE_OCP_RBN5565_n_2346), .o(FE_OCP_RBN5566_n_2346) );
in01s02 FE_OCP_RBC5567_n_2346 ( .a(FE_OCP_RBN5565_n_2346), .o(FE_OCP_RBN5567_n_2346) );
in01m06 FE_OCP_RBC5568_n_2103 ( .a(n_2103), .o(FE_OCP_RBN5568_n_2103) );
in01s01 FE_OCP_RBC5569_n_2103 ( .a(n_2103), .o(FE_OCP_RBN5569_n_2103) );
in01s01 FE_OCP_RBC5574_n_12727 ( .a(n_12727), .o(FE_OCP_RBN5574_n_12727) );
in01m01 FE_OCP_RBC5575_n_12727 ( .a(n_12727), .o(FE_OCP_RBN5575_n_12727) );
in01m02 FE_OCP_RBC5576_n_12727 ( .a(FE_OCP_RBN5575_n_12727), .o(FE_OCP_RBN5576_n_12727) );
in01s10 FE_OCP_RBC5578_n_12753 ( .a(FE_OCP_RBN6564_n_12753), .o(FE_OCP_RBN5578_n_12753) );
in01s01 FE_OCP_RBC5580_n_12753 ( .a(FE_OCP_RBN6565_n_12753), .o(FE_OCP_RBN5580_n_12753) );
in01s08 FE_OCP_RBC5581_n_12753 ( .a(FE_OCP_RBN6565_n_12753), .o(FE_OCP_RBN5581_n_12753) );
in01m01 FE_OCP_RBC5582_n_12802 ( .a(n_12802), .o(FE_OCP_RBN5582_n_12802) );
in01m01 FE_OCP_RBC5583_n_12802 ( .a(n_12802), .o(FE_OCP_RBN5583_n_12802) );
in01m02 FE_OCP_RBC5584_n_12802 ( .a(FE_OCP_RBN5583_n_12802), .o(FE_OCP_RBN5584_n_12802) );
in01s04 FE_OCP_RBC5585_n_33368 ( .a(n_33368), .o(FE_OCP_RBN5585_n_33368) );
in01s03 FE_OCP_RBC5587_FE_RN_1367_0 ( .a(FE_OCP_RBN2490_FE_RN_1367_0), .o(FE_OCP_RBN5587_FE_RN_1367_0) );
in01s03 FE_OCP_RBC5588_FE_RN_1367_0 ( .a(FE_OCP_RBN5587_FE_RN_1367_0), .o(FE_OCP_RBN5588_FE_RN_1367_0) );
in01s01 FE_OCP_RBC5589_FE_RN_1367_0 ( .a(FE_OCP_RBN5587_FE_RN_1367_0), .o(FE_OCP_RBN5589_FE_RN_1367_0) );
in01s03 FE_OCP_RBC5590_FE_RN_1367_0 ( .a(FE_OCP_RBN5588_FE_RN_1367_0), .o(FE_OCP_RBN5590_FE_RN_1367_0) );
in01s01 FE_OCP_RBC5591_FE_RN_1367_0 ( .a(FE_OCP_RBN5589_FE_RN_1367_0), .o(FE_OCP_RBN5591_FE_RN_1367_0) );
in01s01 FE_OCP_RBC5592_FE_RN_1367_0 ( .a(FE_OCP_RBN5590_FE_RN_1367_0), .o(FE_OCP_RBN5592_FE_RN_1367_0) );
in01s02 FE_OCP_RBC5593_FE_RN_1367_0 ( .a(FE_OCP_RBN5592_FE_RN_1367_0), .o(FE_OCP_RBN5593_FE_RN_1367_0) );
in01s01 FE_OCP_RBC5594_n_45903 ( .a(n_45903), .o(FE_OCP_RBN5594_n_45903) );
in01s04 FE_OCP_RBC5595_n_45903 ( .a(n_45903), .o(FE_OCP_RBN5595_n_45903) );
in01m10 FE_OCP_RBC5596_n_45903 ( .a(n_45903), .o(FE_OCP_RBN5596_n_45903) );
in01m10 FE_OCP_RBC5597_n_45903 ( .a(FE_OCP_RBN5596_n_45903), .o(FE_OCP_RBN5597_n_45903) );
in01s01 FE_OCP_RBC5598_n_2100 ( .a(n_2100), .o(FE_OCP_RBN5598_n_2100) );
in01s02 FE_OCP_RBC5599_n_2100 ( .a(n_2100), .o(FE_OCP_RBN5599_n_2100) );
in01s10 FE_OCP_RBC5600_n_44875 ( .a(n_44875), .o(FE_OCP_RBN5600_n_44875) );
in01s01 FE_OCP_RBC5603_n_29056 ( .a(FE_OCP_RBN4900_n_29056), .o(FE_OCP_RBN5603_n_29056) );
in01f02 FE_OCP_RBC5604_n_29056 ( .a(FE_OCP_RBN4900_n_29056), .o(FE_OCP_RBN5604_n_29056) );
in01s02 FE_OCP_RBC5605_n_2430 ( .a(n_2430), .o(FE_OCP_RBN5605_n_2430) );
in01s01 FE_OCP_RBC5606_n_7730 ( .a(n_7730), .o(FE_OCP_RBN5606_n_7730) );
in01s10 FE_OCP_RBC5607_n_7730 ( .a(n_7730), .o(FE_OCP_RBN5607_n_7730) );
in01s02 FE_OCP_RBC5608_n_7730 ( .a(n_7730), .o(FE_OCP_RBN5608_n_7730) );
in01s01 FE_OCP_RBC5609_n_7730 ( .a(FE_OCP_RBN5607_n_7730), .o(FE_OCP_RBN5609_n_7730) );
in01s01 FE_OCP_RBC5610_n_7730 ( .a(FE_OCP_RBN5607_n_7730), .o(FE_OCP_RBN5610_n_7730) );
in01s01 FE_OCP_RBC5611_n_7730 ( .a(FE_OCP_RBN5607_n_7730), .o(FE_OCP_RBN5611_n_7730) );
in01s06 FE_OCP_RBC5612_n_7730 ( .a(FE_OCP_RBN5607_n_7730), .o(FE_OCP_RBN5612_n_7730) );
in01s01 FE_OCP_RBC5613_n_7730 ( .a(FE_OCP_RBN5608_n_7730), .o(FE_OCP_RBN5613_n_7730) );
in01s01 FE_OCP_RBC5614_n_7730 ( .a(FE_OCP_RBN5611_n_7730), .o(FE_OCP_RBN5614_n_7730) );
in01s01 FE_OCP_RBC5615_n_24070 ( .a(n_24070), .o(FE_OCP_RBN5615_n_24070) );
in01s01 FE_OCP_RBC5617_n_18899 ( .a(FE_OCP_RBN4081_n_18899), .o(FE_OCP_RBN5617_n_18899) );
in01s01 FE_OCP_RBC5618_n_18899 ( .a(FE_OCP_RBN4081_n_18899), .o(FE_OCP_RBN5618_n_18899) );
in01s01 FE_OCP_RBC5620_n_18986 ( .a(n_18986), .o(FE_OCP_RBN5620_n_18986) );
in01s04 FE_OCP_RBC5621_n_18986 ( .a(n_18986), .o(FE_OCP_RBN5621_n_18986) );
in01s01 FE_OCP_RBC5622_n_18986 ( .a(FE_OCP_RBN5621_n_18986), .o(FE_OCP_RBN5622_n_18986) );
in01s01 FE_OCP_RBC5625_n_2457 ( .a(n_2457), .o(FE_OCP_RBN5625_n_2457) );
in01s01 FE_OCP_RBC5626_n_2457 ( .a(n_2457), .o(FE_OCP_RBN5626_n_2457) );
in01s02 FE_OCP_RBC5627_n_33976 ( .a(n_33976), .o(FE_OCP_RBN5627_n_33976) );
in01s01 FE_OCP_RBC5628_n_33976 ( .a(FE_OCP_RBN5627_n_33976), .o(FE_OCP_RBN5628_n_33976) );
in01s01 FE_OCP_RBC5629_n_33976 ( .a(FE_OCP_RBN5628_n_33976), .o(FE_OCP_RBN5629_n_33976) );
in01m02 FE_OCP_RBC5630_n_33957 ( .a(n_33957), .o(FE_OCP_RBN5630_n_33957) );
in01s06 FE_OCP_RBC5632_n_7708 ( .a(FE_OCP_RBN6600_n_7708), .o(FE_OCP_RBN5632_n_7708) );
in01s06 FE_OCP_RBC5633_n_7708 ( .a(FE_OCP_RBN5632_n_7708), .o(FE_OCP_RBN5633_n_7708) );
in01s06 FE_OCP_RBC5634_n_7708 ( .a(FE_OCP_RBN5633_n_7708), .o(FE_OCP_RBN5634_n_7708) );
in01s01 FE_OCP_RBC5635_n_7708 ( .a(FE_OCP_RBN5633_n_7708), .o(FE_OCP_RBN5635_n_7708) );
in01s01 FE_OCP_RBC5636_n_7708 ( .a(FE_OCP_RBN5633_n_7708), .o(FE_OCP_RBN5636_n_7708) );
in01s10 FE_OCP_RBC5637_n_41381 ( .a(FE_OCP_RBN4115_n_41381), .o(FE_OCP_RBN5637_n_41381) );
in01s20 FE_OCP_RBC5638_n_41381 ( .a(FE_OCP_RBN5637_n_41381), .o(FE_OCP_RBN5638_n_41381) );
in01s02 FE_OCP_RBC5639_n_41381 ( .a(FE_OCP_RBN5637_n_41381), .o(FE_OCP_RBN5639_n_41381) );
in01m02 FE_OCP_RBC5640_n_19060 ( .a(n_19060), .o(FE_OCP_RBN5640_n_19060) );
in01m06 FE_OCP_RBC5643_n_33977 ( .a(n_33977), .o(FE_OCP_RBN5643_n_33977) );
in01s01 FE_OCP_RBC5644_n_2674 ( .a(n_2674), .o(FE_OCP_RBN5644_n_2674) );
in01s02 FE_OCP_RBC5645_n_29236 ( .a(n_29236), .o(FE_OCP_RBN5645_n_29236) );
in01f04 FE_OCP_RBC5646_n_33785 ( .a(n_33785), .o(FE_OCP_RBN5646_n_33785) );
in01s01 FE_OCP_RBC5647_FE_OCPN855_n_7721 ( .a(FE_OCP_RBN2604_FE_OCPN855_n_7721), .o(FE_OCP_RBN5647_FE_OCPN855_n_7721) );
in01s06 FE_OCP_RBC5648_n_2438 ( .a(FE_OCP_RBN6611_n_2289), .o(FE_OCP_RBN5648_n_2438) );
in01s04 FE_OCP_RBC5649_n_2438 ( .a(FE_OCP_RBN6611_n_2289), .o(FE_OCP_RBN5649_n_2438) );
in01s01 FE_OCP_RBC5650_n_2438 ( .a(FE_OCP_RBN5648_n_2438), .o(FE_OCP_RBN5650_n_2438) );
in01s01 FE_OCP_RBC5651_n_2438 ( .a(FE_OCP_RBN5649_n_2438), .o(FE_OCP_RBN5651_n_2438) );
in01s02 FE_OCP_RBC5652_n_2438 ( .a(FE_OCP_RBN5649_n_2438), .o(FE_OCP_RBN5652_n_2438) );
in01s02 FE_OCP_RBC5653_n_2438 ( .a(FE_OCP_RBN5649_n_2438), .o(FE_OCP_RBN5653_n_2438) );
in01s01 FE_OCP_RBC5654_n_2438 ( .a(FE_OCP_RBN5650_n_2438), .o(FE_OCP_RBN5654_n_2438) );
in01m01 FE_OCP_RBC5655_n_2438 ( .a(FE_OCP_RBN5650_n_2438), .o(FE_OCP_RBN5655_n_2438) );
in01s01 FE_OCP_RBC5656_n_2438 ( .a(FE_OCP_RBN5651_n_2438), .o(FE_OCP_RBN5656_n_2438) );
in01s01 FE_OCP_RBC5657_n_2438 ( .a(FE_OCP_RBN5651_n_2438), .o(FE_OCP_RBN5657_n_2438) );
in01s01 FE_OCP_RBC5658_n_2438 ( .a(FE_OCP_RBN5652_n_2438), .o(FE_OCP_RBN5658_n_2438) );
in01m01 FE_OCP_RBC5659_n_2438 ( .a(FE_OCP_RBN5655_n_2438), .o(FE_OCP_RBN5659_n_2438) );
in01s01 FE_OCP_RBC5660_n_2438 ( .a(FE_OCP_RBN5656_n_2438), .o(FE_OCP_RBN5660_n_2438) );
in01s01 FE_OCP_RBC5661_n_2438 ( .a(FE_OCP_RBN5658_n_2438), .o(FE_OCP_RBN5661_n_2438) );
in01s01 FE_OCP_RBC5662_n_2438 ( .a(FE_OCP_RBN6611_n_2289), .o(FE_OCP_RBN5662_n_2438) );
in01s01 FE_OCP_RBC5663_n_2438 ( .a(FE_OCP_RBN6611_n_2289), .o(FE_OCP_RBN5663_n_2438) );
in01s02 FE_OCP_RBC5664_n_13757 ( .a(n_13757), .o(FE_OCP_RBN5664_n_13757) );
in01m06 FE_OCP_RBC5665_n_19101 ( .a(n_19101), .o(FE_OCP_RBN5665_n_19101) );
in01s01 FE_OCP_RBC5666_n_19101 ( .a(FE_OCP_RBN5665_n_19101), .o(FE_OCP_RBN5666_n_19101) );
in01s01 FE_OCP_RBC5667_n_19101 ( .a(FE_OCP_RBN5666_n_19101), .o(FE_OCP_RBN5667_n_19101) );
in01s01 FE_OCP_RBC5668_n_19101 ( .a(FE_OCP_RBN5666_n_19101), .o(FE_OCP_RBN5668_n_19101) );
in01s01 FE_OCP_RBC5669_n_19101 ( .a(FE_OCP_RBN5666_n_19101), .o(FE_OCP_RBN5669_n_19101) );
in01s01 FE_OCP_RBC5670_n_24288 ( .a(n_24288), .o(FE_OCP_RBN5670_n_24288) );
in01s01 FE_OCP_RBC5671_n_24288 ( .a(n_24288), .o(FE_OCP_RBN5671_n_24288) );
in01m02 FE_OCP_RBC5672_n_29425 ( .a(n_29425), .o(FE_OCP_RBN5672_n_29425) );
in01m20 FE_OCP_RBC5673_n_41420 ( .a(n_41420), .o(FE_OCP_RBN5673_n_41420) );
in01s20 FE_OCP_RBC5674_n_41420 ( .a(n_41420), .o(FE_OCP_RBN5674_n_41420) );
in01m06 FE_OCP_RBC5675_n_41420 ( .a(FE_OCP_RBN5673_n_41420), .o(FE_OCP_RBN5675_n_41420) );
in01s10 FE_OCP_RBC5676_n_41420 ( .a(FE_OCP_RBN5675_n_41420), .o(FE_OCP_RBN5676_n_41420) );
in01s03 FE_OCP_RBC5677_n_19177 ( .a(n_19177), .o(FE_OCP_RBN5677_n_19177) );
in01s02 FE_OCP_RBC5678_n_19177 ( .a(FE_OCP_RBN5677_n_19177), .o(FE_OCP_RBN5678_n_19177) );
in01s01 FE_OCP_RBC5679_n_19177 ( .a(FE_OCP_RBN5678_n_19177), .o(FE_OCP_RBN5679_n_19177) );
in01s01 FE_OCP_RBC5680_n_19177 ( .a(FE_OCP_RBN5678_n_19177), .o(FE_OCP_RBN5680_n_19177) );
in01s02 FE_OCP_RBC5681_n_19177 ( .a(FE_OCP_RBN5678_n_19177), .o(FE_OCP_RBN5681_n_19177) );
in01s01 FE_OCP_RBC5682_n_19177 ( .a(FE_OCP_RBN5678_n_19177), .o(FE_OCP_RBN5682_n_19177) );
in01m06 FE_OCP_RBC5683_n_38474 ( .a(n_38474), .o(FE_OCP_RBN5683_n_38474) );
in01s02 FE_OCP_RBC5684_FE_RN_308_0 ( .a(FE_RN_308_0), .o(FE_OCP_RBN5684_FE_RN_308_0) );
in01s01 FE_OCP_RBC5685_FE_RN_308_0 ( .a(FE_RN_308_0), .o(FE_OCP_RBN5685_FE_RN_308_0) );
in01f04 FE_OCP_RBC5686_FE_RN_308_0 ( .a(FE_RN_308_0), .o(FE_OCP_RBN5686_FE_RN_308_0) );
in01f02 FE_OCP_RBC5687_n_24259 ( .a(n_24259), .o(FE_OCP_RBN5687_n_24259) );
in01s01 FE_OCP_RBC5688_n_24259 ( .a(FE_OCP_RBN5687_n_24259), .o(FE_OCP_RBN5688_n_24259) );
in01m03 FE_OCP_RBC5689_n_38531 ( .a(n_38531), .o(FE_OCP_RBN5689_n_38531) );
in01f02 FE_OCP_RBC5690_n_38515 ( .a(n_38515), .o(FE_OCP_RBN5690_n_38515) );
in01s01 FE_OCP_RBC5691_n_2884 ( .a(n_2884), .o(FE_OCP_RBN5691_n_2884) );
in01m04 FE_OCP_RBC5692_n_2884 ( .a(n_2884), .o(FE_OCP_RBN5692_n_2884) );
in01s01 FE_OCP_RBC5693_n_8138 ( .a(n_8138), .o(FE_OCP_RBN5693_n_8138) );
in01s01 FE_OCP_RBC5695_n_8342 ( .a(FE_OCP_RBN6644_n_8342), .o(FE_OCP_RBN5695_n_8342) );
in01s01 FE_OCP_RBC5697_n_8342 ( .a(FE_OCP_RBN5695_n_8342), .o(FE_OCP_RBN5697_n_8342) );
in01s02 FE_OCP_RBC5698_n_38577 ( .a(n_38577), .o(FE_OCP_RBN5698_n_38577) );
in01f04 FE_OCP_RBC5699_n_42038 ( .a(n_42038), .o(FE_OCP_RBN5699_n_42038) );
in01s01 FE_OCP_RBC5700_n_45828 ( .a(n_45828), .o(FE_OCP_RBN5700_n_45828) );
in01m02 FE_OCP_RBC5701_n_13954 ( .a(n_13954), .o(FE_OCP_RBN5701_n_13954) );
in01m04 FE_OCP_RBC5702_n_29568 ( .a(n_29568), .o(FE_OCP_RBN5702_n_29568) );
in01m02 FE_OCP_RBC5703_n_19663 ( .a(n_19663), .o(FE_OCP_RBN5703_n_19663) );
in01s01 FE_OCP_RBC5704_n_19663 ( .a(n_19663), .o(FE_OCP_RBN5704_n_19663) );
in01s01 FE_OCP_RBC5705_n_19663 ( .a(FE_OCP_RBN5704_n_19663), .o(FE_OCP_RBN5705_n_19663) );
in01s02 FE_OCP_RBC5706_n_24451 ( .a(n_24451), .o(FE_OCP_RBN5706_n_24451) );
in01s01 FE_OCP_RBC5707_n_24451 ( .a(FE_OCP_RBN5706_n_24451), .o(FE_OCP_RBN5707_n_24451) );
in01s01 FE_OCP_RBC5708_n_3055 ( .a(n_3055), .o(FE_OCP_RBN5708_n_3055) );
in01s02 FE_OCP_RBC5709_n_3055 ( .a(n_3055), .o(FE_OCP_RBN5709_n_3055) );
in01s02 FE_OCP_RBC5710_n_13984 ( .a(n_13984), .o(FE_OCP_RBN5710_n_13984) );
in01s01 FE_OCP_RBC5711_n_13984 ( .a(FE_OCP_RBN5710_n_13984), .o(FE_OCP_RBN5711_n_13984) );
in01s06 FE_OCP_RBC5712_n_44102 ( .a(n_44102), .o(FE_OCP_RBN5712_n_44102) );
in01m10 FE_OCP_RBC5713_n_44102 ( .a(n_44102), .o(FE_OCP_RBN5713_n_44102) );
in01s10 FE_OCP_RBC5714_n_44102 ( .a(n_44102), .o(FE_OCP_RBN5714_n_44102) );
in01s01 FE_OCP_RBC5715_n_44102 ( .a(n_44102), .o(FE_OCP_RBN5715_n_44102) );
in01s02 FE_OCP_RBC5716_n_8523 ( .a(n_8523), .o(FE_OCP_RBN5716_n_8523) );
in01m04 FE_OCP_RBC5717_n_24718 ( .a(n_24718), .o(FE_OCP_RBN5717_n_24718) );
in01s01 FE_OCP_RBC5718_n_24718 ( .a(n_24718), .o(FE_OCP_RBN5718_n_24718) );
in01s02 FE_OCP_RBC5719_n_29624 ( .a(n_29624), .o(FE_OCP_RBN5719_n_29624) );
in01s02 FE_OCP_RBC5720_n_29624 ( .a(n_29624), .o(FE_OCP_RBN5720_n_29624) );
in01m04 FE_OCP_RBC5721_n_24506 ( .a(n_24506), .o(FE_OCP_RBN5721_n_24506) );
in01s01 FE_OCP_RBC5722_n_24506 ( .a(n_24506), .o(FE_OCP_RBN5722_n_24506) );
in01s02 FE_OCP_RBC5723_n_47022 ( .a(n_47022), .o(FE_OCP_RBN5723_n_47022) );
in01s01 FE_OCP_RBC5724_n_47022 ( .a(FE_OCP_RBN5723_n_47022), .o(FE_OCP_RBN5724_n_47022) );
in01m02 FE_OCP_RBC5725_n_14120 ( .a(FE_OCP_RBN2071_n_14120), .o(FE_OCP_RBN5725_n_14120) );
in01s01 FE_OCP_RBC5726_n_14120 ( .a(FE_OCP_RBN5725_n_14120), .o(FE_OCP_RBN5726_n_14120) );
in01s01 FE_OCP_RBC5727_n_14120 ( .a(FE_OCP_RBN5726_n_14120), .o(FE_OCP_RBN5727_n_14120) );
in01s01 FE_OCP_RBC5728_n_14120 ( .a(FE_OCP_RBN5726_n_14120), .o(FE_OCP_RBN5728_n_14120) );
in01s02 FE_OCP_RBC5729_n_4211 ( .a(n_4211), .o(FE_OCP_RBN5729_n_4211) );
in01s01 FE_OCP_RBC5730_n_4211 ( .a(n_4211), .o(FE_OCP_RBN5730_n_4211) );
in01s01 FE_OCP_RBC5731_n_4211 ( .a(FE_OCP_RBN5730_n_4211), .o(FE_OCP_RBN5731_n_4211) );
in01s02 FE_OCP_RBC5732_n_19806 ( .a(n_19806), .o(FE_OCP_RBN5732_n_19806) );
in01s02 FE_OCP_RBC5733_n_19806 ( .a(n_19806), .o(FE_OCP_RBN5733_n_19806) );
in01s02 FE_OCP_RBC5734_n_8548 ( .a(n_8548), .o(FE_OCP_RBN5734_n_8548) );
in01f02 FE_OCP_RBC5735_n_38569 ( .a(n_38569), .o(FE_OCP_RBN5735_n_38569) );
in01s01 FE_OCP_RBC5736_n_38569 ( .a(n_38569), .o(FE_OCP_RBN5736_n_38569) );
in01s01 FE_OCP_RBC5737_n_8402 ( .a(FE_OCP_RBN2735_n_8402), .o(FE_OCP_RBN5737_n_8402) );
in01s01 FE_OCP_RBC5738_n_8402 ( .a(FE_OCP_RBN5737_n_8402), .o(FE_OCP_RBN5738_n_8402) );
in01s01 FE_OCP_RBC5739_n_8402 ( .a(FE_OCP_RBN5737_n_8402), .o(FE_OCP_RBN5739_n_8402) );
in01s01 FE_OCP_RBC5740_n_4336 ( .a(n_4336), .o(FE_OCP_RBN5740_n_4336) );
in01s01 FE_OCP_RBC5741_n_4336 ( .a(n_4336), .o(FE_OCP_RBN5741_n_4336) );
in01s02 FE_OCP_RBC5742_n_8540 ( .a(n_8540), .o(FE_OCP_RBN5742_n_8540) );
in01s02 FE_OCP_RBC5743_n_34278 ( .a(n_34278), .o(FE_OCP_RBN5743_n_34278) );
in01m02 FE_OCP_RBC5744_n_42043 ( .a(n_42043), .o(FE_OCP_RBN5744_n_42043) );
in01s02 FE_OCP_RBC5745_n_24618 ( .a(n_24618), .o(FE_OCP_RBN5745_n_24618) );
in01m02 FE_OCP_RBC5746_n_8637 ( .a(n_8637), .o(FE_OCP_RBN5746_n_8637) );
in01s01 FE_OCP_RBC5747_n_8637 ( .a(FE_OCP_RBN5746_n_8637), .o(FE_OCP_RBN5747_n_8637) );
in01s01 FE_OCP_RBC5748_n_8637 ( .a(FE_OCP_RBN5747_n_8637), .o(FE_OCP_RBN5748_n_8637) );
in01m02 FE_OCP_RBC5749_n_8599 ( .a(n_8599), .o(FE_OCP_RBN5749_n_8599) );
in01s01 FE_OCP_RBC5750_n_8599 ( .a(n_8599), .o(FE_OCP_RBN5750_n_8599) );
in01s01 FE_OCP_RBC5751_n_4022 ( .a(n_4022), .o(FE_OCP_RBN5751_n_4022) );
in01s02 FE_OCP_RBC5752_n_4022 ( .a(n_4022), .o(FE_OCP_RBN5752_n_4022) );
in01s01 FE_OCP_RBC5753_n_4022 ( .a(n_4022), .o(FE_OCP_RBN5753_n_4022) );
in01s01 FE_OCP_RBC5754_n_4022 ( .a(FE_OCP_RBN5751_n_4022), .o(FE_OCP_RBN5754_n_4022) );
in01s01 FE_OCP_RBC5756_n_34307 ( .a(n_34307), .o(FE_OCP_RBN5756_n_34307) );
in01m02 FE_OCP_RBC5757_n_14444 ( .a(n_14444), .o(FE_OCP_RBN5757_n_14444) );
in01s01 FE_OCP_RBC5758_n_14444 ( .a(n_14444), .o(FE_OCP_RBN5758_n_14444) );
in01s01 FE_OCP_RBC5759_n_14444 ( .a(FE_OCP_RBN5758_n_14444), .o(FE_OCP_RBN5759_n_14444) );
in01s01 FE_OCP_RBC5760_n_14444 ( .a(FE_OCP_RBN5758_n_14444), .o(FE_OCP_RBN5760_n_14444) );
in01s01 FE_OCP_RBC5762_n_19884 ( .a(n_19884), .o(FE_OCP_RBN5762_n_19884) );
in01m04 FE_OCP_RBC5763_n_19884 ( .a(n_19884), .o(FE_OCP_RBN5763_n_19884) );
in01m06 FE_OCP_RBC5764_n_19884 ( .a(FE_OCP_RBN5763_n_19884), .o(FE_OCP_RBN5764_n_19884) );
in01s01 FE_OCP_RBC5767_n_3498 ( .a(FE_OCP_RBN6688_n_3498), .o(FE_OCP_RBN5767_n_3498) );
in01s01 FE_OCP_RBC5768_n_3498 ( .a(FE_OCP_RBN6688_n_3498), .o(FE_OCP_RBN5768_n_3498) );
in01s01 FE_OCP_RBC5769_n_3338 ( .a(n_3338), .o(FE_OCP_RBN5769_n_3338) );
in01s01 FE_OCP_RBC5770_n_3338 ( .a(FE_OCP_RBN5769_n_3338), .o(FE_OCP_RBN5770_n_3338) );
in01s01 FE_OCP_RBC5771_n_3338 ( .a(FE_OCP_RBN5770_n_3338), .o(FE_OCP_RBN5771_n_3338) );
in01m04 FE_OCP_RBC5772_n_34375 ( .a(n_34375), .o(FE_OCP_RBN5772_n_34375) );
in01m01 FE_OCP_RBC5773_n_34375 ( .a(n_34375), .o(FE_OCP_RBN5773_n_34375) );
in01s02 FE_OCP_RBC5774_n_13796 ( .a(FE_OCP_RBN4203_n_13796), .o(FE_OCP_RBN5774_n_13796) );
in01s06 FE_OCP_RBC5776_n_13796 ( .a(FE_OCP_RBN6692_n_13796), .o(FE_OCP_RBN5776_n_13796) );
in01s01 FE_OCP_RBC5777_n_13796 ( .a(FE_OCP_RBN6692_n_13796), .o(FE_OCP_RBN5777_n_13796) );
in01s01 FE_OCP_RBC5779_n_44570 ( .a(n_44570), .o(FE_OCP_RBN5779_n_44570) );
in01s01 FE_OCP_RBC5780_n_44570 ( .a(n_44570), .o(FE_OCP_RBN5780_n_44570) );
in01s10 FE_OCP_RBC5781_n_44570 ( .a(n_44570), .o(FE_OCP_RBN5781_n_44570) );
in01m02 FE_OCP_RBC5784_n_8657 ( .a(n_8657), .o(FE_OCP_RBN5784_n_8657) );
in01s01 FE_OCP_RBC5785_n_30071 ( .a(n_30071), .o(FE_OCP_RBN5785_n_30071) );
in01s01 FE_OCP_RBC5786_n_3421 ( .a(n_3421), .o(FE_OCP_RBN5786_n_3421) );
in01s01 FE_OCP_RBC5787_n_3421 ( .a(n_3421), .o(FE_OCP_RBN5787_n_3421) );
in01s01 FE_OCP_RBC5790_n_13962 ( .a(FE_OCP_RBN6698_n_13796), .o(FE_OCP_RBN5790_n_13962) );
in01s01 FE_OCP_RBC5791_n_13962 ( .a(FE_OCP_RBN6698_n_13796), .o(FE_OCP_RBN5791_n_13962) );
in01s01 FE_OCP_RBC5792_n_13962 ( .a(FE_OCP_RBN6696_n_13796), .o(FE_OCP_RBN5792_n_13962) );
in01s01 FE_OCP_RBC5793_n_13962 ( .a(FE_OCP_RBN6696_n_13796), .o(FE_OCP_RBN5793_n_13962) );
in01s01 FE_OCP_RBC5794_n_13962 ( .a(FE_OCP_RBN5790_n_13962), .o(FE_OCP_RBN5794_n_13962) );
in01s01 FE_OCP_RBC5795_n_13962 ( .a(FE_OCP_RBN5792_n_13962), .o(FE_OCP_RBN5795_n_13962) );
in01s01 FE_OCP_RBC5796_n_13962 ( .a(FE_OCP_RBN5792_n_13962), .o(FE_OCP_RBN5796_n_13962) );
in01s01 FE_OCP_RBC5797_n_13962 ( .a(FE_OCP_RBN5793_n_13962), .o(FE_OCP_RBN5797_n_13962) );
in01s01 FE_OCP_RBC5798_n_13962 ( .a(FE_OCP_RBN5793_n_13962), .o(FE_OCP_RBN5798_n_13962) );
in01s01 FE_OCP_RBC5799_n_13962 ( .a(FE_OCP_RBN5794_n_13962), .o(FE_OCP_RBN5799_n_13962) );
in01s01 FE_OCP_RBC5800_n_13962 ( .a(FE_OCP_RBN5794_n_13962), .o(FE_OCP_RBN5800_n_13962) );
in01s01 FE_OCP_RBC5801_n_13962 ( .a(FE_OCP_RBN5798_n_13962), .o(FE_OCP_RBN5801_n_13962) );
in01s01 FE_OCP_RBC5802_n_13962 ( .a(FE_OCP_RBN5798_n_13962), .o(FE_OCP_RBN5802_n_13962) );
in01m02 FE_OCP_RBC5803_FE_RN_2224_0 ( .a(FE_RN_2224_0), .o(FE_OCP_RBN5803_FE_RN_2224_0) );
in01s01 FE_OCP_RBC5804_n_47018 ( .a(n_47018), .o(FE_OCP_RBN5804_n_47018) );
in01s01 FE_OCP_RBC5805_n_47018 ( .a(n_47018), .o(FE_OCP_RBN5805_n_47018) );
in01s01 FE_OCP_RBC5806_n_47018 ( .a(FE_OCP_RBN5805_n_47018), .o(FE_OCP_RBN5806_n_47018) );
in01s01 FE_OCP_RBC5807_n_47018 ( .a(FE_OCP_RBN5806_n_47018), .o(FE_OCP_RBN5807_n_47018) );
in01s01 FE_OCP_RBC5808_n_47018 ( .a(FE_OCP_RBN5806_n_47018), .o(FE_OCP_RBN5808_n_47018) );
in01s02 FE_OCP_RBC5809_n_3645 ( .a(n_3645), .o(FE_OCP_RBN5809_n_3645) );
in01s01 FE_OCP_RBC5810_n_3645 ( .a(n_3645), .o(FE_OCP_RBN5810_n_3645) );
in01s01 FE_OCP_RBC5811_n_3645 ( .a(FE_OCP_RBN5810_n_3645), .o(FE_OCP_RBN5811_n_3645) );
in01s01 FE_OCP_RBC5812_n_9014 ( .a(n_9014), .o(FE_OCP_RBN5812_n_9014) );
in01s01 FE_OCP_RBC5813_n_9014 ( .a(FE_OCP_RBN6720_FE_OCP_DRV_N6264_n_9014), .o(FE_OCP_RBN5813_n_9014) );
in01s02 FE_OCP_RBC5814_n_20098 ( .a(n_20098), .o(FE_OCP_RBN5814_n_20098) );
in01m04 FE_OCP_RBC5815_n_24823 ( .a(n_24823), .o(FE_OCP_RBN5815_n_24823) );
in01s02 FE_OCP_RBC5816_n_38678 ( .a(n_38678), .o(FE_OCP_RBN5816_n_38678) );
in01s02 FE_OCP_RBC5817_n_8687 ( .a(n_8687), .o(FE_OCP_RBN5817_n_8687) );
in01s01 FE_OCP_RBC5818_n_8687 ( .a(n_8687), .o(FE_OCP_RBN5818_n_8687) );
in01s01 FE_OCP_RBC5819_n_8651 ( .a(n_8651), .o(FE_OCP_RBN5819_n_8651) );
in01m01 FE_OCP_RBC5820_n_3396 ( .a(n_3396), .o(FE_OCP_RBN5820_n_3396) );
in01s02 FE_OCP_RBC5821_n_3437 ( .a(n_3437), .o(FE_OCP_RBN5821_n_3437) );
in01s02 FE_OCP_RBC5822_n_8985 ( .a(n_8985), .o(FE_OCP_RBN5822_n_8985) );
in01f02 FE_OCP_RBC5823_n_14722 ( .a(n_14722), .o(FE_OCP_RBN5823_n_14722) );
in01f02 FE_OCP_RBC5824_n_14552 ( .a(n_14552), .o(FE_OCP_RBN5824_n_14552) );
in01s01 FE_OCP_RBC5825_n_8692 ( .a(FE_OCP_RBN2854_n_8692), .o(FE_OCP_RBN5825_n_8692) );
in01s02 FE_OCP_RBC5826_n_8692 ( .a(FE_OCP_RBN2854_n_8692), .o(FE_OCP_RBN5826_n_8692) );
in01s01 FE_OCP_RBC5827_n_44579 ( .a(n_44579), .o(FE_OCP_RBN5827_n_44579) );
in01s01 FE_OCP_RBC5828_n_44579 ( .a(n_44579), .o(FE_OCP_RBN5828_n_44579) );
in01s01 FE_OCP_RBC5829_n_44579 ( .a(n_44579), .o(FE_OCP_RBN5829_n_44579) );
in01s01 FE_OCP_RBC5830_n_44579 ( .a(n_44579), .o(FE_OCP_RBN5830_n_44579) );
in01s01 FE_OCP_RBC5833_n_44563 ( .a(FE_OCP_RBN6710_n_44570), .o(FE_OCP_RBN5833_n_44563) );
in01s01 FE_OCP_RBC5834_n_44563 ( .a(FE_OCP_RBN6710_n_44570), .o(FE_OCP_RBN5834_n_44563) );
in01s01 FE_OCP_RBC5835_n_44563 ( .a(FE_OCP_RBN6710_n_44570), .o(FE_OCP_RBN5835_n_44563) );
in01s10 FE_OCP_RBC5836_n_44563 ( .a(FE_OCP_RBN6710_n_44570), .o(FE_OCP_RBN5836_n_44563) );
in01s01 FE_OCP_RBC5837_n_44563 ( .a(FE_OCP_RBN6710_n_44570), .o(FE_OCP_RBN5837_n_44563) );
in01s04 FE_OCP_RBC5838_n_44563 ( .a(FE_OCP_RBN6711_n_44570), .o(FE_OCP_RBN5838_n_44563) );
in01s01 FE_OCP_RBC5842_n_44563 ( .a(FE_OCP_RBN6738_n_44563), .o(FE_OCP_RBN5842_n_44563) );
in01s02 FE_OCP_RBC5843_n_9035 ( .a(n_9035), .o(FE_OCP_RBN5843_n_9035) );
in01m02 FE_OCP_RBC5844_n_42169 ( .a(n_42169), .o(FE_OCP_RBN5844_n_42169) );
in01f02 FE_OCP_RBC5845_n_42169 ( .a(n_42169), .o(FE_OCP_RBN5845_n_42169) );
in01s01 FE_OCP_RBC5846_FE_RN_987_0 ( .a(FE_RN_987_0), .o(FE_OCP_RBN5846_FE_RN_987_0) );
in01s01 FE_OCP_RBC5847_FE_RN_987_0 ( .a(FE_RN_987_0), .o(FE_OCP_RBN5847_FE_RN_987_0) );
in01m02 FE_OCP_RBC5848_FE_RN_2187_0 ( .a(FE_RN_2187_0), .o(FE_OCP_RBN5848_FE_RN_2187_0) );
in01m01 FE_OCP_RBC5849_FE_RN_2187_0 ( .a(FE_OCP_RBN5848_FE_RN_2187_0), .o(FE_OCP_RBN5849_FE_RN_2187_0) );
in01s02 FE_OCP_RBC5850_FE_RN_2187_0 ( .a(FE_OCP_RBN5849_FE_RN_2187_0), .o(FE_OCP_RBN5850_FE_RN_2187_0) );
in01s01 FE_OCP_RBC5851_n_3625 ( .a(n_3625), .o(FE_OCP_RBN5851_n_3625) );
in01s01 FE_OCP_RBC5852_n_3625 ( .a(FE_OCP_RBN5851_n_3625), .o(FE_OCP_RBN5852_n_3625) );
in01s02 FE_OCP_RBC5853_n_14750 ( .a(n_14750), .o(FE_OCP_RBN5853_n_14750) );
in01m04 FE_OCP_RBC5854_n_34908 ( .a(n_34908), .o(FE_OCP_RBN5854_n_34908) );
in01s02 FE_OCP_RBC5855_n_3807 ( .a(n_3807), .o(FE_OCP_RBN5855_n_3807) );
in01s01 FE_OCP_RBC5856_n_3807 ( .a(n_3807), .o(FE_OCP_RBN5856_n_3807) );
in01s01 FE_OCP_RBC5857_FE_RN_998_0 ( .a(FE_RN_998_0), .o(FE_OCP_RBN5857_FE_RN_998_0) );
in01s02 FE_OCP_RBC5858_FE_RN_998_0 ( .a(FE_RN_998_0), .o(FE_OCP_RBN5858_FE_RN_998_0) );
in01s01 FE_OCP_RBC5859_FE_RN_998_0 ( .a(FE_RN_998_0), .o(FE_OCP_RBN5859_FE_RN_998_0) );
in01s02 FE_OCP_RBC5860_FE_RN_998_0 ( .a(FE_OCP_RBN5859_FE_RN_998_0), .o(FE_OCP_RBN5860_FE_RN_998_0) );
in01s01 FE_OCP_RBC5861_n_3718 ( .a(n_3718), .o(FE_OCP_RBN5861_n_3718) );
in01s01 FE_OCP_RBC5862_n_3718 ( .a(n_3718), .o(FE_OCP_RBN5862_n_3718) );
in01s02 FE_OCP_RBC5863_n_3705 ( .a(FE_OCP_RBN4255_n_3705), .o(FE_OCP_RBN5863_n_3705) );
in01s02 FE_OCP_RBC5864_n_3705 ( .a(FE_OCP_RBN5863_n_3705), .o(FE_OCP_RBN5864_n_3705) );
in01s01 FE_OCP_RBC5867_n_3661 ( .a(n_3661), .o(FE_OCP_RBN5867_n_3661) );
in01s01 FE_OCP_RBC5868_n_3704 ( .a(n_3704), .o(FE_OCP_RBN5868_n_3704) );
in01s08 FE_OCP_RBC5869_n_3704 ( .a(n_3704), .o(FE_OCP_RBN5869_n_3704) );
in01s06 FE_OCP_RBC5870_n_3704 ( .a(FE_OCP_RBN5869_n_3704), .o(FE_OCP_RBN5870_n_3704) );
in01m10 FE_OCP_RBC5871_n_3700 ( .a(n_3700), .o(FE_OCP_RBN5871_n_3700) );
in01s10 FE_OCP_RBC5872_n_3700 ( .a(FE_OCP_RBN5871_n_3700), .o(FE_OCP_RBN5872_n_3700) );
in01s04 FE_OCP_RBC5873_n_3700 ( .a(FE_OCP_RBN5871_n_3700), .o(FE_OCP_RBN5873_n_3700) );
in01s01 FE_OCP_RBC5875_n_3700 ( .a(FE_OCP_RBN5873_n_3700), .o(FE_OCP_RBN5875_n_3700) );
in01s01 FE_OCP_RBC5876_n_3848 ( .a(n_3848), .o(FE_OCP_RBN5876_n_3848) );
in01s01 FE_OCP_RBC5877_n_3848 ( .a(n_3848), .o(FE_OCP_RBN5877_n_3848) );
in01s02 FE_OCP_RBC5880_FE_RN_314_0 ( .a(FE_RN_314_0), .o(FE_OCP_RBN5880_FE_RN_314_0) );
in01s01 FE_OCP_RBC5881_FE_RN_314_0 ( .a(FE_RN_314_0), .o(FE_OCP_RBN5881_FE_RN_314_0) );
in01s01 FE_OCP_RBC5882_FE_RN_2220_0 ( .a(FE_RN_2220_0), .o(FE_OCP_RBN5882_FE_RN_2220_0) );
in01m02 FE_OCP_RBC5883_n_9042 ( .a(n_9042), .o(FE_OCP_RBN5883_n_9042) );
in01m02 FE_OCP_RBC5884_n_9306 ( .a(n_9306), .o(FE_OCP_RBN5884_n_9306) );
in01s01 FE_OCP_RBC5885_n_38806 ( .a(n_38806), .o(FE_OCP_RBN5885_n_38806) );
in01f08 FE_OCP_RBC5890_n_38806 ( .a(FE_OCP_RBN6758_n_38806), .o(FE_OCP_RBN5890_n_38806) );
in01s01 FE_OCP_RBC5892_n_38806 ( .a(FE_OCP_RBN6758_n_38806), .o(FE_OCP_RBN5892_n_38806) );
in01s01 FE_OCP_RBC5893_n_38806 ( .a(FE_OCP_RBN6758_n_38806), .o(FE_OCP_RBN5893_n_38806) );
in01s06 FE_OCP_RBC5894_n_38806 ( .a(FE_OCP_RBN6758_n_38806), .o(FE_OCP_RBN5894_n_38806) );
in01f10 FE_OCP_RBC5895_n_38806 ( .a(FE_OCP_RBN5890_n_38806), .o(FE_OCP_RBN5895_n_38806) );
in01m04 FE_OCP_RBC5896_n_38806 ( .a(FE_OCP_RBN5890_n_38806), .o(FE_OCP_RBN5896_n_38806) );
in01s08 FE_OCP_RBC5897_n_38806 ( .a(FE_OCP_RBN5894_n_38806), .o(FE_OCP_RBN5897_n_38806) );
in01m04 FE_OCP_RBC5898_n_35005 ( .a(n_35005), .o(FE_OCP_RBN5898_n_35005) );
in01s01 FE_OCP_RBC5899_n_35005 ( .a(n_35005), .o(FE_OCP_RBN5899_n_35005) );
in01m10 FE_OCP_RBC5900_n_25178 ( .a(FE_OCP_RBN2910_n_25178), .o(FE_OCP_RBN5900_n_25178) );
in01m02 FE_OCP_RBC5901_n_25178 ( .a(FE_OCP_RBN5900_n_25178), .o(FE_OCP_RBN5901_n_25178) );
in01s02 FE_OCP_RBC5902_n_25178 ( .a(FE_OCP_RBN5900_n_25178), .o(FE_OCP_RBN5902_n_25178) );
in01s02 FE_OCP_RBC5903_n_25178 ( .a(FE_OCP_RBN5902_n_25178), .o(FE_OCP_RBN5903_n_25178) );
in01s02 FE_OCP_RBC5904_n_8872 ( .a(FE_OCP_RBN4270_n_8872), .o(FE_OCP_RBN5904_n_8872) );
in01s01 FE_OCP_RBC5905_n_44563 ( .a(FE_OCP_RBN6741_n_44563), .o(FE_OCP_RBN5905_n_44563) );
in01m01 FE_OCP_RBC5906_n_44563 ( .a(FE_OCP_RBN6741_n_44563), .o(FE_OCP_RBN5906_n_44563) );
in01s02 FE_OCP_RBC5907_n_44563 ( .a(FE_OCP_RBN6741_n_44563), .o(FE_OCP_RBN5907_n_44563) );
in01s01 FE_OCP_RBC5908_n_44563 ( .a(FE_OCP_RBN5906_n_44563), .o(FE_OCP_RBN5908_n_44563) );
in01s01 FE_OCP_RBC5909_n_44563 ( .a(FE_OCP_RBN5906_n_44563), .o(FE_OCP_RBN5909_n_44563) );
in01s01 FE_OCP_RBC5910_n_44563 ( .a(FE_OCP_RBN5908_n_44563), .o(FE_OCP_RBN5910_n_44563) );
in01s01 FE_OCP_RBC5911_n_44563 ( .a(FE_OCP_RBN5908_n_44563), .o(FE_OCP_RBN5911_n_44563) );
in01s01 FE_OCP_RBC5912_n_44563 ( .a(FE_OCP_RBN5909_n_44563), .o(FE_OCP_RBN5912_n_44563) );
in01s01 FE_OCP_RBC5913_n_44563 ( .a(FE_OCP_RBN5909_n_44563), .o(FE_OCP_RBN5913_n_44563) );
in01s01 FE_OCP_RBC5914_n_3750 ( .a(n_3750), .o(FE_OCP_RBN5914_n_3750) );
in01s01 FE_OCP_RBC5915_n_3750 ( .a(n_3750), .o(FE_OCP_RBN5915_n_3750) );
in01s02 FE_OCP_RBC5916_n_3875 ( .a(n_3875), .o(FE_OCP_RBN5916_n_3875) );
in01s02 FE_OCP_RBC5917_n_4101 ( .a(n_4101), .o(FE_OCP_RBN5917_n_4101) );
in01s01 FE_OCP_RBC5918_n_4101 ( .a(n_4101), .o(FE_OCP_RBN5918_n_4101) );
in01s02 FE_OCP_RBC5919_n_9456 ( .a(n_9456), .o(FE_OCP_RBN5919_n_9456) );
in01m02 FE_OCP_RBC5920_n_9456 ( .a(n_9456), .o(FE_OCP_RBN5920_n_9456) );
in01m01 FE_OCP_RBC5921_n_20236 ( .a(n_20236), .o(FE_OCP_RBN5921_n_20236) );
in01s02 FE_OCP_RBC5922_n_25211 ( .a(n_25211), .o(FE_OCP_RBN5922_n_25211) );
in01s06 FE_OCP_RBC5923_n_25211 ( .a(n_25211), .o(FE_OCP_RBN5923_n_25211) );
in01s01 FE_OCP_RBC5924_n_25211 ( .a(n_25211), .o(FE_OCP_RBN5924_n_25211) );
in01s10 FE_OCP_RBC5925_n_25211 ( .a(FE_OCP_RBN5923_n_25211), .o(FE_OCP_RBN5925_n_25211) );
in01s02 FE_OCP_RBC5926_n_25211 ( .a(FE_OCP_RBN5925_n_25211), .o(FE_OCP_RBN5926_n_25211) );
in01s06 FE_OCP_RBC5927_n_25211 ( .a(FE_OCP_RBN5925_n_25211), .o(FE_OCP_RBN5927_n_25211) );
in01m02 FE_OCP_RBC5929_n_4158 ( .a(n_4158), .o(FE_OCP_RBN5929_n_4158) );
in01s02 FE_OCP_RBC5930_n_44563 ( .a(FE_OCP_RBN4288_n_44563), .o(FE_OCP_RBN5930_n_44563) );
in01s01 FE_OCP_RBC5931_n_44563 ( .a(FE_OCP_RBN4288_n_44563), .o(FE_OCP_RBN5931_n_44563) );
in01s01 FE_OCP_RBC5932_n_44563 ( .a(FE_OCP_RBN5930_n_44563), .o(FE_OCP_RBN5932_n_44563) );
in01s01 FE_OCP_RBC5933_n_44563 ( .a(FE_OCP_RBN5931_n_44563), .o(FE_OCP_RBN5933_n_44563) );
in01s01 FE_OCP_RBC5934_n_44563 ( .a(FE_OCP_RBN5932_n_44563), .o(FE_OCP_RBN5934_n_44563) );
in01s01 FE_OCP_RBC5935_n_44563 ( .a(FE_OCP_RBN5932_n_44563), .o(FE_OCP_RBN5935_n_44563) );
in01s01 FE_OCP_RBC5936_n_44563 ( .a(FE_OCP_RBN5933_n_44563), .o(FE_OCP_RBN5936_n_44563) );
in01s01 FE_OCP_RBC5937_n_44563 ( .a(FE_OCP_RBN5933_n_44563), .o(FE_OCP_RBN5937_n_44563) );
in01s01 FE_OCP_RBC5938_n_44563 ( .a(FE_OCP_RBN5933_n_44563), .o(FE_OCP_RBN5938_n_44563) );
in01s01 FE_OCP_RBC5939_n_44563 ( .a(FE_OCP_RBN5933_n_44563), .o(FE_OCP_RBN5939_n_44563) );
in01s02 FE_OCP_RBC5940_n_4238 ( .a(n_4238), .o(FE_OCP_RBN5940_n_4238) );
in01m02 FE_OCP_RBC5941_n_9374 ( .a(n_9374), .o(FE_OCP_RBN5941_n_9374) );
in01f03 FE_OCP_RBC5942_n_25544 ( .a(n_25544), .o(FE_OCP_RBN5942_n_25544) );
in01s02 FE_OCP_RBC5943_n_35207 ( .a(n_35207), .o(FE_OCP_RBN5943_n_35207) );
in01s04 FE_OCP_RBC5944_n_35207 ( .a(n_35207), .o(FE_OCP_RBN5944_n_35207) );
in01s04 FE_OCP_RBC5945_FE_RN_1231_0 ( .a(FE_RN_1231_0), .o(FE_OCP_RBN5945_FE_RN_1231_0) );
in01m06 FE_OCP_RBC5946_n_14982 ( .a(n_14982), .o(FE_OCP_RBN5946_n_14982) );
in01m04 FE_OCP_RBC5947_n_14982 ( .a(FE_OCP_RBN5946_n_14982), .o(FE_OCP_RBN5947_n_14982) );
in01s06 FE_OCP_RBC5948_n_14982 ( .a(FE_OCP_RBN5946_n_14982), .o(FE_OCP_RBN5948_n_14982) );
in01s01 FE_OCP_RBC5949_FE_OFN4772_n_44463 ( .a(FE_OFN4772_n_44463), .o(FE_OCP_RBN5949_FE_OFN4772_n_44463) );
in01s01 FE_OCP_RBC5950_FE_OFN4772_n_44463 ( .a(FE_OCP_RBN5949_FE_OFN4772_n_44463), .o(FE_OCP_RBN5950_FE_OFN4772_n_44463) );
in01s01 FE_OCP_RBC5951_FE_OFN4772_n_44463 ( .a(FE_OCP_RBN5949_FE_OFN4772_n_44463), .o(FE_OCP_RBN5951_FE_OFN4772_n_44463) );
in01s01 FE_OCP_RBC5952_FE_OFN4772_n_44463 ( .a(FE_OCP_RBN5950_FE_OFN4772_n_44463), .o(FE_OCP_RBN5952_FE_OFN4772_n_44463) );
in01s01 FE_OCP_RBC5953_FE_OFN4772_n_44463 ( .a(FE_OCP_RBN5950_FE_OFN4772_n_44463), .o(FE_OCP_RBN5953_FE_OFN4772_n_44463) );
in01s01 FE_OCP_RBC5954_FE_OFN4772_n_44463 ( .a(FE_OCP_RBN5951_FE_OFN4772_n_44463), .o(FE_OCP_RBN5954_FE_OFN4772_n_44463) );
in01s02 FE_OCP_RBC5955_FE_OFN4772_n_44463 ( .a(FE_OCP_RBN5951_FE_OFN4772_n_44463), .o(FE_OCP_RBN5955_FE_OFN4772_n_44463) );
in01s01 FE_OCP_RBC5956_n_47012 ( .a(n_47012), .o(FE_OCP_RBN5956_n_47012) );
in01m02 FE_OCP_RBC5957_n_47012 ( .a(n_47012), .o(FE_OCP_RBN5957_n_47012) );
in01s01 FE_OCP_RBC5958_n_4165 ( .a(n_4165), .o(FE_OCP_RBN5958_n_4165) );
in01s02 FE_OCP_RBC5959_n_4165 ( .a(n_4165), .o(FE_OCP_RBN5959_n_4165) );
in01s02 FE_OCP_RBC5960_n_4397 ( .a(n_4397), .o(FE_OCP_RBN5960_n_4397) );
in01s01 FE_OCP_RBC5961_n_20459 ( .a(n_20459), .o(FE_OCP_RBN5961_n_20459) );
in01s01 FE_OCP_RBC5962_n_20459 ( .a(n_20459), .o(FE_OCP_RBN5962_n_20459) );
in01s01 FE_OCP_RBC5963_n_39097 ( .a(n_39097), .o(FE_OCP_RBN5963_n_39097) );
in01s01 FE_OCP_RBC5964_n_39097 ( .a(FE_OCP_RBN5963_n_39097), .o(FE_OCP_RBN5964_n_39097) );
in01s02 FE_OCP_RBC5965_n_39097 ( .a(FE_OCP_RBN5964_n_39097), .o(FE_OCP_RBN5965_n_39097) );
in01s01 FE_OCP_RBC5966_n_39098 ( .a(n_39098), .o(FE_OCP_RBN5966_n_39098) );
in01s02 FE_OCP_RBC5967_n_14905 ( .a(n_14905), .o(FE_OCP_RBN5967_n_14905) );
in01s01 FE_OCP_RBC5968_n_14905 ( .a(n_14905), .o(FE_OCP_RBN5968_n_14905) );
in01m02 FE_OCP_RBC5969_n_9668 ( .a(n_9668), .o(FE_OCP_RBN5969_n_9668) );
in01f02 FE_OCP_RBC5970_n_15235 ( .a(n_15235), .o(FE_OCP_RBN5970_n_15235) );
in01f02 FE_OCP_RBC5971_n_20510 ( .a(n_20510), .o(FE_OCP_RBN5971_n_20510) );
in01f04 FE_OCP_RBC5972_n_9494 ( .a(n_9494), .o(FE_OCP_RBN5972_n_9494) );
in01m02 FE_OCP_RBC5973_n_35231 ( .a(n_35231), .o(FE_OCP_RBN5973_n_35231) );
in01m02 FE_OCP_RBC5974_FE_RN_2033_0 ( .a(FE_RN_2033_0), .o(FE_OCP_RBN5974_FE_RN_2033_0) );
in01s02 FE_OCP_RBC5975_FE_RN_2033_0 ( .a(FE_OCP_RBN5974_FE_RN_2033_0), .o(FE_OCP_RBN5975_FE_RN_2033_0) );
in01s02 FE_OCP_RBC5976_FE_RN_2033_0 ( .a(FE_OCP_RBN5975_FE_RN_2033_0), .o(FE_OCP_RBN5976_FE_RN_2033_0) );
in01s01 FE_OCP_RBC5977_n_4245 ( .a(n_4245), .o(FE_OCP_RBN5977_n_4245) );
in01m01 FE_OCP_RBC5978_n_9682 ( .a(n_9682), .o(FE_OCP_RBN5978_n_9682) );
in01s01 FE_OCP_RBC5979_n_9682 ( .a(n_9682), .o(FE_OCP_RBN5979_n_9682) );
in01s01 FE_OCP_RBC5980_n_9682 ( .a(FE_OCP_RBN5979_n_9682), .o(FE_OCP_RBN5980_n_9682) );
in01s02 FE_OCP_RBC5981_n_9856 ( .a(n_9856), .o(FE_OCP_RBN5981_n_9856) );
in01s01 FE_OCP_RBC5982_n_15160 ( .a(n_15160), .o(FE_OCP_RBN5982_n_15160) );
in01s01 FE_OCP_RBC5983_n_20495 ( .a(n_20495), .o(FE_OCP_RBN5983_n_20495) );
in01f02 FE_OCP_RBC5984_n_15079 ( .a(n_15079), .o(FE_OCP_RBN5984_n_15079) );
in01s01 FE_OCP_RBC5985_n_15079 ( .a(n_15079), .o(FE_OCP_RBN5985_n_15079) );
in01s01 FE_OCP_RBC5987_n_15135 ( .a(FE_OCP_RBN6798_n_15156), .o(FE_OCP_RBN5987_n_15135) );
in01m02 FE_OCP_RBC5988_FE_RN_1865_0 ( .a(FE_RN_1865_0), .o(FE_OCP_RBN5988_FE_RN_1865_0) );
in01m01 FE_OCP_RBC5989_FE_RN_1865_0 ( .a(FE_OCP_RBN5988_FE_RN_1865_0), .o(FE_OCP_RBN5989_FE_RN_1865_0) );
in01s01 FE_OCP_RBC5990_FE_RN_1865_0 ( .a(FE_OCP_RBN5989_FE_RN_1865_0), .o(FE_OCP_RBN5990_FE_RN_1865_0) );
in01s01 FE_OCP_RBC5991_n_4226 ( .a(n_4226), .o(FE_OCP_RBN5991_n_4226) );
in01m02 FE_OCP_RBC5992_n_4376 ( .a(n_4376), .o(FE_OCP_RBN5992_n_4376) );
in01s04 FE_OCP_RBC5993_n_15387 ( .a(n_15387), .o(FE_OCP_RBN5993_n_15387) );
in01f02 FE_OCP_RBC5994_n_15387 ( .a(n_15387), .o(FE_OCP_RBN5994_n_15387) );
in01f02 FE_OCP_RBC5995_n_25702 ( .a(n_25702), .o(FE_OCP_RBN5995_n_25702) );
in01m02 FE_OCP_RBC5996_n_25732 ( .a(n_25732), .o(FE_OCP_RBN5996_n_25732) );
in01s02 FE_OCP_RBC5997_n_25732 ( .a(n_25732), .o(FE_OCP_RBN5997_n_25732) );
in01s02 FE_OCP_RBC5998_n_25732 ( .a(n_25732), .o(FE_OCP_RBN5998_n_25732) );
in01m02 FE_OCP_RBC6000_n_30534 ( .a(n_30534), .o(FE_OCP_RBN6000_n_30534) );
in01s01 FE_OCP_RBC6001_n_30534 ( .a(n_30534), .o(FE_OCP_RBN6001_n_30534) );
in01m02 FE_OCP_RBC6002_n_10015 ( .a(n_10015), .o(FE_OCP_RBN6002_n_10015) );
in01s02 FE_OCP_RBC6003_n_10068 ( .a(n_10068), .o(FE_OCP_RBN6003_n_10068) );
in01s02 FE_OCP_RBC6004_n_10068 ( .a(n_10068), .o(FE_OCP_RBN6004_n_10068) );
in01m02 FE_OCP_RBC6005_n_15704 ( .a(n_15704), .o(FE_OCP_RBN6005_n_15704) );
in01m04 FE_OCP_RBC6006_n_15704 ( .a(n_15704), .o(FE_OCP_RBN6006_n_15704) );
in01s01 FE_OCP_RBC6008_n_30608 ( .a(FE_OCP_RBN6812_n_30608), .o(FE_OCP_RBN6008_n_30608) );
in01s02 FE_OCP_RBC6009_n_4683 ( .a(n_4683), .o(FE_OCP_RBN6009_n_4683) );
in01m01 FE_OCP_RBC6010_n_10277 ( .a(n_10277), .o(FE_OCP_RBN6010_n_10277) );
in01f02 FE_OCP_RBC6011_n_10277 ( .a(FE_OCP_RBN6010_n_10277), .o(FE_OCP_RBN6011_n_10277) );
in01f02 FE_OCP_RBC6012_n_10277 ( .a(FE_OCP_RBN6011_n_10277), .o(FE_OCP_RBN6012_n_10277) );
in01m02 FE_OCP_RBC6013_n_25900 ( .a(n_25900), .o(FE_OCP_RBN6013_n_25900) );
in01m02 FE_OCP_RBC6015_n_10225 ( .a(n_10225), .o(FE_OCP_RBN6015_n_10225) );
in01m02 FE_OCP_RBC6016_n_30625 ( .a(n_30625), .o(FE_OCP_RBN6016_n_30625) );
in01m02 FE_OCP_RBC6017_n_20945 ( .a(n_20945), .o(FE_OCP_RBN6017_n_20945) );
in01m04 FE_OCP_RBC6018_n_25895 ( .a(n_25895), .o(FE_OCP_RBN6018_n_25895) );
in01s03 FE_OCP_RBC6019_n_46959 ( .a(n_46959), .o(FE_OCP_RBN6019_n_46959) );
in01s01 FE_OCP_RBC6020_n_46959 ( .a(FE_OCP_RBN6019_n_46959), .o(FE_OCP_RBN6020_n_46959) );
in01s01 FE_OCP_RBC6021_n_46959 ( .a(FE_OCP_RBN6019_n_46959), .o(FE_OCP_RBN6021_n_46959) );
in01s01 FE_OCP_RBC6022_n_46959 ( .a(FE_OCP_RBN6020_n_46959), .o(FE_OCP_RBN6022_n_46959) );
in01m04 FE_OCP_RBC6023_n_30711 ( .a(n_30711), .o(FE_OCP_RBN6023_n_30711) );
in01s01 FE_OCP_RBC6024_n_30711 ( .a(n_30711), .o(FE_OCP_RBN6024_n_30711) );
in01s02 FE_OCP_RBC6025_n_4858 ( .a(n_4858), .o(FE_OCP_RBN6025_n_4858) );
in01s01 FE_OCP_RBC6026_n_4858 ( .a(n_4858), .o(FE_OCP_RBN6026_n_4858) );
in01s02 FE_OCP_RBC6027_n_10445 ( .a(n_10445), .o(FE_OCP_RBN6027_n_10445) );
in01m04 FE_OCP_RBC6028_n_25928 ( .a(n_25928), .o(FE_OCP_RBN6028_n_25928) );
in01s01 FE_OCP_RBC6029_n_25928 ( .a(n_25928), .o(FE_OCP_RBN6029_n_25928) );
in01s01 FE_OCP_RBC6031_n_25997 ( .a(FE_OCP_RBN6819_n_25997), .o(FE_OCP_RBN6031_n_25997) );
in01f02 FE_OCP_RBC6032_n_30706 ( .a(n_30706), .o(FE_OCP_RBN6032_n_30706) );
in01m04 FE_OCP_RBC6033_n_46962 ( .a(n_46962), .o(FE_OCP_RBN6033_n_46962) );
in01s01 FE_OCP_RBC6034_n_46962 ( .a(n_46962), .o(FE_OCP_RBN6034_n_46962) );
in01f02 FE_OCP_RBC6035_n_30769 ( .a(n_30769), .o(FE_OCP_RBN6035_n_30769) );
in01s02 FE_OCP_RBC6036_n_10399 ( .a(n_10399), .o(FE_OCP_RBN6036_n_10399) );
in01s01 FE_OCP_RBC6037_n_10399 ( .a(n_10399), .o(FE_OCP_RBN6037_n_10399) );
in01s01 FE_OCP_RBC6038_n_30733 ( .a(n_30733), .o(FE_OCP_RBN6038_n_30733) );
in01s02 FE_OCP_RBC6039_n_30733 ( .a(n_30733), .o(FE_OCP_RBN6039_n_30733) );
in01s02 FE_OCP_RBC6040_n_4800 ( .a(n_4800), .o(FE_OCP_RBN6040_n_4800) );
in01s01 FE_OCP_RBC6041_n_10511 ( .a(n_10511), .o(FE_OCP_RBN6041_n_10511) );
in01m10 FE_OCP_RBC6044_n_35487 ( .a(n_35487), .o(FE_OCP_RBN6044_n_35487) );
in01m10 FE_OCP_RBC6045_n_35487 ( .a(FE_OCP_RBN6044_n_35487), .o(FE_OCP_RBN6045_n_35487) );
in01s01 FE_OCP_RBC6046_n_35487 ( .a(FE_OCP_RBN6044_n_35487), .o(FE_OCP_RBN6046_n_35487) );
in01s04 FE_OCP_RBC6047_n_35487 ( .a(FE_OCP_RBN6045_n_35487), .o(FE_OCP_RBN6047_n_35487) );
in01s06 FE_OCP_RBC6048_n_35487 ( .a(FE_OCP_RBN6047_n_35487), .o(FE_OCP_RBN6048_n_35487) );
in01m02 FE_OCP_RBC6049_n_10570 ( .a(n_10570), .o(FE_OCP_RBN6049_n_10570) );
in01s02 FE_OCP_RBC6050_n_21118 ( .a(n_21118), .o(FE_OCP_RBN6050_n_21118) );
in01s01 FE_OCP_RBC6051_n_21118 ( .a(n_21118), .o(FE_OCP_RBN6051_n_21118) );
in01s01 FE_OCP_RBC6053_n_15514 ( .a(FE_OCP_RBN6826_n_15514), .o(FE_OCP_RBN6053_n_15514) );
in01s01 FE_OCP_RBC6055_n_46957 ( .a(n_46957), .o(FE_OCP_RBN6055_n_46957) );
in01s02 FE_OCP_RBC6056_n_46957 ( .a(n_46957), .o(FE_OCP_RBN6056_n_46957) );
in01s04 FE_OCP_RBC6057_n_16011 ( .a(n_16011), .o(FE_OCP_RBN6057_n_16011) );
in01m04 FE_OCP_RBC6058_n_10478 ( .a(n_10478), .o(FE_OCP_RBN6058_n_10478) );
in01s02 FE_OCP_RBC6059_n_15795 ( .a(n_15795), .o(FE_OCP_RBN6059_n_15795) );
in01m02 FE_OCP_RBC6060_n_21194 ( .a(n_21194), .o(FE_OCP_RBN6060_n_21194) );
in01s01 FE_OCP_RBC6061_n_21194 ( .a(n_21194), .o(FE_OCP_RBN6061_n_21194) );
in01s01 FE_OCP_RBC6062_n_21194 ( .a(n_21194), .o(FE_OCP_RBN6062_n_21194) );
in01s01 FE_OCP_RBC6063_n_30908 ( .a(n_30908), .o(FE_OCP_RBN6063_n_30908) );
in01s02 FE_OCP_RBC6064_n_30908 ( .a(n_30908), .o(FE_OCP_RBN6064_n_30908) );
in01s02 FE_OCP_RBC6065_n_26081 ( .a(n_26081), .o(FE_OCP_RBN6065_n_26081) );
in01s01 FE_OCP_RBC6066_n_26081 ( .a(n_26081), .o(FE_OCP_RBN6066_n_26081) );
in01s02 FE_OCP_RBC6067_n_26121 ( .a(n_26121), .o(FE_OCP_RBN6067_n_26121) );
in01f02 FE_OCP_RBC6068_n_26121 ( .a(n_26121), .o(FE_OCP_RBN6068_n_26121) );
in01m02 FE_OCP_RBC6069_n_26140 ( .a(n_26140), .o(FE_OCP_RBN6069_n_26140) );
in01s04 FE_OCP_RBC6070_n_16041 ( .a(n_16041), .o(FE_OCP_RBN6070_n_16041) );
in01s01 FE_OCP_RBC6071_n_16041 ( .a(n_16041), .o(FE_OCP_RBN6071_n_16041) );
in01s06 FE_OCP_RBC6072_n_16086 ( .a(n_16086), .o(FE_OCP_RBN6072_n_16086) );
in01s01 FE_OCP_RBC6073_n_16086 ( .a(n_16086), .o(FE_OCP_RBN6073_n_16086) );
in01m01 FE_OCP_RBC6074_n_44256 ( .a(FE_OCP_RBN4906_n_44256), .o(FE_OCP_RBN6074_n_44256) );
in01s02 FE_OCP_RBC6075_n_44256 ( .a(FE_OCP_RBN4906_n_44256), .o(FE_OCP_RBN6075_n_44256) );
in01s01 FE_OCP_RBC6076_n_44256 ( .a(FE_OCP_RBN4906_n_44256), .o(FE_OCP_RBN6076_n_44256) );
in01s04 FE_OCP_RBC6077_n_16084 ( .a(n_16084), .o(FE_OCP_RBN6077_n_16084) );
in01s01 FE_OCP_RBC6078_n_16084 ( .a(n_16084), .o(FE_OCP_RBN6078_n_16084) );
in01m02 FE_OCP_RBC6079_n_30965 ( .a(n_30965), .o(FE_OCP_RBN6079_n_30965) );
in01s01 FE_OCP_RBC6080_n_5346 ( .a(n_5346), .o(FE_OCP_RBN6080_n_5346) );
in01s02 FE_OCP_RBC6081_n_5486 ( .a(n_5486), .o(FE_OCP_RBN6081_n_5486) );
in01s01 FE_OCP_RBC6082_n_5454 ( .a(n_5454), .o(FE_OCP_RBN6082_n_5454) );
in01s02 FE_OCP_RBC6083_n_5454 ( .a(n_5454), .o(FE_OCP_RBN6083_n_5454) );
in01s01 FE_OCP_RBC6084_n_31010 ( .a(n_31010), .o(FE_OCP_RBN6084_n_31010) );
in01m02 FE_OCP_RBC6085_n_31010 ( .a(n_31010), .o(FE_OCP_RBN6085_n_31010) );
in01s02 FE_OCP_RBC6086_n_10852 ( .a(n_10852), .o(FE_OCP_RBN6086_n_10852) );
in01s01 FE_OCP_RBC6087_n_10852 ( .a(FE_OCP_RBN6086_n_10852), .o(FE_OCP_RBN6087_n_10852) );
in01m02 FE_OCP_RBC6088_n_26181 ( .a(n_26181), .o(FE_OCP_RBN6088_n_26181) );
in01s02 FE_OCP_RBC6089_n_26304 ( .a(n_26304), .o(FE_OCP_RBN6089_n_26304) );
in01m04 FE_OCP_RBC6090_n_26322 ( .a(n_26322), .o(FE_OCP_RBN6090_n_26322) );
in01s02 FE_OCP_RBC6091_n_31153 ( .a(n_31153), .o(FE_OCP_RBN6091_n_31153) );
in01s01 FE_OCP_RBC6092_n_5531 ( .a(n_5531), .o(FE_OCP_RBN6092_n_5531) );
in01m02 FE_OCP_RBC6093_n_10660 ( .a(n_10660), .o(FE_OCP_RBN6093_n_10660) );
in01s02 FE_OCP_RBC6094_n_10946 ( .a(n_10946), .o(FE_OCP_RBN6094_n_10946) );
in01s10 FE_OCP_RBC6095_n_26160 ( .a(FE_OCP_RBN3266_n_26160), .o(FE_OCP_RBN6095_n_26160) );
in01s06 FE_OCP_RBC6096_n_26160 ( .a(FE_OCP_RBN6095_n_26160), .o(FE_OCP_RBN6096_n_26160) );
in01s10 FE_OCP_RBC6097_n_26160 ( .a(FE_OCP_RBN6095_n_26160), .o(FE_OCP_RBN6097_n_26160) );
in01f02 FE_OCP_RBC6098_n_5614 ( .a(n_5614), .o(FE_OCP_RBN6098_n_5614) );
in01s02 FE_OCP_RBC6101_n_21636 ( .a(n_21636), .o(FE_OCP_RBN6101_n_21636) );
in01s02 FE_OCP_RBC6102_n_26358 ( .a(n_26358), .o(FE_OCP_RBN6102_n_26358) );
in01s01 FE_OCP_RBC6104_n_36199 ( .a(n_36199), .o(FE_OCP_RBN6104_n_36199) );
in01m06 FE_OCP_RBC6105_n_39793 ( .a(n_39793), .o(FE_OCP_RBN6105_n_39793) );
in01f04 FE_OCP_RBC6106_n_39793 ( .a(n_39793), .o(FE_OCP_RBN6106_n_39793) );
in01s02 FE_OCP_RBC6108_n_39793 ( .a(FE_OCP_RBN6851_n_39793), .o(FE_OCP_RBN6108_n_39793) );
in01s06 FE_OCP_RBC6109_n_43022 ( .a(n_43022), .o(FE_OCP_RBN6109_n_43022) );
in01s01 FE_OCP_RBC6110_n_43022 ( .a(FE_OCP_RBN6109_n_43022), .o(FE_OCP_RBN6110_n_43022) );
in01s02 FE_OCP_RBC6111_n_5444 ( .a(n_5444), .o(FE_OCP_RBN6111_n_5444) );
in01s01 FE_OCP_RBC6112_n_5444 ( .a(FE_OCP_RBN6111_n_5444), .o(FE_OCP_RBN6112_n_5444) );
in01s01 FE_OCP_RBC6113_n_5444 ( .a(FE_OCP_RBN6112_n_5444), .o(FE_OCP_RBN6113_n_5444) );
in01s01 FE_OCP_RBC6114_n_5444 ( .a(FE_OCP_RBN6112_n_5444), .o(FE_OCP_RBN6114_n_5444) );
in01s01 FE_OCP_RBC6115_n_5444 ( .a(FE_OCP_RBN6112_n_5444), .o(FE_OCP_RBN6115_n_5444) );
in01s02 FE_OCP_RBC6116_n_11004 ( .a(n_11004), .o(FE_OCP_RBN6116_n_11004) );
in01s01 FE_OCP_RBC6117_n_11004 ( .a(n_11004), .o(FE_OCP_RBN6117_n_11004) );
in01s02 FE_OCP_RBC6118_n_5555 ( .a(n_5555), .o(FE_OCP_RBN6118_n_5555) );
in01s01 FE_OCP_RBC6119_n_5555 ( .a(n_5555), .o(FE_OCP_RBN6119_n_5555) );
in01s01 FE_OCP_RBC6120_n_26398 ( .a(n_26398), .o(FE_OCP_RBN6120_n_26398) );
in01m02 FE_OCP_RBC6121_n_26398 ( .a(n_26398), .o(FE_OCP_RBN6121_n_26398) );
in01s02 FE_OCP_RBC6122_n_10904 ( .a(n_10904), .o(FE_OCP_RBN6122_n_10904) );
in01s02 FE_OCP_RBC6123_n_21630 ( .a(n_21630), .o(FE_OCP_RBN6123_n_21630) );
in01s02 FE_OCP_RBC6124_n_5465 ( .a(n_5465), .o(FE_OCP_RBN6124_n_5465) );
in01s02 FE_OCP_RBC6127_n_11026 ( .a(n_11026), .o(FE_OCP_RBN6127_n_11026) );
in01s01 FE_OCP_RBC6128_n_11026 ( .a(n_11026), .o(FE_OCP_RBN6128_n_11026) );
in01m04 FE_OCP_RBC6129_n_21804 ( .a(n_21804), .o(FE_OCP_RBN6129_n_21804) );
in01s01 FE_OCP_RBC6130_n_46424 ( .a(n_46424), .o(FE_OCP_RBN6130_n_46424) );
in01m02 FE_OCP_RBC6131_n_21736 ( .a(n_21736), .o(FE_OCP_RBN6131_n_21736) );
in01s02 FE_OCP_RBC6132_n_26778 ( .a(n_26778), .o(FE_OCP_RBN6132_n_26778) );
in01s02 FE_OCP_RBC6133_n_11169 ( .a(n_11169), .o(FE_OCP_RBN6133_n_11169) );
in01s02 FE_OCP_RBC6134_n_11221 ( .a(n_11221), .o(FE_OCP_RBN6134_n_11221) );
in01f02 FE_OCP_RBC6135_n_16553 ( .a(n_16553), .o(FE_OCP_RBN6135_n_16553) );
in01s02 FE_OCP_RBC6136_n_5816 ( .a(n_5816), .o(FE_OCP_RBN6136_n_5816) );
in01m04 FE_OCP_RBC6137_n_11364 ( .a(n_11364), .o(FE_OCP_RBN6137_n_11364) );
in01s01 FE_OCP_RBC6138_n_31520 ( .a(n_31520), .o(FE_OCP_RBN6138_n_31520) );
in01m04 FE_OCP_RBC6139_n_31520 ( .a(n_31520), .o(FE_OCP_RBN6139_n_31520) );
in01s01 FE_OCP_RBC6144_n_46285 ( .a(n_46285), .o(FE_OCP_RBN6144_n_46285) );
in01m02 FE_OCP_RBC6149_n_5974 ( .a(n_5974), .o(FE_OCP_RBN6149_n_5974) );
in01s02 FE_OCP_RBC6150_n_36501 ( .a(n_36501), .o(FE_OCP_RBN6150_n_36501) );
in01s06 FE_OCP_RBC6151_n_36501 ( .a(n_36501), .o(FE_OCP_RBN6151_n_36501) );
in01m04 FE_OCP_RBC6152_n_39816 ( .a(n_39816), .o(FE_OCP_RBN6152_n_39816) );
in01m06 FE_OCP_RBC6153_n_39816 ( .a(FE_OCP_RBN6152_n_39816), .o(FE_OCP_RBN6153_n_39816) );
in01m20 FE_OCP_RBC6154_n_39816 ( .a(FE_OCP_RBN6153_n_39816), .o(FE_OCP_RBN6154_n_39816) );
in01s01 FE_OCP_RBC6155_n_39816 ( .a(FE_OCP_RBN6153_n_39816), .o(FE_OCP_RBN6155_n_39816) );
in01s02 FE_OCP_RBC6156_n_39816 ( .a(FE_OCP_RBN6154_n_39816), .o(FE_OCP_RBN6156_n_39816) );
in01s10 FE_OCP_RBC6157_n_39816 ( .a(FE_OCP_RBN6154_n_39816), .o(FE_OCP_RBN6157_n_39816) );
in01s01 FE_OCP_RBC6158_n_39816 ( .a(FE_OCP_RBN6156_n_39816), .o(FE_OCP_RBN6158_n_39816) );
in01s02 FE_OCP_RBC6159_n_39816 ( .a(FE_OCP_RBN6156_n_39816), .o(FE_OCP_RBN6159_n_39816) );
in01s06 FE_OCP_RBC6160_n_39816 ( .a(FE_OCP_RBN6157_n_39816), .o(FE_OCP_RBN6160_n_39816) );
in01s06 FE_OCP_RBC6161_n_39816 ( .a(FE_OCP_RBN6160_n_39816), .o(FE_OCP_RBN6161_n_39816) );
in01m08 FE_OCP_RBC6162_FE_RN_1136_0 ( .a(FE_RN_1136_0), .o(FE_OCP_RBN6162_FE_RN_1136_0) );
in01s01 FE_OCP_RBC6163_n_46337 ( .a(n_46337), .o(FE_OCP_RBN6163_n_46337) );
in01s03 FE_OCP_RBC6164_n_46337 ( .a(n_46337), .o(FE_OCP_RBN6164_n_46337) );
in01s08 FE_OCP_RBC6165_n_46337 ( .a(n_46337), .o(FE_OCP_RBN6165_n_46337) );
in01s04 FE_OCP_RBC6166_n_46337 ( .a(FE_OCP_RBN6164_n_46337), .o(FE_OCP_RBN6166_n_46337) );
in01s04 FE_OCP_RBC6167_n_46337 ( .a(FE_OCP_RBN6165_n_46337), .o(FE_OCP_RBN6167_n_46337) );
in01s06 FE_OCP_RBC6168_n_46337 ( .a(FE_OCP_RBN6165_n_46337), .o(FE_OCP_RBN6168_n_46337) );
in01m02 FE_OCP_RBC6169_n_6021 ( .a(n_6021), .o(FE_OCP_RBN6169_n_6021) );
in01s02 FE_OCP_RBC6170_n_6059 ( .a(n_6059), .o(FE_OCP_RBN6170_n_6059) );
in01s02 FE_OCP_RBC6171_n_6059 ( .a(n_6059), .o(FE_OCP_RBN6171_n_6059) );
in01m06 FE_OCP_RBC6172_n_16923 ( .a(n_16923), .o(FE_OCP_RBN6172_n_16923) );
in01s01 FE_OCP_RBC6173_n_16923 ( .a(n_16923), .o(FE_OCP_RBN6173_n_16923) );
in01m01 FE_OCP_RBC6174_n_16923 ( .a(n_16923), .o(FE_OCP_RBN6174_n_16923) );
in01m08 FE_OCP_RBC6175_n_16923 ( .a(FE_OCP_RBN6172_n_16923), .o(FE_OCP_RBN6175_n_16923) );
in01s01 FE_OCP_RBC6176_n_16923 ( .a(FE_OCP_RBN6175_n_16923), .o(FE_OCP_RBN6176_n_16923) );
in01s04 FE_OCP_RBC6177_n_36444 ( .a(n_36444), .o(FE_OCP_RBN6177_n_36444) );
in01s02 FE_OCP_RBC6178_n_22106 ( .a(n_22106), .o(FE_OCP_RBN6178_n_22106) );
in01s01 FE_OCP_RBC6179_n_22106 ( .a(n_22106), .o(FE_OCP_RBN6179_n_22106) );
in01s02 FE_OCP_RBC6182_n_44267 ( .a(n_44267), .o(FE_OCP_RBN6182_n_44267) );
in01m08 FE_OCP_RBC6183_n_44267 ( .a(n_44267), .o(FE_OCP_RBN6183_n_44267) );
in01f08 FE_OCP_RBC6184_n_44267 ( .a(FE_OCP_RBN6183_n_44267), .o(FE_OCP_RBN6184_n_44267) );
in01s01 FE_OCP_RBC6185_n_44267 ( .a(FE_OCP_RBN6183_n_44267), .o(FE_OCP_RBN6185_n_44267) );
in01m02 FE_OCP_RBC6186_n_16824 ( .a(n_16824), .o(FE_OCP_RBN6186_n_16824) );
in01s01 FE_OCP_RBC6187_n_31916 ( .a(n_31916), .o(FE_OCP_RBN6187_n_31916) );
in01s02 FE_OCP_RBC6188_n_11403 ( .a(n_11403), .o(FE_OCP_RBN6188_n_11403) );
in01s02 FE_OCP_RBC6189_n_11403 ( .a(n_11403), .o(FE_OCP_RBN6189_n_11403) );
in01m10 FE_OCP_RBC6190_n_43103 ( .a(FE_OCP_RBN4457_n_43103), .o(FE_OCP_RBN6190_n_43103) );
in01s20 FE_OCP_RBC6191_n_43103 ( .a(FE_OCP_RBN6190_n_43103), .o(FE_OCP_RBN6191_n_43103) );
in01s06 FE_OCP_RBC6192_n_43103 ( .a(FE_OCP_RBN6190_n_43103), .o(FE_OCP_RBN6192_n_43103) );
in01s01 FE_OCP_RBC6193_n_10636 ( .a(n_10636), .o(FE_OCP_RBN6193_n_10636) );
in01s01 FE_OCP_RBC6194_n_10636 ( .a(FE_OCP_RBN6193_n_10636), .o(FE_OCP_RBN6194_n_10636) );
in01m10 FE_OCP_RBC6195_FE_OFN789_n_46195 ( .a(FE_OFN789_n_46195), .o(FE_OCP_RBN6195_FE_OFN789_n_46195) );
in01s02 FE_OCP_RBC6196_FE_OFN789_n_46195 ( .a(FE_OFN789_n_46195), .o(FE_OCP_RBN6196_FE_OFN789_n_46195) );
in01m06 FE_OCP_RBC6197_FE_OFN789_n_46195 ( .a(FE_OCP_RBN6195_FE_OFN789_n_46195), .o(FE_OCP_RBN6197_FE_OFN789_n_46195) );
in01s01 FE_OCP_RBC6198_FE_OFN789_n_46195 ( .a(FE_OCP_RBN6197_FE_OFN789_n_46195), .o(FE_OCP_RBN6198_FE_OFN789_n_46195) );
in01s02 FE_OCP_RBC6199_FE_OFN789_n_46195 ( .a(FE_OCP_RBN6197_FE_OFN789_n_46195), .o(FE_OCP_RBN6199_FE_OFN789_n_46195) );
in01s02 FE_OCP_RBC6200_FE_OFN789_n_46195 ( .a(FE_OCP_RBN6197_FE_OFN789_n_46195), .o(FE_OCP_RBN6200_FE_OFN789_n_46195) );
in01s02 FE_OCP_RBC6201_FE_OFN789_n_46195 ( .a(FE_OCP_RBN6197_FE_OFN789_n_46195), .o(FE_OCP_RBN6201_FE_OFN789_n_46195) );
in01s06 FE_OCP_RBC6202_n_31819 ( .a(FE_OCP_RBN3390_n_31819), .o(FE_OCP_RBN6202_n_31819) );
in01s04 FE_OCP_RBC6203_n_31819 ( .a(FE_OCP_RBN3390_n_31819), .o(FE_OCP_RBN6203_n_31819) );
in01s01 FE_OCP_RBC6204_n_31819 ( .a(FE_OCP_RBN6202_n_31819), .o(FE_OCP_RBN6204_n_31819) );
in01s02 FE_OCP_RBC6207_n_11486 ( .a(n_11486), .o(FE_OCP_RBN6207_n_11486) );
in01s02 FE_OCP_RBC6208_n_11486 ( .a(n_11486), .o(FE_OCP_RBN6208_n_11486) );
in01s06 FE_OCP_RBC6209_n_11486 ( .a(n_11486), .o(FE_OCP_RBN6209_n_11486) );
in01f02 FE_OCP_RBC6211_n_22421 ( .a(n_22421), .o(FE_OCP_RBN6211_n_22421) );
in01s01 FE_OCP_RBC6212_n_16962 ( .a(n_16962), .o(FE_OCP_RBN6212_n_16962) );
in01s02 FE_OCP_RBC6213_n_27086 ( .a(n_27086), .o(FE_OCP_RBN6213_n_27086) );
in01s02 FE_OCP_RBC6214_n_27086 ( .a(n_27086), .o(FE_OCP_RBN6214_n_27086) );
in01s03 FE_OCP_RBC6216_n_27086 ( .a(n_27086), .o(FE_OCP_RBN6216_n_27086) );
in01m08 FE_OCP_RBC6217_n_27110 ( .a(n_27110), .o(FE_OCP_RBN6217_n_27110) );
in01s06 FE_OCP_RBC6218_n_27110 ( .a(FE_OCP_RBN6217_n_27110), .o(FE_OCP_RBN6218_n_27110) );
in01f03 FE_OCP_RBC6219_n_27110 ( .a(FE_OCP_RBN6217_n_27110), .o(FE_OCP_RBN6219_n_27110) );
in01s01 FE_OCP_RBC6220_n_27110 ( .a(FE_OCP_RBN6217_n_27110), .o(FE_OCP_RBN6220_n_27110) );
in01s01 FE_OCP_RBC6221_n_27110 ( .a(FE_OCP_RBN6217_n_27110), .o(FE_OCP_RBN6221_n_27110) );
in01s01 FE_OCP_RBC6222_n_27110 ( .a(FE_OCP_RBN6220_n_27110), .o(FE_OCP_RBN6222_n_27110) );
in01s01 FE_OCP_RBC6223_n_27110 ( .a(FE_OCP_RBN6220_n_27110), .o(FE_OCP_RBN6223_n_27110) );
in01s01 FE_OCP_RBC6224_n_32061 ( .a(n_32061), .o(FE_OCP_RBN6224_n_32061) );
in01s01 FE_OCP_RBC6225_n_11713 ( .a(n_11713), .o(FE_OCP_RBN6225_n_11713) );
in01s01 FE_OCP_RBC6226_n_32178 ( .a(n_32178), .o(FE_OCP_RBN6226_n_32178) );
in01s01 FE_OCP_RBC6227_n_32216 ( .a(n_32216), .o(FE_OCP_RBN6227_n_32216) );
in01f02 FE_OCP_RBC6228_n_40565 ( .a(n_40565), .o(FE_OCP_RBN6228_n_40565) );
in01m02 FE_OCP_RBC6229_n_36693 ( .a(n_36693), .o(FE_OCP_RBN6229_n_36693) );
in01f02 FE_OCP_RBC6230_n_43882 ( .a(n_43882), .o(FE_OCP_RBN6230_n_43882) );
in01s02 FE_OCP_RBC6231_n_22639 ( .a(n_22639), .o(FE_OCP_RBN6231_n_22639) );
in01s04 FE_OCP_RBC6232_n_22639 ( .a(n_22639), .o(FE_OCP_RBN6232_n_22639) );
in01s01 FE_OCP_RBC6233_n_27504 ( .a(n_27504), .o(FE_OCP_RBN6233_n_27504) );
in01s01 FE_OCP_RBC6234_n_36778 ( .a(n_36778), .o(FE_OCP_RBN6234_n_36778) );
in01s01 FE_OCP_RBC6235_n_36780 ( .a(n_36780), .o(FE_OCP_RBN6235_n_36780) );
in01f02 FE_OCP_RBC6236_n_40586 ( .a(n_40586), .o(FE_OCP_RBN6236_n_40586) );
in01m06 FE_OCP_RBC6237_n_11853 ( .a(n_11853), .o(FE_OCP_RBN6237_n_11853) );
in01s02 FE_OCP_RBC6238_n_22718 ( .a(n_22718), .o(FE_OCP_RBN6238_n_22718) );
in01s02 FE_OCP_RBC6239_n_6456 ( .a(n_6456), .o(FE_OCP_RBN6239_n_6456) );
in01s01 FE_OCP_RBC6240_n_6438 ( .a(n_6438), .o(FE_OCP_RBN6240_n_6438) );
in01f02 FE_OCP_RBC6241_n_22622 ( .a(n_22622), .o(FE_OCP_RBN6241_n_22622) );
in01m02 FE_OCP_RBC6242_n_27436 ( .a(n_27436), .o(FE_OCP_RBN6242_n_27436) );
in01s02 FE_OCP_RBC6243_n_32305 ( .a(n_32305), .o(FE_OCP_RBN6243_n_32305) );
in01f02 FE_OCP_RBC6244_n_6535 ( .a(n_6535), .o(FE_OCP_RBN6244_n_6535) );
in01s02 FE_OCP_RBC6245_n_17587 ( .a(n_17587), .o(FE_OCP_RBN6245_n_17587) );
in01s01 FE_OCP_RBC6246_n_17587 ( .a(n_17587), .o(FE_OCP_RBN6246_n_17587) );
in01s01 FE_OCP_RBC6247_n_6477 ( .a(n_6477), .o(FE_OCP_RBN6247_n_6477) );
in01m02 FE_OCP_RBC6248_n_6477 ( .a(n_6477), .o(FE_OCP_RBN6248_n_6477) );
in01s01 FE_OCP_RBC6249_n_6567 ( .a(n_6567), .o(FE_OCP_RBN6249_n_6567) );
in01s01 FE_OCP_RBC6250_n_6567 ( .a(n_6567), .o(FE_OCP_RBN6250_n_6567) );
in01s02 FE_OCP_RBC6251_n_12067 ( .a(n_12067), .o(FE_OCP_RBN6251_n_12067) );
in01s01 FE_OCP_RBC6252_n_12067 ( .a(n_12067), .o(FE_OCP_RBN6252_n_12067) );
in01m02 FE_OCP_RBC6253_n_12117 ( .a(n_12117), .o(FE_OCP_RBN6253_n_12117) );
in01s01 FE_OCP_RBC6254_n_17723 ( .a(n_17723), .o(FE_OCP_RBN6254_n_17723) );
in01m02 FE_OCP_RBC6255_FE_RN_1283_0 ( .a(FE_RN_1283_0), .o(FE_OCP_RBN6255_FE_RN_1283_0) );
in01m02 FE_OCP_RBC6256_FE_RN_2452_0 ( .a(FE_RN_2452_0), .o(FE_OCP_RBN6256_FE_RN_2452_0) );
in01s02 FE_OCP_RBC6257_n_43842 ( .a(n_43842), .o(FE_OCP_RBN6257_n_43842) );
in01s02 FE_OCP_RBC6258_n_27743 ( .a(n_27743), .o(FE_OCP_RBN6258_n_27743) );
in01m02 FE_OCP_RBC6259_n_27726 ( .a(n_27726), .o(FE_OCP_RBN6259_n_27726) );
in01m10 FE_OCP_RBC6307_n_45224 ( .a(n_45224), .o(FE_OCP_RBN6307_n_45224) );
in01s10 FE_OCP_RBC6308_n_45224 ( .a(n_45224), .o(FE_OCP_RBN6308_n_45224) );
in01s10 FE_OCP_RBC6309_n_45224 ( .a(FE_OCP_RBN6311_n_45224), .o(FE_OCP_RBN6309_n_45224) );
in01s20 FE_OCP_RBC6310_n_45224 ( .a(FE_OCP_RBN6311_n_45224), .o(FE_OCP_RBN6310_n_45224) );
in01s20 FE_OCP_RBC6311_n_45224 ( .a(n_45224), .o(FE_OCP_RBN6311_n_45224) );
in01s06 FE_OCP_RBC6312_n_45224 ( .a(n_45224), .o(FE_OCP_RBN6312_n_45224) );
in01s06 FE_OCP_RBC6313_n_45224 ( .a(FE_OCP_RBN6315_n_45224), .o(FE_OCP_RBN6313_n_45224) );
in01s20 FE_OCP_RBC6314_n_45224 ( .a(FE_OCP_RBN6315_n_45224), .o(FE_OCP_RBN6314_n_45224) );
in01s20 FE_OCP_RBC6315_n_45224 ( .a(n_45224), .o(FE_OCP_RBN6315_n_45224) );
in01s10 FE_OCP_RBC6316_n_45224 ( .a(n_45224), .o(FE_OCP_RBN6316_n_45224) );
in01s08 FE_OCP_RBC6317_n_45224 ( .a(n_45224), .o(FE_OCP_RBN6317_n_45224) );
in01s10 FE_OCP_RBC6318_n_45224 ( .a(n_45224), .o(FE_OCP_RBN6318_n_45224) );
in01m08 FE_OCP_RBC6319_n_45224 ( .a(n_45224), .o(FE_OCP_RBN6319_n_45224) );
in01s10 FE_OCP_RBC6320_n_45224 ( .a(n_45224), .o(FE_OCP_RBN6320_n_45224) );
in01s04 FE_OCP_RBC6321_n_45224 ( .a(n_45224), .o(FE_OCP_RBN6321_n_45224) );
in01s01 FE_OCP_RBC6369_n_27773 ( .a(n_27773), .o(FE_OCP_RBN6369_n_27773) );
in01s04 FE_OCP_RBC6370_n_17582 ( .a(n_17582), .o(FE_OCP_RBN6370_n_17582) );
in01s02 FE_OCP_RBC6371_FE_RN_1425_0 ( .a(FE_RN_1425_0), .o(FE_OCP_RBN6371_FE_RN_1425_0) );
in01f02 FE_OCP_RBC6372_FE_RN_1425_0 ( .a(FE_RN_1425_0), .o(FE_OCP_RBN6372_FE_RN_1425_0) );
in01s01 FE_OCP_RBC6373_n_19701 ( .a(n_19701), .o(FE_OCP_RBN6373_n_19701) );
in01m01 FE_OCP_RBC6374_n_19722 ( .a(n_19722), .o(FE_OCP_RBN6374_n_19722) );
in01s02 FE_OCP_RBC6375_n_14154 ( .a(n_14154), .o(FE_OCP_RBN6375_n_14154) );
in01s02 FE_OCP_RBC6376_n_14154 ( .a(n_14154), .o(FE_OCP_RBN6376_n_14154) );
in01m02 FE_OCP_RBC6377_n_14380 ( .a(n_14380), .o(FE_OCP_RBN6377_n_14380) );
in01m02 FE_OCP_RBC6378_n_14380 ( .a(n_14380), .o(FE_OCP_RBN6378_n_14380) );
in01m04 FE_OCP_RBC6379_n_14380 ( .a(FE_OCP_RBN6377_n_14380), .o(FE_OCP_RBN6379_n_14380) );
in01s02 FE_OCP_RBC6380_n_20125 ( .a(n_20125), .o(FE_OCP_RBN6380_n_20125) );
in01m02 FE_OCP_RBC6381_n_30824 ( .a(n_30824), .o(FE_OCP_RBN6381_n_30824) );
in01f02 FE_OCP_RBC6382_n_21087 ( .a(n_21087), .o(FE_OCP_RBN6382_n_21087) );
in01s01 FE_OCP_RBC6383_n_21087 ( .a(n_21087), .o(FE_OCP_RBN6383_n_21087) );
in01s01 FE_OCP_RBC6384_n_21087 ( .a(FE_OCP_RBN6383_n_21087), .o(FE_OCP_RBN6384_n_21087) );
in01s04 FE_OCP_RBC6385_n_21429 ( .a(n_21429), .o(FE_OCP_RBN6385_n_21429) );
in01m04 FE_OCP_RBC6386_n_21429 ( .a(FE_OCP_RBN6385_n_21429), .o(FE_OCP_RBN6386_n_21429) );
in01m10 FE_OCP_RBC6387_n_32238 ( .a(n_32238), .o(FE_OCP_RBN6387_n_32238) );
in01s03 FE_OCP_RBC6388_n_32238 ( .a(n_32238), .o(FE_OCP_RBN6388_n_32238) );
in01m06 FE_OCP_RBC6407_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN6407_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s40 FE_OCP_RBC6408_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN6408_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01m06 FE_OCP_RBC6409_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN6409_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s03 FE_OCP_RBC6410_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN6410_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s06 FE_OCP_RBC6413_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN6413_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s20 FE_OCP_RBC6435_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN6435_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01m10 FE_OCP_RBC6438_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN6438_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01s06 FE_OCP_RBC6439_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN6439_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01s20 FE_OCP_RBC6440_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN6440_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01s40 FE_OCP_RBC6442_delay_sub_ln23_unr9_stage4_stallmux_q_3_ ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(FE_OCP_RBN6442_delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
in01s40 FE_OCP_RBC6444_delay_xor_ln21_unr9_stage4_stallmux_q_1_ ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_1_), .o(FE_OCP_RBN6444_delay_xor_ln21_unr9_stage4_stallmux_q_1_) );
in01s10 FE_OCP_RBC6463_n_44061 ( .a(n_44061), .o(FE_OCP_RBN6463_n_44061) );
in01s03 FE_OCP_RBC6464_n_44061 ( .a(FE_OCP_RBN6465_n_44061), .o(FE_OCP_RBN6464_n_44061) );
in01s03 FE_OCP_RBC6465_n_44061 ( .a(n_44061), .o(FE_OCP_RBN6465_n_44061) );
in01s10 FE_OCP_RBC6466_n_44061 ( .a(n_44061), .o(FE_OCP_RBN6466_n_44061) );
in01s80 FE_OCP_RBC6467_n_44061 ( .a(FE_OCP_RBN6468_n_44061), .o(FE_OCP_RBN6467_n_44061) );
in01s40 FE_OCP_RBC6468_n_44061 ( .a(n_44061), .o(FE_OCP_RBN6468_n_44061) );
in01m40 FE_OCP_RBC6471_delay_xor_ln21_unr15_stage6_stallmux_q_3_ ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_3_), .o(FE_OCP_RBN6471_delay_xor_ln21_unr15_stage6_stallmux_q_3_) );
in01s06 FE_OCP_RBC6499_n_44610 ( .a(n_44610), .o(FE_OCP_RBN6499_n_44610) );
in01s06 FE_OCP_RBC6500_n_44610 ( .a(n_44610), .o(FE_OCP_RBN6500_n_44610) );
in01s06 FE_OCP_RBC6501_n_44610 ( .a(n_44610), .o(FE_OCP_RBN6501_n_44610) );
in01s06 FE_OCP_RBC6502_n_44610 ( .a(FE_OCP_RBN6501_n_44610), .o(FE_OCP_RBN6502_n_44610) );
in01s10 FE_OCP_RBC6503_n_44610 ( .a(FE_OCP_RBN6502_n_44610), .o(FE_OCP_RBN6503_n_44610) );
in01s40 FE_OCP_RBC6506_delay_add_ln22_unr23_stage9_stallmux_q_24_ ( .a(delay_add_ln22_unr23_stage9_stallmux_q_24_), .o(FE_OCP_RBN6506_delay_add_ln22_unr23_stage9_stallmux_q_24_) );
in01s10 FE_OCP_RBC6507_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN6438_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN6507_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01s20 FE_OCP_RBC6508_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN6507_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN6508_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01s10 FE_OCP_RBC6509_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN6508_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN6509_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01s20 FE_OCP_RBC6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN6509_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01s02 FE_OCP_RBC6511_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN6511_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01s02 FE_OCP_RBC6512_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN6511_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN6512_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01s01 FE_OCP_RBC6513_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN6413_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN6513_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s01 FE_OCP_RBC6514_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN6413_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN6514_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s06 FE_OCP_RBC6515_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN6413_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN6515_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01s06 FE_OCP_RBC6516_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN6515_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN6516_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01m03 FE_OCP_RBC6517_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN6515_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN6517_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01m10 FE_OCP_RBC6518_n_32706 ( .a(n_32706), .o(FE_OCP_RBN6518_n_32706) );
in01s10 FE_OCP_RBC6519_n_32706 ( .a(n_32706), .o(FE_OCP_RBN6519_n_32706) );
in01s10 FE_OCP_RBC6520_n_32706 ( .a(FE_OCP_RBN6519_n_32706), .o(FE_OCP_RBN6520_n_32706) );
in01s01 FE_OCP_RBC6521_n_32706 ( .a(FE_OCP_RBN6520_n_32706), .o(FE_OCP_RBN6521_n_32706) );
in01m06 FE_OCP_RBC6523_n_45224 ( .a(FE_OCP_RBN6310_n_45224), .o(FE_OCP_RBN6523_n_45224) );
in01s01 FE_OCP_RBC6524_n_6649 ( .a(n_6649), .o(FE_OCP_RBN6524_n_6649) );
in01s06 FE_OCP_RBC6525_n_11829 ( .a(n_11829), .o(FE_OCP_RBN6525_n_11829) );
in01s20 FE_OCP_RBC6526_n_44962 ( .a(FE_OCP_RBN4630_n_44962), .o(FE_OCP_RBN6526_n_44962) );
in01s40 FE_OCP_RBC6527_n_44962 ( .a(FE_OCP_RBN4630_n_44962), .o(FE_OCP_RBN6527_n_44962) );
in01s02 FE_OCP_RBC6528_n_6745 ( .a(n_6745), .o(FE_OCP_RBN6528_n_6745) );
in01s01 FE_OCP_RBC6529_n_6745 ( .a(n_6745), .o(FE_OCP_RBN6529_n_6745) );
in01m10 FE_OCP_RBC6530_n_22822 ( .a(n_22822), .o(FE_OCP_RBN6530_n_22822) );
in01s06 FE_OCP_RBC6531_n_11780 ( .a(n_11780), .o(FE_OCP_RBN6531_n_11780) );
in01m20 FE_OCP_RBC6532_n_32791 ( .a(n_32791), .o(FE_OCP_RBN6532_n_32791) );
in01s02 FE_OCP_RBC6533_n_32436 ( .a(FE_OCP_RBN5517_n_32436), .o(FE_OCP_RBN6533_n_32436) );
in01s01 FE_OCP_RBC6534_n_1577 ( .a(n_1577), .o(FE_OCP_RBN6534_n_1577) );
in01m08 FE_OCP_RBC6535_n_1602 ( .a(n_1602), .o(FE_OCP_RBN6535_n_1602) );
in01s01 FE_OCP_RBC6536_n_1602 ( .a(n_1602), .o(FE_OCP_RBN6536_n_1602) );
in01s01 FE_OCP_RBC6537_n_1614 ( .a(n_1614), .o(FE_OCP_RBN6537_n_1614) );
in01m10 FE_OCP_RBC6538_n_1614 ( .a(n_1614), .o(FE_OCP_RBN6538_n_1614) );
in01s80 FE_OCP_RBC6539_n_44083 ( .a(FE_OCP_RBN5537_n_44083), .o(FE_OCP_RBN6539_n_44083) );
in01s80 FE_OCP_RBC6540_n_44083 ( .a(FE_OCP_RBN6539_n_44083), .o(FE_OCP_RBN6540_n_44083) );
in01s40 FE_OCP_RBC6541_n_44083 ( .a(FE_OCP_RBN6539_n_44083), .o(FE_OCP_RBN6541_n_44083) );
in01f04 FE_OCP_RBC6542_n_23186 ( .a(n_23186), .o(FE_OCP_RBN6542_n_23186) );
in01s10 FE_OCP_RBC6543_n_45145 ( .a(FE_OCP_RBN5546_n_45145), .o(FE_OCP_RBN6543_n_45145) );
in01s10 FE_OCP_RBC6544_n_45145 ( .a(FE_OCP_RBN5546_n_45145), .o(FE_OCP_RBN6544_n_45145) );
in01m08 FE_OCP_RBC6545_n_1672 ( .a(n_1672), .o(FE_OCP_RBN6545_n_1672) );
in01s01 FE_OCP_RBC6546_n_1672 ( .a(n_1672), .o(FE_OCP_RBN6546_n_1672) );
in01m04 FE_OCP_RBC6547_n_1725 ( .a(n_1725), .o(FE_OCP_RBN6547_n_1725) );
in01s01 FE_OCP_RBC6548_n_1725 ( .a(n_1725), .o(FE_OCP_RBN6548_n_1725) );
in01m02 FE_OCP_RBC6549_n_37377 ( .a(n_37377), .o(FE_OCP_RBN6549_n_37377) );
in01m06 FE_OCP_RBC6550_n_37377 ( .a(n_37377), .o(FE_OCP_RBN6550_n_37377) );
in01s01 FE_OCP_RBC6551_n_1905 ( .a(n_1905), .o(FE_OCP_RBN6551_n_1905) );
in01s01 FE_OCP_RBC6552_n_28458 ( .a(FE_OCP_RBN4028_n_28458), .o(FE_OCP_RBN6552_n_28458) );
in01s20 FE_OCP_RBC6553_n_28458 ( .a(FE_OCP_RBN4028_n_28458), .o(FE_OCP_RBN6553_n_28458) );
in01s20 FE_OCP_RBC6554_n_28458 ( .a(FE_OCP_RBN6553_n_28458), .o(FE_OCP_RBN6554_n_28458) );
in01s02 FE_OCP_RBC6555_n_28458 ( .a(FE_OCP_RBN6553_n_28458), .o(FE_OCP_RBN6555_n_28458) );
in01s02 FE_OCP_RBC6556_n_28458 ( .a(FE_OCP_RBN6553_n_28458), .o(FE_OCP_RBN6556_n_28458) );
in01m08 FE_OCP_RBC6557_n_23572 ( .a(n_23572), .o(FE_OCP_RBN6557_n_23572) );
in01m02 FE_OCP_RBC6558_n_23572 ( .a(FE_OCP_RBN6557_n_23572), .o(FE_OCP_RBN6558_n_23572) );
in01s01 FE_OCP_RBC6559_n_23572 ( .a(FE_OCP_RBN6557_n_23572), .o(FE_OCP_RBN6559_n_23572) );
in01s06 FE_OCP_RBC6560_n_23572 ( .a(FE_OCP_RBN6558_n_23572), .o(FE_OCP_RBN6560_n_23572) );
in01s06 FE_OCP_RBC6561_n_33208 ( .a(n_33208), .o(FE_OCP_RBN6561_n_33208) );
in01s06 FE_OCP_RBC6562_n_33208 ( .a(FE_OCP_RBN6561_n_33208), .o(FE_OCP_RBN6562_n_33208) );
in01s01 FE_OCP_RBC6563_n_12753 ( .a(n_12753), .o(FE_OCP_RBN6563_n_12753) );
in01f10 FE_OCP_RBC6564_n_12753 ( .a(n_12753), .o(FE_OCP_RBN6564_n_12753) );
in01f08 FE_OCP_RBC6565_n_12753 ( .a(FE_OCP_RBN6564_n_12753), .o(FE_OCP_RBN6565_n_12753) );
in01s02 FE_OCP_RBC6566_n_33368 ( .a(n_33368), .o(FE_OCP_RBN6566_n_33368) );
in01m02 FE_OCP_RBC6567_n_12714 ( .a(n_12714), .o(FE_OCP_RBN6567_n_12714) );
in01s01 FE_OCP_RBC6568_n_33803 ( .a(n_33803), .o(FE_OCP_RBN6568_n_33803) );
in01f02 FE_OCP_RBC6569_n_33803 ( .a(n_33803), .o(FE_OCP_RBN6569_n_33803) );
in01s01 FE_OCP_RBC6570_n_44875 ( .a(FE_OCP_RBN5600_n_44875), .o(FE_OCP_RBN6570_n_44875) );
in01s10 FE_OCP_RBC6571_n_44875 ( .a(FE_OCP_RBN5600_n_44875), .o(FE_OCP_RBN6571_n_44875) );
in01s06 FE_OCP_RBC6572_n_44875 ( .a(FE_OCP_RBN5600_n_44875), .o(FE_OCP_RBN6572_n_44875) );
in01s03 FE_OCP_RBC6573_n_44875 ( .a(FE_OCP_RBN6572_n_44875), .o(FE_OCP_RBN6573_n_44875) );
in01s01 FE_OCP_RBC6574_n_44875 ( .a(FE_OCP_RBN6572_n_44875), .o(FE_OCP_RBN6574_n_44875) );
in01s06 FE_OCP_RBC6575_n_44875 ( .a(FE_OCP_RBN6573_n_44875), .o(FE_OCP_RBN6575_n_44875) );
in01m02 FE_OCP_RBC6576_n_13011 ( .a(n_13011), .o(FE_OCP_RBN6576_n_13011) );
in01f04 FE_OCP_RBC6577_n_13011 ( .a(n_13011), .o(FE_OCP_RBN6577_n_13011) );
in01s01 FE_OCP_RBC6578_n_8676 ( .a(n_8676), .o(FE_OCP_RBN6578_n_8676) );
in01s01 FE_OCP_RBC6579_n_8676 ( .a(n_8676), .o(FE_OCP_RBN6579_n_8676) );
in01s01 FE_OCP_RBC6580_n_8676 ( .a(FE_OCP_RBN6578_n_8676), .o(FE_OCP_RBN6580_n_8676) );
in01s01 FE_OCP_RBC6581_n_8021 ( .a(n_8021), .o(FE_OCP_RBN6581_n_8021) );
in01s01 FE_OCP_RBC6582_n_8021 ( .a(FE_OCP_RBN6581_n_8021), .o(FE_OCP_RBN6582_n_8021) );
in01s01 FE_OCP_RBC6583_n_8021 ( .a(FE_OCP_RBN6581_n_8021), .o(FE_OCP_RBN6583_n_8021) );
in01s03 FE_OCP_RBC6584_n_41491 ( .a(n_41491), .o(FE_OCP_RBN6584_n_41491) );
in01s01 FE_OCP_RBC6585_n_41491 ( .a(n_41491), .o(FE_OCP_RBN6585_n_41491) );
in01s02 FE_OCP_RBC6586_n_41491 ( .a(n_41491), .o(FE_OCP_RBN6586_n_41491) );
in01s02 FE_OCP_RBC6587_n_41491 ( .a(n_41491), .o(FE_OCP_RBN6587_n_41491) );
in01s04 FE_OCP_RBC6588_n_41491 ( .a(n_41491), .o(FE_OCP_RBN6588_n_41491) );
in01s02 FE_OCP_RBC6589_n_41491 ( .a(n_41491), .o(FE_OCP_RBN6589_n_41491) );
in01s03 FE_OCP_RBC6590_n_41491 ( .a(FE_OCP_RBN6584_n_41491), .o(FE_OCP_RBN6590_n_41491) );
in01s02 FE_OCP_RBC6591_n_41491 ( .a(FE_OCP_RBN6584_n_41491), .o(FE_OCP_RBN6591_n_41491) );
in01s06 FE_OCP_RBC6592_n_41491 ( .a(FE_OCP_RBN6588_n_41491), .o(FE_OCP_RBN6592_n_41491) );
in01s01 FE_OCP_RBC6593_n_41491 ( .a(FE_OCP_RBN6589_n_41491), .o(FE_OCP_RBN6593_n_41491) );
in01s01 FE_OCP_RBC6594_n_41491 ( .a(FE_OCP_RBN6593_n_41491), .o(FE_OCP_RBN6594_n_41491) );
in01s01 FE_OCP_RBC6595_n_41491 ( .a(FE_OCP_RBN6593_n_41491), .o(FE_OCP_RBN6595_n_41491) );
in01s01 FE_OCP_RBC6596_n_7708 ( .a(FE_OCP_RBN4075_n_7708), .o(FE_OCP_RBN6596_n_7708) );
in01s06 FE_OCP_RBC6597_n_7708 ( .a(FE_OCP_RBN4075_n_7708), .o(FE_OCP_RBN6597_n_7708) );
in01s01 FE_OCP_RBC6598_n_7708 ( .a(FE_OCP_RBN4075_n_7708), .o(FE_OCP_RBN6598_n_7708) );
in01m02 FE_OCP_RBC6599_n_7708 ( .a(FE_OCP_RBN4075_n_7708), .o(FE_OCP_RBN6599_n_7708) );
in01s10 FE_OCP_RBC6600_n_7708 ( .a(FE_OCP_RBN6597_n_7708), .o(FE_OCP_RBN6600_n_7708) );
in01s06 FE_OCP_RBC6601_n_7708 ( .a(FE_OCP_RBN6599_n_7708), .o(FE_OCP_RBN6601_n_7708) );
in01s01 FE_OCP_RBC6602_n_7881 ( .a(n_7881), .o(FE_OCP_RBN6602_n_7881) );
in01s01 FE_OCP_RBC6603_n_7881 ( .a(FE_OCP_RBN6602_n_7881), .o(FE_OCP_RBN6603_n_7881) );
in01s01 FE_OCP_RBC6604_n_7881 ( .a(FE_OCP_RBN6602_n_7881), .o(FE_OCP_RBN6604_n_7881) );
in01s01 FE_OCP_RBC6605_n_7881 ( .a(FE_OCP_RBN6603_n_7881), .o(FE_OCP_RBN6605_n_7881) );
in01s06 FE_OCP_RBC6606_n_2289 ( .a(FE_OCP_RBN4073_n_2289), .o(FE_OCP_RBN6606_n_2289) );
in01s10 FE_OCP_RBC6607_n_2289 ( .a(FE_OCP_RBN4073_n_2289), .o(FE_OCP_RBN6607_n_2289) );
in01s01 FE_OCP_RBC6608_n_2289 ( .a(FE_OCP_RBN6606_n_2289), .o(FE_OCP_RBN6608_n_2289) );
in01s01 FE_OCP_RBC6609_n_2289 ( .a(FE_OCP_RBN6606_n_2289), .o(FE_OCP_RBN6609_n_2289) );
in01s06 FE_OCP_RBC6610_n_2289 ( .a(FE_OCP_RBN6607_n_2289), .o(FE_OCP_RBN6610_n_2289) );
in01s10 FE_OCP_RBC6611_n_2289 ( .a(FE_OCP_RBN6607_n_2289), .o(FE_OCP_RBN6611_n_2289) );
in01s01 FE_OCP_RBC6612_n_2289 ( .a(FE_OCP_RBN6608_n_2289), .o(FE_OCP_RBN6612_n_2289) );
in01s01 FE_OCP_RBC6613_n_2289 ( .a(FE_OCP_RBN6608_n_2289), .o(FE_OCP_RBN6613_n_2289) );
in01s01 FE_OCP_RBC6614_n_2289 ( .a(FE_OCP_RBN6608_n_2289), .o(FE_OCP_RBN6614_n_2289) );
in01s01 FE_OCP_RBC6615_n_2289 ( .a(FE_OCP_RBN6609_n_2289), .o(FE_OCP_RBN6615_n_2289) );
in01s01 FE_OCP_RBC6616_n_2289 ( .a(FE_OCP_RBN6609_n_2289), .o(FE_OCP_RBN6616_n_2289) );
in01s01 FE_OCP_RBC6617_n_2289 ( .a(FE_OCP_RBN6609_n_2289), .o(FE_OCP_RBN6617_n_2289) );
in01s02 FE_OCP_RBC6618_n_41381 ( .a(FE_OCP_RBN4115_n_41381), .o(FE_OCP_RBN6618_n_41381) );
in01s02 FE_OCP_RBC6619_n_41381 ( .a(FE_OCP_RBN4115_n_41381), .o(FE_OCP_RBN6619_n_41381) );
in01s01 FE_OCP_RBC6620_n_41381 ( .a(FE_OCP_RBN4115_n_41381), .o(FE_OCP_RBN6620_n_41381) );
in01s01 FE_OCP_RBC6621_n_7821 ( .a(n_7821), .o(FE_OCP_RBN6621_n_7821) );
in01s01 FE_OCP_RBC6622_n_7943 ( .a(n_7943), .o(FE_OCP_RBN6622_n_7943) );
in01s02 FE_OCP_RBC6623_n_24175 ( .a(FE_OCP_RBN1007_n_24175), .o(FE_OCP_RBN6623_n_24175) );
in01s01 FE_OCP_RBC6624_n_24175 ( .a(FE_OCP_RBN1007_n_24175), .o(FE_OCP_RBN6624_n_24175) );
in01m04 FE_OCP_RBC6625_n_2537 ( .a(n_2537), .o(FE_OCP_RBN6625_n_2537) );
in01s01 FE_OCP_RBC6626_n_2537 ( .a(n_2537), .o(FE_OCP_RBN6626_n_2537) );
in01s01 FE_OCP_RBC6627_n_7832 ( .a(n_7832), .o(FE_OCP_RBN6627_n_7832) );
in01s02 FE_OCP_RBC6628_n_8269 ( .a(n_8269), .o(FE_OCP_RBN6628_n_8269) );
in01s01 FE_OCP_RBC6629_n_8269 ( .a(n_8269), .o(FE_OCP_RBN6629_n_8269) );
in01s01 FE_OCP_RBC6630_n_8269 ( .a(n_8269), .o(FE_OCP_RBN6630_n_8269) );
in01m02 FE_OCP_RBC6631_n_8111 ( .a(n_8111), .o(FE_OCP_RBN6631_n_8111) );
in01m04 FE_OCP_RBC6632_n_2633 ( .a(n_2633), .o(FE_OCP_RBN6632_n_2633) );
in01s01 FE_OCP_RBC6633_n_2633 ( .a(n_2633), .o(FE_OCP_RBN6633_n_2633) );
in01s01 FE_OCP_RBC6634_n_9304 ( .a(n_9304), .o(FE_OCP_RBN6634_n_9304) );
in01s01 FE_OCP_RBC6635_n_9304 ( .a(n_9304), .o(FE_OCP_RBN6635_n_9304) );
in01s01 FE_OCP_RBC6636_n_33983 ( .a(n_33983), .o(FE_OCP_RBN6636_n_33983) );
in01f06 FE_OCP_RBC6637_n_33983 ( .a(n_33983), .o(FE_OCP_RBN6637_n_33983) );
in01s02 FE_OCP_RBC6638_n_13726 ( .a(FE_OCP_RBN5019_n_13726), .o(FE_OCP_RBN6638_n_13726) );
in01s01 FE_OCP_RBC6639_n_13726 ( .a(FE_OCP_RBN5019_n_13726), .o(FE_OCP_RBN6639_n_13726) );
in01s06 FE_OCP_RBC6640_n_24268 ( .a(n_24268), .o(FE_OCP_RBN6640_n_24268) );
in01s01 FE_OCP_RBC6641_n_3502 ( .a(n_3502), .o(FE_OCP_RBN6641_n_3502) );
in01s02 FE_OCP_RBC6642_n_3502 ( .a(n_3502), .o(FE_OCP_RBN6642_n_3502) );
in01s02 FE_OCP_RBC6643_n_8342 ( .a(n_8342), .o(FE_OCP_RBN6643_n_8342) );
in01s01 FE_OCP_RBC6644_n_8342 ( .a(n_8342), .o(FE_OCP_RBN6644_n_8342) );
in01s01 FE_OCP_RBC6645_n_8342 ( .a(FE_OCP_RBN6644_n_8342), .o(FE_OCP_RBN6645_n_8342) );
in01s02 FE_OCP_RBC6646_n_13818 ( .a(FE_OCP_RBN2684_n_13818), .o(FE_OCP_RBN6646_n_13818) );
in01s01 FE_OCP_RBC6647_n_13818 ( .a(FE_OCP_RBN2684_n_13818), .o(FE_OCP_RBN6647_n_13818) );
in01s01 FE_OCP_RBC6648_n_13818 ( .a(FE_OCP_RBN6646_n_13818), .o(FE_OCP_RBN6648_n_13818) );
in01s01 FE_OCP_RBC6649_n_13818 ( .a(FE_OCP_RBN6647_n_13818), .o(FE_OCP_RBN6649_n_13818) );
in01s01 FE_OCP_RBC6650_n_13818 ( .a(FE_OCP_RBN6648_n_13818), .o(FE_OCP_RBN6650_n_13818) );
in01s01 FE_OCP_RBC6651_n_13818 ( .a(FE_OCP_RBN6648_n_13818), .o(FE_OCP_RBN6651_n_13818) );
in01s01 FE_OCP_RBC6652_n_29494 ( .a(n_29494), .o(FE_OCP_RBN6652_n_29494) );
in01f04 FE_OCP_RBC6653_n_29494 ( .a(n_29494), .o(FE_OCP_RBN6653_n_29494) );
in01s02 FE_OCP_RBC6654_n_8187 ( .a(n_8187), .o(FE_OCP_RBN6654_n_8187) );
in01s01 FE_OCP_RBC6655_n_8187 ( .a(n_8187), .o(FE_OCP_RBN6655_n_8187) );
in01s01 FE_OCP_RBC6656_n_8187 ( .a(FE_OCP_RBN6655_n_8187), .o(FE_OCP_RBN6656_n_8187) );
in01s02 FE_OCP_RBC6657_n_44352 ( .a(n_44352), .o(FE_OCP_RBN6657_n_44352) );
in01s02 FE_OCP_RBC6658_n_44352 ( .a(n_44352), .o(FE_OCP_RBN6658_n_44352) );
in01s01 FE_OCP_RBC6659_n_2829 ( .a(n_2829), .o(FE_OCP_RBN6659_n_2829) );
in01s02 FE_OCP_RBC6660_n_13884 ( .a(n_13884), .o(FE_OCP_RBN6660_n_13884) );
in01m02 FE_OCP_RBC6661_n_13702 ( .a(n_13702), .o(FE_OCP_RBN6661_n_13702) );
in01f04 FE_OCP_RBC6662_n_13702 ( .a(n_13702), .o(FE_OCP_RBN6662_n_13702) );
in01s02 FE_OCP_RBC6663_n_8355 ( .a(n_8355), .o(FE_OCP_RBN6663_n_8355) );
in01s08 FE_OCP_RBC6664_n_34297 ( .a(n_34297), .o(FE_OCP_RBN6664_n_34297) );
in01m04 FE_OCP_RBC6665_n_34297 ( .a(n_34297), .o(FE_OCP_RBN6665_n_34297) );
in01s03 FE_OCP_RBC6666_n_34297 ( .a(n_34297), .o(FE_OCP_RBN6666_n_34297) );
in01s01 FE_OCP_RBC6667_n_34297 ( .a(FE_OCP_RBN6664_n_34297), .o(FE_OCP_RBN6667_n_34297) );
in01s10 FE_OCP_RBC6668_n_34297 ( .a(FE_OCP_RBN6664_n_34297), .o(FE_OCP_RBN6668_n_34297) );
in01s02 FE_OCP_RBC6669_n_34297 ( .a(FE_OCP_RBN6665_n_34297), .o(FE_OCP_RBN6669_n_34297) );
in01s01 FE_OCP_RBC6670_n_34297 ( .a(FE_OCP_RBN6666_n_34297), .o(FE_OCP_RBN6670_n_34297) );
in01s02 FE_OCP_RBC6671_n_34297 ( .a(FE_OCP_RBN6669_n_34297), .o(FE_OCP_RBN6671_n_34297) );
in01s01 FE_OCP_RBC6672_n_34297 ( .a(FE_OCP_RBN6670_n_34297), .o(FE_OCP_RBN6672_n_34297) );
in01s01 FE_OCP_RBC6673_n_34297 ( .a(FE_OCP_RBN6670_n_34297), .o(FE_OCP_RBN6673_n_34297) );
in01f02 FE_OCP_RBC6674_n_38519 ( .a(n_38519), .o(FE_OCP_RBN6674_n_38519) );
in01s01 FE_OCP_RBC6675_n_8288 ( .a(FE_OCP_RBN4186_n_8288), .o(FE_OCP_RBN6675_n_8288) );
in01s01 FE_OCP_RBC6676_n_8288 ( .a(FE_OCP_RBN4186_n_8288), .o(FE_OCP_RBN6676_n_8288) );
in01s01 FE_OCP_RBC6677_n_8288 ( .a(FE_OCP_RBN6676_n_8288), .o(FE_OCP_RBN6677_n_8288) );
in01s01 FE_OCP_RBC6678_n_8288 ( .a(FE_OCP_RBN6677_n_8288), .o(FE_OCP_RBN6678_n_8288) );
in01s01 FE_OCP_RBC6679_n_8288 ( .a(FE_OCP_RBN6677_n_8288), .o(FE_OCP_RBN6679_n_8288) );
in01f02 FE_OCP_RBC6680_n_8448 ( .a(n_8448), .o(FE_OCP_RBN6680_n_8448) );
in01m06 FE_OCP_RBC6681_n_24648 ( .a(n_24648), .o(FE_OCP_RBN6681_n_24648) );
in01s01 FE_OCP_RBC6682_FE_OCPN4529_FE_OCP_RBN2748_n_8474 ( .a(FE_OCPN4529_FE_OCP_RBN2748_n_8474), .o(FE_OCP_RBN6682_FE_OCPN4529_FE_OCP_RBN2748_n_8474) );
in01s01 FE_OCP_RBC6683_FE_OCPN4529_FE_OCP_RBN2748_n_8474 ( .a(FE_OCPN4529_FE_OCP_RBN2748_n_8474), .o(FE_OCP_RBN6683_FE_OCPN4529_FE_OCP_RBN2748_n_8474) );
in01s01 FE_OCP_RBC6684_FE_OCPN4529_FE_OCP_RBN2748_n_8474 ( .a(FE_OCP_RBN6682_FE_OCPN4529_FE_OCP_RBN2748_n_8474), .o(FE_OCP_RBN6684_FE_OCPN4529_FE_OCP_RBN2748_n_8474) );
in01s01 FE_OCP_RBC6685_FE_OCPN4529_FE_OCP_RBN2748_n_8474 ( .a(FE_OCP_RBN6684_FE_OCPN4529_FE_OCP_RBN2748_n_8474), .o(FE_OCP_RBN6685_FE_OCPN4529_FE_OCP_RBN2748_n_8474) );
in01s02 FE_OCP_RBC6686_n_3498 ( .a(n_3498), .o(FE_OCP_RBN6686_n_3498) );
in01s01 FE_OCP_RBC6687_n_3498 ( .a(n_3498), .o(FE_OCP_RBN6687_n_3498) );
in01s01 FE_OCP_RBC6688_n_3498 ( .a(FE_OCP_RBN6687_n_3498), .o(FE_OCP_RBN6688_n_3498) );
in01s03 FE_OCP_RBC6689_n_38655 ( .a(n_38655), .o(FE_OCP_RBN6689_n_38655) );
in01m02 FE_OCP_RBC6690_n_38655 ( .a(n_38655), .o(FE_OCP_RBN6690_n_38655) );
in01s01 FE_OCP_RBC6691_n_8629 ( .a(n_8629), .o(FE_OCP_RBN6691_n_8629) );
in01m06 FE_OCP_RBC6692_n_13796 ( .a(FE_OCP_RBN4203_n_13796), .o(FE_OCP_RBN6692_n_13796) );
in01s40 FE_OCP_RBC6693_n_13796 ( .a(FE_OCP_RBN6692_n_13796), .o(FE_OCP_RBN6693_n_13796) );
in01s01 FE_OCP_RBC6694_n_13796 ( .a(FE_OCP_RBN4205_n_13796), .o(FE_OCP_RBN6694_n_13796) );
in01m10 FE_OCP_RBC6695_n_13796 ( .a(FE_OCP_RBN4205_n_13796), .o(FE_OCP_RBN6695_n_13796) );
in01s10 FE_OCP_RBC6696_n_13796 ( .a(FE_OCP_RBN6695_n_13796), .o(FE_OCP_RBN6696_n_13796) );
in01s01 FE_OCP_RBC6697_n_13796 ( .a(FE_OCP_RBN6695_n_13796), .o(FE_OCP_RBN6697_n_13796) );
in01s01 FE_OCP_RBC6698_n_13796 ( .a(FE_OCP_RBN6695_n_13796), .o(FE_OCP_RBN6698_n_13796) );
in01s01 FE_OCP_RBC6699_n_13796 ( .a(FE_OCP_RBN6697_n_13796), .o(FE_OCP_RBN6699_n_13796) );
in01s01 FE_OCP_RBC6700_n_13796 ( .a(FE_OCP_RBN6698_n_13796), .o(FE_OCP_RBN6700_n_13796) );
in01s02 FE_OCP_RBC6701_n_14444 ( .a(FE_OCP_RBN5760_n_14444), .o(FE_OCP_RBN6701_n_14444) );
in01s01 FE_OCP_RBC6702_n_14444 ( .a(FE_OCP_RBN5760_n_14444), .o(FE_OCP_RBN6702_n_14444) );
in01s02 FE_OCP_RBC6703_n_14444 ( .a(FE_OCP_RBN6701_n_14444), .o(FE_OCP_RBN6703_n_14444) );
in01m02 FE_OCP_RBC6704_n_8762 ( .a(n_8762), .o(FE_OCP_RBN6704_n_8762) );
in01s01 FE_OCP_RBC6705_n_8762 ( .a(n_8762), .o(FE_OCP_RBN6705_n_8762) );
in01f04 FE_OCP_RBC6706_n_29787 ( .a(n_29787), .o(FE_OCP_RBN6706_n_29787) );
in01s01 FE_OCP_RBC6707_n_8719 ( .a(n_8719), .o(FE_OCP_RBN6707_n_8719) );
in01s01 FE_OCP_RBC6708_n_44570 ( .a(FE_OCP_RBN5781_n_44570), .o(FE_OCP_RBN6708_n_44570) );
in01s10 FE_OCP_RBC6709_n_44570 ( .a(FE_OCP_RBN5781_n_44570), .o(FE_OCP_RBN6709_n_44570) );
in01s10 FE_OCP_RBC6710_n_44570 ( .a(FE_OCP_RBN6709_n_44570), .o(FE_OCP_RBN6710_n_44570) );
in01s02 FE_OCP_RBC6711_n_44570 ( .a(FE_OCP_RBN6709_n_44570), .o(FE_OCP_RBN6711_n_44570) );
in01s01 FE_OCP_RBC6712_n_44570 ( .a(FE_OCP_RBN6709_n_44570), .o(FE_OCP_RBN6712_n_44570) );
in01f02 FE_OCP_RBC6713_n_8800 ( .a(n_8800), .o(FE_OCP_RBN6713_n_8800) );
in01s01 FE_OCP_RBC6714_n_3604 ( .a(n_3604), .o(FE_OCP_RBN6714_n_3604) );
in01s02 FE_OCP_RBC6715_n_3604 ( .a(n_3604), .o(FE_OCP_RBN6715_n_3604) );
in01s06 FE_OCP_RBC6716_n_3604 ( .a(n_3604), .o(FE_OCP_RBN6716_n_3604) );
in01s04 FE_OCP_RBC6717_n_3604 ( .a(FE_OCP_RBN6716_n_3604), .o(FE_OCP_RBN6717_n_3604) );
in01s01 FE_OCP_RBC6718_n_3604 ( .a(FE_OCP_RBN6716_n_3604), .o(FE_OCP_RBN6718_n_3604) );
in01s01 FE_OCP_RBC6719_n_3604 ( .a(FE_OCP_RBN6716_n_3604), .o(FE_OCP_RBN6719_n_3604) );
in01s01 FE_OCP_RBC6720_FE_OCP_DRV_N6264_n_9014 ( .a(FE_OCP_DRV_N6264_n_9014), .o(FE_OCP_RBN6720_FE_OCP_DRV_N6264_n_9014) );
in01s01 FE_OCP_RBC6721_FE_OCP_DRV_N6264_n_9014 ( .a(FE_OCP_DRV_N6264_n_9014), .o(FE_OCP_RBN6721_FE_OCP_DRV_N6264_n_9014) );
in01s02 FE_OCP_RBC6722_n_9034 ( .a(n_9034), .o(FE_OCP_RBN6722_n_9034) );
in01m02 FE_OCP_RBC6723_n_44055 ( .a(n_44055), .o(FE_OCP_RBN6723_n_44055) );
in01s01 FE_OCP_RBC6724_n_44055 ( .a(n_44055), .o(FE_OCP_RBN6724_n_44055) );
in01s01 FE_OCP_RBC6725_n_34388 ( .a(n_34388), .o(FE_OCP_RBN6725_n_34388) );
in01s04 FE_OCP_RBC6726_n_34388 ( .a(n_34388), .o(FE_OCP_RBN6726_n_34388) );
in01s01 FE_OCP_RBC6727_n_34388 ( .a(FE_OCP_RBN6726_n_34388), .o(FE_OCP_RBN6727_n_34388) );
in01s01 FE_OCP_RBC6728_n_34388 ( .a(FE_OCP_RBN6727_n_34388), .o(FE_OCP_RBN6728_n_34388) );
in01s01 FE_OCP_RBC6729_n_44579 ( .a(FE_OCP_RBN5829_n_44579), .o(FE_OCP_RBN6729_n_44579) );
in01s01 FE_OCP_RBC6730_n_44579 ( .a(FE_OCP_RBN6729_n_44579), .o(FE_OCP_RBN6730_n_44579) );
in01s02 FE_OCP_RBC6731_n_44579 ( .a(FE_OCP_RBN6729_n_44579), .o(FE_OCP_RBN6731_n_44579) );
in01s01 FE_OCP_RBC6732_n_44579 ( .a(FE_OCP_RBN6729_n_44579), .o(FE_OCP_RBN6732_n_44579) );
in01s01 FE_OCP_RBC6733_n_44579 ( .a(FE_OCP_RBN5830_n_44579), .o(FE_OCP_RBN6733_n_44579) );
in01s01 FE_OCP_RBC6734_n_44579 ( .a(FE_OCP_RBN5830_n_44579), .o(FE_OCP_RBN6734_n_44579) );
in01s01 FE_OCP_RBC6735_n_44579 ( .a(FE_OCP_RBN5830_n_44579), .o(FE_OCP_RBN6735_n_44579) );
in01s01 FE_OCP_RBC6736_n_44579 ( .a(FE_OCP_RBN6735_n_44579), .o(FE_OCP_RBN6736_n_44579) );
in01s02 FE_OCP_RBC6737_n_44563 ( .a(FE_OCP_RBN5836_n_44563), .o(FE_OCP_RBN6737_n_44563) );
in01s02 FE_OCP_RBC6738_n_44563 ( .a(FE_OCP_RBN5836_n_44563), .o(FE_OCP_RBN6738_n_44563) );
in01m10 FE_OCP_RBC6739_n_44563 ( .a(FE_OCP_RBN5836_n_44563), .o(FE_OCP_RBN6739_n_44563) );
in01s10 FE_OCP_RBC6740_n_44563 ( .a(FE_OCP_RBN6739_n_44563), .o(FE_OCP_RBN6740_n_44563) );
in01s02 FE_OCP_RBC6741_n_44563 ( .a(FE_OCP_RBN6739_n_44563), .o(FE_OCP_RBN6741_n_44563) );
in01s02 FE_OCP_RBC6742_n_3746 ( .a(n_3746), .o(FE_OCP_RBN6742_n_3746) );
in01s01 FE_OCP_RBC6743_n_3746 ( .a(n_3746), .o(FE_OCP_RBN6743_n_3746) );
in01s01 FE_OCP_RBC6744_n_3746 ( .a(FE_OCP_RBN6743_n_3746), .o(FE_OCP_RBN6744_n_3746) );
in01s01 FE_OCP_RBC6745_n_3746 ( .a(FE_OCP_RBN6744_n_3746), .o(FE_OCP_RBN6745_n_3746) );
in01s01 FE_OCP_RBC6746_n_30170 ( .a(n_30170), .o(FE_OCP_RBN6746_n_30170) );
in01s01 FE_OCP_RBC6747_n_30170 ( .a(FE_OCP_RBN6746_n_30170), .o(FE_OCP_RBN6747_n_30170) );
in01s01 FE_OCP_RBC6748_n_30170 ( .a(FE_OCP_RBN6747_n_30170), .o(FE_OCP_RBN6748_n_30170) );
in01m02 FE_OCP_RBC6749_n_9198 ( .a(n_9198), .o(FE_OCP_RBN6749_n_9198) );
in01s01 FE_OCP_RBC6750_n_9198 ( .a(FE_OCP_RBN6749_n_9198), .o(FE_OCP_RBN6750_n_9198) );
in01s02 FE_OCP_RBC6751_n_9185 ( .a(n_9185), .o(FE_OCP_RBN6751_n_9185) );
in01s01 FE_OCP_RBC6752_n_30273 ( .a(n_30273), .o(FE_OCP_RBN6752_n_30273) );
in01m02 FE_OCP_RBC6753_n_35049 ( .a(n_35049), .o(FE_OCP_RBN6753_n_35049) );
in01m04 FE_OCP_RBC6754_n_38806 ( .a(n_38806), .o(FE_OCP_RBN6754_n_38806) );
in01m06 FE_OCP_RBC6755_n_38806 ( .a(n_38806), .o(FE_OCP_RBN6755_n_38806) );
in01s02 FE_OCP_RBC6756_n_38806 ( .a(FE_OCP_RBN6755_n_38806), .o(FE_OCP_RBN6756_n_38806) );
in01m04 FE_OCP_RBC6757_n_38806 ( .a(FE_OCP_RBN6755_n_38806), .o(FE_OCP_RBN6757_n_38806) );
in01f08 FE_OCP_RBC6758_n_38806 ( .a(FE_OCP_RBN6755_n_38806), .o(FE_OCP_RBN6758_n_38806) );
in01s01 FE_OCP_RBC6759_n_9075 ( .a(n_9075), .o(FE_OCP_RBN6759_n_9075) );
in01m02 FE_OCP_RBC6760_n_9075 ( .a(n_9075), .o(FE_OCP_RBN6760_n_9075) );
in01s02 FE_OCP_RBC6761_n_3705 ( .a(FE_OCP_RBN5864_n_3705), .o(FE_OCP_RBN6761_n_3705) );
in01s01 FE_OCP_RBC6762_n_3790 ( .a(n_3790), .o(FE_OCP_RBN6762_n_3790) );
in01m06 FE_OCP_RBC6763_FE_RN_2259_0 ( .a(FE_RN_2259_0), .o(FE_OCP_RBN6763_FE_RN_2259_0) );
in01m01 FE_OCP_RBC6764_FE_RN_2259_0 ( .a(FE_RN_2259_0), .o(FE_OCP_RBN6764_FE_RN_2259_0) );
in01s02 FE_OCP_RBC6765_n_3704 ( .a(FE_OCP_RBN5870_n_3704), .o(FE_OCP_RBN6765_n_3704) );
in01s01 FE_OCP_RBC6766_n_3704 ( .a(FE_OCP_RBN6765_n_3704), .o(FE_OCP_RBN6766_n_3704) );
in01s01 FE_OCP_RBC6767_n_3704 ( .a(FE_OCP_RBN6765_n_3704), .o(FE_OCP_RBN6767_n_3704) );
in01s04 FE_OCP_RBC6768_n_3700 ( .a(FE_OCP_RBN5873_n_3700), .o(FE_OCP_RBN6768_n_3700) );
in01s01 FE_OCP_RBC6769_n_3700 ( .a(FE_OCP_RBN6768_n_3700), .o(FE_OCP_RBN6769_n_3700) );
in01s01 FE_OCP_RBC6770_n_3700 ( .a(FE_OCP_RBN6769_n_3700), .o(FE_OCP_RBN6770_n_3700) );
in01s01 FE_OCP_RBC6771_n_3700 ( .a(FE_OCP_RBN6769_n_3700), .o(FE_OCP_RBN6771_n_3700) );
in01s01 FE_OCP_RBC6772_n_3700 ( .a(FE_OCP_RBN6769_n_3700), .o(FE_OCP_RBN6772_n_3700) );
in01s01 FE_OCP_RBC6773_n_4046 ( .a(n_4046), .o(FE_OCP_RBN6773_n_4046) );
in01s10 FE_OCP_RBC6774_n_4046 ( .a(n_4046), .o(FE_OCP_RBN6774_n_4046) );
in01s01 FE_OCP_RBC6775_n_4046 ( .a(FE_OCP_RBN6773_n_4046), .o(FE_OCP_RBN6775_n_4046) );
in01s01 FE_OCP_RBC6776_n_4046 ( .a(FE_OCP_RBN6773_n_4046), .o(FE_OCP_RBN6776_n_4046) );
in01s10 FE_OCP_RBC6777_n_4046 ( .a(FE_OCP_RBN6774_n_4046), .o(FE_OCP_RBN6777_n_4046) );
in01s01 FE_OCP_RBC6778_n_4046 ( .a(FE_OCP_RBN6774_n_4046), .o(FE_OCP_RBN6778_n_4046) );
in01s01 FE_OCP_RBC6779_n_4046 ( .a(FE_OCP_RBN6775_n_4046), .o(FE_OCP_RBN6779_n_4046) );
in01s06 FE_OCP_RBC6780_n_4046 ( .a(FE_OCP_RBN6777_n_4046), .o(FE_OCP_RBN6780_n_4046) );
in01s01 FE_OCP_RBC6781_n_4046 ( .a(FE_OCP_RBN6777_n_4046), .o(FE_OCP_RBN6781_n_4046) );
in01s01 FE_OCP_RBC6782_n_4046 ( .a(FE_OCP_RBN6778_n_4046), .o(FE_OCP_RBN6782_n_4046) );
in01s01 FE_OCP_RBC6783_n_4046 ( .a(FE_OCP_RBN6779_n_4046), .o(FE_OCP_RBN6783_n_4046) );
in01s06 FE_OCP_RBC6784_n_4046 ( .a(FE_OCP_RBN6780_n_4046), .o(FE_OCP_RBN6784_n_4046) );
in01f02 FE_OCP_RBC6785_n_14704 ( .a(n_14704), .o(FE_OCP_RBN6785_n_14704) );
in01m02 FE_OCP_RBC6786_n_9410 ( .a(n_9410), .o(FE_OCP_RBN6786_n_9410) );
in01s01 FE_OCP_RBC6787_n_35130 ( .a(n_35130), .o(FE_OCP_RBN6787_n_35130) );
in01m02 FE_OCP_RBC6788_n_35130 ( .a(n_35130), .o(FE_OCP_RBN6788_n_35130) );
in01m04 FE_OCP_RBC6789_n_20242 ( .a(FE_OCP_RBN2943_n_20242), .o(FE_OCP_RBN6789_n_20242) );
in01s04 FE_OCP_RBC6790_n_20242 ( .a(FE_OCP_RBN6789_n_20242), .o(FE_OCP_RBN6790_n_20242) );
in01s06 FE_OCP_RBC6791_n_20242 ( .a(FE_OCP_RBN6789_n_20242), .o(FE_OCP_RBN6791_n_20242) );
in01s01 FE_OCP_RBC6792_n_9510 ( .a(n_9510), .o(FE_OCP_RBN6792_n_9510) );
in01s01 FE_OCP_RBC6793_n_25211 ( .a(FE_OCP_RBN5927_n_25211), .o(FE_OCP_RBN6793_n_25211) );
in01s01 FE_OCP_RBC6794_n_25211 ( .a(FE_OCP_RBN5927_n_25211), .o(FE_OCP_RBN6794_n_25211) );
in01m03 FE_OCP_RBC6795_n_25211 ( .a(FE_OCP_RBN5927_n_25211), .o(FE_OCP_RBN6795_n_25211) );
in01m03 FE_OCP_RBC6796_n_25211 ( .a(FE_OCP_RBN6795_n_25211), .o(FE_OCP_RBN6796_n_25211) );
in01s01 FE_OCP_RBC6797_n_25211 ( .a(FE_OCP_RBN6795_n_25211), .o(FE_OCP_RBN6797_n_25211) );
in01s02 FE_OCP_RBC6798_n_15156 ( .a(FE_OCP_RBN4323_n_15156), .o(FE_OCP_RBN6798_n_15156) );
in01s01 FE_OCP_RBC6799_n_15156 ( .a(FE_OCP_RBN4323_n_15156), .o(FE_OCP_RBN6799_n_15156) );
in01s03 FE_OCP_RBC6800_n_15156 ( .a(FE_OCP_RBN4323_n_15156), .o(FE_OCP_RBN6800_n_15156) );
in01s06 FE_OCP_RBC6801_n_15156 ( .a(FE_OCP_RBN4323_n_15156), .o(FE_OCP_RBN6801_n_15156) );
in01s06 FE_OCP_RBC6802_n_15156 ( .a(FE_OCP_RBN6800_n_15156), .o(FE_OCP_RBN6802_n_15156) );
in01s01 FE_OCP_RBC6803_n_20565 ( .a(n_20565), .o(FE_OCP_RBN6803_n_20565) );
in01s02 FE_OCP_RBC6804_n_9742 ( .a(n_9742), .o(FE_OCP_RBN6804_n_9742) );
in01s01 FE_OCP_RBC6805_n_9742 ( .a(n_9742), .o(FE_OCP_RBN6805_n_9742) );
in01s01 FE_OCP_RBC6806_n_4411 ( .a(n_4411), .o(FE_OCP_RBN6806_n_4411) );
in01f02 FE_OCP_RBC6807_n_15110 ( .a(n_15110), .o(FE_OCP_RBN6807_n_15110) );
in01s02 FE_OCP_RBC6808_n_20667 ( .a(n_20667), .o(FE_OCP_RBN6808_n_20667) );
in01s02 FE_OCP_RBC6809_n_4563 ( .a(n_4563), .o(FE_OCP_RBN6809_n_4563) );
in01m04 FE_OCP_RBC6810_n_39551 ( .a(n_39551), .o(FE_OCP_RBN6810_n_39551) );
in01s01 FE_OCP_RBC6811_n_39551 ( .a(n_39551), .o(FE_OCP_RBN6811_n_39551) );
in01s01 FE_OCP_RBC6812_n_30608 ( .a(n_30608), .o(FE_OCP_RBN6812_n_30608) );
in01s02 FE_OCP_RBC6813_n_30608 ( .a(n_30608), .o(FE_OCP_RBN6813_n_30608) );
in01s02 FE_OCP_RBC6814_n_9893 ( .a(n_9893), .o(FE_OCP_RBN6814_n_9893) );
in01s02 FE_OCP_RBC6815_n_25753 ( .a(n_25753), .o(FE_OCP_RBN6815_n_25753) );
in01s02 FE_OCP_RBC6816_n_4654 ( .a(n_4654), .o(FE_OCP_RBN6816_n_4654) );
in01m02 FE_OCP_RBC6817_n_20889 ( .a(n_20889), .o(FE_OCP_RBN6817_n_20889) );
in01m02 FE_OCP_RBC6818_n_25997 ( .a(n_25997), .o(FE_OCP_RBN6818_n_25997) );
in01s01 FE_OCP_RBC6819_n_25997 ( .a(FE_OCP_RBN6818_n_25997), .o(FE_OCP_RBN6819_n_25997) );
in01s01 FE_OCP_RBC6820_n_5152 ( .a(n_5152), .o(FE_OCP_RBN6820_n_5152) );
in01m02 FE_OCP_RBC6821_n_45319 ( .a(n_45319), .o(FE_OCP_RBN6821_n_45319) );
in01m02 FE_OCP_RBC6822_FE_RN_592_0 ( .a(FE_RN_592_0), .o(FE_OCP_RBN6822_FE_RN_592_0) );
in01m01 FE_OCP_RBC6823_FE_RN_592_0 ( .a(FE_RN_592_0), .o(FE_OCP_RBN6823_FE_RN_592_0) );
in01s01 FE_OCP_RBC6824_n_39542 ( .a(n_39542), .o(FE_OCP_RBN6824_n_39542) );
in01f02 FE_OCP_RBC6825_n_39542 ( .a(n_39542), .o(FE_OCP_RBN6825_n_39542) );
in01s01 FE_OCP_RBC6826_n_15514 ( .a(FE_OCP_RBN4375_n_15514), .o(FE_OCP_RBN6826_n_15514) );
in01s02 FE_OCP_RBC6827_n_15514 ( .a(FE_OCP_RBN4375_n_15514), .o(FE_OCP_RBN6827_n_15514) );
in01s02 FE_OCP_RBC6828_n_15514 ( .a(FE_OCP_RBN6827_n_15514), .o(FE_OCP_RBN6828_n_15514) );
in01s01 FE_OCP_RBC6829_n_15514 ( .a(FE_OCP_RBN6827_n_15514), .o(FE_OCP_RBN6829_n_15514) );
in01m02 FE_OCP_RBC6830_n_45484 ( .a(n_45484), .o(FE_OCP_RBN6830_n_45484) );
in01f02 FE_OCP_RBC6831_n_15676 ( .a(n_15676), .o(FE_OCP_RBN6831_n_15676) );
in01s01 FE_OCP_RBC6832_n_31073 ( .a(n_31073), .o(FE_OCP_RBN6832_n_31073) );
in01s02 FE_OCP_RBC6833_n_31073 ( .a(n_31073), .o(FE_OCP_RBN6833_n_31073) );
in01s01 FE_OCP_RBC6834_n_31073 ( .a(n_31073), .o(FE_OCP_RBN6834_n_31073) );
in01s01 FE_OCP_RBC6835_n_39577 ( .a(n_39577), .o(FE_OCP_RBN6835_n_39577) );
in01m04 FE_OCP_RBC6836_n_39577 ( .a(n_39577), .o(FE_OCP_RBN6836_n_39577) );
in01f02 FE_OCP_RBC6837_FE_RN_586_0 ( .a(FE_RN_586_0), .o(FE_OCP_RBN6837_FE_RN_586_0) );
in01s04 FE_OCP_RBC6838_FE_RN_586_0 ( .a(FE_RN_586_0), .o(FE_OCP_RBN6838_FE_RN_586_0) );
in01m02 FE_OCP_RBC6839_FE_RN_2660_0 ( .a(FE_RN_2660_0), .o(FE_OCP_RBN6839_FE_RN_2660_0) );
in01s02 FE_OCP_RBC6840_FE_RN_2660_0 ( .a(FE_RN_2660_0), .o(FE_OCP_RBN6840_FE_RN_2660_0) );
in01s02 FE_OCP_RBC6841_n_31023 ( .a(n_31023), .o(FE_OCP_RBN6841_n_31023) );
in01s02 FE_OCP_RBC6842_n_5397 ( .a(n_5397), .o(FE_OCP_RBN6842_n_5397) );
in01s02 FE_OCP_RBC6843_n_31194 ( .a(n_31194), .o(FE_OCP_RBN6843_n_31194) );
in01s01 FE_OCP_RBC6844_n_15599 ( .a(FE_OCP_RBN3186_n_15599), .o(FE_OCP_RBN6844_n_15599) );
in01s02 FE_OCP_RBC6845_n_15599 ( .a(FE_OCP_RBN3186_n_15599), .o(FE_OCP_RBN6845_n_15599) );
in01s01 FE_OCP_RBC6846_n_15599 ( .a(FE_OCP_RBN3186_n_15599), .o(FE_OCP_RBN6846_n_15599) );
in01s01 FE_OCP_RBC6847_n_15599 ( .a(FE_OCP_RBN6845_n_15599), .o(FE_OCP_RBN6847_n_15599) );
in01s01 FE_OCP_RBC6848_n_15599 ( .a(FE_OCP_RBN6846_n_15599), .o(FE_OCP_RBN6848_n_15599) );
in01s04 FE_OCP_RBC6849_n_26358 ( .a(n_26358), .o(FE_OCP_RBN6849_n_26358) );
in01m01 FE_OCP_RBC6850_n_26504 ( .a(n_26504), .o(FE_OCP_RBN6850_n_26504) );
in01m10 FE_OCP_RBC6851_n_39793 ( .a(FE_OCP_RBN6105_n_39793), .o(FE_OCP_RBN6851_n_39793) );
in01m10 FE_OCP_RBC6852_n_39793 ( .a(FE_OCP_RBN6851_n_39793), .o(FE_OCP_RBN6852_n_39793) );
in01s08 FE_OCP_RBC6853_n_39793 ( .a(FE_OCP_RBN6851_n_39793), .o(FE_OCP_RBN6853_n_39793) );
in01s01 FE_OCP_RBC6854_n_5735 ( .a(n_5735), .o(FE_OCP_RBN6854_n_5735) );
in01s01 FE_OCP_RBC6855_n_5735 ( .a(n_5735), .o(FE_OCP_RBN6855_n_5735) );
in01s06 FE_OCP_RBC6856_n_26160 ( .a(FE_OCP_RBN4405_n_26160), .o(FE_OCP_RBN6856_n_26160) );
in01s06 FE_OCP_RBC6857_n_26160 ( .a(FE_OCP_RBN6856_n_26160), .o(FE_OCP_RBN6857_n_26160) );
in01s06 FE_OCP_RBC6858_n_26160 ( .a(FE_OCP_RBN6856_n_26160), .o(FE_OCP_RBN6858_n_26160) );
in01s01 FE_OCP_RBC6859_n_26160 ( .a(FE_OCP_RBN6857_n_26160), .o(FE_OCP_RBN6859_n_26160) );
in01s01 FE_OCP_RBC6860_n_26160 ( .a(FE_OCP_RBN6859_n_26160), .o(FE_OCP_RBN6860_n_26160) );
in01s06 FE_OCP_RBC6861_n_46285 ( .a(n_46285), .o(FE_OCP_RBN6861_n_46285) );
in01s04 FE_OCP_RBC6862_n_46285 ( .a(FE_OCP_RBN6861_n_46285), .o(FE_OCP_RBN6862_n_46285) );
in01s06 FE_OCP_RBC6863_n_46285 ( .a(FE_OCP_RBN6861_n_46285), .o(FE_OCP_RBN6863_n_46285) );
in01s06 FE_OCP_RBC6864_n_46285 ( .a(FE_OCP_RBN6861_n_46285), .o(FE_OCP_RBN6864_n_46285) );
in01s02 FE_OCP_RBC6865_n_46285 ( .a(FE_OCP_RBN6861_n_46285), .o(FE_OCP_RBN6865_n_46285) );
in01m02 FE_OCP_RBC6866_n_5743 ( .a(n_5743), .o(FE_OCP_RBN6866_n_5743) );
in01s01 FE_OCP_RBC6867_n_16392 ( .a(n_16392), .o(FE_OCP_RBN6867_n_16392) );
in01f04 FE_OCP_RBC6868_n_16392 ( .a(n_16392), .o(FE_OCP_RBN6868_n_16392) );
in01m02 FE_OCP_RBC6869_n_5751 ( .a(n_5751), .o(FE_OCP_RBN6869_n_5751) );
in01m02 FE_OCP_RBC6870_FE_RN_2289_0 ( .a(FE_RN_2289_0), .o(FE_OCP_RBN6870_FE_RN_2289_0) );
in01s04 FE_OCP_RBC6871_FE_RN_2289_0 ( .a(FE_RN_2289_0), .o(FE_OCP_RBN6871_FE_RN_2289_0) );
in01s01 FE_OCP_RBC6872_n_31520 ( .a(FE_OCP_RBN6138_n_31520), .o(FE_OCP_RBN6872_n_31520) );
in01s01 FE_OCP_RBC6873_n_31520 ( .a(FE_OCP_RBN6138_n_31520), .o(FE_OCP_RBN6873_n_31520) );
in01s01 FE_OCP_RBC6874_n_31520 ( .a(FE_OCP_RBN6873_n_31520), .o(FE_OCP_RBN6874_n_31520) );
in01s02 FE_OCP_RBC6875_n_31520 ( .a(FE_OCP_RBN6873_n_31520), .o(FE_OCP_RBN6875_n_31520) );
in01s01 FE_OCP_RBC6876_n_16920 ( .a(n_16920), .o(FE_OCP_RBN6876_n_16920) );
in01s02 FE_OCP_RBC6877_n_16920 ( .a(n_16920), .o(FE_OCP_RBN6877_n_16920) );
in01f08 FE_OCP_RBC6878_n_44267 ( .a(FE_OCP_RBN6184_n_44267), .o(FE_OCP_RBN6878_n_44267) );
in01s06 FE_OCP_RBC6879_n_31819 ( .a(FE_OCP_RBN6202_n_31819), .o(FE_OCP_RBN6879_n_31819) );
in01s02 FE_OCP_RBC6880_n_31819 ( .a(FE_OCP_RBN6202_n_31819), .o(FE_OCP_RBN6880_n_31819) );
in01s01 FE_OCP_RBC6881_n_31819 ( .a(FE_OCP_RBN6879_n_31819), .o(FE_OCP_RBN6881_n_31819) );
in01s02 FE_OCP_RBC6882_n_11486 ( .a(FE_OCP_RBN6209_n_11486), .o(FE_OCP_RBN6882_n_11486) );
in01s04 FE_OCP_RBC6883_n_11486 ( .a(FE_OCP_RBN6209_n_11486), .o(FE_OCP_RBN6883_n_11486) );
in01s40 FE_OCP_RBC7005_n_44962 ( .a(n_44962), .o(FE_OCP_RBN7005_n_44962) );
in01s06 FE_OCP_RBC7006_n_44962 ( .a(FE_OCP_RBN7007_n_44962), .o(FE_OCP_RBN7006_n_44962) );
in01s01 FE_OCP_RBC7007_n_44962 ( .a(n_44962), .o(FE_OCP_RBN7007_n_44962) );
in01s40 FE_OCP_RBC7008_n_44962 ( .a(n_44962), .o(FE_OCP_RBN7008_n_44962) );
in01m03 FE_OCP_RBC7009_n_44962 ( .a(FE_OCP_RBN7011_n_44962), .o(FE_OCP_RBN7009_n_44962) );
in01s02 FE_OCP_RBC7010_n_44962 ( .a(FE_OCP_RBN7011_n_44962), .o(FE_OCP_RBN7010_n_44962) );
in01m01 FE_OCP_RBC7011_n_44962 ( .a(n_44962), .o(FE_OCP_RBN7011_n_44962) );
in01s40 FE_OCP_RBC7012_n_44962 ( .a(FE_OCP_RBN7014_n_44962), .o(FE_OCP_RBN7012_n_44962) );
in01s06 FE_OCP_RBC7013_n_44962 ( .a(FE_OCP_RBN7014_n_44962), .o(FE_OCP_RBN7013_n_44962) );
in01s06 FE_OCP_RBC7014_n_44962 ( .a(n_44962), .o(FE_OCP_RBN7014_n_44962) );
in01s40 FE_OCP_RBC7015_n_44962 ( .a(n_44962), .o(FE_OCP_RBN7015_n_44962) );
in01m10 FE_OCP_RBC7016_n_32687 ( .a(n_32687), .o(FE_OCP_RBN7016_n_32687) );
in01m08 FE_OCP_RBC7017_n_32687 ( .a(FE_OCP_RBN7016_n_32687), .o(FE_OCP_RBN7017_n_32687) );
in01s10 FE_OCP_RBC7018_n_32649 ( .a(n_32649), .o(FE_OCP_RBN7018_n_32649) );
in01s01 FE_OCP_RBC7019_n_28166 ( .a(n_28166), .o(FE_OCP_RBN7019_n_28166) );
in01s01 FE_OCP_RBC7020_n_17717 ( .a(n_17717), .o(FE_OCP_RBN7020_n_17717) );
in01s01 FE_OCP_RBC7021_n_33330 ( .a(n_33330), .o(FE_OCP_RBN7021_n_33330) );
in01s01 FE_OCP_RBC7022_n_18248 ( .a(n_18248), .o(FE_OCP_RBN7022_n_18248) );
in01s06 FE_OCP_RBC7023_n_18650 ( .a(n_18650), .o(FE_OCP_RBN7023_n_18650) );
in01f03 FE_OCP_RBC7024_FE_RN_1738_0 ( .a(FE_RN_1738_0), .o(FE_OCP_RBN7024_FE_RN_1738_0) );
in01s02 FE_OCP_RBC7025_n_18873 ( .a(n_18873), .o(FE_OCP_RBN7025_n_18873) );
in01s01 FE_OCP_RBC7026_n_18866 ( .a(n_18866), .o(FE_OCP_RBN7026_n_18866) );
in01s01 FE_OCP_RBC7027_n_18866 ( .a(FE_OCP_RBN7026_n_18866), .o(FE_OCP_RBN7027_n_18866) );
in01s01 FE_OCP_RBC7028_n_18866 ( .a(FE_OCP_RBN7027_n_18866), .o(FE_OCP_RBN7028_n_18866) );
in01f03 FE_OCP_RBC7029_n_44259 ( .a(n_44259), .o(FE_OCP_RBN7029_n_44259) );
in01s06 FE_OCP_RBC7030_n_44259 ( .a(n_44259), .o(FE_OCP_RBN7030_n_44259) );
in01f02 FE_OCP_RBC7031_n_18981 ( .a(n_18981), .o(FE_OCP_RBN7031_n_18981) );
in01s01 FE_OCP_RBC7032_n_18981 ( .a(n_18981), .o(FE_OCP_RBN7032_n_18981) );
in01s02 FE_OCP_RBC7033_n_18981 ( .a(FE_OCP_RBN7032_n_18981), .o(FE_OCP_RBN7033_n_18981) );
in01s01 FE_OCP_RBC7034_n_18981 ( .a(FE_OCP_RBN7033_n_18981), .o(FE_OCP_RBN7034_n_18981) );
in01s01 FE_OCP_RBC7035_n_18981 ( .a(FE_OCP_RBN7033_n_18981), .o(FE_OCP_RBN7035_n_18981) );
in01s04 FE_OCP_RBC7036_n_18982 ( .a(n_18982), .o(FE_OCP_RBN7036_n_18982) );
in01m08 FE_OCP_RBC7037_n_18982 ( .a(n_18982), .o(FE_OCP_RBN7037_n_18982) );
in01s01 FE_OCP_RBC7038_n_34903 ( .a(n_34903), .o(FE_OCP_RBN7038_n_34903) );
in01s04 FE_OCP_RBC7039_n_34903 ( .a(n_34903), .o(FE_OCP_RBN7039_n_34903) );
in01m02 FE_OCP_RBC7040_n_20167 ( .a(n_20167), .o(FE_OCP_RBN7040_n_20167) );
in01s01 FE_OCP_RBC7041_n_20336 ( .a(n_20336), .o(FE_OCP_RBN7041_n_20336) );
in01f02 FE_OCP_RBC7042_n_20336 ( .a(n_20336), .o(FE_OCP_RBN7042_n_20336) );
in01s01 FE_OCP_RBC7043_n_20336 ( .a(FE_OCP_RBN7041_n_20336), .o(FE_OCP_RBN7043_n_20336) );
in01f01 FE_OCP_RBC7044_FE_RN_1462_0 ( .a(FE_RN_1462_0), .o(FE_OCP_RBN7044_FE_RN_1462_0) );
in01s02 FE_OCP_RBC7045_FE_RN_1462_0 ( .a(FE_RN_1462_0), .o(FE_OCP_RBN7045_FE_RN_1462_0) );
in01s01 FE_OCP_RBC7046_n_20941 ( .a(n_20941), .o(FE_OCP_RBN7046_n_20941) );
in01m02 FE_OCP_RBC7047_n_20941 ( .a(n_20941), .o(FE_OCP_RBN7047_n_20941) );
in01s01 FE_OCP_RBC7048_n_20941 ( .a(n_20941), .o(FE_OCP_RBN7048_n_20941) );
in01s01 FE_OCP_RBC7049_n_20941 ( .a(FE_OCP_RBN7046_n_20941), .o(FE_OCP_RBN7049_n_20941) );
in01s01 FE_OCP_RBC7050_n_20941 ( .a(FE_OCP_RBN7048_n_20941), .o(FE_OCP_RBN7050_n_20941) );
in01s01 FE_OCP_RBC7051_n_20941 ( .a(FE_OCP_RBN7050_n_20941), .o(FE_OCP_RBN7051_n_20941) );
in01s01 FE_OCP_RBC7052_n_20941 ( .a(FE_OCP_RBN7050_n_20941), .o(FE_OCP_RBN7052_n_20941) );
in01m02 FE_OCP_RBC7053_n_30867 ( .a(n_30867), .o(FE_OCP_RBN7053_n_30867) );
in01s02 FE_OCP_RBC7055_FE_OCPN1068_n_21973 ( .a(FE_OCPN1068_n_21973), .o(FE_OCP_RBN7055_FE_OCPN1068_n_21973) );
in01s02 FE_OCP_RBC7056_FE_OCPN1068_n_21973 ( .a(FE_OCPN1068_n_21973), .o(FE_OCP_RBN7056_FE_OCPN1068_n_21973) );
in01m06 FE_OCP_RBC7057_n_36677 ( .a(n_36677), .o(FE_OCP_RBN7057_n_36677) );
in01s10 FE_OCP_RBC7101_n_44365 ( .a(n_44365), .o(FE_OCP_RBN7101_n_44365) );
in01s40 FE_OCP_RBC7102_n_44365 ( .a(FE_OCP_RBN7104_n_44365), .o(FE_OCP_RBN7102_n_44365) );
in01s06 FE_OCP_RBC7103_n_44365 ( .a(FE_OCP_RBN7104_n_44365), .o(FE_OCP_RBN7103_n_44365) );
in01m20 FE_OCP_RBC7104_n_44365 ( .a(n_44365), .o(FE_OCP_RBN7104_n_44365) );
in01s06 FE_OCP_RBC7105_n_44365 ( .a(n_44365), .o(FE_OCP_RBN7105_n_44365) );
in01s20 FE_OCP_RBC7106_n_44365 ( .a(FE_OCP_RBN7107_n_44365), .o(FE_OCP_RBN7106_n_44365) );
in01s20 FE_OCP_RBC7107_n_44365 ( .a(n_44365), .o(FE_OCP_RBN7107_n_44365) );
in01s10 FE_OCP_RBC7108_n_44365 ( .a(FE_OCP_RBN7110_n_44365), .o(FE_OCP_RBN7108_n_44365) );
in01s40 FE_OCP_RBC7109_n_44365 ( .a(FE_OCP_RBN7110_n_44365), .o(FE_OCP_RBN7109_n_44365) );
in01s40 FE_OCP_RBC7110_n_44365 ( .a(n_44365), .o(FE_OCP_RBN7110_n_44365) );
in01s08 FE_OCP_RBC7111_n_44365 ( .a(n_44365), .o(FE_OCP_RBN7111_n_44365) );
in01s20 FE_OCP_RBC7112_n_44365 ( .a(n_44365), .o(FE_OCP_RBN7112_n_44365) );
in01s10 FE_OCP_RBC7113_n_44365 ( .a(n_44365), .o(FE_OCP_RBN7113_n_44365) );
in01m10 FE_OCP_RBC7114_n_44365 ( .a(n_44365), .o(FE_OCP_RBN7114_n_44365) );
in01m01 FE_OCP_RBC7117_delay_xor_ln22_unr12_stage5_stallmux_q_0_ ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_0_), .o(FE_OCP_RBN7117_delay_xor_ln22_unr12_stage5_stallmux_q_0_) );
in01s06 FE_OCP_RBC7118_delay_xor_ln22_unr12_stage5_stallmux_q_0_ ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_0_), .o(FE_OCP_RBN7118_delay_xor_ln22_unr12_stage5_stallmux_q_0_) );
in01s80 FE_OCP_RBC7127_n_44722 ( .a(FE_OCP_RBN7129_n_44722), .o(FE_OCP_RBN7127_n_44722) );
in01s80 FE_OCP_RBC7128_n_44722 ( .a(FE_OCP_RBN7129_n_44722), .o(FE_OCP_RBN7128_n_44722) );
in01s80 FE_OCP_RBC7129_n_44722 ( .a(n_44722), .o(FE_OCP_RBN7129_n_44722) );
in01s02 FE_OCP_RBC7130_n_29262 ( .a(n_29262), .o(FE_OCP_RBN7130_n_29262) );
in01s02 FE_OCP_RBC7131_n_29262 ( .a(FE_OCP_RBN7130_n_29262), .o(FE_OCP_RBN7131_n_29262) );
in01f02 FE_OCP_RBC983_n_24262 ( .a(n_24262), .o(FE_OCP_RBN983_n_24262) );
in01s03 FE_OCP_RBC984_n_22822 ( .a(n_22822), .o(FE_OCP_RBN984_n_22822) );
in01s01 FE_OFC0_n_43918 ( .a(n_43918), .o(FE_OFN0_n_43918) );
in01s01 FE_OFC1178_n_916 ( .a(FE_OFN4810_n_916), .o(FE_OFN1178_n_916) );
in01s01 FE_OFC1180_n_13195 ( .a(FE_OFN4790_n_13195), .o(FE_OFN1180_n_13195) );
in01s01 FE_OFC1181_n_13195 ( .a(FE_OFN4790_n_13195), .o(FE_OFN1181_n_13195) );
in01s01 FE_OFC1182_n_24059 ( .a(n_24059), .o(FE_OFN1182_n_24059) );
in01s02 FE_OFC1183_n_24059 ( .a(FE_OFN1182_n_24059), .o(FE_OFN1183_n_24059) );
in01s01 FE_OFC1185_n_19801 ( .a(FE_OFN4805_n_19801), .o(FE_OFN1185_n_19801) );
in01s01 FE_OFC1194_n_27014 ( .a(n_27014), .o(FE_OFN1194_n_27014) );
in01s02 FE_OFC1196_n_27014 ( .a(FE_RN_1461_0), .o(FE_OFN1196_n_27014) );
in01s01 FE_OFC1198_n_27014 ( .a(FE_OFN1194_n_27014), .o(FE_OFN1198_n_27014) );
in01s01 FE_OFC1199_n_27014 ( .a(FE_OFN1194_n_27014), .o(FE_OFN1199_n_27014) );
in01s03 FE_OFC1_n_43918 ( .a(FE_OFN0_n_43918), .o(FE_OFN1_n_43918) );
in01s01 FE_OFC230_n_35655 ( .a(n_35655), .o(FE_OFN230_n_35655) );
in01s01 FE_OFC231_n_35655 ( .a(FE_OFN230_n_35655), .o(FE_OFN231_n_35655) );
in01s01 FE_OFC2_n_43918 ( .a(FE_OFN0_n_43918), .o(TIMEBOOST_net_2323) );
in01s01 FE_OFC321_n_2929 ( .a(FE_OFN794_n_2929), .o(FE_OFN321_n_2929) );
in01s01 FE_OFC380_n_9391 ( .a(n_9391), .o(FE_OFN380_n_9391) );
in01s01 FE_OFC381_n_9391 ( .a(FE_OFN380_n_9391), .o(FE_OFN381_n_9391) );
in01s01 FE_OFC3_n_43918 ( .a(FE_OFN4653_n_43918), .o(FE_OFN3_n_43918) );
in01s01 FE_OFC4650_n_43918 ( .a(FE_OFN5_n_43918), .o(FE_OFN4650_n_43918) );
in01s02 FE_OFC4651_n_43918 ( .a(FE_OFN4650_n_43918), .o(FE_OFN4651_n_43918) );
in01s01 FE_OFC4652_n_43918 ( .a(FE_OFN1_n_43918), .o(FE_OFN4652_n_43918) );
in01s02 FE_OFC4653_n_43918 ( .a(FE_OFN4652_n_43918), .o(FE_OFN4653_n_43918) );
in01f02 FE_OFC4669_n_16873 ( .a(FE_OFN4812_n_16873), .o(FE_OFN4669_n_16873) );
in01s01 FE_OFC4701_n_7702 ( .a(FE_OFN4806_n_7702), .o(FE_OFN4701_n_7702) );
in01s01 FE_OFC4714_n_18642 ( .a(n_18642), .o(FE_OFN4714_n_18642) );
in01s01 FE_OFC4715_n_18642 ( .a(FE_OFN4714_n_18642), .o(FE_OFN4715_n_18642) );
in01s01 FE_OFC4730_n_31403 ( .a(n_31403), .o(FE_OFN4730_n_31403) );
in01s01 FE_OFC4731_n_31403 ( .a(FE_OFN4730_n_31403), .o(FE_OFN4731_n_31403) );
in01s01 FE_OFC4732_n_29677 ( .a(n_29677), .o(FE_OFN4732_n_29677) );
in01s01 FE_OFC4733_n_29677 ( .a(FE_OFN4732_n_29677), .o(FE_OFN4733_n_29677) );
in01s01 FE_OFC4755_n_41563 ( .a(FE_OFN4809_n_41563), .o(FE_OFN4755_n_41563) );
in01s06 FE_OFC4762_n_3029 ( .a(n_3029), .o(FE_OFN4762_n_3029) );
in01s06 FE_OFC4763_n_3029 ( .a(FE_OFN4762_n_3029), .o(FE_OFN4763_n_3029) );
in01s03 FE_OFC4764_n_3029 ( .a(FE_OFN4762_n_3029), .o(FE_OFN4764_n_3029) );
in01s03 FE_OFC4765_n_3029 ( .a(FE_OFN4762_n_3029), .o(FE_OFN4765_n_3029) );
in01s01 FE_OFC4766_n_8309 ( .a(n_8309), .o(FE_OFN4766_n_8309) );
in01s01 FE_OFC4767_n_8309 ( .a(FE_OFN4766_n_8309), .o(FE_OFN4767_n_8309) );
in01s01 FE_OFC4768_n_8309 ( .a(FE_OFN4766_n_8309), .o(FE_OFN4768_n_8309) );
in01s01 FE_OFC4769_n_8309 ( .a(n_8309), .o(FE_OFN4769_n_8309) );
in01s01 FE_OFC4770_n_8309 ( .a(FE_OFN4769_n_8309), .o(FE_OFN4770_n_8309) );
in01s01 FE_OFC4771_n_8309 ( .a(FE_OFN4769_n_8309), .o(FE_OFN4771_n_8309) );
in01s10 FE_OFC4772_n_44463 ( .a(FE_OCP_RBN6740_n_44563), .o(FE_OFN4772_n_44463) );
in01s01 FE_OFC4774_n_44463 ( .a(FE_OCP_RBN6740_n_44563), .o(FE_OFN4774_n_44463) );
in01s02 FE_OFC4775_n_44463 ( .a(FE_OFN4774_n_44463), .o(FE_OFN4775_n_44463) );
in01s01 FE_OFC4776_n_44463 ( .a(FE_OFN4774_n_44463), .o(FE_OFN4776_n_44463) );
in01m20 FE_OFC4777_n_44490 ( .a(n_44490), .o(FE_OFN4777_n_44490) );
in01s02 FE_OFC4778_n_44490 ( .a(FE_OFN4777_n_44490), .o(FE_OFN4778_n_44490) );
in01m20 FE_OFC4779_n_44490 ( .a(FE_OFN4777_n_44490), .o(FE_OFN4779_n_44490) );
in01s01 FE_OFC4780_n_45813 ( .a(FE_OFN758_n_45813), .o(FE_OFN4780_n_45813) );
in01s01 FE_OFC4781_n_45813 ( .a(FE_OFN758_n_45813), .o(FE_OFN4781_n_45813) );
in01s02 FE_OFC4782_n_45813 ( .a(FE_OFN758_n_45813), .o(FE_OFN4782_n_45813) );
in01s01 FE_OFC4783_n_45813 ( .a(FE_OFN758_n_45813), .o(FE_OFN4783_n_45813) );
in01s01 FE_OFC4784_n_45813 ( .a(FE_OFN758_n_45813), .o(FE_OFN4784_n_45813) );
in01s01 FE_OFC4785_n_45813 ( .a(FE_OFN758_n_45813), .o(FE_OFN4785_n_45813) );
in01s01 FE_OFC4786_n_45813 ( .a(FE_OFN758_n_45813), .o(FE_OFN4786_n_45813) );
in01f02 FE_OFC4787_n_46137 ( .a(FE_OFN767_n_46137), .o(FE_OFN4787_n_46137) );
in01m08 FE_OFC4788_n_46137 ( .a(FE_OFN767_n_46137), .o(FE_OFN4788_n_46137) );
in01m10 FE_OFC4789_n_46137 ( .a(FE_OFN767_n_46137), .o(FE_OFN4789_n_46137) );
in01s01 FE_OFC4790_n_13195 ( .a(n_13195), .o(FE_OFN4790_n_13195) );
in01s01 FE_OFC4791_n_13195 ( .a(n_13195), .o(FE_OFN4791_n_13195) );
in01s01 FE_OFC4792_n_13195 ( .a(FE_OFN4791_n_13195), .o(FE_OFN4792_n_13195) );
in01s02 FE_OFC4793_n_13195 ( .a(FE_OFN4791_n_13195), .o(FE_OFN4793_n_13195) );
in01s03 FE_OFC4794_n_13195 ( .a(n_13195), .o(FE_OFN4794_n_13195) );
in01s06 FE_OFC4795_n_13195 ( .a(FE_OFN4794_n_13195), .o(FE_OFN4795_n_13195) );
in01s01 FE_OFC4796_n_13195 ( .a(FE_OFN4794_n_13195), .o(FE_OFN4796_n_13195) );
in01s01 FE_OFC4797_n_44498 ( .a(n_44498), .o(FE_OFN4797_n_44498) );
in01s02 FE_OFC4798_n_44498 ( .a(n_44498), .o(FE_OFN4798_n_44498) );
in01s06 FE_OFC4799_n_44498 ( .a(FE_OFN4797_n_44498), .o(FE_OFN4799_n_44498) );
in01m01 FE_OFC4800_n_44498 ( .a(FE_OFN4797_n_44498), .o(FE_OFN4800_n_44498) );
in01s01 FE_OFC4801_n_44498 ( .a(FE_OFN4798_n_44498), .o(FE_OFN4801_n_44498) );
in01s01 FE_OFC4802_n_44498 ( .a(FE_OFN4798_n_44498), .o(FE_OFN4802_n_44498) );
in01s01 FE_OFC4804_n_19384 ( .a(FE_OFN4813_n_19384), .o(FE_OFN4804_n_19384) );
in01s01 FE_OFC4805_n_19801 ( .a(n_19801), .o(FE_OFN4805_n_19801) );
in01s01 FE_OFC4806_n_7702 ( .a(n_7702), .o(FE_OFN4806_n_7702) );
in01s01 FE_OFC4807_n_2432 ( .a(FE_OFN4814_n_2432), .o(FE_OFN4807_n_2432) );
in01s01 FE_OFC4808_n_28820 ( .a(n_28820), .o(FE_OFN4808_n_28820) );
in01s01 FE_OFC4809_n_41563 ( .a(n_41563), .o(FE_OFN4809_n_41563) );
in01s01 FE_OFC4810_n_916 ( .a(n_916), .o(FE_OFN4810_n_916) );
in01s01 FE_OFC4811_n_902 ( .a(FE_OFN812_n_902), .o(FE_OFN4811_n_902) );
in01f02 FE_OFC4812_n_16873 ( .a(n_16873), .o(FE_OFN4812_n_16873) );
in01s01 FE_OFC4813_n_19384 ( .a(n_19384), .o(FE_OFN4813_n_19384) );
in01s01 FE_OFC4814_n_2432 ( .a(n_2432), .o(FE_OFN4814_n_2432) );
in01s01 FE_OFC4815_n_4018 ( .a(FE_OFN805_n_4018), .o(FE_OFN4815_n_4018) );
in01s01 FE_OFC4816_n_47017 ( .a(FE_OFN781_n_47017), .o(FE_OFN4816_n_47017) );
in01s01 FE_OFC4817_n_920 ( .a(n_920), .o(FE_OFN4817_n_920) );
in01s01 FE_OFC4818_n_920 ( .a(n_920), .o(FE_OFN4818_n_920) );
in01s03 FE_OFC4_n_43918 ( .a(FE_OFN3_n_43918), .o(FE_OFN4_n_43918) );
in01s01 FE_OFC5063_n_1545 ( .a(n_1545), .o(FE_OFN5063_n_1545) );
in01s01 FE_OFC5064_n_1545 ( .a(FE_OFN5063_n_1545), .o(FE_OFN5064_n_1545) );
in01f02 FE_OFC5065_n_8904 ( .a(n_8904), .o(FE_OFN5065_n_8904) );
in01f04 FE_OFC5066_n_8904 ( .a(FE_OFN5065_n_8904), .o(FE_OFN5066_n_8904) );
in01s01 FE_OFC5069_n_13646 ( .a(n_13646), .o(FE_OFN5069_n_13646) );
in01s01 FE_OFC5070_n_13646 ( .a(FE_OFN5069_n_13646), .o(FE_OFN5070_n_13646) );
in01s01 FE_OFC5071_n_18287 ( .a(n_18287), .o(FE_OFN5071_n_18287) );
in01s01 FE_OFC5072_n_18287 ( .a(FE_OFN5071_n_18287), .o(FE_OFN5072_n_18287) );
in01m01 FE_OFC5073_delay_sub_ln23_0_unr15_stage6_stallmux_q ( .a(FE_OFN742_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_OFN5073_delay_sub_ln23_0_unr15_stage6_stallmux_q) );
in01s01 FE_OFC5074_delay_sub_ln23_0_unr15_stage6_stallmux_q ( .a(FE_OFN5073_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_OFN5074_delay_sub_ln23_0_unr15_stage6_stallmux_q) );
in01s06 FE_OFC5075_delay_sub_ln23_0_unr15_stage6_stallmux_q ( .a(FE_OFN5073_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q) );
in01s01 FE_OFC5076_n_31435 ( .a(n_31435), .o(FE_OFN5076_n_31435) );
in01s01 FE_OFC5077_n_31435 ( .a(FE_OFN5076_n_31435), .o(FE_OFN5077_n_31435) );
in01s01 FE_OFC5078_n_29014 ( .a(n_29014), .o(FE_OFN5078_n_29014) );
in01s01 FE_OFC5079_n_29014 ( .a(FE_OFN5078_n_29014), .o(FE_OFN5079_n_29014) );
in01s01 FE_OFC5080_n_36439 ( .a(n_36439), .o(FE_OFN5080_n_36439) );
in01s01 FE_OFC5081_n_36439 ( .a(FE_OFN5080_n_36439), .o(FE_OFN5081_n_36439) );
in01s01 FE_OFC5082_n_36750 ( .a(n_36750), .o(FE_OFN5082_n_36750) );
in01s02 FE_OFC5083_n_36750 ( .a(FE_OFN5082_n_36750), .o(FE_OFN5083_n_36750) );
in01s02 FE_OFC5084_n_36750 ( .a(FE_OFN5082_n_36750), .o(FE_OFN5084_n_36750) );
in01s01 FE_OFC5085_delay_sub_ln23_0_unr22_stage8_stallmux_q ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(FE_OFN5085_delay_sub_ln23_0_unr22_stage8_stallmux_q) );
in01s04 FE_OFC5086_delay_sub_ln23_0_unr22_stage8_stallmux_q ( .a(FE_OFN5085_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q) );
in01s01 FE_OFC5087_delay_sub_ln23_0_unr22_stage8_stallmux_q ( .a(FE_OFN5085_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(FE_OFN5087_delay_sub_ln23_0_unr22_stage8_stallmux_q) );
in01s01 FE_OFC5088_delay_sub_ln23_0_unr25_stage9_stallmux_q ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(FE_OFN5088_delay_sub_ln23_0_unr25_stage9_stallmux_q) );
in01s01 FE_OFC5089_delay_sub_ln23_0_unr25_stage9_stallmux_q ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(FE_OFN5089_delay_sub_ln23_0_unr25_stage9_stallmux_q) );
in01s01 FE_OFC5090_delay_sub_ln23_0_unr25_stage9_stallmux_q ( .a(FE_OFN5088_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(FE_OFN5090_delay_sub_ln23_0_unr25_stage9_stallmux_q) );
in01s01 FE_OFC5091_delay_sub_ln23_0_unr25_stage9_stallmux_q ( .a(FE_OFN5088_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(FE_OFN5091_delay_sub_ln23_0_unr25_stage9_stallmux_q) );
in01s06 FE_OFC5092_delay_sub_ln23_0_unr25_stage9_stallmux_q ( .a(FE_OFN5089_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(FE_OFN5092_delay_sub_ln23_0_unr25_stage9_stallmux_q) );
in01s01 FE_OFC5093_delay_sub_ln23_0_unr25_stage9_stallmux_q ( .a(FE_OFN5089_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(FE_OFN5093_delay_sub_ln23_0_unr25_stage9_stallmux_q) );
in01s03 FE_OFC5_n_43918 ( .a(FE_OFN3_n_43918), .o(FE_OFN5_n_43918) );
in01s01 FE_OFC620_n_28336 ( .a(n_28336), .o(FE_OFN620_n_28336) );
in01s02 FE_OFC621_n_28336 ( .a(FE_OFN620_n_28336), .o(FE_OFN621_n_28336) );
in01s01 FE_OFC622_n_28336 ( .a(FE_OFN620_n_28336), .o(FE_OFN622_n_28336) );
in01s80 FE_OFC735_n_17093 ( .a(n_17093), .o(FE_OFN735_n_17093) );
in01s20 FE_OFC736_n_17093 ( .a(FE_OFN735_n_17093), .o(FE_OFN736_n_17093) );
in01s03 FE_OFC737_n_17093 ( .a(FE_OFN735_n_17093), .o(FE_OFN737_n_17093) );
in01f03 FE_OFC738_n_17093 ( .a(FE_OFN735_n_17093), .o(FE_OFN738_n_17093) );
in01s02 FE_OFC739_n_17093 ( .a(FE_OFN735_n_17093), .o(FE_OFN739_n_17093) );
in01s06 FE_OFC740_delay_sub_ln23_0_unr15_stage6_stallmux_q ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_OFN740_delay_sub_ln23_0_unr15_stage6_stallmux_q) );
in01s02 FE_OFC741_delay_sub_ln23_0_unr15_stage6_stallmux_q ( .a(FE_OFN740_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_OFN741_delay_sub_ln23_0_unr15_stage6_stallmux_q) );
in01s03 FE_OFC742_delay_sub_ln23_0_unr15_stage6_stallmux_q ( .a(FE_OFN740_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_OFN742_delay_sub_ln23_0_unr15_stage6_stallmux_q) );
in01s04 FE_OFC743_delay_sub_ln23_0_unr15_stage6_stallmux_q ( .a(FE_OFN740_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_OFN743_delay_sub_ln23_0_unr15_stage6_stallmux_q) );
in01s06 FE_OFC744_n_22641 ( .a(n_22641), .o(FE_OFN744_n_22641) );
in01s02 FE_OFC745_n_22641 ( .a(FE_OFN744_n_22641), .o(FE_OFN745_n_22641) );
in01s03 FE_OFC747_n_22641 ( .a(FE_OFN744_n_22641), .o(FE_OFN747_n_22641) );
in01s06 FE_OFC748_n_22641 ( .a(FE_OFN744_n_22641), .o(FE_OFN748_n_22641) );
in01m02 FE_OFC752_n_13889 ( .a(n_13889), .o(FE_OFN752_n_13889) );
in01s01 FE_OFC753_n_13889 ( .a(FE_OFN752_n_13889), .o(FE_OFN753_n_13889) );
in01m04 FE_OFC754_n_13889 ( .a(FE_OFN752_n_13889), .o(FE_OFN754_n_13889) );
in01s10 FE_OFC755_n_44464 ( .a(FE_OFN4772_n_44463), .o(FE_OFN755_n_44464) );
in01s20 FE_OFC756_n_44464 ( .a(FE_OFN755_n_44464), .o(FE_OFN756_n_44464) );
in01s02 FE_OFC757_n_44464 ( .a(FE_OFN755_n_44464), .o(FE_OFN757_n_44464) );
in01s02 FE_OFC758_n_45813 ( .a(n_45813), .o(FE_OFN758_n_45813) );
in01s02 FE_OFC759_n_45813 ( .a(FE_OFN758_n_45813), .o(FE_OFN759_n_45813) );
in01s02 FE_OFC765_n_46337 ( .a(FE_OCP_RBN6163_n_46337), .o(FE_OFN765_n_46337) );
in01s01 FE_OFC766_n_46137 ( .a(n_46137), .o(FE_OFN766_n_46137) );
in01f08 FE_OFC767_n_46137 ( .a(n_46137), .o(FE_OFN767_n_46137) );
in01s02 FE_OFC768_n_46137 ( .a(FE_OFN766_n_46137), .o(FE_OFN768_n_46137) );
in01s02 FE_OFC769_n_46196 ( .a(n_46195), .o(FE_OFN769_n_46196) );
in01s03 FE_OFC770_n_46196 ( .a(FE_OFN769_n_46196), .o(FE_OFN770_n_46196) );
in01s04 FE_OFC771_n_46196 ( .a(FE_OFN769_n_46196), .o(FE_OFN771_n_46196) );
in01s06 FE_OFC772_n_25834 ( .a(n_25834), .o(FE_OFN772_n_25834) );
in01f03 FE_OFC773_n_25834 ( .a(FE_OFN772_n_25834), .o(FE_OFN773_n_25834) );
in01s40 FE_OFC774_n_25834 ( .a(FE_OFN772_n_25834), .o(FE_OFN774_n_25834) );
in01s01 FE_OFC775_n_25834 ( .a(FE_OFN772_n_25834), .o(FE_RN_2448_0) );
in01m06 FE_OFC776_n_18268 ( .a(n_18268), .o(FE_OFN776_n_18268) );
in01m10 FE_OFC777_n_18268 ( .a(FE_OFN776_n_18268), .o(FE_OFN777_n_18268) );
in01s02 FE_OFC778_n_23803 ( .a(n_23803), .o(FE_OFN778_n_23803) );
in01s02 FE_OFC779_n_23803 ( .a(FE_OFN778_n_23803), .o(FE_OFN779_n_23803) );
in01s04 FE_OFC780_n_23803 ( .a(FE_OFN778_n_23803), .o(FE_OFN780_n_23803) );
in01s01 FE_OFC781_n_47017 ( .a(n_47017), .o(FE_OFN781_n_47017) );
in01s02 FE_OFC787_n_46285 ( .a(FE_OCP_RBN6144_n_46285), .o(FE_OFN787_n_46285) );
in01m06 FE_OFC789_n_46195 ( .a(n_46195), .o(FE_OFN789_n_46195) );
in01s01 FE_OFC792_n_1909 ( .a(FE_OFN813_n_1909), .o(FE_OFN792_n_1909) );
in01s01 FE_OFC793_n_2056 ( .a(FE_OFN814_n_2056), .o(FE_OFN793_n_2056) );
in01s01 FE_OFC794_n_2929 ( .a(n_2929), .o(FE_OFN794_n_2929) );
in01s01 FE_OFC795_n_19885 ( .a(FE_OFN815_n_19885), .o(FE_OFN795_n_19885) );
in01s01 FE_OFC796_n_2719 ( .a(FE_OFN816_n_2719), .o(FE_OFN796_n_2719) );
in01s01 FE_OFC797_n_2285 ( .a(FE_OFN819_n_2285), .o(FE_OFN797_n_2285) );
in01s01 FE_OFC798_n_2620 ( .a(FE_OFN818_n_2620), .o(FE_OFN798_n_2620) );
in01s01 FE_OFC799_n_2644 ( .a(FE_OFN817_n_2644), .o(FE_OFN799_n_2644) );
in01s01 FE_OFC800_n_3771 ( .a(FE_OFN820_n_3771), .o(FE_OFN800_n_3771) );
in01s01 FE_OFC801_n_3902 ( .a(FE_OFN821_n_3902), .o(FE_OFN801_n_3902) );
in01s01 FE_OFC802_n_3911 ( .a(FE_OFN825_n_3911), .o(FE_OFN802_n_3911) );
in01s01 FE_OFC803_n_4142 ( .a(FE_OFN826_n_4142), .o(FE_OFN803_n_4142) );
in01s01 FE_OFC804_n_4575 ( .a(FE_OFN827_n_4575), .o(FE_OFN804_n_4575) );
in01s01 FE_OFC805_n_4018 ( .a(n_4018), .o(FE_OFN805_n_4018) );
in01s01 FE_OFC806_n_13742 ( .a(FE_OFN829_n_13742), .o(FE_OFN806_n_13742) );
in01s01 FE_OFC807_n_4686 ( .a(FE_OFN828_n_4686), .o(FE_OFN807_n_4686) );
in01s01 FE_OFC808_n_3264 ( .a(FE_OFN830_n_3264), .o(FE_OFN808_n_3264) );
in01s01 FE_OFC809_n_9939 ( .a(FE_OFN831_n_9939), .o(FE_OFN809_n_9939) );
in01s01 FE_OFC810_n_9028 ( .a(FE_OFN832_n_9028), .o(FE_OFN810_n_9028) );
in01s01 FE_OFC812_n_902 ( .a(n_902), .o(FE_OFN812_n_902) );
in01s01 FE_OFC813_n_1909 ( .a(n_1909), .o(FE_OFN813_n_1909) );
in01s01 FE_OFC814_n_2056 ( .a(n_2056), .o(FE_OFN814_n_2056) );
in01s01 FE_OFC815_n_19885 ( .a(n_19885), .o(FE_OFN815_n_19885) );
in01s01 FE_OFC816_n_2719 ( .a(n_2719), .o(FE_OFN816_n_2719) );
in01s01 FE_OFC817_n_2644 ( .a(n_2644), .o(FE_OFN817_n_2644) );
in01s01 FE_OFC818_n_2620 ( .a(n_2620), .o(FE_OFN818_n_2620) );
in01s01 FE_OFC819_n_2285 ( .a(n_2285), .o(FE_OFN819_n_2285) );
in01s01 FE_OFC81_n_4117 ( .a(n_4117), .o(FE_OFN81_n_4117) );
in01s01 FE_OFC820_n_3771 ( .a(n_3771), .o(FE_OFN820_n_3771) );
in01s01 FE_OFC821_n_3902 ( .a(n_3902), .o(FE_OFN821_n_3902) );
in01s01 FE_OFC822_n_1045 ( .a(n_1045), .o(FE_OFN822_n_1045) );
in01s01 FE_OFC823_n_1045 ( .a(FE_OFN822_n_1045), .o(FE_OFN823_n_1045) );
in01s01 FE_OFC824_n_1045 ( .a(FE_OFN822_n_1045), .o(FE_OFN824_n_1045) );
in01s01 FE_OFC825_n_3911 ( .a(n_3911), .o(FE_OFN825_n_3911) );
in01s01 FE_OFC826_n_4142 ( .a(n_4142), .o(FE_OFN826_n_4142) );
in01s01 FE_OFC827_n_4575 ( .a(n_4575), .o(FE_OFN827_n_4575) );
in01s01 FE_OFC828_n_4686 ( .a(n_4686), .o(FE_OFN828_n_4686) );
in01s01 FE_OFC829_n_13742 ( .a(n_13742), .o(FE_OFN829_n_13742) );
in01s01 FE_OFC82_n_4117 ( .a(FE_OFN81_n_4117), .o(FE_OFN82_n_4117) );
in01s01 FE_OFC830_n_3264 ( .a(n_3264), .o(FE_OFN830_n_3264) );
in01s01 FE_OFC831_n_9939 ( .a(n_9939), .o(FE_OFN831_n_9939) );
in01s01 FE_OFC832_n_9028 ( .a(n_9028), .o(FE_OFN832_n_9028) );
oa22m02 FE_RC_0_0 ( .a(n_18128), .b(n_18283), .c(n_18129), .d(n_18282), .o(n_18405) );
na02f08 FE_RC_1001_0 ( .a(FE_RN_306_0), .b(FE_RN_307_0), .o(FE_RN_308_0) );
ao22f04 FE_RC_1005_0 ( .a(n_13418), .b(n_14072), .c(n_13514), .d(FE_OCP_RBN2728_n_14072), .o(n_14177) );
oa22f02 FE_RC_1006_0 ( .a(FE_OCPN935_n_7802), .b(n_8548), .c(FE_OCP_RBN4138_n_7743), .d(FE_OCP_RBN5734_n_8548), .o(n_8696) );
ao22m04 FE_RC_1007_0 ( .a(n_2913), .b(n_3385), .c(FE_OCP_RBN2629_n_2737), .d(n_4228), .o(n_3481) );
oa22m06 FE_RC_1008_0 ( .a(n_33404), .b(n_33875), .c(n_33900), .d(n_33405), .o(n_33976) );
oa22m02 FE_RC_1009_0 ( .a(n_8376), .b(n_7498), .c(n_7499), .d(n_8386), .o(n_8474) );
oa22s06 FE_RC_1010_0 ( .a(n_14021), .b(n_13420), .c(n_14022), .d(n_13419), .o(n_14157) );
oa22s06 FE_RC_1011_0 ( .a(FE_OFN1180_n_13195), .b(n_14157), .c(n_13469), .d(FE_OCP_RBN2749_n_14157), .o(n_14323) );
oa22s02 FE_RC_1019_0 ( .a(n_17177), .b(n_17487), .c(n_17176), .d(n_17512), .o(n_17688) );
oa22f04 FE_RC_1022_0 ( .a(n_14367), .b(FE_OCP_RBN2727_n_14018), .c(n_14366), .d(FE_OCP_RBN2726_n_14018), .o(n_14544) );
no02s01 TIMEBOOST_cell_6157 ( .a(n_26512), .b(FE_OCP_RBN6097_n_26160), .o(TIMEBOOST_net_1930) );
in01s02 FE_RC_1024_0 ( .a(n_8196), .o(FE_RN_310_0) );
in01m02 FE_RC_1025_0 ( .a(FE_RN_311_0), .o(n_8271) );
no02s01 TIMEBOOST_cell_6158 ( .a(TIMEBOOST_net_1930), .b(n_26486), .o(n_26611) );
ao22s04 FE_RC_1028_0 ( .a(n_3641), .b(n_2913), .c(FE_OFN4764_n_3029), .d(n_4528), .o(n_3720) );
oa22m04 FE_RC_1029_0 ( .a(FE_OCP_RBN4190_n_14279), .b(n_13207), .c(n_13206), .d(n_14279), .o(n_14444) );
ao22m04 FE_RC_1036_0 ( .a(n_2905), .b(n_3595), .c(n_2904), .d(n_3636), .o(n_3807) );
ao22m06 FE_RC_1037_0 ( .a(n_23964), .b(n_24563), .c(n_23965), .d(n_24562), .o(n_24684) );
oa22f04 FE_RC_1038_0 ( .a(n_28824), .b(n_29343), .c(n_28825), .d(n_29344), .o(n_29485) );
ao22f04 FE_RC_103_0 ( .a(n_20506), .b(n_20310), .c(n_20505), .d(n_20312), .o(n_20640) );
ao22s04 FE_RC_1043_0 ( .a(n_28822), .b(n_29384), .c(n_28823), .d(n_29383), .o(n_29479) );
oa22f06 FE_RC_1047_0 ( .a(n_42155), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .c(n_42196), .d(n_42154), .o(n_42182) );
oa22m04 FE_RC_1049_0 ( .a(n_9527), .b(FE_OCP_RBN3011_n_9565), .c(n_9565), .d(n_9528), .o(n_9742) );
no02m06 TIMEBOOST_cell_8877 ( .a(TIMEBOOST_net_2925), .b(n_27124), .o(TIMEBOOST_net_2687) );
oa22f06 FE_RC_1055_0 ( .a(delay_sub_ln23_0_unr29_stage10_stallmux_q), .b(n_42128), .c(n_42196), .d(n_42129), .o(n_42156) );
oa22m04 FE_RC_1057_0 ( .a(n_38198), .b(FE_OCP_RBN5689_n_38531), .c(n_38197), .d(n_38531), .o(n_38586) );
ao22s02 FE_RC_1061_0 ( .a(FE_OCP_RBN6770_n_3700), .b(n_47014), .c(FE_OCP_RBN5870_n_3704), .d(FE_OCP_RBN4289_n_47014), .o(n_4030) );
in01s01 FE_RC_1062_0 ( .a(n_25859), .o(FE_RN_315_0) );
na02s02 TIMEBOOST_cell_4937 ( .a(TIMEBOOST_net_1416), .b(n_7160), .o(n_7244) );
in01m04 FE_RC_1064_0 ( .a(FE_RN_317_0), .o(n_29533) );
no02m06 TIMEBOOST_cell_4947 ( .a(TIMEBOOST_net_1421), .b(TIMEBOOST_net_140), .o(n_12469) );
ao22m04 FE_RC_1066_0 ( .a(n_40139), .b(n_40521), .c(n_40140), .d(n_40531), .o(n_40568) );
no02m06 TIMEBOOST_cell_3115 ( .a(n_10720), .b(TIMEBOOST_net_848), .o(n_10869) );
in01f02 FE_RC_1068_0 ( .a(n_9556), .o(FE_RN_319_0) );
in01f04 FE_RC_1069_0 ( .a(FE_RN_320_0), .o(n_9926) );
no02s06 TIMEBOOST_cell_3116 ( .a(FE_RN_678_0), .b(FE_RN_677_0), .o(TIMEBOOST_net_849) );
oa22f04 FE_RC_1071_0 ( .a(n_22393), .b(n_24932), .c(FE_OCPN1354_n_22484), .d(n_24933), .o(n_25036) );
oa22s04 FE_RC_1072_0 ( .a(n_24684), .b(n_24870), .c(n_24717), .d(n_24850), .o(n_24934) );
na02m06 TIMEBOOST_cell_5983 ( .a(n_12207), .b(n_12401), .o(TIMEBOOST_net_1843) );
in01m08 FE_RC_1075_0 ( .a(FE_RN_323_0), .o(n_25453) );
no02m08 TIMEBOOST_cell_4297 ( .a(TIMEBOOST_net_807), .b(FE_RN_1051_0), .o(TIMEBOOST_net_1239) );
ao22m02 FE_RC_1080_0 ( .a(n_7632), .b(n_8700), .c(n_45503), .d(n_7631), .o(n_8767) );
oa22s01 FE_RC_1083_0 ( .a(FE_OCP_RBN6715_n_3604), .b(n_5109), .c(n_3381), .d(FE_OCP_RBN4255_n_3705), .o(n_3929) );
in01s01 FE_RC_1086_0 ( .a(n_4416), .o(FE_RN_324_0) );
in01s02 FE_RC_1087_0 ( .a(n_4363), .o(FE_RN_325_0) );
no02s04 FE_RC_1088_0 ( .a(FE_RN_324_0), .b(FE_RN_325_0), .o(FE_RN_326_0) );
no02s01 TIMEBOOST_cell_6129 ( .a(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n_22089), .o(TIMEBOOST_net_1916) );
oa22m02 FE_RC_1090_0 ( .a(n_8536), .b(n_8654), .c(n_8570), .d(n_8653), .o(n_8781) );
oa22f02 FE_RC_1091_0 ( .a(n_38624), .b(n_38673), .c(n_38637), .d(n_38674), .o(n_38747) );
ao22f04 FE_RC_1092_0 ( .a(FE_OCP_RBN2890_n_14460), .b(FE_OCP_RBN4205_n_13796), .c(n_14460), .d(FE_OCP_RBN6695_n_13796), .o(n_14591) );
ao22m04 FE_RC_1093_0 ( .a(n_38778), .b(n_38606), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .d(n_38605), .o(n_38669) );
oa22f02 FE_RC_1095_0 ( .a(FE_OCP_RBN6707_n_8719), .b(n_8859), .c(n_8719), .d(n_8836), .o(n_9009) );
ao22f02 FE_RC_1096_0 ( .a(n_8934), .b(n_8899), .c(n_8891), .d(n_8898), .o(n_9075) );
in01m03 FE_RC_10_0 ( .a(n_18051), .o(FE_RN_4_0) );
ao22f04 FE_RC_1101_0 ( .a(FE_OCP_RBN2926_n_14684), .b(FE_OCP_RBN2834_n_13962), .c(FE_OCP_RBN6700_n_13796), .d(n_14684), .o(n_14785) );
oa22f04 FE_RC_1102_0 ( .a(n_33643), .b(FE_OCP_RBN2543_n_33584), .c(n_33584), .d(n_33660), .o(n_33757) );
oa22f02 FE_RC_1105_0 ( .a(FE_OCP_RBN6732_n_44579), .b(FE_OCP_RBN6749_n_9198), .c(FE_OCP_RBN6738_n_44563), .d(n_9198), .o(n_9410) );
in01s01 FE_RC_110_0 ( .a(n_17572), .o(FE_RN_21_0) );
oa22m06 FE_RC_1111_0 ( .a(FE_OCP_RBN6731_n_44579), .b(FE_OCP_RBN5972_n_9494), .c(FE_OCP_RBN6738_n_44563), .d(n_9494), .o(n_9666) );
ao22m06 FE_RC_1115_0 ( .a(n_34423), .b(n_34908), .c(n_34424), .d(FE_OCP_RBN5854_n_34908), .o(n_35005) );
oa22f04 FE_RC_1116_0 ( .a(n_14618), .b(n_46982), .c(FE_OCP_RBN4369_n_46982), .d(n_14452), .o(n_15761) );
ao22m08 FE_RC_1118_0 ( .a(n_34703), .b(n_35026), .c(n_34702), .d(n_35048), .o(n_35132) );
in01s01 FE_RC_1119_0 ( .a(n_15636), .o(FE_RN_327_0) );
in01s02 FE_RC_111_0 ( .a(n_17613), .o(FE_RN_22_0) );
in01s03 FE_RC_1120_0 ( .a(n_15857), .o(FE_RN_328_0) );
no02s06 FE_RC_1121_0 ( .a(FE_RN_328_0), .b(FE_RN_327_0), .o(FE_RN_329_0) );
oa22m04 FE_RC_1123_0 ( .a(FE_OCP_RBN5939_n_44563), .b(FE_OCP_RBN3091_n_10023), .c(FE_OCP_RBN5911_n_44563), .d(n_10023), .o(n_10192) );
oa22m06 FE_RC_1124_0 ( .a(n_15908), .b(n_15601), .c(n_15602), .d(n_15909), .o(n_16088) );
oa22f04 FE_RC_1126_0 ( .a(n_15453), .b(n_15858), .c(n_15454), .d(n_15815), .o(n_16053) );
oa22f02 FE_RC_1129_0 ( .a(n_5098), .b(n_45322), .c(n_5099), .d(n_45321), .o(n_5444) );
na02s03 FE_RC_112_0 ( .a(FE_RN_22_0), .b(FE_RN_21_0), .o(FE_RN_23_0) );
oa22m06 FE_RC_1130_0 ( .a(n_25583), .b(n_25925), .c(FE_OCP_RBN3150_n_25925), .d(n_25584), .o(n_26045) );
oa22m04 FE_RC_1134_0 ( .a(n_10494), .b(n_10880), .c(n_10881), .d(n_10495), .o(n_11004) );
in01s01 FE_RC_1136_0 ( .a(n_30292), .o(FE_RN_330_0) );
in01s04 FE_RC_1137_0 ( .a(n_30535), .o(FE_RN_331_0) );
na02m08 TIMEBOOST_cell_1091 ( .a(FE_RN_1716_0), .b(n_32919), .o(TIMEBOOST_net_160) );
na02f08 TIMEBOOST_cell_1092 ( .a(FE_RN_1715_0), .b(TIMEBOOST_net_160), .o(n_33207) );
ao22m06 FE_RC_1140_0 ( .a(n_30316), .b(n_30610), .c(n_30317), .d(n_30609), .o(n_30711) );
na03m04 FE_RC_1141_0 ( .a(n_6162), .b(n_6187), .c(n_6188), .o(n_6189) );
in01s01 FE_RC_1153_0 ( .a(n_30281), .o(FE_RN_336_0) );
in01m04 FE_RC_1154_0 ( .a(n_30644), .o(FE_RN_337_0) );
na02m08 FE_RC_1155_0 ( .a(FE_RN_337_0), .b(FE_RN_336_0), .o(FE_RN_338_0) );
na02m08 FE_RC_1156_0 ( .a(FE_RN_338_0), .b(n_30675), .o(n_46958) );
ao22m06 FE_RC_1157_0 ( .a(n_21197), .b(FE_OCP_RBN3118_n_20812), .c(n_20812), .d(n_21198), .o(n_21360) );
ao22m04 FE_RC_1158_0 ( .a(n_45024), .b(n_21194), .c(n_45026), .d(FE_OCP_RBN6060_n_21194), .o(n_21361) );
ao22m04 FE_RC_1159_0 ( .a(n_26324), .b(n_25722), .c(FE_OCPN1675_n_25721), .d(n_26376), .o(n_26464) );
oa22f04 FE_RC_1161_0 ( .a(n_16390), .b(n_16530), .c(n_16391), .d(n_16531), .o(n_16622) );
oa22s04 FE_RC_1164_0 ( .a(n_46956), .b(FE_OCP_DRV_N6897_FE_OCPN1679_n_27315), .c(n_27366), .d(n_31017), .o(n_31101) );
oa22m04 FE_RC_1165_0 ( .a(n_21636), .b(n_21492), .c(n_21491), .d(FE_OCP_RBN6101_n_21636), .o(n_21789) );
oa22f08 FE_RC_1168_0 ( .a(n_26456), .b(n_27008), .c(n_26487), .d(n_27017), .o(n_27083) );
oa22s02 FE_RC_1170_0 ( .a(FE_OFN787_n_46285), .b(n_12196), .c(FE_OCP_RBN3352_FE_OFN760_n_46337), .d(FE_OCP_RBN3458_n_12196), .o(n_46347) );
oa22s02 FE_RC_1171_0 ( .a(FE_OFN787_n_46285), .b(n_12197), .c(FE_OCP_RBN3352_FE_OFN760_n_46337), .d(n_12116), .o(n_46350) );
ao22s04 FE_RC_1172_0 ( .a(n_36139), .b(FE_OCP_RBN6177_n_36444), .c(n_36140), .d(n_36444), .o(n_36515) );
oa22s02 FE_RC_1173_0 ( .a(FE_OFN787_n_46285), .b(n_12217), .c(FE_OCP_RBN3352_FE_OFN760_n_46337), .d(n_12190), .o(n_46344) );
oa22s01 FE_RC_1181_0 ( .a(n_36754), .b(n_36778), .c(n_36753), .d(FE_OCP_RBN6234_n_36778), .o(n_36830) );
oa22s02 FE_RC_1182_0 ( .a(n_17584), .b(n_17725), .c(n_17753), .d(n_17674), .o(n_17769) );
oa22m02 FE_RC_1183_0 ( .a(n_17336), .b(n_17686), .c(FE_OCP_RBN3196_n_15599), .d(n_44153), .o(n_17755) );
oa22f02 FE_RC_1184_0 ( .a(FE_OCP_RBN3199_n_15599), .b(n_17685), .c(n_17753), .d(n_44147), .o(n_17754) );
oa22s02 FE_RC_1185_0 ( .a(n_17584), .b(n_17723), .c(n_17753), .d(FE_OCP_RBN6254_n_17723), .o(n_17770) );
oa22f02 FE_RC_1186_0 ( .a(n_17336), .b(n_17697), .c(n_16339), .d(FE_OCP_RBN3450_n_17697), .o(n_17776) );
oa22f02 FE_RC_1194_0 ( .a(FE_OCPN1394_n_22801), .b(FE_OCP_RBN6241_n_22622), .c(n_22580), .d(n_22622), .o(n_22742) );
oa22f02 FE_RC_1195_0 ( .a(n_22961), .b(n_22631), .c(n_20252), .d(n_22611), .o(n_22704) );
oa22m02 FE_RC_1197_0 ( .a(n_20231), .b(n_22774), .c(n_22751), .d(n_22580), .o(n_22826) );
oa22m02 FE_RC_1199_0 ( .a(n_17336), .b(n_17630), .c(FE_OCP_RBN3196_n_15599), .d(n_17628), .o(n_17731) );
in01s06 FE_RC_119_0 ( .a(n_17970), .o(FE_RN_27_0) );
na02s10 FE_RC_11_0 ( .a(FE_RN_3_0), .b(FE_RN_4_0), .o(FE_RN_5_0) );
no03s02 TIMEBOOST_cell_7728 ( .a(n_26549), .b(n_26510), .c(FE_OCP_RBN6097_n_26160), .o(TIMEBOOST_net_2495) );
in01s02 FE_RC_1202_0 ( .a(n_17391), .o(FE_RN_340_0) );
in01m02 FE_RC_1203_0 ( .a(FE_RN_341_0), .o(n_17495) );
na02m08 TIMEBOOST_cell_7455 ( .a(TIMEBOOST_net_2358), .b(n_11984), .o(n_12137) );
oa22s02 FE_RC_1207_0 ( .a(n_17387), .b(n_17657), .c(n_17386), .d(n_17629), .o(n_17811) );
oa22s02 FE_RC_1208_0 ( .a(n_17378), .b(n_17627), .c(n_17379), .d(n_17601), .o(n_17759) );
in01s06 FE_RC_120_0 ( .a(n_17971), .o(FE_RN_28_0) );
oa22f02 FE_RC_1210_0 ( .a(FE_OFN621_n_28336), .b(n_44216), .c(n_32287), .d(n_32290), .o(n_32337) );
oa22s01 FE_RC_1212_0 ( .a(n_17336), .b(n_17759), .c(n_17753), .d(n_44334), .o(n_17832) );
no02s01 TIMEBOOST_cell_7665 ( .a(TIMEBOOST_net_2463), .b(FE_OCP_RBN6626_n_2537), .o(n_2718) );
in01s01 FE_RC_1215_0 ( .a(FE_RN_344_0), .o(n_17600) );
no03f08 TIMEBOOST_cell_3498 ( .a(n_32697), .b(FE_OCP_RBN2434_n_32702), .c(FE_RN_1631_0), .o(n_32722) );
oa22m02 FE_RC_1219_0 ( .a(n_32287), .b(n_32338), .c(FE_OFN621_n_28336), .d(n_44432), .o(n_32373) );
na03m20 TIMEBOOST_cell_2154 ( .a(FE_RN_2103_0), .b(n_44061), .c(n_22634), .o(TIMEBOOST_net_15) );
oa22s06 FE_RC_1220_0 ( .a(n_17382), .b(n_17689), .c(n_17383), .d(FE_OCP_RBN1875_n_17689), .o(n_17834) );
oa22m02 FE_RC_1223_0 ( .a(n_32287), .b(FE_OCP_RBN3441_n_32266), .c(FE_OFN621_n_28336), .d(n_32266), .o(n_32334) );
oa22m02 FE_RC_1224_0 ( .a(n_32566), .b(n_32340), .c(FE_OFN621_n_28336), .d(FE_OCP_RBN5055_n_32340), .o(n_32374) );
ao22s02 FE_RC_1229_0 ( .a(n_27501), .b(n_27648), .c(n_27649), .d(n_27500), .o(n_27729) );
na03f10 TIMEBOOST_cell_6435 ( .a(n_23412), .b(n_23144), .c(n_23396), .o(n_23502) );
in01s01 FE_RC_1233_0 ( .a(n_27373), .o(FE_RN_345_0) );
na03m08 TIMEBOOST_cell_3519 ( .a(FE_RN_2718_0), .b(FE_RN_2719_0), .c(FE_RN_2721_0), .o(TIMEBOOST_net_741) );
in01s01 FE_RC_1235_0 ( .a(FE_RN_347_0), .o(n_27690) );
na02s01 TIMEBOOST_cell_4858 ( .a(FE_OCP_RBN6410_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(n_1369), .o(TIMEBOOST_net_1377) );
oa22s01 FE_RC_1237_0 ( .a(n_32566), .b(n_32518), .c(n_28336), .d(FE_OCP_RBN5349_n_32518), .o(n_32571) );
oa22s02 FE_RC_1238_0 ( .a(n_32287), .b(n_32468), .c(n_28336), .d(n_32395), .o(n_32515) );
oa22f01 FE_RC_1239_0 ( .a(n_28336), .b(n_32466), .c(n_32566), .d(n_32517), .o(n_32565) );
oa22s01 FE_RC_1241_0 ( .a(n_24350), .b(n_27781), .c(n_27796), .d(n_27752), .o(n_27838) );
oa22m01 FE_RC_1242_0 ( .a(n_24350), .b(n_27768), .c(n_27796), .d(n_27736), .o(n_27797) );
oa22s01 FE_RC_1243_0 ( .a(n_24350), .b(n_27782), .c(n_27845), .d(n_45309), .o(n_27836) );
oa22s01 FE_RC_1244_0 ( .a(n_24350), .b(n_27755), .c(n_27845), .d(n_27729), .o(n_27780) );
oa22s01 FE_RC_1245_0 ( .a(FE_OFN1183_n_24059), .b(n_27784), .c(n_27845), .d(n_27757), .o(n_27846) );
oa22s01 FE_RC_1246_0 ( .a(n_24350), .b(n_27783), .c(n_27845), .d(n_27756), .o(n_27844) );
oa22s01 FE_RC_1247_0 ( .a(FE_OFN1183_n_24059), .b(n_27785), .c(n_27796), .d(n_27758), .o(n_27843) );
no02s04 TIMEBOOST_cell_1636 ( .a(TIMEBOOST_net_432), .b(n_30578), .o(n_30623) );
oa22m01 FE_RC_1250_0 ( .a(n_32287), .b(FE_OCP_RBN5058_n_32427), .c(n_28336), .d(n_32427), .o(n_32541) );
oa22f02 FE_RC_1251_0 ( .a(FE_OCPN1394_n_22801), .b(n_22684), .c(n_22833), .d(n_22637), .o(n_22758) );
oa22s01 FE_RC_1252_0 ( .a(n_32287), .b(n_32519), .c(n_28336), .d(n_32469), .o(n_32569) );
oa22f02 FE_RC_1254_0 ( .a(n_22961), .b(n_22778), .c(n_22580), .d(n_22757), .o(n_22832) );
ao22m02 FE_RC_1256_0 ( .a(n_45496), .b(n_22309), .c(n_45497), .d(n_22272), .o(n_22710) );
oa22s06 FE_RC_1257_0 ( .a(n_22379), .b(n_22618), .c(n_22380), .d(n_22636), .o(n_22806) );
oa22m02 FE_RC_1258_0 ( .a(FE_OCPN1394_n_22801), .b(FE_OCP_RBN3451_n_22710), .c(n_22833), .d(n_22710), .o(n_22802) );
in01s03 FE_RC_125_0 ( .a(n_17765), .o(FE_RN_30_0) );
oa22s02 FE_RC_1260_0 ( .a(n_20231), .b(n_22875), .c(n_22833), .d(n_44329), .o(n_22949) );
oa22m02 FE_RC_1261_0 ( .a(n_22961), .b(FE_OCP_RBN4492_n_22755), .c(n_22833), .d(n_22755), .o(n_22834) );
oa22m02 FE_RC_1262_0 ( .a(n_20231), .b(n_22914), .c(n_22793), .d(n_22871), .o(n_22973) );
oa22s02 FE_RC_1263_0 ( .a(n_20231), .b(n_22835), .c(n_22580), .d(n_22804), .o(n_22913) );
oa22s02 FE_RC_1264_0 ( .a(FE_OFN1183_n_24059), .b(n_27799), .c(n_27796), .d(n_27766), .o(n_27855) );
oa22f01 FE_RC_1265_0 ( .a(n_24350), .b(n_27835), .c(n_27796), .d(n_27795), .o(n_27894) );
oa22s02 FE_RC_1266_0 ( .a(n_24350), .b(n_27800), .c(n_27796), .d(n_27767), .o(n_27858) );
oa22s01 FE_RC_1267_0 ( .a(n_24350), .b(n_27771), .c(n_27845), .d(n_27744), .o(n_27819) );
oa22s02 FE_RC_1269_0 ( .a(n_24350), .b(n_27772), .c(n_27796), .d(n_27745), .o(n_27818) );
in01s06 FE_RC_126_0 ( .a(n_17885), .o(FE_RN_31_0) );
no02s06 TIMEBOOST_cell_1892 ( .a(TIMEBOOST_net_560), .b(n_40059), .o(n_40104) );
no02s10 TIMEBOOST_cell_7417 ( .a(TIMEBOOST_net_2339), .b(n_17341), .o(n_17507) );
na02m06 FE_RC_127_0 ( .a(FE_RN_31_0), .b(FE_RN_30_0), .o(FE_RN_32_0) );
oa22f10 FE_RC_1281_0 ( .a(delay_xor_ln23_unr6_stage3_stallmux_q), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(n_6505), .d(FE_OCP_RBN6440_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6528) );
na03s01 TIMEBOOST_cell_4676 ( .a(n_2878), .b(n_2877), .c(n_2913), .o(FE_RN_899_0) );
in01s02 FE_RC_1283_0 ( .a(n_17973), .o(FE_RN_348_0) );
in01s01 FE_RC_1284_0 ( .a(n_18113), .o(FE_RN_349_0) );
no02s04 TIMEBOOST_cell_5091 ( .a(TIMEBOOST_net_1493), .b(n_2361), .o(n_2511) );
in01s01 TIMEBOOST_cell_8911 ( .a(TIMEBOOST_net_2954), .o(TIMEBOOST_net_2955) );
in01m01 FE_RC_1293_0 ( .a(n_18133), .o(FE_RN_354_0) );
in01s02 FE_RC_1294_0 ( .a(n_18135), .o(FE_RN_355_0) );
na02s08 TIMEBOOST_cell_4923 ( .a(n_7144), .b(TIMEBOOST_net_1409), .o(n_7222) );
na02f04 TIMEBOOST_cell_6238 ( .a(TIMEBOOST_net_1970), .b(n_36222), .o(n_35681) );
oa22f04 FE_RC_1298_0 ( .a(n_27632), .b(n_27497), .c(n_27496), .d(FE_OCP_RBN3453_n_27632), .o(n_27728) );
oa22f02 FE_RC_1299_0 ( .a(FE_OFN1183_n_24059), .b(n_27728), .c(n_27796), .d(n_27706), .o(n_27750) );
no02s04 TIMEBOOST_cell_1664 ( .a(TIMEBOOST_net_446), .b(n_20137), .o(n_20181) );
oa22m06 FE_RC_1300_0 ( .a(n_38109), .b(n_38449), .c(n_38108), .d(n_38448), .o(n_38530) );
ao22m02 FE_RC_1303_0 ( .a(FE_OCP_RBN5753_n_4022), .b(n_3405), .c(n_4022), .d(n_3373), .o(n_3495) );
na02m04 TIMEBOOST_cell_2141 ( .a(FE_OCP_RBN1871_n_36489), .b(n_36750), .o(TIMEBOOST_net_685) );
ao22m04 FE_RC_1307_0 ( .a(n_3015), .b(n_3935), .c(n_3014), .d(n_3859), .o(n_4158) );
no02f02 TIMEBOOST_cell_1607 ( .a(FE_OCP_RBN6754_n_38806), .b(n_38882), .o(TIMEBOOST_net_418) );
oa22m02 FE_RC_1315_0 ( .a(FE_OCP_RBN3193_n_15599), .b(FE_OCP_RBN6245_n_17587), .c(n_17753), .d(n_17587), .o(n_17677) );
ao22f04 FE_RC_1316_0 ( .a(n_4880), .b(n_4816), .c(n_4815), .d(n_4881), .o(n_5049) );
oa22m02 FE_RC_1317_0 ( .a(FE_OCP_RBN2962_n_4046), .b(n_4784), .c(FE_OCP_RBN2966_n_4046), .d(FE_OCP_RBN3123_n_4784), .o(n_4959) );
in01f10 FE_RC_1318_0 ( .a(n_27839), .o(FE_RN_360_0) );
in01s08 FE_RC_1319_0 ( .a(n_27919), .o(FE_RN_361_0) );
no03f08 TIMEBOOST_cell_2367 ( .a(n_33621), .b(n_33581), .c(n_33644), .o(n_33715) );
no02f02 TIMEBOOST_cell_8667 ( .a(TIMEBOOST_net_2820), .b(n_31097), .o(TIMEBOOST_net_1718) );
oa22f02 FE_RC_1323_0 ( .a(FE_OFN787_n_46285), .b(n_12211), .c(FE_OFN765_n_46337), .d(n_12151), .o(n_46342) );
oa22s02 FE_RC_1324_0 ( .a(FE_OFN787_n_46285), .b(FE_OCP_RBN6251_n_12067), .c(FE_OFN765_n_46337), .d(n_12067), .o(n_46358) );
oa22s01 FE_RC_1326_0 ( .a(n_17336), .b(n_44447), .c(n_16339), .d(n_17729), .o(n_17808) );
oa22m04 FE_RC_1328_0 ( .a(n_12027), .b(n_11806), .c(n_11807), .d(n_12028), .o(n_12240) );
oa22m02 FE_RC_1329_0 ( .a(FE_OFN787_n_46285), .b(n_12240), .c(FE_OFN765_n_46337), .d(n_12189), .o(n_46340) );
oa22m02 FE_RC_1330_0 ( .a(FE_OCPN931_n_7817), .b(FE_OCP_RBN2781_n_8664), .c(FE_OCP_RBN2599_n_7743), .d(n_8664), .o(n_8803) );
in01s01 FE_RC_1331_0 ( .a(n_39426), .o(FE_RN_363_0) );
in01s01 FE_RC_1332_0 ( .a(n_39840), .o(FE_RN_364_0) );
no02s01 FE_RC_1333_0 ( .a(FE_RN_363_0), .b(FE_RN_364_0), .o(FE_RN_365_0) );
no02f08 FE_RC_1334_0 ( .a(n_39812), .b(FE_RN_365_0), .o(n_39907) );
oa22m04 FE_RC_1335_0 ( .a(FE_OCP_RBN6683_FE_OCPN4529_FE_OCP_RBN2748_n_8474), .b(FE_OCP_RBN2856_n_8755), .c(FE_OCP_RBN6684_FE_OCPN4529_FE_OCP_RBN2748_n_8474), .d(n_8755), .o(n_8889) );
oa22f02 FE_RC_1339_0 ( .a(n_17584), .b(n_17550), .c(n_17753), .d(n_17475), .o(n_17585) );
oa22f02 FE_RC_1343_0 ( .a(n_40598), .b(n_40577), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .d(n_44690), .o(n_40589) );
ao22m02 FE_RC_1345_0 ( .a(n_7591), .b(n_8788), .c(n_7590), .d(n_8769), .o(n_8915) );
oa22m02 FE_RC_1347_0 ( .a(n_11588), .b(n_11652), .c(n_11587), .d(n_11702), .o(n_11873) );
oa22s02 FE_RC_1348_0 ( .a(FE_OCP_RBN6865_n_46285), .b(n_11873), .c(FE_OCP_RBN4448_FE_OFN760_n_46337), .d(n_11841), .o(n_46359) );
ao22m06 FE_RC_1354_0 ( .a(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n_24366), .c(n_22089), .d(n_24395), .o(n_24465) );
in01s01 FE_RC_1355_0 ( .a(n_19438), .o(FE_RN_366_0) );
na02m04 FE_RC_1356_0 ( .a(n_19707), .b(n_19505), .o(FE_RN_367_0) );
na02m06 FE_RC_1358_0 ( .a(FE_RN_367_0), .b(FE_OCPN5274_FE_RN_366_0), .o(FE_RN_368_0) );
oa22s01 FE_RC_1361_0 ( .a(n_24350), .b(n_27804), .c(n_27845), .d(FE_OCP_RBN1878_n_27804), .o(n_27862) );
ao22f06 FE_RC_1363_0 ( .a(FE_OCPN3578_n_23354), .b(n_25928), .c(n_23317), .d(FE_OCP_RBN6028_n_25928), .o(n_26039) );
oa22f04 FE_RC_1364_0 ( .a(n_22295), .b(n_22444), .c(n_22296), .d(n_22475), .o(n_22596) );
ao22f02 FE_RC_1366_0 ( .a(n_14741), .b(n_14790), .c(n_14720), .d(n_14791), .o(n_14905) );
oa22f02 FE_RC_1368_0 ( .a(n_14928), .b(n_15055), .c(n_14953), .d(FE_OCP_RBN3014_n_15055), .o(n_15200) );
ao22m04 FE_RC_1369_0 ( .a(n_25395), .b(n_25634), .c(n_25394), .d(n_25655), .o(n_25763) );
oa22m04 FE_RC_1373_0 ( .a(n_20836), .b(n_21091), .c(n_20837), .d(n_21090), .o(n_21236) );
ao22f04 FE_RC_1375_0 ( .a(n_30875), .b(n_30950), .c(n_30876), .d(n_30949), .o(n_31056) );
ao22f04 FE_RC_1379_0 ( .a(n_31802), .b(FE_OCP_RBN5053_n_32169), .c(n_31803), .d(n_32169), .o(n_32254) );
oa22f02 FE_RC_1380_0 ( .a(n_32287), .b(FE_OCP_RBN3432_n_32239), .c(FE_OFN621_n_28336), .d(n_32239), .o(n_32288) );
in01s02 FE_RC_1381_0 ( .a(n_31821), .o(FE_RN_369_0) );
na02m02 TIMEBOOST_cell_5624 ( .a(n_26664), .b(FE_OCP_DRV_N6899_FE_OCPN5276_n_23590), .o(TIMEBOOST_net_1760) );
in01s04 FE_RC_1383_0 ( .a(FE_RN_371_0), .o(n_32172) );
oa22m06 FE_RC_1385_0 ( .a(n_31829), .b(n_32244), .c(n_31830), .d(n_32226), .o(n_32340) );
oa22m04 FE_RC_1387_0 ( .a(FE_OFN747_n_22641), .b(n_25890), .c(n_23259), .d(n_25891), .o(n_25983) );
in01s01 FE_RC_1388_0 ( .a(n_31738), .o(FE_RN_372_0) );
no02f04 TIMEBOOST_cell_6703 ( .a(n_14955), .b(FE_OCP_RBN6695_n_13796), .o(TIMEBOOST_net_2109) );
ao22m04 FE_RC_138_0 ( .a(n_19477), .b(n_18670), .c(n_19476), .d(n_18669), .o(n_19599) );
in01s02 FE_RC_1390_0 ( .a(FE_RN_374_0), .o(n_32224) );
no02m08 TIMEBOOST_cell_8583 ( .a(TIMEBOOST_net_2778), .b(TIMEBOOST_net_881), .o(n_35154) );
oa22s02 FE_RC_1394_0 ( .a(n_27675), .b(n_27526), .c(n_27525), .d(n_27697), .o(n_27785) );
oa22s02 FE_RC_1399_0 ( .a(n_17336), .b(n_17834), .c(n_17753), .d(n_17803), .o(n_17878) );
oa22m04 FE_RC_139_0 ( .a(n_18630), .b(n_19539), .c(n_18629), .d(n_19519), .o(n_19663) );
ao22f04 FE_RC_1402_0 ( .a(n_30640), .b(FE_OCP_RBN5336_n_30865), .c(n_30621), .d(n_30865), .o(n_31046) );
oa22m02 FE_RC_1403_0 ( .a(FE_OCP_RBN3061_n_30575), .b(FE_OFN1196_n_27014), .c(FE_OCPN1677_n_27062), .d(n_30575), .o(n_30692) );
oa22f02 FE_RC_1404_0 ( .a(n_26068), .b(n_26061), .c(n_26028), .d(n_26062), .o(n_26184) );
oa22m02 FE_RC_1406_0 ( .a(n_22907), .b(n_22806), .c(n_20252), .d(n_22776), .o(n_22872) );
in01s01 FE_RC_1407_0 ( .a(n_32052), .o(FE_RN_375_0) );
oa22m06 FE_RC_140_0 ( .a(n_17881), .b(n_19342), .c(n_19418), .d(n_19372), .o(n_19450) );
oa22f02 FE_RC_1412_0 ( .a(n_22801), .b(n_22818), .c(n_22793), .d(FE_OCP_RBN5350_n_22818), .o(n_22894) );
no02s01 FE_RC_1421_0 ( .a(n_17360), .b(n_17359), .o(FE_RN_382_0) );
na02s06 FE_RC_1422_0 ( .a(n_17499), .b(FE_RN_382_0), .o(FE_RN_383_0) );
no02f08 FE_RC_1423_0 ( .a(n_17863), .b(FE_RN_383_0), .o(n_17939) );
na02s01 FE_RC_1427_0 ( .a(n_42358), .b(n_42562), .o(FE_RN_386_0) );
na02s01 FE_RC_1428_0 ( .a(FE_RN_386_0), .b(n_42285), .o(FE_RN_387_0) );
na02f08 FE_RC_1429_0 ( .a(FE_RN_387_0), .b(n_42600), .o(n_42652) );
na02s03 FE_RC_1430_0 ( .a(n_42332), .b(n_42402), .o(FE_RN_388_0) );
no02f08 FE_RC_1431_0 ( .a(FE_RN_388_0), .b(n_42652), .o(n_42705) );
no02s02 FE_RC_1432_0 ( .a(n_35740), .b(n_35739), .o(FE_RN_389_0) );
na02m08 FE_RC_1433_0 ( .a(n_36280), .b(FE_RN_389_0), .o(n_36352) );
na02f04 FE_RC_1436_0 ( .a(n_10111), .b(n_10107), .o(FE_RN_391_0) );
no02m04 FE_RC_1437_0 ( .a(n_10092), .b(n_10050), .o(FE_RN_392_0) );
na02f06 FE_RC_1438_0 ( .a(FE_RN_391_0), .b(FE_RN_392_0), .o(n_10355) );
na02m03 FE_RC_1441_0 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_1_), .b(FE_OCP_RBN5434_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_RN_394_0) );
na02s06 FE_RC_1442_0 ( .a(FE_RN_394_0), .b(n_6619), .o(n_6637) );
in01s02 FE_RC_1443_0 ( .a(delay_xor_ln23_unr3_stage2_stallmux_q), .o(FE_RN_395_0) );
na03f06 TIMEBOOST_cell_8390 ( .a(FE_OCP_RBN6059_n_15795), .b(n_15758), .c(n_15850), .o(n_16071) );
no02s06 TIMEBOOST_cell_5016 ( .a(n_18323), .b(FE_OCP_RBN5031_n_18951), .o(TIMEBOOST_net_1456) );
no02m06 TIMEBOOST_cell_4944 ( .a(FE_RN_130_0), .b(FE_RN_129_0), .o(TIMEBOOST_net_1420) );
no03s02 TIMEBOOST_cell_8227 ( .a(FE_RN_1550_0), .b(FE_OCP_RBN6555_n_28458), .c(FE_RN_1553_0), .o(TIMEBOOST_net_1452) );
in01s01 FE_RC_1448_0 ( .a(n_1494), .o(FE_RN_398_0) );
in01s01 FE_RC_1449_0 ( .a(n_1491), .o(FE_RN_399_0) );
in01s01 FE_RC_1451_0 ( .a(n_12275), .o(FE_RN_400_0) );
in01m04 FE_RC_1452_0 ( .a(n_12294), .o(FE_RN_401_0) );
in01m06 FE_RC_1453_0 ( .a(n_12309), .o(FE_RN_402_0) );
no02m08 FE_RC_1454_0 ( .a(FE_RN_401_0), .b(FE_RN_402_0), .o(FE_RN_403_0) );
na02m04 TIMEBOOST_cell_8799 ( .a(TIMEBOOST_net_2886), .b(n_24783), .o(n_24868) );
na02f04 TIMEBOOST_cell_8794 ( .a(n_24231), .b(n_24319), .o(TIMEBOOST_net_2884) );
na02m08 FE_RC_1457_0 ( .a(FE_RN_400_0), .b(FE_RN_405_0), .o(n_44426) );
na02m08 TIMEBOOST_cell_8841 ( .a(TIMEBOOST_net_2907), .b(n_10782), .o(n_10922) );
no02f02 TIMEBOOST_cell_3969 ( .a(n_19377), .b(FE_OFN738_n_17093), .o(TIMEBOOST_net_1075) );
ao22f02 FE_RC_1479_0 ( .a(n_45319), .b(n_5106), .c(FE_OCP_RBN6821_n_45319), .d(n_5105), .o(n_5284) );
no02f08 FE_RC_1480_0 ( .a(n_23613), .b(n_23580), .o(FE_RN_424_0) );
na02s01 TIMEBOOST_cell_6753 ( .a(n_39144), .b(n_39260), .o(TIMEBOOST_net_2134) );
na02f08 FE_RC_1482_0 ( .a(n_23586), .b(n_23584), .o(FE_RN_426_0) );
na02m80 TIMEBOOST_cell_2791 ( .a(TIMEBOOST_net_686), .b(n_32687), .o(n_32754) );
no02s01 TIMEBOOST_cell_2792 ( .a(n_6512), .b(FE_OCP_RBN5504_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(TIMEBOOST_net_687) );
na02m10 FE_RC_1486_0 ( .a(n_33331), .b(FE_RN_428_0), .o(n_33388) );
in01s06 FE_RC_1487_0 ( .a(n_17897), .o(FE_RN_429_0) );
na02s06 FE_RC_1488_0 ( .a(FE_RN_429_0), .b(n_17954), .o(FE_RN_430_0) );
oa12s06 FE_RC_1490_0 ( .a(FE_RN_430_0), .b(FE_RN_429_0), .c(n_17954), .o(n_18056) );
na02s01 TIMEBOOST_cell_5170 ( .a(n_44102), .b(FE_OCP_RBN1812_n_33750), .o(TIMEBOOST_net_1533) );
no03m10 TIMEBOOST_cell_6430 ( .a(n_37596), .b(TIMEBOOST_net_1442), .c(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37702) );
in01s01 FE_RC_14_0 ( .a(n_18018), .o(FE_RN_6_0) );
in01f04 FE_RC_1502_0 ( .a(n_19501), .o(FE_RN_437_0) );
in01f04 FE_RC_1503_0 ( .a(n_19556), .o(FE_RN_438_0) );
na02f08 FE_RC_1504_0 ( .a(FE_RN_437_0), .b(FE_RN_438_0), .o(FE_RN_439_0) );
in01f06 FE_RC_1505_0 ( .a(FE_RN_440_0), .o(n_19860) );
no02f08 FE_RC_1506_0 ( .a(n_19726), .b(FE_RN_439_0), .o(FE_RN_440_0) );
oa22m04 FE_RC_150_0 ( .a(n_20673), .b(FE_OCP_RBN6017_n_20945), .c(n_20945), .d(n_20672), .o(n_21087) );
in01s01 FE_RC_1510_0 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_), .o(FE_RN_443_0) );
no02s06 FE_RC_1511_0 ( .a(n_32525), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .o(FE_RN_444_0) );
no02m06 FE_RC_1519_0 ( .a(n_12619), .b(n_13270), .o(FE_RN_448_0) );
no02f08 FE_RC_1520_0 ( .a(FE_RN_448_0), .b(n_12620), .o(n_13413) );
na02s01 FE_RC_1521_0 ( .a(n_27416), .b(n_25781), .o(FE_RN_449_0) );
na02s06 FE_RC_1522_0 ( .a(FE_RN_449_0), .b(n_27110), .o(FE_RN_450_0) );
na02f08 FE_RC_1523_0 ( .a(n_27404), .b(FE_RN_450_0), .o(n_27476) );
na02s02 FE_RC_1528_0 ( .a(n_28652), .b(n_28533), .o(FE_RN_453_0) );
no02f04 FE_RC_1529_0 ( .a(n_28976), .b(FE_RN_453_0), .o(n_28997) );
in01s01 FE_RC_1533_0 ( .a(n_23714), .o(FE_RN_456_0) );
no02s04 FE_RC_1534_0 ( .a(FE_RN_456_0), .b(n_24139), .o(FE_RN_457_0) );
in01m04 FE_RC_1537_0 ( .a(n_45327), .o(FE_RN_459_0) );
in01m04 FE_RC_1538_0 ( .a(n_35237), .o(FE_RN_460_0) );
oa22f06 FE_RC_1539_0 ( .a(FE_RN_460_0), .b(FE_RN_459_0), .c(n_35237), .d(n_45327), .o(n_35368) );
na02s02 FE_RC_1541_0 ( .a(n_12836), .b(FE_RN_464_0), .o(FE_RN_462_0) );
no02s10 TIMEBOOST_cell_8825 ( .a(TIMEBOOST_net_2899), .b(FE_OCP_RBN6072_n_16086), .o(n_16330) );
in01s01 FE_RC_1543_0 ( .a(n_12766), .o(FE_RN_464_0) );
in01s02 FE_RC_1546_0 ( .a(n_17339), .o(FE_RN_466_0) );
na02s08 FE_RC_1547_0 ( .a(FE_RN_466_0), .b(n_17401), .o(n_17582) );
na03s06 TIMEBOOST_cell_6454 ( .a(n_2492), .b(n_2520), .c(FE_OCP_RBN5625_n_2457), .o(n_2559) );
in01s01 FE_RC_1550_0 ( .a(n_28628), .o(FE_RN_469_0) );
na02s04 FE_RC_1553_0 ( .a(n_13913), .b(FE_OCP_RBN2056_n_13784), .o(FE_RN_471_0) );
oa22f02 FE_RC_1555_0 ( .a(n_12899), .b(n_13694), .c(n_12898), .d(FE_OCP_RBN2050_n_13694), .o(n_13756) );
na02s06 FE_RC_1560_0 ( .a(n_14510), .b(n_14508), .o(FE_RN_474_0) );
na02m08 FE_RC_1563_0 ( .a(n_14587), .b(FE_RN_476_0), .o(n_14673) );
no02f08 FE_RC_1566_0 ( .a(FE_OCP_RBN2074_n_29603), .b(FE_OCP_RBN6653_n_29494), .o(FE_RN_479_0) );
no02f08 FE_RC_1567_0 ( .a(FE_RN_479_0), .b(n_29586), .o(n_29663) );
no02f08 TIMEBOOST_cell_3247 ( .a(TIMEBOOST_net_914), .b(n_15917), .o(n_16122) );
in01s01 FE_RC_1570_0 ( .a(FE_OCP_RBN5039_n_13927), .o(FE_RN_480_0) );
na02f02 FE_RC_1571_0 ( .a(n_14201), .b(FE_RN_480_0), .o(FE_RN_481_0) );
na02f06 FE_RC_1573_0 ( .a(n_24553), .b(n_24556), .o(FE_RN_482_0) );
na02f08 FE_RC_1574_0 ( .a(FE_RN_482_0), .b(n_24592), .o(n_24779) );
in01s08 FE_RC_1578_0 ( .a(n_16984), .o(FE_RN_485_0) );
no02s10 FE_RC_1579_0 ( .a(n_16936), .b(n_16893), .o(FE_RN_486_0) );
in01f04 FE_RC_158_0 ( .a(FE_RN_35_0), .o(n_21195) );
in01s03 FE_RC_1595_0 ( .a(n_27057), .o(FE_RN_495_0) );
no02f06 FE_RC_1596_0 ( .a(n_27073), .b(n_27024), .o(FE_RN_496_0) );
na02f06 FE_RC_1597_0 ( .a(n_27057), .b(n_27068), .o(FE_RN_497_0) );
no02s02 FE_RC_1599_0 ( .a(n_18758), .b(n_18264), .o(n_18864) );
no02s02 TIMEBOOST_cell_3248 ( .a(n_45072), .b(n_21218), .o(TIMEBOOST_net_915) );
in01s02 FE_RC_15_0 ( .a(n_18020), .o(FE_RN_7_0) );
na02s02 FE_RC_1611_0 ( .a(n_18864), .b(n_18336), .o(n_18947) );
no02s02 FE_RC_1618_0 ( .a(n_23848), .b(n_24251), .o(FE_RN_510_0) );
no02s10 FE_RC_1621_0 ( .a(FE_OCP_RBN6216_n_27086), .b(FE_OCP_RBN5204_n_25729), .o(n_27150) );
no02s01 FE_RC_1627_0 ( .a(n_18461), .b(n_18462), .o(FE_RN_516_0) );
na02s06 FE_RC_1628_0 ( .a(FE_RN_516_0), .b(n_19284), .o(n_19333) );
no02m04 FE_RC_1629_0 ( .a(n_17732), .b(n_18986), .o(FE_RN_517_0) );
no02f08 FE_RC_1630_0 ( .a(n_19112), .b(FE_RN_517_0), .o(n_19213) );
na02s02 FE_RC_1633_0 ( .a(FE_RN_519_0), .b(n_18947), .o(n_19055) );
in01s01 FE_RC_1643_0 ( .a(n_30145), .o(FE_RN_525_0) );
no02f06 FE_RC_1646_0 ( .a(n_26186), .b(n_26293), .o(FE_RN_526_0) );
no02f08 FE_RC_1647_0 ( .a(FE_RN_526_0), .b(n_26212), .o(n_26425) );
in01s01 FE_RC_1648_0 ( .a(n_20124), .o(FE_RN_527_0) );
na02m04 TIMEBOOST_cell_2002 ( .a(n_33610), .b(TIMEBOOST_net_615), .o(n_33636) );
in01s01 FE_RC_1650_0 ( .a(n_19497), .o(FE_RN_529_0) );
in01s02 FE_RC_1651_0 ( .a(n_19653), .o(FE_RN_530_0) );
no02f08 TIMEBOOST_cell_3900 ( .a(n_23826), .b(TIMEBOOST_net_1040), .o(n_24000) );
no02s04 TIMEBOOST_cell_3901 ( .a(n_18893), .b(n_17783), .o(TIMEBOOST_net_1041) );
na02s08 FE_RC_1654_0 ( .a(FE_RN_528_0), .b(FE_RN_532_0), .o(n_20167) );
na02f04 FE_RC_1657_0 ( .a(n_19774), .b(n_19704), .o(FE_RN_533_0) );
no02f04 FE_RC_1659_0 ( .a(FE_OCP_RBN1151_FE_RN_533_0), .b(n_19695), .o(n_19890) );
oa22f04 FE_RC_1660_0 ( .a(n_22508), .b(n_22511), .c(n_22531), .d(n_22469), .o(n_22631) );
in01s02 FE_RC_1661_0 ( .a(n_31103), .o(FE_RN_535_0) );
na02m06 FE_RC_1662_0 ( .a(n_31246), .b(FE_RN_535_0), .o(FE_RN_536_0) );
in01s02 FE_RC_1663_0 ( .a(n_31103), .o(FE_RN_537_0) );
oa12m06 FE_RC_1664_0 ( .a(FE_RN_536_0), .b(n_31246), .c(FE_RN_537_0), .o(n_31404) );
in01m02 FE_RC_1665_0 ( .a(n_31305), .o(FE_RN_538_0) );
in01s02 FE_RC_1666_0 ( .a(n_31156), .o(FE_RN_539_0) );
na02m02 FE_RC_1669_0 ( .a(n_19325), .b(FE_OCP_RBN1133_n_19077), .o(FE_RN_541_0) );
na02f06 FE_RC_1679_0 ( .a(n_19318), .b(n_19152), .o(FE_RN_546_0) );
na02f08 FE_RC_1680_0 ( .a(FE_RN_546_0), .b(n_19348), .o(n_19514) );
na02m06 FE_RC_1681_0 ( .a(n_26069), .b(n_25624), .o(FE_RN_547_0) );
na02f06 FE_RC_1682_0 ( .a(FE_RN_547_0), .b(n_25625), .o(n_26153) );
in01m01 FE_RC_1689_0 ( .a(n_25457), .o(FE_RN_552_0) );
na02m02 FE_RC_1690_0 ( .a(n_25383), .b(FE_RN_552_0), .o(FE_RN_553_0) );
no02m04 FE_RC_1691_0 ( .a(n_25726), .b(FE_RN_553_0), .o(n_25753) );
in01f06 FE_RC_1693_0 ( .a(FE_RN_555_0), .o(n_26963) );
no02f04 FE_RC_1697_0 ( .a(n_25920), .b(FE_RN_1106_0), .o(FE_RN_557_0) );
no02s01 TIMEBOOST_cell_6802 ( .a(TIMEBOOST_net_2158), .b(n_6304), .o(TIMEBOOST_net_921) );
no03m04 TIMEBOOST_cell_3487 ( .a(n_23047), .b(TIMEBOOST_net_591), .c(n_45311), .o(n_23194) );
no03m20 TIMEBOOST_cell_7122 ( .a(FE_RN_32_0), .b(n_17845), .c(n_17884), .o(n_17914) );
no02f02 FE_RC_1701_0 ( .a(n_20504), .b(n_45101), .o(FE_RN_559_0) );
in01s01 FE_RC_1702_0 ( .a(FE_OCPN869_n_45003), .o(FE_RN_560_0) );
ao12f02 FE_RC_1703_0 ( .a(FE_RN_559_0), .b(FE_RN_560_0), .c(n_20504), .o(n_20727) );
ao22m04 FE_RC_1706_0 ( .a(n_31842), .b(n_32150), .c(n_31843), .d(n_32145), .o(n_32239) );
in01s01 FE_RC_1711_0 ( .a(n_20289), .o(FE_RN_563_0) );
na02s03 FE_RC_1712_0 ( .a(FE_RN_563_0), .b(FE_OCP_RBN3001_n_20400), .o(FE_RN_564_0) );
in01s01 FE_RC_1713_0 ( .a(n_20305), .o(FE_RN_565_0) );
no02f06 FE_RC_1714_0 ( .a(n_20616), .b(FE_RN_565_0), .o(FE_RN_566_0) );
na02s02 FE_RC_1715_0 ( .a(n_47257), .b(n_20305), .o(FE_RN_567_0) );
na02m02 FE_RC_1716_0 ( .a(n_20400), .b(FE_RN_567_0), .o(FE_RN_568_0) );
oa12f04 FE_RC_1717_0 ( .a(FE_RN_564_0), .b(FE_RN_566_0), .c(FE_RN_568_0), .o(FE_RN_569_0) );
in01s01 FE_RC_1718_0 ( .a(n_47257), .o(FE_RN_570_0) );
na02s02 TIMEBOOST_cell_5424 ( .a(FE_OCP_RBN3215_n_5003), .b(FE_OCP_RBN2962_n_4046), .o(TIMEBOOST_net_1660) );
na02f04 FE_RC_1721_0 ( .a(FE_RN_569_0), .b(FE_RN_572_0), .o(n_20848) );
in01s02 FE_RC_1724_0 ( .a(n_20570), .o(FE_RN_574_0) );
no02s01 TIMEBOOST_cell_4878 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_30_), .o(TIMEBOOST_net_1387) );
na02s02 FE_RC_1731_0 ( .a(n_45091), .b(n_21118), .o(FE_RN_579_0) );
no02s01 TIMEBOOST_cell_4498 ( .a(TIMEBOOST_net_1339), .b(n_27110), .o(n_27226) );
no02s01 TIMEBOOST_cell_4499 ( .a(FE_OCP_RBN3386_n_11439), .b(n_10613), .o(TIMEBOOST_net_1340) );
in01f02 FE_RC_173_0 ( .a(n_20963), .o(FE_RN_42_0) );
no02s04 FE_RC_1744_0 ( .a(n_30619), .b(FE_OCPN1676_n_27062), .o(FE_RN_588_0) );
in01s01 FE_RC_1749_0 ( .a(n_45023), .o(FE_RN_591_0) );
in01m02 FE_RC_174_0 ( .a(n_20991), .o(FE_RN_43_0) );
na02m02 FE_RC_1751_0 ( .a(FE_RN_591_0), .b(n_21084), .o(FE_RN_592_0) );
na02s06 FE_RC_1755_0 ( .a(n_30824), .b(FE_OCPN5286_n_30708), .o(FE_RN_595_0) );
na02m08 FE_RC_1756_0 ( .a(n_31018), .b(FE_RN_595_0), .o(n_31079) );
na02s02 TIMEBOOST_cell_5400 ( .a(n_42856), .b(n_43103), .o(TIMEBOOST_net_1648) );
no02m06 TIMEBOOST_cell_7719 ( .a(TIMEBOOST_net_2490), .b(FE_OCP_RBN2929_n_34971), .o(n_35075) );
na02f06 TIMEBOOST_cell_5403 ( .a(TIMEBOOST_net_1649), .b(n_43193), .o(n_43334) );
no02s06 TIMEBOOST_cell_8518 ( .a(n_13260), .b(n_13778), .o(TIMEBOOST_net_2746) );
na02m10 FE_RC_1771_0 ( .a(FE_RN_604_0), .b(n_31971), .o(n_32026) );
no02s04 FE_RC_1774_0 ( .a(n_21540), .b(FE_OCP_RBN1170_n_21318), .o(n_21573) );
no02m04 FE_RC_1776_0 ( .a(n_22066), .b(FE_OCP_RBN4645_n_20420), .o(FE_RN_606_0) );
oa22s01 FE_RC_1781_0 ( .a(n_24350), .b(n_27805), .c(n_27796), .d(n_45132), .o(n_27863) );
na02s02 TIMEBOOST_cell_8664 ( .a(n_40028), .b(FE_OCP_RBN4431_n_39942), .o(TIMEBOOST_net_2819) );
in01s01 FE_RC_1783_0 ( .a(n_27470), .o(FE_RN_611_0) );
in01s01 FE_RC_1784_0 ( .a(FE_RN_612_0), .o(n_27531) );
na03m02 TIMEBOOST_cell_8430 ( .a(FE_OCP_RBN4440_n_5891), .b(n_47270), .c(FE_OCP_RBN4444_n_5849), .o(TIMEBOOST_net_564) );
na02s04 FE_RC_1788_0 ( .a(n_31463), .b(n_31234), .o(FE_RN_614_0) );
in01s01 FE_RC_1793_0 ( .a(FE_OCPN5113_n_22249), .o(FE_RN_617_0) );
in01s01 FE_RC_1794_0 ( .a(FE_OCP_RBN3259_n_21360), .o(FE_RN_618_0) );
na02s02 FE_RC_1796_0 ( .a(FE_RN_618_0), .b(FE_OCP_RBN4484_n_22667), .o(FE_RN_620_0) );
na02s02 FE_RC_1797_0 ( .a(FE_RN_617_0), .b(FE_RN_620_0), .o(FE_RN_621_0) );
na02s02 FE_RC_1798_0 ( .a(n_22470), .b(FE_RN_621_0), .o(FE_RN_622_0) );
no02s06 TIMEBOOST_cell_8722 ( .a(n_37417), .b(n_37151), .o(TIMEBOOST_net_2848) );
in01s01 FE_RC_1800_0 ( .a(n_22413), .o(FE_RN_624_0) );
na02s02 FE_RC_1801_0 ( .a(FE_OCP_RBN4487_n_22438), .b(FE_RN_624_0), .o(FE_RN_625_0) );
no02s02 FE_RC_1805_0 ( .a(n_22233), .b(n_22235), .o(FE_RN_628_0) );
in01s01 FE_RC_1806_0 ( .a(n_22273), .o(FE_RN_629_0) );
na02m06 FE_RC_1807_0 ( .a(n_45498), .b(FE_RN_629_0), .o(FE_RN_630_0) );
na02m08 FE_RC_1808_0 ( .a(FE_RN_630_0), .b(FE_RN_628_0), .o(n_22720) );
ao22f04 FE_RC_180_0 ( .a(n_22502), .b(FE_OCP_RBN5345_n_22476), .c(FE_OCP_RBN1173_n_22476), .d(n_22503), .o(n_22622) );
in01s06 FE_RC_1810_0 ( .a(n_37205), .o(FE_RN_631_0) );
na02s08 FE_RC_1811_0 ( .a(FE_RN_631_0), .b(n_37157), .o(FE_RN_632_0) );
no02m08 FE_RC_1812_0 ( .a(n_37092), .b(FE_RN_632_0), .o(FE_RN_633_0) );
in01s06 FE_RC_1813_0 ( .a(n_37279), .o(FE_RN_634_0) );
no02s06 FE_RC_1814_0 ( .a(FE_RN_634_0), .b(n_37034), .o(FE_RN_635_0) );
no02m01 TIMEBOOST_cell_8060 ( .a(FE_OCP_RBN3333_n_39942), .b(FE_OCP_RBN6824_n_39542), .o(TIMEBOOST_net_2661) );
in01m01 FE_RC_1816_0 ( .a(n_37161), .o(FE_RN_637_0) );
no02s06 TIMEBOOST_cell_1625 ( .a(n_19148), .b(n_17881), .o(TIMEBOOST_net_427) );
no02m06 TIMEBOOST_cell_5061 ( .a(TIMEBOOST_net_1478), .b(FE_OCP_RBN5677_n_19177), .o(n_19360) );
in01m08 FE_RC_1819_0 ( .a(n_37253), .o(FE_RN_640_0) );
no02m10 FE_RC_1820_0 ( .a(FE_RN_640_0), .b(FE_RN_639_0), .o(FE_RN_641_0) );
na02f10 FE_RC_1821_0 ( .a(FE_RN_641_0), .b(FE_RN_636_0), .o(n_37353) );
in01s20 FE_RC_1824_0 ( .a(n_22944), .o(FE_RN_643_0) );
no02s20 FE_RC_1825_0 ( .a(FE_RN_643_0), .b(n_22823), .o(FE_RN_644_0) );
no02s06 FE_RC_1827_0 ( .a(n_32949), .b(n_32914), .o(FE_RN_645_0) );
na02s06 FE_RC_1828_0 ( .a(FE_RN_645_0), .b(n_33274), .o(FE_RN_646_0) );
no02s01 TIMEBOOST_cell_3213 ( .a(TIMEBOOST_net_897), .b(n_5994), .o(n_6051) );
na02s02 TIMEBOOST_cell_3214 ( .a(FE_RN_570_0), .b(FE_OCP_RBN3002_n_20400), .o(TIMEBOOST_net_898) );
na02f04 TIMEBOOST_cell_8812 ( .a(n_14764), .b(FE_OCP_RBN5776_n_13796), .o(TIMEBOOST_net_2893) );
no03s06 TIMEBOOST_cell_7176 ( .a(n_2461), .b(n_2475), .c(FE_OCP_RBN5605_n_2430), .o(n_2517) );
no03s08 FE_RC_1833_0 ( .a(n_33159), .b(n_33380), .c(n_33160), .o(FE_RN_650_0) );
no02s01 TIMEBOOST_cell_1783 ( .a(n_15806), .b(n_15293), .o(TIMEBOOST_net_506) );
no02s04 TIMEBOOST_cell_1784 ( .a(TIMEBOOST_net_506), .b(n_15808), .o(n_15906) );
no02s06 FE_RC_1842_0 ( .a(n_33083), .b(FE_RN_656_0), .o(FE_RN_657_0) );
no02s06 FE_RC_1843_0 ( .a(n_42260), .b(n_42288), .o(FE_RN_658_0) );
na02f08 FE_RC_1844_0 ( .a(FE_RN_658_0), .b(n_42541), .o(n_42554) );
no02s01 FE_RC_1845_0 ( .a(n_22695), .b(n_22692), .o(FE_RN_659_0) );
na02s02 FE_RC_1846_0 ( .a(n_22763), .b(FE_RN_659_0), .o(FE_RN_660_0) );
no02m06 FE_RC_1847_0 ( .a(n_23221), .b(FE_RN_660_0), .o(n_23242) );
ao22s04 FE_RC_184_0 ( .a(n_22505), .b(n_22589), .c(n_22504), .d(FE_OCP_RBN4647_n_22553), .o(n_22739) );
in01s01 FE_RC_1851_0 ( .a(FE_OCPN873_n_42202), .o(FE_RN_663_0) );
in01s01 FE_RC_1852_0 ( .a(n_42304), .o(FE_RN_664_0) );
in01s01 FE_RC_1853_0 ( .a(n_42327), .o(FE_RN_665_0) );
no02f10 TIMEBOOST_cell_3027 ( .a(n_8733), .b(TIMEBOOST_net_804), .o(n_8875) );
in01s01 TIMEBOOST_cell_5919 ( .a(FE_OFN1_n_43918), .o(TIMEBOOST_net_1808) );
no02f08 TIMEBOOST_cell_6066 ( .a(TIMEBOOST_net_1884), .b(n_12977), .o(n_13011) );
na02m04 FE_RC_1857_0 ( .a(FE_RN_668_0), .b(n_42428), .o(FE_RN_669_0) );
na03s02 FE_RC_1858_0 ( .a(n_42359), .b(n_42328), .c(n_42360), .o(FE_RN_670_0) );
na02f08 TIMEBOOST_cell_853 ( .a(FE_RN_173_0), .b(n_37175), .o(TIMEBOOST_net_41) );
na02f08 TIMEBOOST_cell_854 ( .a(TIMEBOOST_net_41), .b(n_37033), .o(n_37193) );
in01s01 FE_RC_1861_0 ( .a(n_42285), .o(FE_RN_672_0) );
in01s01 FE_RC_1862_0 ( .a(n_42423), .o(FE_RN_673_0) );
in01s01 FE_RC_1863_0 ( .a(n_42443), .o(FE_RN_674_0) );
no02f06 TIMEBOOST_cell_2961 ( .a(TIMEBOOST_net_771), .b(n_24598), .o(n_24720) );
no02m02 TIMEBOOST_cell_2962 ( .a(FE_OCP_RBN1829_n_19528), .b(FE_OCPN1665_FE_OCP_RBN1138_n_19270), .o(TIMEBOOST_net_772) );
na02s02 FE_RC_1866_0 ( .a(FE_RN_676_0), .b(n_42434), .o(FE_RN_677_0) );
na03s02 FE_RC_1867_0 ( .a(n_42397), .b(n_42451), .c(n_42395), .o(FE_RN_678_0) );
na02m06 TIMEBOOST_cell_6776 ( .a(TIMEBOOST_net_2145), .b(n_9457), .o(n_9623) );
na02f02 TIMEBOOST_cell_6010 ( .a(n_41155), .b(TIMEBOOST_net_1856), .o(n_41233) );
in01m04 FE_RC_1872_0 ( .a(FE_RN_681_0), .o(n_44996) );
no02m04 FE_RC_1873_0 ( .a(n_23494), .b(n_23053), .o(FE_RN_681_0) );
in01s01 FE_RC_1874_0 ( .a(n_17308), .o(FE_RN_682_0) );
in01f04 FE_RC_1875_0 ( .a(FE_RN_683_0), .o(n_18104) );
na02f06 FE_RC_1876_0 ( .a(n_18013), .b(FE_RN_682_0), .o(FE_RN_683_0) );
no03m02 TIMEBOOST_cell_8321 ( .a(TIMEBOOST_net_1583), .b(n_9261), .c(FE_OCP_RBN6720_FE_OCP_DRV_N6264_n_9014), .o(TIMEBOOST_net_2507) );
na02s04 FE_RC_1881_0 ( .a(FE_RN_686_0), .b(n_42492), .o(FE_RN_687_0) );
no02f08 FE_RC_1882_0 ( .a(FE_RN_687_0), .b(n_42790), .o(n_42834) );
in01s01 FE_RC_1883_0 ( .a(n_25053), .o(FE_RN_688_0) );
na02s01 FE_RC_1884_0 ( .a(FE_RN_688_0), .b(n_25548), .o(FE_RN_689_0) );
no02f04 FE_RC_1885_0 ( .a(FE_RN_689_0), .b(n_25470), .o(n_25528) );
in01s04 FE_RC_1886_0 ( .a(n_17665), .o(FE_RN_690_0) );
na02m08 TIMEBOOST_cell_7704 ( .a(n_22089), .b(FE_OCP_RBN5721_n_24506), .o(TIMEBOOST_net_2483) );
no02s08 FE_RC_1889_0 ( .a(FE_RN_692_0), .b(n_17734), .o(FE_RN_693_0) );
in01s02 FE_RC_1890_0 ( .a(n_17611), .o(FE_RN_694_0) );
no02s06 FE_RC_1891_0 ( .a(FE_RN_694_0), .b(n_17663), .o(FE_RN_695_0) );
na02f08 FE_RC_1892_0 ( .a(n_45524), .b(FE_RN_695_0), .o(FE_RN_696_0) );
na02f10 FE_RC_1893_0 ( .a(FE_RN_696_0), .b(FE_RN_693_0), .o(n_18421) );
in01s01 FE_RC_1894_0 ( .a(n_25189), .o(FE_RN_697_0) );
no02s06 TIMEBOOST_cell_6777 ( .a(n_24310), .b(n_24386), .o(TIMEBOOST_net_2146) );
in01s01 FE_RC_1896_0 ( .a(n_25160), .o(FE_RN_699_0) );
na03m08 TIMEBOOST_cell_2214 ( .a(n_40790), .b(n_40702), .c(n_45149), .o(n_40795) );
no02f06 TIMEBOOST_cell_7681 ( .a(TIMEBOOST_net_2471), .b(TIMEBOOST_net_1467), .o(n_37944) );
na02s06 TIMEBOOST_cell_8665 ( .a(TIMEBOOST_net_2819), .b(n_40030), .o(n_40134) );
oa22m04 FE_RC_18_0 ( .a(n_18333), .b(n_18520), .c(n_18519), .d(n_18334), .o(n_18682) );
no02s06 TIMEBOOST_cell_5603 ( .a(TIMEBOOST_net_1749), .b(FE_OCP_RBN3369_n_31520), .o(n_31831) );
no03f08 TIMEBOOST_cell_7335 ( .a(n_28291), .b(n_28290), .c(FE_RN_127_0), .o(FE_RN_128_0) );
na02s08 FE_RC_1902_0 ( .a(n_34380), .b(n_34381), .o(FE_RN_704_0) );
no02m08 FE_RC_1903_0 ( .a(FE_RN_704_0), .b(n_34406), .o(n_34459) );
no02s01 TIMEBOOST_cell_2875 ( .a(TIMEBOOST_net_728), .b(n_37858), .o(n_38022) );
na02m02 TIMEBOOST_cell_2876 ( .a(n_37756), .b(n_37700), .o(TIMEBOOST_net_729) );
na02f08 FE_RC_1906_0 ( .a(FE_RN_706_0), .b(n_34342), .o(n_34375) );
no03m08 TIMEBOOST_cell_3533 ( .a(n_37945), .b(FE_RN_952_0), .c(n_37980), .o(FE_RN_954_0) );
ao22f06 FE_RC_1908_0 ( .a(n_41783), .b(n_42038), .c(n_41782), .d(FE_OCP_RBN5699_n_42038), .o(n_42100) );
no02s01 FE_RC_1909_0 ( .a(n_27878), .b(n_27990), .o(FE_RN_707_0) );
na02m04 FE_RC_1910_0 ( .a(n_28138), .b(FE_RN_707_0), .o(n_28205) );
na02s01 FE_RC_1911_0 ( .a(n_1580), .b(n_1441), .o(FE_RN_708_0) );
no02s01 FE_RC_1912_0 ( .a(FE_RN_708_0), .b(n_1630), .o(FE_RN_709_0) );
na02f06 FE_RC_1913_0 ( .a(FE_RN_709_0), .b(n_1869), .o(FE_RN_710_0) );
na02f06 FE_RC_1914_0 ( .a(FE_RN_710_0), .b(n_1442), .o(n_1958) );
no02s06 TIMEBOOST_cell_2966 ( .a(n_41293), .b(FE_OCPN3555_n_40986), .o(TIMEBOOST_net_774) );
in01s01 FE_RC_1931_0 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_), .o(FE_RN_724_0) );
in01s01 FE_RC_1932_0 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_), .o(FE_RN_725_0) );
no02s03 TIMEBOOST_cell_1557 ( .a(n_30098), .b(n_30066), .o(TIMEBOOST_net_393) );
na02s06 TIMEBOOST_cell_2922 ( .a(FE_RN_2399_0), .b(n_12954), .o(TIMEBOOST_net_752) );
no02m04 FE_RC_1935_0 ( .a(n_28401), .b(FE_RN_727_0), .o(n_28399) );
in01s01 FE_RC_1936_0 ( .a(n_28016), .o(FE_RN_728_0) );
no02s01 TIMEBOOST_cell_6681 ( .a(FE_OCP_RBN4143_n_7743), .b(FE_OCP_RBN4138_n_7743), .o(TIMEBOOST_net_2098) );
no02m04 TIMEBOOST_cell_1667 ( .a(n_25932), .b(FE_OFN748_n_22641), .o(TIMEBOOST_net_448) );
na02s04 TIMEBOOST_cell_4339 ( .a(n_7968), .b(n_7832), .o(TIMEBOOST_net_1260) );
no02s01 FE_RC_1940_0 ( .a(n_28050), .b(n_28018), .o(FE_RN_732_0) );
na02s01 TIMEBOOST_cell_4880 ( .a(FE_RN_737_0), .b(FE_RN_738_0), .o(TIMEBOOST_net_1388) );
na02s02 TIMEBOOST_cell_1883 ( .a(n_36091), .b(n_35613), .o(TIMEBOOST_net_556) );
no02s01 FE_RC_1944_0 ( .a(n_28108), .b(n_28109), .o(FE_RN_735_0) );
na02s01 FE_RC_1945_0 ( .a(FE_RN_735_0), .b(n_28154), .o(FE_RN_736_0) );
no02s08 FE_RC_1946_0 ( .a(FE_OCP_RBN2480_FE_RN_734_0), .b(FE_RN_736_0), .o(n_28539) );
in01s01 FE_RC_1947_0 ( .a(n_27923), .o(FE_RN_737_0) );
in01s01 FE_RC_1948_0 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_30_), .o(FE_RN_738_0) );
in01s01 FE_RC_1949_0 ( .a(n_28152), .o(FE_RN_739_0) );
in01s03 FE_RC_194_0 ( .a(n_23391), .o(FE_RN_45_0) );
no02s06 TIMEBOOST_cell_3028 ( .a(n_34427), .b(n_34037), .o(TIMEBOOST_net_805) );
no02s02 TIMEBOOST_cell_1656 ( .a(TIMEBOOST_net_442), .b(n_3612), .o(n_3755) );
na02s06 FE_RC_1952_0 ( .a(n_28261), .b(FE_RN_741_0), .o(FE_RN_742_0) );
in01s01 FE_RC_1953_0 ( .a(n_28214), .o(FE_RN_743_0) );
no02f04 TIMEBOOST_cell_6327 ( .a(n_16434), .b(n_16444), .o(TIMEBOOST_net_2015) );
no02m06 TIMEBOOST_cell_8723 ( .a(TIMEBOOST_net_2848), .b(TIMEBOOST_net_1025), .o(n_37527) );
no03s02 TIMEBOOST_cell_7131 ( .a(n_23606), .b(n_23605), .c(n_23679), .o(n_23714) );
na02s06 TIMEBOOST_cell_8669 ( .a(TIMEBOOST_net_2821), .b(FE_OCP_RBN3169_n_44211), .o(n_35691) );
in01m20 FE_RC_1959_0 ( .a(n_23308), .o(FE_RN_747_0) );
in01s10 FE_RC_195_0 ( .a(n_23390), .o(FE_RN_46_0) );
na02m20 FE_RC_1960_0 ( .a(FE_OCP_RBN5540_n_23307), .b(FE_RN_747_0), .o(FE_RN_748_0) );
in01m20 FE_RC_1963_0 ( .a(n_23015), .o(FE_RN_749_0) );
no02m40 FE_RC_1965_0 ( .a(FE_RN_749_0), .b(n_22889), .o(FE_RN_751_0) );
na02m20 FE_RC_1966_0 ( .a(FE_RN_751_0), .b(n_23040), .o(n_23064) );
in01s01 FE_RC_1967_0 ( .a(n_37913), .o(FE_RN_752_0) );
in01s02 FE_RC_1968_0 ( .a(n_37981), .o(FE_RN_753_0) );
in01s01 FE_RC_1969_0 ( .a(n_37912), .o(FE_RN_754_0) );
na02s10 FE_RC_196_0 ( .a(FE_RN_46_0), .b(FE_RN_45_0), .o(FE_RN_47_0) );
na02s10 TIMEBOOST_cell_8695 ( .a(TIMEBOOST_net_2834), .b(n_32690), .o(n_32732) );
no02s06 TIMEBOOST_cell_8724 ( .a(n_28090), .b(FE_OCP_RBN5549_n_28319), .o(TIMEBOOST_net_2849) );
no03m04 TIMEBOOST_cell_8231 ( .a(n_37605), .b(n_37659), .c(n_37579), .o(n_37717) );
na02s06 TIMEBOOST_cell_1957 ( .a(n_37366), .b(n_37219), .o(TIMEBOOST_net_593) );
na02f06 FE_RC_1975_0 ( .a(FE_RN_759_0), .b(n_38122), .o(FE_RN_760_0) );
no02s04 FE_RC_1976_0 ( .a(n_37939), .b(n_37946), .o(FE_RN_761_0) );
na02m06 FE_RC_1977_0 ( .a(n_37975), .b(FE_RN_761_0), .o(FE_RN_762_0) );
no02s01 TIMEBOOST_cell_3895 ( .a(n_37732), .b(n_37529), .o(TIMEBOOST_net_1038) );
no02s04 TIMEBOOST_cell_3946 ( .a(TIMEBOOST_net_1063), .b(FE_OCP_RBN2800_n_8817), .o(n_8951) );
in01s01 FE_RC_1980_0 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_), .o(FE_RN_764_0) );
in01s01 FE_RC_1981_0 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_), .o(FE_RN_765_0) );
no02s01 TIMEBOOST_cell_1563 ( .a(n_2976), .b(n_4073), .o(TIMEBOOST_net_396) );
no02m04 TIMEBOOST_cell_4265 ( .a(n_33771), .b(n_34037), .o(TIMEBOOST_net_1223) );
no02f08 FE_RC_1984_0 ( .a(FE_RN_767_0), .b(n_12418), .o(n_12413) );
na02s02 FE_RC_1985_0 ( .a(n_6569), .b(n_6540), .o(FE_RN_768_0) );
na02s06 TIMEBOOST_cell_8639 ( .a(TIMEBOOST_net_2806), .b(n_30851), .o(n_30991) );
no02f06 TIMEBOOST_cell_6732 ( .a(TIMEBOOST_net_2123), .b(FE_OCP_RBN2101_n_15083), .o(n_15281) );
na02m20 FE_RC_1989_0 ( .a(FE_RN_770_0), .b(delay_xor_ln21_unr21_stage8_stallmux_q_10_), .o(n_32863) );
no02f04 TIMEBOOST_cell_1708 ( .a(n_20270), .b(TIMEBOOST_net_468), .o(n_20376) );
in01s01 FE_RC_1993_0 ( .a(n_1936), .o(FE_RN_773_0) );
no03m06 TIMEBOOST_cell_8209 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_11_), .b(FE_RN_204_0), .c(n_32879), .o(FE_RN_206_0) );
na02s06 TIMEBOOST_cell_8668 ( .a(TIMEBOOST_net_556), .b(FE_OCP_RBN3168_n_44211), .o(TIMEBOOST_net_2821) );
in01s01 FE_RC_1996_0 ( .a(n_11896), .o(FE_RN_775_0) );
na02s06 FE_RC_1997_0 ( .a(n_12050), .b(FE_RN_775_0), .o(FE_RN_776_0) );
no02f10 FE_RC_1998_0 ( .a(FE_RN_776_0), .b(n_12514), .o(n_12535) );
no02s06 TIMEBOOST_cell_4926 ( .a(n_40681), .b(n_45153), .o(TIMEBOOST_net_1411) );
no02m08 TIMEBOOST_cell_4927 ( .a(n_40914), .b(TIMEBOOST_net_1411), .o(n_40943) );
in01s01 FE_RC_2001_0 ( .a(n_2005), .o(FE_RN_778_0) );
na02s01 TIMEBOOST_cell_6815 ( .a(n_36062), .b(n_36096), .o(TIMEBOOST_net_2165) );
in01m06 FE_RC_2003_0 ( .a(FE_RN_780_0), .o(n_45488) );
no03f04 TIMEBOOST_cell_2764 ( .a(n_39702), .b(n_39685), .c(n_39712), .o(n_39739) );
in01s02 FE_RC_2005_0 ( .a(n_12170), .o(FE_RN_781_0) );
in01s01 FE_RC_2006_0 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_22_), .o(FE_RN_782_0) );
in01s01 FE_RC_2007_0 ( .a(n_11973), .o(FE_RN_783_0) );
no02m10 TIMEBOOST_cell_4895 ( .a(TIMEBOOST_net_1395), .b(FE_OCP_RBN6538_n_1614), .o(n_1672) );
no02m08 TIMEBOOST_cell_1722 ( .a(TIMEBOOST_net_475), .b(n_20441), .o(n_20472) );
in01s01 FE_RC_2010_0 ( .a(n_12051), .o(FE_RN_786_0) );
na02s06 FE_RC_2011_0 ( .a(FE_RN_786_0), .b(FE_RN_785_0), .o(FE_RN_787_0) );
in01s02 FE_RC_2012_0 ( .a(n_12170), .o(FE_RN_788_0) );
ao22f10 FE_RC_2013_0 ( .a(FE_RN_787_0), .b(FE_RN_781_0), .c(FE_RN_788_0), .d(n_12535), .o(n_12623) );
oa22f04 FE_RC_2014_0 ( .a(n_40306), .b(n_40563), .c(FE_OCP_RBN3430_n_40563), .d(n_45306), .o(n_40593) );
no02s06 FE_RC_2015_0 ( .a(n_43435), .b(n_43387), .o(FE_RN_789_0) );
na02s06 FE_RC_2016_0 ( .a(FE_RN_789_0), .b(n_43523), .o(FE_RN_790_0) );
no02m10 FE_RC_2017_0 ( .a(n_43768), .b(FE_RN_790_0), .o(n_43822) );
in01s01 FE_RC_2018_0 ( .a(n_12278), .o(FE_RN_791_0) );
in01s01 FE_RC_2019_0 ( .a(n_12279), .o(FE_RN_792_0) );
na02s02 FE_RC_2020_0 ( .a(FE_RN_791_0), .b(FE_RN_792_0), .o(FE_RN_793_0) );
in01s01 FE_RC_2021_0 ( .a(n_12119), .o(FE_RN_794_0) );
no02s03 FE_RC_2022_0 ( .a(FE_RN_793_0), .b(FE_RN_794_0), .o(FE_RN_795_0) );
in01s01 FE_RC_2023_0 ( .a(FE_OCP_RBN2394_n_45697), .o(FE_RN_796_0) );
in01s01 FE_RC_2024_0 ( .a(n_12168), .o(FE_RN_797_0) );
no02m06 TIMEBOOST_cell_1717 ( .a(FE_OCP_RBN2861_n_44921), .b(n_38973), .o(TIMEBOOST_net_473) );
na03s10 TIMEBOOST_cell_5697 ( .a(n_32578), .b(n_32577), .c(n_32582), .o(n_32625) );
na02m06 TIMEBOOST_cell_5062 ( .a(n_13515), .b(FE_OCP_RBN5757_n_14444), .o(TIMEBOOST_net_1479) );
na02s08 TIMEBOOST_cell_4896 ( .a(n_11867), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_14_), .o(TIMEBOOST_net_1396) );
oa22f02 FE_RC_2040_0 ( .a(n_40598), .b(n_40593), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .d(n_40584), .o(n_40599) );
in01s01 FE_RC_2041_0 ( .a(n_43522), .o(FE_RN_811_0) );
in01s02 FE_RC_2042_0 ( .a(n_43822), .o(FE_RN_812_0) );
no02s06 FE_RC_2043_0 ( .a(FE_RN_811_0), .b(FE_RN_812_0), .o(FE_RN_813_0) );
no02s06 FE_RC_2044_0 ( .a(FE_RN_813_0), .b(n_43681), .o(n_43842) );
in01s01 FE_RC_2047_0 ( .a(n_6940), .o(FE_RN_816_0) );
in01s02 FE_RC_204_0 ( .a(n_23461), .o(FE_RN_51_0) );
na02s06 FE_RC_2050_0 ( .a(n_39980), .b(n_40013), .o(FE_RN_818_0) );
no02f08 FE_RC_2051_0 ( .a(FE_RN_818_0), .b(n_40406), .o(n_40422) );
na02m06 FE_RC_2056_0 ( .a(n_3000), .b(n_2231), .o(FE_RN_821_0) );
na02m08 FE_RC_2057_0 ( .a(FE_RN_821_0), .b(n_2232), .o(n_3092) );
na02s01 TIMEBOOST_cell_5522 ( .a(n_11007), .b(FE_OCP_RBN4483_n_11439), .o(TIMEBOOST_net_1709) );
in01s06 FE_RC_205_0 ( .a(n_23462), .o(FE_RN_52_0) );
no02s02 TIMEBOOST_cell_8827 ( .a(TIMEBOOST_net_2900), .b(n_4692), .o(TIMEBOOST_net_1309) );
in01s01 FE_RC_2061_0 ( .a(n_2149), .o(FE_RN_824_0) );
no02s04 TIMEBOOST_cell_4110 ( .a(TIMEBOOST_net_1145), .b(n_10619), .o(n_10742) );
no02s01 TIMEBOOST_cell_4111 ( .a(FE_OCP_RBN6076_n_44256), .b(n_35005), .o(TIMEBOOST_net_1146) );
no02s02 FE_RC_2065_0 ( .a(n_35616), .b(n_35617), .o(FE_RN_826_0) );
na02s06 FE_RC_2066_0 ( .a(FE_RN_826_0), .b(n_35640), .o(FE_RN_827_0) );
no02f08 FE_RC_2067_0 ( .a(n_36208), .b(FE_RN_827_0), .o(n_36280) );
no02f10 FE_RC_2068_0 ( .a(n_39347), .b(n_39278), .o(FE_RN_828_0) );
na02m10 FE_RC_2069_0 ( .a(n_39254), .b(n_39253), .o(FE_RN_829_0) );
na02m08 FE_RC_206_0 ( .a(FE_RN_51_0), .b(FE_RN_52_0), .o(FE_RN_53_0) );
no02f20 FE_RC_2070_0 ( .a(FE_RN_828_0), .b(FE_RN_829_0), .o(n_39493) );
no02f06 FE_RC_2074_0 ( .a(n_39187), .b(n_39446), .o(FE_RN_832_0) );
ao12f04 FE_RC_2075_0 ( .a(FE_RN_832_0), .b(n_39187), .c(n_39446), .o(n_39542) );
na02m06 FE_RC_2076_0 ( .a(n_1795), .b(n_1667), .o(FE_RN_833_0) );
na02m08 FE_RC_2077_0 ( .a(FE_RN_833_0), .b(n_1666), .o(n_1847) );
no02m08 TIMEBOOST_cell_3884 ( .a(n_28634), .b(TIMEBOOST_net_1032), .o(n_28749) );
na02m02 TIMEBOOST_cell_3885 ( .a(n_18148), .b(n_17948), .o(TIMEBOOST_net_1033) );
in01m08 FE_RC_2080_0 ( .a(FE_RN_835_0), .o(n_45740) );
na02f08 FE_RC_2081_0 ( .a(n_39652), .b(n_39637), .o(FE_RN_835_0) );
in01s01 FE_RC_2084_0 ( .a(n_7095), .o(FE_RN_837_0) );
no02s03 TIMEBOOST_cell_8094 ( .a(n_36553), .b(n_36750), .o(TIMEBOOST_net_2678) );
no02s02 TIMEBOOST_cell_8520 ( .a(TIMEBOOST_net_2215), .b(FE_OCP_RBN4131_n_24077), .o(TIMEBOOST_net_2747) );
in01s01 FE_RC_2087_0 ( .a(n_7132), .o(FE_RN_839_0) );
no03s08 TIMEBOOST_cell_8188 ( .a(FE_OCPN937_n_17684), .b(n_17683), .c(n_17726), .o(n_17727) );
na03s02 TIMEBOOST_cell_7972 ( .a(n_4430), .b(n_4431), .c(n_4144), .o(TIMEBOOST_net_2617) );
no02s02 FE_RC_2090_0 ( .a(n_40130), .b(n_40128), .o(FE_RN_841_0) );
na02f08 FE_RC_2091_0 ( .a(n_40495), .b(FE_RN_841_0), .o(n_40511) );
in01s01 FE_RC_2092_0 ( .a(n_18524), .o(FE_RN_842_0) );
na02s02 FE_RC_2093_0 ( .a(n_18620), .b(FE_RN_842_0), .o(FE_RN_843_0) );
no02s03 FE_RC_2094_0 ( .a(n_18661), .b(FE_RN_843_0), .o(FE_RN_844_0) );
na02m04 FE_RC_2095_0 ( .a(n_18966), .b(n_18612), .o(FE_RN_845_0) );
na02m06 FE_RC_2096_0 ( .a(FE_RN_845_0), .b(FE_RN_844_0), .o(n_19097) );
na02s04 TIMEBOOST_cell_1690 ( .a(TIMEBOOST_net_459), .b(n_20024), .o(FE_RN_528_0) );
na02s01 FE_RC_2098_0 ( .a(n_18658), .b(n_18659), .o(FE_RN_846_0) );
no02s02 FE_RC_2099_0 ( .a(n_18696), .b(FE_RN_846_0), .o(FE_RN_847_0) );
na02m06 FE_RC_2100_0 ( .a(n_19097), .b(FE_RN_847_0), .o(n_19125) );
oa22s02 FE_RC_2101_0 ( .a(n_1496), .b(n_1461), .c(n_1495), .d(n_1460), .o(n_1571) );
na02s01 FE_RC_2104_0 ( .a(n_18810), .b(n_18722), .o(FE_RN_849_0) );
in01m02 FE_RC_2105_0 ( .a(n_18884), .o(FE_RN_850_0) );
no02s04 FE_RC_2106_0 ( .a(FE_RN_850_0), .b(FE_RN_849_0), .o(FE_RN_851_0) );
no02s01 FE_RC_2107_0 ( .a(n_18769), .b(n_18724), .o(FE_RN_852_0) );
no02f08 TIMEBOOST_cell_5145 ( .a(TIMEBOOST_net_1520), .b(n_14616), .o(n_14721) );
no02s01 TIMEBOOST_cell_8480 ( .a(n_6610), .b(n_6802), .o(TIMEBOOST_net_2727) );
no02s02 FE_RC_2110_0 ( .a(n_41687), .b(n_41527), .o(FE_RN_854_0) );
no02s02 FE_RC_2111_0 ( .a(n_41529), .b(n_41530), .o(FE_RN_855_0) );
in01m02 FE_RC_2113_0 ( .a(FE_RN_857_0), .o(n_41941) );
no02m02 TIMEBOOST_cell_7937 ( .a(TIMEBOOST_net_2599), .b(n_5231), .o(n_5461) );
no02s02 TIMEBOOST_cell_7520 ( .a(n_13312), .b(n_13110), .o(TIMEBOOST_net_2391) );
in01s01 FE_RC_2116_0 ( .a(n_18843), .o(FE_RN_859_0) );
no02s04 FE_RC_2117_0 ( .a(n_18964), .b(FE_RN_859_0), .o(FE_RN_860_0) );
no03m06 TIMEBOOST_cell_8842 ( .a(n_10339), .b(n_10338), .c(n_10354), .o(TIMEBOOST_net_2908) );
na02s04 TIMEBOOST_cell_8645 ( .a(TIMEBOOST_net_2809), .b(n_31105), .o(n_31194) );
na02s06 TIMEBOOST_cell_6789 ( .a(FE_OCP_RBN4457_n_43103), .b(n_43140), .o(TIMEBOOST_net_2152) );
na02s02 TIMEBOOST_cell_7618 ( .a(n_2697), .b(n_2393), .o(TIMEBOOST_net_2440) );
in01s01 FE_RC_2122_0 ( .a(n_7768), .o(FE_RN_864_0) );
in01s01 FE_RC_2123_0 ( .a(FE_OCP_RBN5608_n_7730), .o(FE_RN_865_0) );
no02s01 FE_RC_2124_0 ( .a(FE_RN_865_0), .b(FE_RN_864_0), .o(FE_RN_866_0) );
na02f06 FE_RC_2126_0 ( .a(FE_RN_867_0), .b(n_7815), .o(n_8215) );
no02s03 TIMEBOOST_cell_7747 ( .a(TIMEBOOST_net_2504), .b(FE_RN_1916_0), .o(n_47005) );
in01s01 FE_RC_2132_0 ( .a(n_37654), .o(FE_RN_871_0) );
in01s02 FE_RC_2133_0 ( .a(n_38185), .o(FE_RN_872_0) );
na02s06 FE_RC_2134_0 ( .a(FE_RN_871_0), .b(FE_RN_872_0), .o(FE_RN_873_0) );
no02s03 FE_RC_2135_0 ( .a(n_38164), .b(n_38131), .o(FE_RN_874_0) );
ao22f08 FE_RC_2136_0 ( .a(FE_OCP_RBN4058_n_44875), .b(FE_RN_873_0), .c(FE_RN_874_0), .d(n_38420), .o(n_38474) );
na02s01 FE_RC_2137_0 ( .a(n_8059), .b(n_8018), .o(FE_RN_875_0) );
in01s01 FE_RC_2138_0 ( .a(n_8048), .o(FE_RN_876_0) );
no02s01 FE_RC_2139_0 ( .a(FE_RN_875_0), .b(FE_RN_876_0), .o(FE_RN_877_0) );
in01s02 FE_RC_213_0 ( .a(n_23043), .o(FE_RN_57_0) );
na02f08 FE_RC_2140_0 ( .a(n_8684), .b(FE_RN_877_0), .o(n_8733) );
na02s06 FE_RC_2141_0 ( .a(FE_OCPN1354_n_22484), .b(n_24964), .o(FE_RN_878_0) );
no02s06 FE_RC_2142_0 ( .a(n_24986), .b(FE_RN_878_0), .o(n_25067) );
oa22s02 FE_RC_2143_0 ( .a(n_6639), .b(n_6665), .c(n_6640), .d(n_6666), .o(n_6832) );
in01s06 FE_RC_2144_0 ( .a(FE_RN_879_0), .o(n_36887) );
no02f03 FE_RC_2145_0 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_2_), .b(delay_add_ln22_unr23_stage9_stallmux_q_2_), .o(FE_RN_879_0) );
in01s06 FE_RC_2146_0 ( .a(n_12039), .o(FE_RN_880_0) );
in01s06 FE_RC_2147_0 ( .a(n_12038), .o(FE_RN_881_0) );
in01m06 FE_RC_214_0 ( .a(n_23046), .o(FE_RN_58_0) );
in01s06 FE_RC_2150_0 ( .a(n_12056), .o(FE_RN_882_0) );
na02s08 FE_RC_2151_0 ( .a(n_12423), .b(FE_RN_882_0), .o(n_12492) );
in01s01 FE_RC_2155_0 ( .a(n_2817), .o(FE_RN_885_0) );
no02s01 FE_RC_2156_0 ( .a(FE_RN_885_0), .b(n_2838), .o(FE_RN_886_0) );
na02f08 FE_RC_2157_0 ( .a(FE_RN_886_0), .b(n_3326), .o(n_3365) );
no02s02 FE_RC_2158_0 ( .a(n_2935), .b(n_2900), .o(FE_RN_887_0) );
in01s01 FE_RC_2159_0 ( .a(FE_OFN797_n_2285), .o(FE_RN_888_0) );
no02f08 FE_RC_215_0 ( .a(FE_RN_58_0), .b(FE_RN_57_0), .o(FE_RN_59_0) );
in01s01 FE_RC_2160_0 ( .a(n_2814), .o(FE_RN_889_0) );
na02f08 TIMEBOOST_cell_2071 ( .a(n_34186), .b(FE_RN_2094_0), .o(TIMEBOOST_net_650) );
in01s01 FE_RC_2162_0 ( .a(n_2913), .o(FE_RN_891_0) );
no02f04 TIMEBOOST_cell_2068 ( .a(TIMEBOOST_net_648), .b(n_8741), .o(n_8835) );
in01s01 FE_RC_2164_0 ( .a(n_2880), .o(FE_RN_893_0) );
na02s06 TIMEBOOST_cell_2846 ( .a(FE_RN_800_0), .b(FE_RN_795_0), .o(TIMEBOOST_net_714) );
na02f08 FE_RC_2166_0 ( .a(n_3365), .b(FE_RN_894_0), .o(FE_RN_895_0) );
na02f10 FE_RC_2167_0 ( .a(FE_RN_895_0), .b(FE_RN_887_0), .o(n_3456) );
in01s01 FE_RC_2168_0 ( .a(n_2882), .o(FE_RN_896_0) );
no02s01 FE_RC_2169_0 ( .a(FE_RN_896_0), .b(n_2937), .o(FE_RN_897_0) );
na02m40 TIMEBOOST_cell_7401 ( .a(n_32577), .b(TIMEBOOST_net_2331), .o(n_32575) );
no02s08 TIMEBOOST_cell_8483 ( .a(TIMEBOOST_net_2728), .b(TIMEBOOST_net_2195), .o(n_12128) );
no02m10 TIMEBOOST_cell_3001 ( .a(n_29258), .b(TIMEBOOST_net_791), .o(n_29316) );
na02m06 TIMEBOOST_cell_3002 ( .a(n_41978), .b(n_41860), .o(TIMEBOOST_net_792) );
na02f06 FE_RC_2174_0 ( .a(n_2009), .b(n_1844), .o(FE_RN_901_0) );
na02f08 FE_RC_2175_0 ( .a(FE_RN_901_0), .b(n_1845), .o(n_2063) );
in01s02 FE_RC_2176_0 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_21_), .o(FE_RN_902_0) );
na02s01 TIMEBOOST_cell_7596 ( .a(FE_OCP_RBN2570_n_33735), .b(FE_OCP_RBN6668_n_34297), .o(TIMEBOOST_net_2429) );
no03s04 TIMEBOOST_cell_3572 ( .a(FE_RN_942_0), .b(FE_RN_943_0), .c(n_3032), .o(n_47022) );
na02m06 FE_RC_2179_0 ( .a(FE_RN_904_0), .b(n_40894), .o(n_40942) );
in01m08 FE_RC_217_0 ( .a(FE_OCP_RBN2388_n_23227), .o(FE_RN_60_0) );
no02m08 FE_RC_2180_0 ( .a(n_40777), .b(n_40811), .o(FE_RN_905_0) );
na02f08 FE_RC_2181_0 ( .a(FE_RN_905_0), .b(n_40866), .o(n_41084) );
in01m40 FE_RC_2187_0 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_2_), .o(FE_RN_909_0) );
na02m80 FE_RC_2188_0 ( .a(FE_RN_909_0), .b(n_44962), .o(n_32577) );
in01m08 FE_RC_218_0 ( .a(n_23226), .o(FE_RN_61_0) );
na02s06 FE_RC_2191_0 ( .a(n_12810), .b(n_12841), .o(FE_RN_911_0) );
no02f08 FE_RC_2192_0 ( .a(FE_RN_911_0), .b(n_13100), .o(n_13136) );
in01s01 FE_RC_2193_0 ( .a(n_18171), .o(FE_RN_912_0) );
na02m02 FE_RC_2194_0 ( .a(n_18202), .b(FE_RN_912_0), .o(n_18218) );
oa22m04 FE_RC_2195_0 ( .a(FE_OCP_RBN4221_n_8732), .b(n_44576), .c(n_8732), .d(FE_OCP_RBN6712_n_44570), .o(n_9020) );
na02m08 FE_RC_219_0 ( .a(FE_RN_60_0), .b(FE_RN_61_0), .o(FE_RN_62_0) );
oa22m02 FE_RC_2201_0 ( .a(n_36706), .b(n_36772), .c(n_36771), .d(FE_OCP_RBN3410_n_36706), .o(n_36800) );
in01s02 FE_RC_2202_0 ( .a(n_11991), .o(FE_RN_916_0) );
in01s01 FE_RC_2203_0 ( .a(n_11882), .o(FE_RN_917_0) );
na02s06 FE_RC_2204_0 ( .a(FE_RN_916_0), .b(FE_RN_917_0), .o(FE_RN_918_0) );
no02s01 TIMEBOOST_cell_8856 ( .a(n_16977), .b(FE_OCP_RBN6073_n_16086), .o(TIMEBOOST_net_2915) );
ao22s02 FE_RC_2206_0 ( .a(n_3639), .b(n_4642), .c(n_3638), .d(n_3025), .o(n_3677) );
in01s01 FE_RC_2207_0 ( .a(n_2871), .o(FE_RN_919_0) );
na02s02 FE_RC_2208_0 ( .a(FE_OCP_RBN5566_n_2346), .b(n_2799), .o(FE_RN_920_0) );
no02m04 FE_RC_2209_0 ( .a(n_3063), .b(FE_RN_920_0), .o(FE_RN_921_0) );
in01s01 FE_RC_2210_0 ( .a(n_2870), .o(FE_RN_922_0) );
no02m04 FE_RC_2211_0 ( .a(n_3034), .b(n_3063), .o(FE_RN_923_0) );
oa22m04 FE_RC_2212_0 ( .a(FE_RN_919_0), .b(FE_RN_921_0), .c(FE_RN_922_0), .d(FE_RN_923_0), .o(n_3149) );
na02s06 TIMEBOOST_cell_6007 ( .a(n_28544), .b(n_28542), .o(TIMEBOOST_net_1855) );
no02s02 TIMEBOOST_cell_5662 ( .a(FE_OCPN900_n_16923), .b(FE_OCP_RBN4396_n_16146), .o(TIMEBOOST_net_1779) );
no02f06 FE_RC_2215_0 ( .a(n_4927), .b(n_4371), .o(FE_RN_925_0) );
na02s02 FE_RC_2216_0 ( .a(n_4261), .b(n_4215), .o(FE_RN_926_0) );
in01s01 FE_RC_2217_0 ( .a(n_4371), .o(FE_RN_927_0) );
ao12f06 FE_RC_2218_0 ( .a(FE_RN_925_0), .b(FE_RN_926_0), .c(FE_RN_927_0), .o(n_5144) );
in01s01 FE_RC_2219_0 ( .a(n_37068), .o(FE_RN_928_0) );
no02m02 TIMEBOOST_cell_1647 ( .a(n_14979), .b(FE_OCP_RBN2834_n_13962), .o(TIMEBOOST_net_438) );
in01s02 FE_RC_2220_0 ( .a(n_37290), .o(FE_RN_929_0) );
no02s02 FE_RC_2221_0 ( .a(FE_RN_929_0), .b(FE_RN_928_0), .o(FE_RN_930_0) );
in01s01 FE_RC_2222_0 ( .a(n_36955), .o(FE_RN_931_0) );
no02s01 TIMEBOOST_cell_4535 ( .a(FE_OCP_RBN6875_n_31520), .b(FE_OCPN908_n_46956), .o(TIMEBOOST_net_1358) );
in01m08 FE_RC_2224_0 ( .a(FE_RN_933_0), .o(n_37694) );
na02f06 TIMEBOOST_cell_8739 ( .a(TIMEBOOST_net_2856), .b(n_13860), .o(TIMEBOOST_net_2408) );
no02s01 TIMEBOOST_cell_4885 ( .a(TIMEBOOST_net_1390), .b(n_44042), .o(TIMEBOOST_net_163) );
na02s04 TIMEBOOST_cell_8644 ( .a(FE_OCP_RBN6833_n_31073), .b(FE_OCPN1340_n_27246), .o(TIMEBOOST_net_2809) );
no02s02 TIMEBOOST_cell_1257 ( .a(n_37850), .b(n_37849), .o(TIMEBOOST_net_243) );
no02f06 TIMEBOOST_cell_1258 ( .a(TIMEBOOST_net_243), .b(n_37892), .o(n_38010) );
no02f08 FE_RC_2232_0 ( .a(FE_RN_938_0), .b(n_22172), .o(FE_RN_939_0) );
in01s06 FE_RC_2233_0 ( .a(n_22041), .o(FE_RN_940_0) );
oa22f08 FE_RC_2234_0 ( .a(FE_RN_940_0), .b(FE_RN_939_0), .c(FE_RN_940_0), .d(n_22356), .o(n_22450) );
na02s02 FE_RC_2235_0 ( .a(n_3958), .b(n_4035), .o(FE_RN_941_0) );
no02s04 FE_RC_2236_0 ( .a(FE_RN_941_0), .b(n_4075), .o(n_4235) );
in01s01 FE_RC_2237_0 ( .a(n_2333), .o(FE_RN_942_0) );
in01s01 FE_RC_2238_0 ( .a(n_3031), .o(FE_RN_943_0) );
no02f08 TIMEBOOST_cell_4142 ( .a(n_35673), .b(TIMEBOOST_net_1161), .o(n_35878) );
no02s01 TIMEBOOST_cell_4143 ( .a(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(FE_OFN5084_n_36750), .o(TIMEBOOST_net_1162) );
in01s08 FE_RC_2241_0 ( .a(n_22927), .o(FE_RN_945_0) );
in01s06 FE_RC_2242_0 ( .a(n_22748), .o(FE_RN_946_0) );
na03s08 TIMEBOOST_cell_8190 ( .a(n_11917), .b(n_11765), .c(n_11957), .o(n_12098) );
na02s04 TIMEBOOST_cell_5641 ( .a(TIMEBOOST_net_1768), .b(n_6133), .o(n_6233) );
in01s20 FE_RC_2245_0 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_8_), .o(FE_RN_948_0) );
no02s40 FE_RC_2246_0 ( .a(FE_RN_948_0), .b(FE_OCP_RBN2039_n_44722), .o(n_28032) );
ao22m10 FE_RC_2249_0 ( .a(n_45224), .b(n_11696), .c(FE_OCP_RBN6317_n_45224), .d(delay_xor_ln22_unr9_stage4_stallmux_q_2_), .o(n_11734) );
in01s02 FE_RC_224_0 ( .a(FE_OCPN1906_n_23322), .o(FE_RN_63_0) );
oa22s06 FE_RC_2250_0 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_0_), .b(n_45224), .c(n_11593), .d(FE_OCP_RBN6321_n_45224), .o(n_11761) );
in01s01 FE_RC_2254_0 ( .a(n_37894), .o(FE_RN_952_0) );
na02s06 TIMEBOOST_cell_6606 ( .a(TIMEBOOST_net_2060), .b(FE_RN_179_0), .o(n_17667) );
no02f04 TIMEBOOST_cell_8120 ( .a(FE_RN_42_0), .b(FE_RN_43_0), .o(TIMEBOOST_net_2691) );
no02f06 FE_RC_2257_0 ( .a(FE_RN_954_0), .b(n_38062), .o(n_38122) );
in01s01 FE_RC_225_0 ( .a(n_23229), .o(FE_RN_64_0) );
na02f04 FE_RC_2265_0 ( .a(n_20070), .b(FE_OCP_RBN3706_n_18716), .o(FE_RN_959_0) );
in01s02 FE_RC_2266_0 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_9_), .o(FE_RN_960_0) );
in01m02 FE_RC_2267_0 ( .a(n_23266), .o(FE_RN_961_0) );
na02f04 TIMEBOOST_cell_7956 ( .a(n_10598), .b(n_10624), .o(TIMEBOOST_net_2609) );
no02m02 TIMEBOOST_cell_8753 ( .a(TIMEBOOST_net_2863), .b(FE_RN_310_0), .o(FE_RN_311_0) );
na02s04 FE_RC_226_0 ( .a(FE_RN_63_0), .b(FE_RN_64_0), .o(FE_RN_65_0) );
in01s02 FE_RC_2273_0 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_3_), .o(FE_RN_964_0) );
no02s06 FE_RC_2275_0 ( .a(FE_RN_964_0), .b(FE_OCP_RBN6514_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_RN_966_0) );
no02s06 FE_RC_2276_0 ( .a(n_1542), .b(FE_RN_966_0), .o(n_1436) );
no02m06 TIMEBOOST_cell_1674 ( .a(TIMEBOOST_net_451), .b(n_34830), .o(n_34903) );
in01s01 FE_RC_2278_0 ( .a(n_38279), .o(FE_RN_967_0) );
no02s01 FE_RC_2279_0 ( .a(FE_RN_967_0), .b(n_37569), .o(FE_RN_968_0) );
no02s01 TIMEBOOST_cell_1635 ( .a(FE_OCPN1270_n_30577), .b(n_30244), .o(TIMEBOOST_net_432) );
no02s06 FE_RC_2280_0 ( .a(n_38007), .b(FE_RN_968_0), .o(n_38121) );
in01s10 FE_RC_2281_0 ( .a(n_17617), .o(FE_RN_969_0) );
na03s04 TIMEBOOST_cell_8290 ( .a(n_9271), .b(FE_OFN4768_n_8309), .c(FE_OCP_RBN4236_n_9089), .o(FE_RN_314_0) );
no02s02 TIMEBOOST_cell_6761 ( .a(n_15810), .b(n_15516), .o(TIMEBOOST_net_2138) );
na02m04 TIMEBOOST_cell_7989 ( .a(n_26140), .b(TIMEBOOST_net_2625), .o(n_26180) );
oa22m02 FE_RC_2287_0 ( .a(n_8657), .b(FE_OCP_RBN5739_n_8402), .c(FE_OCP_RBN5737_n_8402), .d(FE_OCP_RBN5784_n_8657), .o(n_8776) );
no02s01 TIMEBOOST_cell_3823 ( .a(n_6504), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(TIMEBOOST_net_1002) );
in01m02 FE_RC_2289_0 ( .a(n_8251), .o(FE_RN_974_0) );
no02s03 TIMEBOOST_cell_1661 ( .a(n_19732), .b(n_20058), .o(TIMEBOOST_net_445) );
no03f10 TIMEBOOST_cell_2218 ( .a(n_40825), .b(n_40826), .c(n_40725), .o(n_40866) );
in01s02 FE_RC_2291_0 ( .a(n_8208), .o(FE_RN_976_0) );
no02m04 FE_RC_2292_0 ( .a(FE_RN_975_0), .b(FE_RN_976_0), .o(FE_RN_977_0) );
no02m06 FE_RC_2293_0 ( .a(n_8234), .b(FE_RN_977_0), .o(n_8403) );
oa22m04 FE_RC_2294_0 ( .a(n_38201), .b(n_38506), .c(n_38202), .d(n_38460), .o(n_38537) );
oa22f04 FE_RC_2295_0 ( .a(n_38778), .b(n_38545), .c(FE_OCP_RBN4172_n_38545), .d(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38594) );
oa22f04 FE_RC_2296_0 ( .a(n_38214), .b(FE_OCP_RBN6674_n_38519), .c(n_38215), .d(n_38519), .o(n_38583) );
na02m04 FE_RC_2297_0 ( .a(n_38778), .b(n_38537), .o(FE_RN_978_0) );
no02m08 TIMEBOOST_cell_4206 ( .a(TIMEBOOST_net_1193), .b(n_32741), .o(n_32788) );
na02s01 TIMEBOOST_cell_8832 ( .a(n_4316), .b(FE_OCP_RBN2966_n_4046), .o(TIMEBOOST_net_2903) );
in01s01 FE_RC_2300_0 ( .a(n_8437), .o(FE_RN_980_0) );
in01f02 FE_RC_2301_0 ( .a(FE_RN_981_0), .o(n_8626) );
na02f02 FE_RC_2302_0 ( .a(FE_RN_980_0), .b(n_8515), .o(FE_RN_981_0) );
in01s01 FE_RC_2303_0 ( .a(n_2526), .o(FE_RN_982_0) );
no02m08 TIMEBOOST_cell_3005 ( .a(TIMEBOOST_net_793), .b(n_24561), .o(n_24718) );
no02f08 TIMEBOOST_cell_3006 ( .a(FE_RN_2375_0), .b(FE_OCPN939_n_23577), .o(TIMEBOOST_net_794) );
in01s01 FE_RC_2307_0 ( .a(n_41121), .o(FE_RN_985_0) );
na02s04 FE_RC_2308_0 ( .a(n_41435), .b(FE_RN_985_0), .o(n_41577) );
oa22f06 FE_RC_230_0 ( .a(n_25380), .b(n_25632), .c(n_25354), .d(n_25600), .o(n_25731) );
ao22m04 FE_RC_2311_0 ( .a(n_23717), .b(n_24094), .c(n_23716), .d(FE_OCP_RBN1006_n_24094), .o(n_24175) );
na02m06 FE_RC_2312_0 ( .a(n_3204), .b(n_2385), .o(FE_RN_986_0) );
na02m08 FE_RC_2313_0 ( .a(FE_RN_986_0), .b(FE_OCPN3560_n_2386), .o(n_3318) );
no02m02 FE_RC_2315_0 ( .a(FE_OCP_RBN6583_n_8021), .b(n_8776), .o(FE_RN_987_0) );
na02m02 FE_RC_2316_0 ( .a(FE_OCPN931_n_7817), .b(n_8803), .o(FE_RN_988_0) );
na02m04 FE_RC_2317_0 ( .a(FE_RN_988_0), .b(n_8799), .o(n_8968) );
in01s01 FE_RC_2319_0 ( .a(n_37587), .o(FE_RN_989_0) );
na02s06 FE_RC_2320_0 ( .a(n_38007), .b(FE_RN_989_0), .o(n_38089) );
in01m04 FE_RC_2321_0 ( .a(n_22998), .o(FE_RN_990_0) );
no02m06 FE_RC_2322_0 ( .a(n_23110), .b(FE_RN_990_0), .o(n_23176) );
na02s02 FE_RC_2324_0 ( .a(FE_OCP_RBN2598_n_7743), .b(n_8915), .o(FE_RN_991_0) );
in01s01 FE_RC_2325_0 ( .a(FE_OFN4770_n_8309), .o(FE_RN_992_0) );
oa12m02 FE_RC_2326_0 ( .a(FE_RN_991_0), .b(FE_RN_992_0), .c(n_8915), .o(n_9080) );
in01s01 FE_RC_2327_0 ( .a(n_9012), .o(FE_RN_993_0) );
in01m04 FE_RC_2328_0 ( .a(FE_RN_994_0), .o(n_9347) );
na02m02 FE_RC_2329_0 ( .a(FE_RN_993_0), .b(n_9080), .o(FE_RN_994_0) );
ao22s02 FE_RC_2330_0 ( .a(n_2912), .b(n_3812), .c(n_2911), .d(n_3736), .o(n_3981) );
ao22m04 FE_RC_2332_0 ( .a(n_7574), .b(n_8910), .c(n_7575), .d(n_8864), .o(n_9044) );
no02f02 FE_RC_2333_0 ( .a(FE_OCPN1073_n_12638), .b(n_12983), .o(FE_RN_995_0) );
no02f06 FE_RC_2335_0 ( .a(n_42199), .b(n_42234), .o(FE_RN_996_0) );
no02f08 FE_RC_2336_0 ( .a(FE_RN_996_0), .b(n_42207), .o(n_42240) );
in01s01 FE_RC_2337_0 ( .a(n_2947), .o(FE_RN_997_0) );
no02s01 FE_RC_2339_0 ( .a(FE_RN_997_0), .b(n_3830), .o(FE_RN_998_0) );
no02s06 FE_RC_2343_0 ( .a(n_11608), .b(n_11596), .o(FE_RN_1000_0) );
na02m08 FE_RC_2344_0 ( .a(n_11777), .b(FE_RN_1000_0), .o(n_11853) );
ao22s03 FE_RC_2345_0 ( .a(n_3635), .b(n_2810), .c(n_2809), .d(n_3579), .o(n_3718) );
oa22m02 FE_RC_2353_0 ( .a(n_3106), .b(FE_OCP_RBN4292_n_4080), .c(n_3082), .d(n_4080), .o(n_4313) );
oa22m04 FE_RC_2354_0 ( .a(n_3807), .b(FE_OFN4763_n_3029), .c(n_3615), .d(FE_OCP_RBN5855_n_3807), .o(n_3963) );
oa22s02 FE_RC_2358_0 ( .a(n_4057), .b(n_2998), .c(n_2997), .d(n_4131), .o(n_4238) );
no02m06 FE_RC_2359_0 ( .a(n_34037), .b(n_33825), .o(FE_RN_1005_0) );
no02m08 FE_RC_2360_0 ( .a(FE_RN_1005_0), .b(FE_OCP_RBN1815_n_33873), .o(n_33957) );
no02f06 FE_RC_2363_0 ( .a(n_29349), .b(n_28737), .o(FE_RN_1007_0) );
ao12f04 FE_RC_2364_0 ( .a(FE_RN_1007_0), .b(n_28737), .c(n_29349), .o(n_29450) );
ao22m04 FE_RC_2365_0 ( .a(n_23917), .b(n_24424), .c(n_23918), .d(n_24423), .o(n_24518) );
na02f02 FE_RC_2366_0 ( .a(n_29450), .b(FE_OFN774_n_25834), .o(FE_RN_1008_0) );
in01s01 FE_RC_2367_0 ( .a(n_29561), .o(FE_RN_1009_0) );
oa12f02 FE_RC_2368_0 ( .a(FE_RN_1008_0), .b(FE_RN_1009_0), .c(n_29450), .o(n_29566) );
in01s02 FE_RC_2369_0 ( .a(n_9351), .o(FE_RN_1010_0) );
oa22f04 FE_RC_236_0 ( .a(n_25670), .b(n_26154), .c(n_25671), .d(n_26153), .o(n_26291) );
no02s04 FE_RC_2370_0 ( .a(FE_RN_1010_0), .b(n_9552), .o(FE_RN_1011_0) );
na02m04 FE_RC_2371_0 ( .a(FE_RN_1011_0), .b(n_9424), .o(FE_RN_1012_0) );
no02f06 FE_RC_2373_0 ( .a(FE_RN_1013_0), .b(FE_RN_1012_0), .o(n_9764) );
in01f04 FE_RC_2375_0 ( .a(n_13689), .o(FE_RN_1015_0) );
na02f08 FE_RC_2376_0 ( .a(FE_OCP_RBN2540_n_12880), .b(FE_RN_1015_0), .o(FE_RN_1016_0) );
na02f08 FE_RC_2377_0 ( .a(n_47253), .b(FE_RN_1016_0), .o(n_13702) );
in01s01 FE_RC_2378_0 ( .a(FE_RN_1018_0), .o(FE_RN_1017_0) );
no02s01 FE_RC_2379_0 ( .a(FE_RN_1017_0), .b(n_23124), .o(n_23235) );
in01m04 FE_RC_2380_0 ( .a(n_23124), .o(FE_RN_1019_0) );
na02f06 FE_RC_2381_0 ( .a(n_23191), .b(n_23187), .o(FE_RN_1018_0) );
na02m06 FE_RC_2385_0 ( .a(delay_sub_ln23_0_unr21_stage8_stallmux_q), .b(n_33872), .o(FE_RN_1021_0) );
na02m08 FE_RC_2386_0 ( .a(FE_RN_1021_0), .b(n_33957), .o(n_33977) );
oa22m02 FE_RC_2389_0 ( .a(n_13016), .b(n_13633), .c(n_13044), .d(n_13594), .o(n_13667) );
no02s01 TIMEBOOST_cell_5218 ( .a(FE_OCP_RBN2078_n_14149), .b(n_15142), .o(TIMEBOOST_net_1557) );
in01f04 FE_RC_2390_0 ( .a(FE_RN_1023_0), .o(n_23196) );
no02f06 FE_RC_2391_0 ( .a(n_23069), .b(delay_add_ln22_unr14_stage6_stallmux_q_4_), .o(FE_RN_1023_0) );
ao22s02 FE_RC_2392_0 ( .a(n_4690), .b(n_4754), .c(n_4753), .d(n_4624), .o(n_4925) );
in01s01 FE_RC_2394_0 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_23_), .o(FE_RN_1025_0) );
na02s06 FE_RC_2395_0 ( .a(n_13213), .b(FE_RN_1025_0), .o(FE_RN_1026_0) );
no02s03 FE_RC_2396_0 ( .a(n_46414), .b(n_13173), .o(FE_RN_1027_0) );
na02f08 FE_RC_2398_0 ( .a(n_15035), .b(n_15124), .o(FE_RN_1028_0) );
na02f08 FE_RC_2399_0 ( .a(n_15036), .b(FE_RN_1028_0), .o(n_15321) );
in01s02 FE_RC_239_0 ( .a(n_23077), .o(FE_RN_67_0) );
na02s06 FE_RC_2400_0 ( .a(n_29417), .b(n_29630), .o(FE_RN_1029_0) );
na02f08 FE_RC_2401_0 ( .a(FE_RN_1029_0), .b(n_29697), .o(n_29730) );
na02s01 TIMEBOOST_cell_8762 ( .a(n_14376), .b(n_13515), .o(TIMEBOOST_net_2868) );
no02s01 TIMEBOOST_cell_3878 ( .a(TIMEBOOST_net_1029), .b(n_521), .o(n_1045) );
na02f06 FE_RC_2406_0 ( .a(n_19104), .b(FE_RN_1032_0), .o(n_19168) );
no02s02 TIMEBOOST_cell_5598 ( .a(FE_OCPN5122_n_44438), .b(n_31931), .o(TIMEBOOST_net_1747) );
in01m10 FE_RC_2408_0 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_3_), .o(FE_RN_1034_0) );
na03m04 TIMEBOOST_cell_7309 ( .a(n_31365), .b(n_31244), .c(n_31383), .o(n_31474) );
in01s02 FE_RC_240_0 ( .a(FE_RN_68_0), .o(n_23107) );
no02s02 TIMEBOOST_cell_5599 ( .a(TIMEBOOST_net_1747), .b(FE_OCP_RBN6203_n_31819), .o(n_32132) );
no02s02 FE_RC_2413_0 ( .a(FE_OCP_RBN5960_n_4397), .b(n_4403), .o(FE_RN_1038_0) );
oa22m04 FE_RC_2415_0 ( .a(FE_RN_1038_0), .b(n_4592), .c(FE_OCP_RBN3026_n_4699), .d(n_4630), .o(n_4906) );
na02s01 FE_RC_2416_0 ( .a(sin_out_20), .b(FE_OFN5_n_43918), .o(FE_RN_1040_0) );
in01s01 FE_RC_2417_0 ( .a(n_43398), .o(FE_RN_1041_0) );
no02s02 FE_RC_2418_0 ( .a(FE_RN_1041_0), .b(n_43809), .o(FE_RN_1042_0) );
in01s01 FE_RC_2419_0 ( .a(n_43398), .o(FE_RN_1043_0) );
no02s01 TIMEBOOST_cell_3949 ( .a(n_20036), .b(n_19787), .o(TIMEBOOST_net_1065) );
ao12s02 FE_RC_2420_0 ( .a(FE_RN_1042_0), .b(FE_RN_1043_0), .c(n_43809), .o(FE_RN_1044_0) );
oa12s02 FE_RC_2421_0 ( .a(FE_RN_1040_0), .b(FE_OFN5_n_43918), .c(FE_RN_1044_0), .o(n_43888) );
na02m04 FE_RC_2423_0 ( .a(n_33648), .b(FE_OCPN1630_n_33196), .o(FE_RN_1045_0) );
no02s02 FE_RC_2425_0 ( .a(n_43349), .b(n_43646), .o(FE_RN_1046_0) );
in01s01 FE_RC_2426_0 ( .a(n_43359), .o(FE_RN_1047_0) );
na02f04 FE_RC_2427_0 ( .a(n_43833), .b(FE_RN_1047_0), .o(FE_RN_1048_0) );
na02f04 FE_RC_2428_0 ( .a(FE_RN_1048_0), .b(FE_RN_1046_0), .o(n_43874) );
ao22m02 FE_RC_2429_0 ( .a(n_4968), .b(n_5083), .c(n_5082), .d(n_4969), .o(n_5221) );
ao22s10 FE_RC_242_0 ( .a(FE_OCP_RBN1109_n_44061), .b(delay_xor_ln21_unr15_stage6_stallmux_q_4_), .c(FE_OCP_RBN5179_n_44061), .d(n_22939), .o(n_22992) );
no02s06 FE_RC_2434_0 ( .a(n_34224), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(FE_RN_1051_0) );
no02m06 TIMEBOOST_cell_2092 ( .a(TIMEBOOST_net_660), .b(n_30576), .o(n_30643) );
na02s01 TIMEBOOST_cell_8492 ( .a(n_7250), .b(n_7348), .o(TIMEBOOST_net_2733) );
no02m02 TIMEBOOST_cell_4159 ( .a(n_26664), .b(n_26663), .o(TIMEBOOST_net_1170) );
in01s01 FE_RC_2439_0 ( .a(n_13204), .o(FE_RN_1054_0) );
in01m04 FE_RC_243_0 ( .a(n_363), .o(FE_RN_69_0) );
na02s01 FE_RC_2440_0 ( .a(FE_RN_1054_0), .b(n_13777), .o(FE_RN_1055_0) );
no02m06 FE_RC_2441_0 ( .a(n_13732), .b(FE_RN_1055_0), .o(n_13774) );
na02m04 FE_RC_2442_0 ( .a(n_7844), .b(n_7938), .o(FE_RN_1056_0) );
na02m06 FE_RC_2443_0 ( .a(n_7847), .b(FE_RN_1056_0), .o(n_8066) );
na02s06 FE_RC_2447_0 ( .a(n_39009), .b(n_39010), .o(FE_RN_1059_0) );
no02s06 FE_RC_2448_0 ( .a(FE_RN_1059_0), .b(n_38987), .o(n_39139) );
in01s01 FE_RC_2449_0 ( .a(n_29630), .o(FE_RN_1060_0) );
no02m03 TIMEBOOST_cell_4890 ( .a(n_12071), .b(n_11796), .o(TIMEBOOST_net_1393) );
no02s06 FE_RC_2450_0 ( .a(n_29628), .b(FE_RN_1060_0), .o(FE_RN_522_0) );
oa22m06 FE_RC_2451_0 ( .a(n_9297), .b(n_9438), .c(n_9368), .d(n_9357), .o(n_9629) );
in01s01 FE_RC_2452_0 ( .a(n_38060), .o(FE_RN_1061_0) );
na02m04 FE_RC_2453_0 ( .a(FE_RN_1061_0), .b(FE_OCP_RBN5885_n_38806), .o(n_38864) );
oa22m06 FE_RC_2455_0 ( .a(n_17783), .b(FE_OCP_RBN1131_n_19077), .c(n_17900), .d(n_19077), .o(n_19278) );
ao22m04 FE_RC_2456_0 ( .a(n_18032), .b(FE_OCP_RBN1826_n_19513), .c(n_19418), .d(n_19513), .o(n_19633) );
na02f02 FE_RC_2458_0 ( .a(n_5477), .b(n_5472), .o(FE_RN_1062_0) );
no02m02 FE_RC_2459_0 ( .a(n_5476), .b(n_5512), .o(FE_RN_1063_0) );
in01f06 FE_RC_245_0 ( .a(FE_RN_71_0), .o(n_386) );
na02f02 FE_RC_2460_0 ( .a(FE_RN_1062_0), .b(FE_RN_1063_0), .o(n_5608) );
in01s01 FE_RC_2463_0 ( .a(n_18631), .o(FE_RN_1065_0) );
no02s06 TIMEBOOST_cell_1945 ( .a(n_32600), .b(n_32602), .o(TIMEBOOST_net_587) );
no02f06 TIMEBOOST_cell_8646 ( .a(FE_RN_1873_0), .b(n_39596), .o(TIMEBOOST_net_2810) );
no02s04 TIMEBOOST_cell_8562 ( .a(n_44872), .b(n_37909), .o(TIMEBOOST_net_2768) );
in01s01 FE_RC_2470_0 ( .a(n_33613), .o(FE_RN_1069_0) );
no02s06 FE_RC_2471_0 ( .a(n_44102), .b(FE_RN_1069_0), .o(n_34162) );
in01s01 FE_RC_2472_0 ( .a(n_23914), .o(FE_RN_1070_0) );
na02s04 FE_RC_2473_0 ( .a(FE_RN_1070_0), .b(n_24323), .o(FE_RN_1071_0) );
in01s01 FE_RC_2476_0 ( .a(FE_OCP_RBN4087_n_12880), .o(FE_RN_1073_0) );
in01m02 FE_RC_2477_0 ( .a(FE_RN_1074_0), .o(n_14203) );
no02f02 FE_RC_2478_0 ( .a(FE_RN_1073_0), .b(n_14096), .o(FE_RN_1074_0) );
no02m02 TIMEBOOST_cell_1975 ( .a(n_37602), .b(n_37579), .o(TIMEBOOST_net_602) );
in01m04 FE_RC_247_0 ( .a(n_23208), .o(FE_RN_72_0) );
no02s01 TIMEBOOST_cell_8500 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_), .b(FE_RN_216_0), .o(TIMEBOOST_net_2737) );
oa22f04 FE_RC_2481_0 ( .a(n_27605), .b(n_27499), .c(n_27604), .d(n_27498), .o(n_27686) );
na02f10 FE_RC_2482_0 ( .a(n_27554), .b(n_27189), .o(n_27568) );
no02f04 FE_RC_2486_0 ( .a(n_38698), .b(n_38766), .o(FE_RN_1077_0) );
na02f04 FE_RC_2487_0 ( .a(n_38698), .b(n_38766), .o(FE_RN_1078_0) );
ao12f04 FE_RC_2488_0 ( .a(FE_RN_1077_0), .b(FE_RN_1078_0), .c(n_38747), .o(n_38780) );
na02f08 TIMEBOOST_cell_6918 ( .a(TIMEBOOST_net_2217), .b(n_24262), .o(n_24359) );
oa22f04 FE_RC_2494_0 ( .a(n_13332), .b(n_13293), .c(n_13245), .d(n_13294), .o(n_13398) );
na02s02 FE_RC_2495_0 ( .a(n_10270), .b(FE_OCP_RBN5906_n_44563), .o(FE_RN_1082_0) );
na02m04 FE_RC_2496_0 ( .a(n_10503), .b(FE_RN_1082_0), .o(FE_RN_1083_0) );
no02f04 FE_RC_2497_0 ( .a(FE_RN_1083_0), .b(n_10377), .o(n_10624) );
in01f03 FE_RC_249_0 ( .a(FE_RN_74_0), .o(n_23365) );
no02s06 FE_RC_2502_0 ( .a(n_19222), .b(n_19223), .o(FE_RN_1086_0) );
no02f06 FE_RC_2503_0 ( .a(n_19516), .b(FE_RN_1086_0), .o(n_19603) );
oa22s02 FE_RC_2504_0 ( .a(n_17330), .b(FE_OCP_RBN1026_n_17417), .c(FE_OCP_RBN1028_n_17417), .d(n_17327), .o(n_17728) );
no03f08 TIMEBOOST_cell_5799 ( .a(n_44946), .b(n_38993), .c(n_38890), .o(TIMEBOOST_net_1577) );
oa22s01 FE_RC_2507_0 ( .a(n_17336), .b(n_17728), .c(FE_OCP_RBN3196_n_15599), .d(n_17682), .o(n_17777) );
no02f04 FE_RC_2508_0 ( .a(n_13290), .b(n_13183), .o(FE_RN_1088_0) );
no02f08 FE_RC_2509_0 ( .a(n_13224), .b(FE_RN_1088_0), .o(n_13394) );
na03s02 TIMEBOOST_cell_2544 ( .a(n_4016), .b(FE_OCP_RBN6744_n_3746), .c(n_4068), .o(n_4360) );
oa22m02 FE_RC_2512_0 ( .a(n_9229), .b(n_9306), .c(n_9230), .d(FE_OCP_RBN5884_n_9306), .o(n_9506) );
na02s01 TIMEBOOST_cell_8588 ( .a(n_29113), .b(n_30364), .o(TIMEBOOST_net_2781) );
in01f04 FE_RC_2517_0 ( .a(n_39907), .o(FE_RN_1093_0) );
na02m04 TIMEBOOST_cell_8510 ( .a(n_13362), .b(n_13365), .o(TIMEBOOST_net_2742) );
no02f06 FE_RC_251_0 ( .a(FE_RN_75_0), .b(n_355), .o(n_379) );
oa22f04 FE_RC_2522_0 ( .a(n_10089), .b(FE_OCP_RBN6011_n_10277), .c(n_10090), .d(FE_OCP_RBN6012_n_10277), .o(n_10477) );
no02s01 FE_RC_2523_0 ( .a(n_34564), .b(n_34565), .o(FE_RN_1095_0) );
in01s02 FE_RC_2524_0 ( .a(n_34511), .o(FE_RN_1096_0) );
na02s06 FE_RC_2525_0 ( .a(FE_RN_1096_0), .b(FE_RN_1095_0), .o(FE_RN_1097_0) );
no02m10 FE_RC_2526_0 ( .a(n_34872), .b(FE_RN_1097_0), .o(n_34927) );
na02f08 FE_RC_2527_0 ( .a(n_25206), .b(n_25205), .o(FE_RN_1098_0) );
no02f10 FE_RC_2528_0 ( .a(n_25513), .b(FE_RN_1098_0), .o(n_25601) );
no02s01 FE_RC_252_0 ( .a(FE_RN_77_0), .b(FE_RN_76_0), .o(FE_RN_75_0) );
na02s02 TIMEBOOST_cell_5544 ( .a(n_6077), .b(n_5966), .o(TIMEBOOST_net_1720) );
na03m08 TIMEBOOST_cell_574 ( .a(n_6288), .b(n_6298), .c(n_6386), .o(n_6387) );
no02s01 TIMEBOOST_cell_4195 ( .a(n_36750), .b(FE_OCPN1950_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_1188) );
ao22m02 FE_RC_2535_0 ( .a(n_10511), .b(n_10322), .c(n_10323), .d(FE_OCP_RBN6041_n_10511), .o(n_10644) );
ao22m02 FE_RC_2537_0 ( .a(n_25662), .b(n_26016), .c(n_25956), .d(n_25661), .o(n_26081) );
no02f04 FE_RC_2538_0 ( .a(n_10399), .b(FE_OCP_RBN5936_n_44563), .o(FE_RN_1104_0) );
na02f08 TIMEBOOST_cell_6928 ( .a(n_29110), .b(TIMEBOOST_net_2222), .o(n_29154) );
in01s01 FE_RC_253_0 ( .a(beta_0), .o(FE_RN_76_0) );
in01s01 TIMEBOOST_cell_8910 ( .a(n_1317), .o(TIMEBOOST_net_2954) );
in01s01 FE_RC_2542_0 ( .a(n_23271), .o(FE_RN_1106_0) );
ao22s04 FE_RC_2545_0 ( .a(n_24830), .b(n_24922), .c(n_24921), .d(n_24831), .o(n_25045) );
in01s01 FE_RC_254_0 ( .a(beta_1), .o(FE_RN_77_0) );
in01s06 FE_RC_2553_0 ( .a(n_25301), .o(FE_RN_1112_0) );
no03m08 TIMEBOOST_cell_8200 ( .a(FE_RN_1977_0), .b(n_32672), .c(n_32761), .o(n_32822) );
na02m02 TIMEBOOST_cell_8654 ( .a(n_36668), .b(FE_OFN5084_n_36750), .o(TIMEBOOST_net_2814) );
in01s01 FE_RC_2561_0 ( .a(n_23447), .o(FE_RN_1116_0) );
in01s03 FE_RC_2562_0 ( .a(FE_RN_1117_0), .o(n_26473) );
no02s02 FE_RC_2563_0 ( .a(FE_RN_1116_0), .b(n_26320), .o(FE_RN_1117_0) );
no02s02 FE_RC_2567_0 ( .a(FE_OCPN1238_n_30470), .b(n_30198), .o(FE_RN_1120_0) );
na02s08 FE_RC_2568_0 ( .a(FE_RN_1120_0), .b(n_30452), .o(n_30467) );
in01s01 FE_RC_256_0 ( .a(n_353), .o(FE_RN_78_0) );
na02m06 FE_RC_2570_0 ( .a(n_10995), .b(n_10957), .o(FE_RN_1121_0) );
no02f06 TIMEBOOST_cell_8121 ( .a(TIMEBOOST_net_2691), .b(n_21034), .o(n_46968) );
na02s06 TIMEBOOST_cell_6612 ( .a(TIMEBOOST_net_2063), .b(n_12161), .o(n_12336) );
in01s01 FE_RC_2573_0 ( .a(n_30369), .o(FE_RN_1123_0) );
in01s01 FE_RC_2574_0 ( .a(n_30601), .o(FE_RN_1124_0) );
ao22f02 FE_RC_2576_0 ( .a(n_14959), .b(n_14871), .c(n_14846), .d(n_14960), .o(n_15079) );
in01s02 FE_RC_2578_0 ( .a(n_10654), .o(FE_RN_1126_0) );
no02m02 TIMEBOOST_cell_5507 ( .a(TIMEBOOST_net_1701), .b(n_5395), .o(n_5549) );
in01s01 FE_RC_257_0 ( .a(n_50), .o(FE_RN_79_0) );
na03s03 TIMEBOOST_cell_8369 ( .a(n_3897), .b(n_3980), .c(n_4010), .o(n_4281) );
na02s02 FE_RC_2581_0 ( .a(FE_OCPN1679_n_27315), .b(n_30733), .o(FE_RN_1128_0) );
na02m06 TIMEBOOST_cell_7804 ( .a(FE_OCP_RBN5954_FE_OFN4772_n_44463), .b(FE_OCP_RBN3288_n_10915), .o(TIMEBOOST_net_2533) );
no02s02 TIMEBOOST_cell_8575 ( .a(TIMEBOOST_net_2774), .b(n_3913), .o(TIMEBOOST_net_1585) );
in01s01 FE_RC_2587_0 ( .a(n_30401), .o(FE_RN_1132_0) );
na02s02 FE_RC_2588_0 ( .a(FE_RN_1132_0), .b(n_30885), .o(FE_RN_1133_0) );
no02s01 FE_RC_258_0 ( .a(FE_RN_78_0), .b(FE_RN_79_0), .o(FE_RN_80_0) );
na02s03 FE_RC_2591_0 ( .a(FE_OFN4799_n_44498), .b(n_11223), .o(FE_RN_1135_0) );
na02m08 FE_RC_2593_0 ( .a(n_11299), .b(FE_RN_1135_0), .o(FE_RN_1136_0) );
oa22f02 FE_RC_2595_0 ( .a(n_40598), .b(n_40578), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .d(n_44687), .o(n_40588) );
na02f08 TIMEBOOST_cell_2989 ( .a(n_13494), .b(TIMEBOOST_net_785), .o(n_13587) );
no02m02 TIMEBOOST_cell_5283 ( .a(TIMEBOOST_net_1589), .b(n_4243), .o(n_4529) );
no02f06 FE_RC_259_0 ( .a(n_354), .b(FE_RN_80_0), .o(n_355) );
no02s06 TIMEBOOST_cell_2990 ( .a(n_19246), .b(n_18849), .o(TIMEBOOST_net_786) );
in01f02 FE_RC_2603_0 ( .a(n_15196), .o(FE_RN_1141_0) );
ao22s03 FE_RC_2606_0 ( .a(n_20745), .b(n_21068), .c(n_20744), .d(n_21067), .o(n_21218) );
oa22f04 FE_RC_2607_0 ( .a(n_45066), .b(FE_OCP_RBN5971_n_20510), .c(n_20510), .d(n_45101), .o(n_20650) );
na02m06 FE_RC_2613_0 ( .a(n_20628), .b(n_20997), .o(FE_RN_1146_0) );
na02m08 FE_RC_2614_0 ( .a(FE_RN_1146_0), .b(FE_OCP_RBN6803_n_20565), .o(n_21149) );
ao22m02 FE_RC_2615_0 ( .a(n_45024), .b(FE_OCP_RBN3211_n_21203), .c(n_45023), .d(n_21203), .o(n_21390) );
ao22f04 FE_RC_2616_0 ( .a(n_14452), .b(FE_OCP_RBN3202_n_15900), .c(n_14419), .d(n_15900), .o(n_16074) );
na02m08 TIMEBOOST_cell_4254 ( .a(TIMEBOOST_net_1217), .b(n_13436), .o(n_13529) );
na02s02 TIMEBOOST_cell_4091 ( .a(n_31021), .b(n_27518), .o(TIMEBOOST_net_1136) );
in01s01 FE_RC_2619_0 ( .a(FE_OCP_RBN2744_n_14114), .o(FE_RN_1149_0) );
oa22f02 FE_RC_2622_0 ( .a(n_45010), .b(FE_OCP_RBN3718_n_20621), .c(n_45012), .d(n_20621), .o(n_20771) );
in01m04 FE_RC_2623_0 ( .a(FE_RN_1151_0), .o(n_16333) );
no02s02 FE_RC_2627_0 ( .a(FE_OCPN1733_n_14524), .b(n_16197), .o(FE_RN_1152_0) );
no02s06 FE_RC_2628_0 ( .a(FE_RN_1152_0), .b(n_16446), .o(n_16495) );
no02s01 FE_RC_2631_0 ( .a(n_19461), .b(n_20429), .o(FE_RN_1154_0) );
in01s01 FE_RC_2632_0 ( .a(n_19461), .o(FE_RN_1155_0) );
no02s02 FE_RC_2633_0 ( .a(FE_RN_1155_0), .b(FE_OCP_RBN4351_n_20456), .o(FE_RN_1156_0) );
no02s02 FE_RC_2634_0 ( .a(FE_RN_1154_0), .b(FE_RN_1156_0), .o(n_20672) );
in01s01 FE_RC_2637_0 ( .a(FE_OCP_DRV_N5161_n_30322), .o(FE_RN_1158_0) );
na02s06 FE_RC_2638_0 ( .a(n_31476), .b(FE_RN_1158_0), .o(n_31501) );
na02s02 TIMEBOOST_cell_5035 ( .a(TIMEBOOST_net_1465), .b(FE_OCP_RBN4133_n_38028), .o(n_38201) );
no02m02 FE_RC_2642_0 ( .a(n_25401), .b(n_25358), .o(FE_RN_1161_0) );
na02m02 FE_RC_2643_0 ( .a(n_25635), .b(n_25399), .o(FE_RN_1162_0) );
na02f04 FE_RC_2644_0 ( .a(FE_RN_1162_0), .b(FE_RN_1161_0), .o(n_25702) );
na02s04 FE_RC_2645_0 ( .a(n_31502), .b(n_31475), .o(FE_RN_1163_0) );
na02s08 FE_RC_2646_0 ( .a(n_31520), .b(FE_RN_1163_0), .o(FE_RN_1164_0) );
na02s10 FE_RC_2647_0 ( .a(FE_RN_1164_0), .b(n_31548), .o(n_31746) );
na02s01 FE_RC_2648_0 ( .a(n_30224), .b(n_30324), .o(FE_RN_1165_0) );
na02s06 FE_RC_2649_0 ( .a(n_31466), .b(FE_RN_1165_0), .o(n_31751) );
in01m02 FE_RC_264_0 ( .a(n_22560), .o(FE_RN_82_0) );
na02s01 TIMEBOOST_cell_3139 ( .a(n_35717), .b(TIMEBOOST_net_860), .o(n_35853) );
na02s01 TIMEBOOST_cell_3140 ( .a(n_35884), .b(FE_OCP_RBN3299_n_35539), .o(TIMEBOOST_net_861) );
no02m10 FE_RC_2657_0 ( .a(n_25732), .b(FE_RN_1171_0), .o(n_25786) );
in01m04 FE_RC_265_0 ( .a(FE_RN_83_0), .o(n_22632) );
no02s03 FE_RC_2660_0 ( .a(n_20891), .b(n_20526), .o(FE_RN_1172_0) );
ao12m04 FE_RC_2661_0 ( .a(FE_RN_1172_0), .b(n_20526), .c(n_20891), .o(n_21004) );
no02m02 FE_RC_2662_0 ( .a(n_30890), .b(n_30887), .o(FE_RN_1173_0) );
na02f06 FE_RC_2663_0 ( .a(n_31061), .b(FE_RN_1173_0), .o(n_31058) );
no02s02 TIMEBOOST_cell_8857 ( .a(TIMEBOOST_net_2915), .b(n_17117), .o(n_17313) );
na02m06 TIMEBOOST_cell_8627 ( .a(TIMEBOOST_net_2800), .b(n_10719), .o(n_46989) );
na02m06 TIMEBOOST_cell_5036 ( .a(FE_OCP_RBN5703_n_19663), .b(FE_OCPN1727_n_18099), .o(TIMEBOOST_net_1466) );
in01f02 FE_RC_2672_0 ( .a(n_16466), .o(FE_RN_1179_0) );
in01s02 FE_RC_2673_0 ( .a(n_16567), .o(FE_RN_1180_0) );
na02f06 TIMEBOOST_cell_5543 ( .a(TIMEBOOST_net_1719), .b(n_36652), .o(n_36715) );
no03s04 TIMEBOOST_cell_5782 ( .a(n_9495), .b(FE_OCP_RBN2887_n_9492), .c(FE_RN_2220_0), .o(FE_RN_1013_0) );
no02m04 TIMEBOOST_cell_7753 ( .a(TIMEBOOST_net_2507), .b(n_9299), .o(n_9514) );
in01f04 FE_RC_2677_0 ( .a(n_21603), .o(FE_RN_1183_0) );
no03f06 TIMEBOOST_cell_4636 ( .a(n_24263), .b(n_24246), .c(FE_OCP_RBN6623_n_24175), .o(n_24362) );
in01s01 FE_RC_2680_0 ( .a(n_23486), .o(FE_RN_1185_0) );
na02f04 FE_RC_2689_0 ( .a(FE_OCP_RBN2086_n_14911), .b(n_16622), .o(FE_RN_1190_0) );
oa22f06 FE_RC_2690_0 ( .a(n_30766), .b(n_30864), .c(n_30767), .d(n_30863), .o(n_31013) );
in01m02 FE_RC_2691_0 ( .a(n_26872), .o(FE_RN_1191_0) );
no02m06 FE_RC_2692_0 ( .a(n_26824), .b(FE_RN_1191_0), .o(FE_RN_555_0) );
no02f04 FE_RC_2693_0 ( .a(n_30944), .b(n_30703), .o(FE_RN_1192_0) );
na02m04 FE_RC_2694_0 ( .a(n_30944), .b(n_30703), .o(FE_RN_1193_0) );
ao12f04 FE_RC_2695_0 ( .a(FE_RN_1192_0), .b(FE_RN_1193_0), .c(n_30862), .o(n_31003) );
in01f02 FE_RC_2696_0 ( .a(n_15175), .o(FE_RN_1194_0) );
in01f02 FE_RC_2697_0 ( .a(n_15231), .o(FE_RN_1195_0) );
oa22f04 FE_RC_2698_0 ( .a(FE_RN_1194_0), .b(n_15231), .c(n_15175), .d(FE_RN_1195_0), .o(n_15459) );
no02f04 FE_RC_2700_0 ( .a(n_21736), .b(FE_OCP_RBN3361_n_21847), .o(FE_RN_1197_0) );
na02s01 TIMEBOOST_cell_1237 ( .a(FE_RN_1330_0), .b(FE_OCPN1610_n_23503), .o(TIMEBOOST_net_233) );
na02s01 TIMEBOOST_cell_1238 ( .a(TIMEBOOST_net_233), .b(FE_RN_1329_0), .o(FE_RN_1334_0) );
na02m02 TIMEBOOST_cell_6100 ( .a(TIMEBOOST_net_1901), .b(n_8951), .o(TIMEBOOST_net_1535) );
oa22f02 FE_RC_2712_0 ( .a(n_32287), .b(n_32311), .c(FE_OFN621_n_28336), .d(n_32286), .o(n_32352) );
oa22f02 FE_RC_2713_0 ( .a(n_32287), .b(FE_OCP_RBN3421_n_32254), .c(FE_OFN621_n_28336), .d(n_32254), .o(n_32304) );
oa22s02 FE_RC_2716_0 ( .a(n_32566), .b(n_32310), .c(FE_OFN621_n_28336), .d(n_32285), .o(n_32353) );
oa22m06 FE_RC_2718_0 ( .a(n_31825), .b(n_32172), .c(n_31826), .d(n_32195), .o(n_32290) );
oa22s02 FE_RC_2719_0 ( .a(n_32287), .b(n_32339), .c(FE_OFN621_n_28336), .d(n_44434), .o(n_32370) );
in01f04 FE_RC_271_0 ( .a(n_24099), .o(FE_RN_85_0) );
oa22m02 FE_RC_2720_0 ( .a(n_24059), .b(n_27655), .c(n_27845), .d(n_27641), .o(n_27700) );
in01s01 FE_RC_2721_0 ( .a(n_26797), .o(FE_RN_1203_0) );
no02s04 FE_RC_2722_0 ( .a(n_26920), .b(FE_RN_1203_0), .o(n_26879) );
oa22s02 FE_RC_2723_0 ( .a(FE_OFN1183_n_24059), .b(n_27720), .c(n_27796), .d(n_27698), .o(n_27741) );
oa22s01 FE_RC_2724_0 ( .a(n_24350), .b(n_27739), .c(n_27796), .d(n_27730), .o(n_27779) );
in01m02 FE_RC_2725_0 ( .a(n_31025), .o(FE_RN_1204_0) );
na02m04 FE_RC_2726_0 ( .a(n_31050), .b(FE_RN_1204_0), .o(n_31070) );
in01s02 FE_RC_2729_0 ( .a(n_21240), .o(FE_RN_1205_0) );
in01f04 FE_RC_272_0 ( .a(FE_RN_86_0), .o(n_24269) );
no02m04 FE_RC_2730_0 ( .a(n_21399), .b(FE_RN_1205_0), .o(n_21442) );
ao22f06 FE_RC_2731_0 ( .a(n_30799), .b(n_31046), .c(n_31045), .d(n_31122), .o(n_31148) );
in01s01 FE_RC_2732_0 ( .a(n_22793), .o(FE_RN_1206_0) );
na02f02 FE_RC_2733_0 ( .a(n_22750), .b(FE_RN_1206_0), .o(FE_RN_1207_0) );
oa12f02 FE_RC_2734_0 ( .a(FE_RN_1207_0), .b(FE_OCPN1394_n_22801), .c(n_22750), .o(n_22794) );
oa22f02 FE_RC_2735_0 ( .a(n_14901), .b(n_14881), .c(FE_OCP_RBN4315_n_14881), .d(n_14902), .o(n_15001) );
ao22f04 FE_RC_2737_0 ( .a(n_32101), .b(n_32296), .c(n_32102), .d(n_32300), .o(n_32380) );
no03s02 TIMEBOOST_cell_8240 ( .a(n_2503), .b(n_2504), .c(n_3222), .o(TIMEBOOST_net_2090) );
no02f04 FE_RC_2740_0 ( .a(n_26369), .b(FE_OCPN5290_n_26125), .o(FE_RN_1209_0) );
na02f04 FE_RC_2741_0 ( .a(n_26369), .b(n_26125), .o(FE_RN_1210_0) );
ao12f04 FE_RC_2742_0 ( .a(FE_RN_1209_0), .b(FE_RN_1210_0), .c(n_26267), .o(n_26412) );
na02s01 FE_RC_2746_0 ( .a(n_26171), .b(n_27222), .o(FE_RN_1213_0) );
na02s01 FE_RC_2747_0 ( .a(n_27204), .b(FE_RN_1213_0), .o(n_27400) );
no02s02 TIMEBOOST_cell_1601 ( .a(FE_OCPN1244_n_13992), .b(n_15103), .o(TIMEBOOST_net_415) );
in01s02 FE_RC_275_0 ( .a(n_24182), .o(FE_RN_87_0) );
no02s04 TIMEBOOST_cell_1618 ( .a(n_34714), .b(TIMEBOOST_net_423), .o(n_34729) );
oa22f04 FE_RC_2762_0 ( .a(n_7769), .b(FE_RN_866_0), .c(n_7767), .d(n_8093), .o(FE_RN_867_0) );
oa22f04 FE_RC_2765_0 ( .a(n_19738), .b(n_19920), .c(n_19737), .d(n_19890), .o(n_20020) );
oa22s02 FE_RC_2767_0 ( .a(FE_RN_1220_0), .b(FE_OCP_RBN5527_n_6760), .c(n_6760), .d(FE_RN_1221_0), .o(n_6874) );
in01s01 FE_RC_2768_0 ( .a(n_6601), .o(FE_RN_1221_0) );
in01s01 FE_RC_2769_0 ( .a(FE_RN_1221_0), .o(FE_RN_1220_0) );
in01s02 FE_RC_276_0 ( .a(n_23772), .o(FE_RN_88_0) );
oa22s01 FE_RC_2770_0 ( .a(n_1188), .b(n_44652), .c(n_1186), .d(n_44637), .o(n_1329) );
oa22s01 FE_RC_2771_0 ( .a(n_1142), .b(n_44652), .c(n_1130), .d(n_44661), .o(n_1299) );
oa22m04 FE_RC_2773_0 ( .a(n_8534), .b(n_8366), .c(FE_OCPN3568_n_8348), .d(n_8533), .o(n_8677) );
oa22f02 FE_RC_2774_0 ( .a(FE_OCP_RBN2751_FE_RN_1223_0), .b(FE_OCP_RBN2797_n_8530), .c(n_8530), .d(FE_OCP_RBN2719_n_8242), .o(n_8580) );
in01s01 FE_RC_2775_0 ( .a(FE_OCP_RBN2717_n_8242), .o(FE_RN_1223_0) );
oa22m04 FE_RC_2777_0 ( .a(n_10263), .b(n_10441), .c(n_10440), .d(n_10262), .o(n_10570) );
na02s06 FE_RC_277_0 ( .a(FE_RN_87_0), .b(FE_RN_88_0), .o(FE_RN_89_0) );
oa22m04 FE_RC_2780_0 ( .a(n_10521), .b(n_10946), .c(n_10522), .d(FE_OCP_RBN6094_n_10946), .o(n_11087) );
na03m06 FE_RC_2782_0 ( .a(n_11076), .b(n_11195), .c(n_11110), .o(n_11196) );
ao22s04 FE_RC_2783_0 ( .a(n_7589), .b(n_9011), .c(n_7588), .d(n_9010), .o(n_9188) );
oa22s02 FE_RC_2784_0 ( .a(n_7693), .b(FE_OCPN6919_n_7726), .c(n_7725), .d(n_7675), .o(n_7747) );
oa22m04 FE_RC_2786_0 ( .a(n_8806), .b(n_8815), .c(n_8825), .d(FE_OCP_RBN2885_n_8806), .o(n_8981) );
ao22m02 FE_RC_2788_0 ( .a(n_9764), .b(FE_OCP_RBN2970_n_9676), .c(n_9676), .d(n_9712), .o(n_9904) );
ao22m02 FE_RC_2789_0 ( .a(n_44575), .b(FE_OCP_RBN2937_n_8981), .c(FE_OCP_RBN5834_n_44563), .d(n_8981), .o(n_9102) );
ao22s02 FE_RC_2791_0 ( .a(n_44355), .b(FE_OCP_RBN6225_n_11713), .c(n_11713), .d(n_44354), .o(n_12058) );
oa22f04 FE_RC_2793_0 ( .a(FE_OCP_RBN7033_n_18981), .b(n_19249), .c(FE_OCP_RBN7034_n_18981), .d(n_19271), .o(n_19437) );
oa22s02 FE_RC_2794_0 ( .a(n_7764), .b(n_8942), .c(n_7765), .d(n_8941), .o(n_9090) );
ao22m02 FE_RC_2795_0 ( .a(n_9083), .b(n_8967), .c(n_9084), .d(n_8966), .o(n_9292) );
oa22m04 FE_RC_2796_0 ( .a(FE_OCP_RBN4270_n_8872), .b(n_8998), .c(FE_OCP_RBN5904_n_8872), .d(n_8999), .o(n_9182) );
in01s01 FE_RC_2797_0 ( .a(FE_OFN4768_n_8309), .o(FE_RN_1224_0) );
in01s02 FE_RC_2798_0 ( .a(n_9271), .o(FE_RN_1225_0) );
na02s04 FE_RC_2799_0 ( .a(FE_RN_1225_0), .b(FE_RN_1224_0), .o(FE_RN_1226_0) );
na02m06 FE_RC_2800_0 ( .a(n_9261), .b(FE_RN_1226_0), .o(n_9362) );
oa22m04 FE_RC_2801_0 ( .a(n_9718), .b(FE_OCP_RBN5969_n_9668), .c(n_9668), .d(n_9719), .o(n_9859) );
in01f04 FE_RC_2803_0 ( .a(n_9293), .o(FE_RN_1227_0) );
in01m02 FE_RC_2804_0 ( .a(n_9170), .o(FE_RN_1228_0) );
no02m08 FE_RC_2805_0 ( .a(FE_RN_1227_0), .b(FE_RN_1228_0), .o(FE_RN_1229_0) );
ao12m08 FE_RC_2806_0 ( .a(FE_RN_1229_0), .b(n_9215), .c(FE_OCP_RBN5945_FE_RN_1231_0), .o(n_9494) );
in01m02 FE_RC_2807_0 ( .a(n_9242), .o(FE_RN_1231_0) );
ao22m04 FE_RC_2809_0 ( .a(FE_OCP_RBN4305_n_44579), .b(n_9584), .c(FE_OCP_RBN5930_n_44563), .d(FE_OCP_RBN3028_n_9584), .o(n_9747) );
in01s02 FE_RC_2811_0 ( .a(FE_RN_574_0), .o(FE_RN_1232_0) );
in01s02 FE_RC_2812_0 ( .a(n_20973), .o(FE_RN_1233_0) );
na02m04 FE_RC_2813_0 ( .a(FE_RN_1232_0), .b(FE_RN_1233_0), .o(FE_RN_1234_0) );
na02s04 TIMEBOOST_cell_8850 ( .a(n_10014), .b(FE_OCP_RBN6814_n_9893), .o(TIMEBOOST_net_2912) );
ao22m02 FE_RC_2816_0 ( .a(n_9701), .b(n_9714), .c(n_9713), .d(n_9660), .o(n_9892) );
in01s01 TIMEBOOST_cell_5904 ( .a(TIMEBOOST_net_1792), .o(TIMEBOOST_net_1793) );
ao22m04 FE_RC_281_0 ( .a(n_24010), .b(n_24399), .c(n_24398), .d(n_24009), .o(n_24501) );
in01m02 FE_RC_2821_0 ( .a(n_21535), .o(FE_RN_1236_0) );
na02m04 FE_RC_2822_0 ( .a(FE_OCP_RBN3244_n_21269), .b(FE_RN_1236_0), .o(FE_RN_1237_0) );
na02m04 FE_RC_2823_0 ( .a(FE_RN_1237_0), .b(n_21576), .o(n_46966) );
ao22f02 FE_RC_2824_0 ( .a(n_21273), .b(n_21464), .c(n_21272), .d(n_21420), .o(n_21640) );
oa22f06 FE_RC_2825_0 ( .a(n_21306), .b(FE_OCP_RBN5340_n_21261), .c(n_21261), .d(n_21307), .o(n_21494) );
oa22f04 FE_RC_2827_0 ( .a(n_22381), .b(n_22518), .c(n_22382), .d(n_22538), .o(n_22640) );
oa22f02 FE_RC_2828_0 ( .a(n_22961), .b(n_46965), .c(n_22580), .d(n_22594), .o(n_22671) );
no03m08 TIMEBOOST_cell_8233 ( .a(n_29533), .b(n_29502), .c(n_29630), .o(TIMEBOOST_net_1505) );
ao22f02 FE_RC_2831_0 ( .a(n_21619), .b(n_21686), .c(n_21588), .d(n_21710), .o(n_21816) );
oa22s02 FE_RC_2833_0 ( .a(FE_OFN787_n_46285), .b(n_12144), .c(FE_OCP_RBN3352_FE_OFN760_n_46337), .d(n_12112), .o(n_46351) );
oa22s02 FE_RC_2834_0 ( .a(FE_OFN787_n_46285), .b(n_12150), .c(FE_OCP_RBN3352_FE_OFN760_n_46337), .d(n_12058), .o(n_46356) );
oa22s04 FE_RC_2836_0 ( .a(n_11922), .b(n_11799), .c(n_11800), .d(n_11923), .o(n_12068) );
ao22m02 FE_RC_2838_0 ( .a(FE_OCP_RBN3426_n_11810), .b(n_11870), .c(n_11810), .d(n_11850), .o(n_12060) );
ao22m02 FE_RC_283_0 ( .a(n_22089), .b(FE_OCP_RBN2712_n_24501), .c(n_22280), .d(n_24501), .o(n_24618) );
oa22s02 FE_RC_2840_0 ( .a(FE_OCPN1394_n_22801), .b(n_22718), .c(n_22833), .d(FE_OCP_RBN6238_n_22718), .o(n_22777) );
oa22f02 FE_RC_2841_0 ( .a(n_22961), .b(n_22635), .c(n_22580), .d(n_22614), .o(n_22712) );
oa22f08 FE_RC_2847_0 ( .a(n_40643), .b(n_40659), .c(n_40664), .d(n_40644), .o(n_40715) );
ao22m04 FE_RC_284_0 ( .a(n_24327), .b(FE_OCPN1368_n_23923), .c(n_23924), .d(n_24348), .o(n_24451) );
in01s06 FE_RC_2853_0 ( .a(n_40732), .o(FE_RN_1244_0) );
in01f04 FE_RC_2854_0 ( .a(n_40743), .o(FE_RN_1245_0) );
no02f08 FE_RC_2855_0 ( .a(FE_RN_1244_0), .b(FE_RN_1245_0), .o(FE_RN_1246_0) );
no03s20 TIMEBOOST_cell_5698 ( .a(n_32706), .b(n_32440), .c(FE_OCP_RBN7010_n_44962), .o(n_32597) );
in01s01 FE_RC_2857_0 ( .a(n_40572), .o(FE_RN_1247_0) );
in01m02 FE_RC_2858_0 ( .a(n_40822), .o(FE_RN_1248_0) );
no02m04 FE_RC_2859_0 ( .a(FE_RN_1247_0), .b(FE_RN_1248_0), .o(FE_RN_1249_0) );
no02m06 FE_RC_2860_0 ( .a(FE_OCP_RBN2441_n_44798), .b(FE_RN_1249_0), .o(n_40963) );
in01s01 TIMEBOOST_cell_8912 ( .a(n_1299), .o(TIMEBOOST_net_2956) );
no02f10 TIMEBOOST_cell_1750 ( .a(n_39293), .b(TIMEBOOST_net_489), .o(n_39450) );
no02m04 TIMEBOOST_cell_1817 ( .a(n_16233), .b(n_16236), .o(TIMEBOOST_net_523) );
ao22f04 FE_RC_2864_0 ( .a(n_42166), .b(n_42157), .c(n_42156), .d(n_42173), .o(n_42179) );
ao22f04 FE_RC_2865_0 ( .a(n_42178), .b(n_42176), .c(n_42175), .d(n_42177), .o(n_42194) );
ao22s02 FE_RC_2866_0 ( .a(n_43617), .b(FE_OCP_RBN3412_n_43829), .c(n_43618), .d(n_43829), .o(n_43864) );
ao22s02 FE_RC_2867_0 ( .a(n_43258), .b(n_43765), .c(n_43259), .d(n_43764), .o(n_43815) );
ao22s02 FE_RC_2868_0 ( .a(n_43348), .b(n_43782), .c(n_43347), .d(n_43781), .o(n_43839) );
ao22f02 FE_RC_2869_0 ( .a(n_43609), .b(n_43893), .c(n_43610), .d(n_43892), .o(n_43911) );
ao22f02 FE_RC_2870_0 ( .a(n_43534), .b(FE_OCP_RBN3431_n_43880), .c(n_43533), .d(n_43880), .o(n_43907) );
ao22f02 FE_RC_2871_0 ( .a(n_43428), .b(n_43877), .c(n_43427), .d(n_43876), .o(n_43901) );
ao22f02 FE_RC_2872_0 ( .a(n_43559), .b(n_43872), .c(n_43871), .d(n_43558), .o(n_43900) );
ao22m02 FE_RC_2873_0 ( .a(n_43834), .b(n_43463), .c(n_43462), .d(n_43819), .o(n_43878) );
ao22s02 FE_RC_2874_0 ( .a(n_43635), .b(n_43842), .c(n_43634), .d(FE_OCP_RBN6257_n_43842), .o(n_43866) );
ao22m08 FE_RC_2878_0 ( .a(n_11816), .b(n_47212), .c(n_11815), .d(n_47213), .o(n_12261) );
oa22m04 FE_RC_2880_0 ( .a(FE_RN_1250_0), .b(n_31001), .c(n_30368), .d(FE_OCP_RBN3175_n_31001), .o(n_31107) );
in01s01 FE_RC_2881_0 ( .a(n_30367), .o(FE_RN_1251_0) );
in01s01 FE_RC_2882_0 ( .a(FE_RN_1251_0), .o(FE_RN_1250_0) );
oa22f02 FE_RC_2883_0 ( .a(FE_OFN1183_n_24059), .b(n_27686), .c(n_27845), .d(n_27662), .o(n_27725) );
na02s01 TIMEBOOST_cell_8768 ( .a(FE_OCP_RBN2757_n_13796), .b(FE_OCP_RBN6694_n_13796), .o(TIMEBOOST_net_2871) );
oa22m01 FE_RC_2889_0 ( .a(n_36846), .b(n_36723), .c(n_36722), .d(n_36889), .o(n_36890) );
in01s20 FE_RC_2890_0 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_12_), .o(FE_RN_1255_0) );
in01s03 FE_RC_2891_0 ( .a(FE_OCP_RBN6540_n_44083), .o(FE_RN_1256_0) );
no02f02 TIMEBOOST_cell_1735 ( .a(n_26139), .b(n_23414), .o(TIMEBOOST_net_482) );
no02s02 TIMEBOOST_cell_1737 ( .a(n_26240), .b(n_23564), .o(TIMEBOOST_net_483) );
na03m10 TIMEBOOST_cell_2157 ( .a(n_36931), .b(n_36917), .c(n_36932), .o(n_37033) );
ao22m08 FE_RC_2896_0 ( .a(FE_OCP_RBN6525_n_11829), .b(n_11819), .c(n_11829), .d(n_11881), .o(n_11978) );
in01m10 FE_RC_2897_0 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_7_), .o(FE_RN_1258_0) );
in01s03 FE_RC_2898_0 ( .a(FE_OCP_RBN5529_n_44061), .o(FE_RN_1259_0) );
na02s02 TIMEBOOST_cell_8526 ( .a(n_13440), .b(n_14024), .o(TIMEBOOST_net_2750) );
ao22f06 FE_RC_289_0 ( .a(FE_OCP_RBN2709_n_24505), .b(n_25017), .c(n_25104), .d(n_25016), .o(n_25127) );
ao22f04 FE_RC_2904_0 ( .a(n_12688), .b(n_12527), .c(n_12526), .d(n_12689), .o(n_12800) );
ao22f04 FE_RC_290_0 ( .a(n_24868), .b(n_25071), .c(n_24869), .d(n_25072), .o(n_25149) );
oa22m10 FE_RC_2912_0 ( .a(n_32664), .b(FE_OCP_RBN7018_n_32649), .c(n_32663), .d(n_32649), .o(n_32773) );
oa22f08 FE_RC_2917_0 ( .a(n_22945), .b(n_22966), .c(n_22965), .d(n_22900), .o(n_23069) );
ao22m10 FE_RC_2918_0 ( .a(n_32625), .b(n_32473), .c(n_32596), .d(n_32472), .o(n_32667) );
ao22f04 FE_RC_2923_0 ( .a(n_28572), .b(n_28951), .c(n_28573), .d(n_28950), .o(n_29033) );
ao22m08 FE_RC_2930_0 ( .a(n_44061), .b(FE_OCP_RBN2270_delay_xor_ln22_unr15_stage6_stallmux_q_2_), .c(delay_xor_ln22_unr15_stage6_stallmux_q_2_), .d(FE_OCP_RBN6466_n_44061), .o(n_22771) );
oa22m04 FE_RC_2935_0 ( .a(n_22458), .b(n_22745), .c(n_22457), .d(n_22707), .o(n_22901) );
in01s01 FE_RC_2938_0 ( .a(n_23823), .o(FE_RN_1267_0) );
in01s04 FE_RC_2939_0 ( .a(FE_RN_89_0), .o(FE_RN_1268_0) );
na02m08 FE_RC_2940_0 ( .a(FE_RN_1268_0), .b(FE_RN_1267_0), .o(FE_RN_1269_0) );
na02s02 TIMEBOOST_cell_8763 ( .a(TIMEBOOST_net_2868), .b(n_14362), .o(TIMEBOOST_net_2444) );
oa22s06 FE_RC_2943_0 ( .a(n_23787), .b(n_24148), .c(n_23786), .d(n_24166), .o(n_24254) );
oa22f04 FE_RC_2949_0 ( .a(n_35201), .b(n_35475), .c(n_35228), .d(n_35443), .o(n_35505) );
oa22m04 FE_RC_294_0 ( .a(FE_OCP_RBN2665_n_24372), .b(n_24787), .c(n_24529), .d(n_24836), .o(n_24944) );
oa22f04 FE_RC_2951_0 ( .a(n_14722), .b(n_14665), .c(n_14693), .d(FE_OCP_RBN5823_n_14722), .o(n_14823) );
oa22f06 FE_RC_2953_0 ( .a(n_25831), .b(n_25816), .c(FE_OCP_RBN3076_n_25816), .d(n_25829), .o(n_25912) );
in01m02 FE_RC_2956_0 ( .a(n_36069), .o(FE_RN_1271_0) );
in01s02 FE_RC_2957_0 ( .a(FE_RN_1271_0), .o(FE_RN_1270_0) );
oa22m02 FE_RC_2959_0 ( .a(n_15076), .b(n_15164), .c(n_15075), .d(n_15163), .o(n_15319) );
na03m08 FE_RC_2964_0 ( .a(n_15410), .b(FE_OCP_RBN3015_n_15300), .c(n_15407), .o(n_15492) );
in01f02 FE_RC_2966_0 ( .a(n_26555), .o(FE_RN_1273_0) );
no02f04 FE_RC_2967_0 ( .a(n_26394), .b(FE_RN_1273_0), .o(FE_RN_1274_0) );
no03s10 TIMEBOOST_cell_3424 ( .a(n_1427), .b(n_1435), .c(n_1494), .o(n_1513) );
na02f02 TIMEBOOST_cell_1900 ( .a(TIMEBOOST_net_564), .b(n_5842), .o(FE_RN_2273_0) );
in01s01 FE_RC_296_0 ( .a(n_24502), .o(FE_RN_90_0) );
in01s01 FE_RC_2971_0 ( .a(FE_RN_1149_0), .o(FE_RN_1275_0) );
in01s01 FE_RC_2972_0 ( .a(FE_OCP_RBN6802_n_15156), .o(FE_RN_1276_0) );
na02f03 TIMEBOOST_cell_5255 ( .a(TIMEBOOST_net_1575), .b(n_3530), .o(n_3674) );
na02s03 TIMEBOOST_cell_3080 ( .a(n_8108), .b(FE_OCP_RBN4162_FE_OCPN857_n_7802), .o(TIMEBOOST_net_831) );
oa22m02 FE_RC_2975_0 ( .a(n_36657), .b(FE_OCP_RBN6229_n_36693), .c(n_36631), .d(n_36693), .o(n_36741) );
in01s02 FE_RC_2981_0 ( .a(n_30882), .o(FE_RN_1279_0) );
na03s02 TIMEBOOST_cell_8384 ( .a(n_4831), .b(n_4515), .c(n_4876), .o(n_5063) );
na02f04 TIMEBOOST_cell_5627 ( .a(TIMEBOOST_net_1761), .b(n_16826), .o(n_17128) );
ao22f04 FE_RC_2984_0 ( .a(n_25935), .b(n_45329), .c(n_25919), .d(n_25964), .o(n_26085) );
oa22s04 FE_RC_2985_0 ( .a(n_27521), .b(n_27670), .c(n_27522), .d(n_27690), .o(n_27782) );
ao22m02 FE_RC_2987_0 ( .a(n_26276), .b(n_23414), .c(n_23466), .d(FE_OCP_RBN3252_n_26276), .o(n_26424) );
oa22s02 FE_RC_2989_0 ( .a(n_32566), .b(n_32305), .c(FE_OFN621_n_28336), .d(FE_OCP_RBN6243_n_32305), .o(n_32350) );
no02s01 TIMEBOOST_cell_6151 ( .a(FE_OCP_RBN2837_n_13962), .b(FE_OCP_RBN5800_n_13962), .o(TIMEBOOST_net_1927) );
ao22m06 FE_RC_2990_0 ( .a(n_31800), .b(n_45518), .c(n_31801), .d(n_45516), .o(n_32266) );
ao22m02 FE_RC_2991_0 ( .a(n_47187), .b(n_21578), .c(n_21543), .d(n_47186), .o(n_21791) );
oa22s02 FE_RC_2993_0 ( .a(n_27520), .b(n_27674), .c(n_27519), .d(n_27696), .o(n_27784) );
oa22s02 FE_RC_2998_0 ( .a(n_22961), .b(n_22789), .c(n_22580), .d(n_22739), .o(n_22815) );
na02s06 TIMEBOOST_cell_2862 ( .a(n_37351), .b(n_37101), .o(TIMEBOOST_net_722) );
oa22s01 FE_RC_3004_0 ( .a(n_17584), .b(n_17687), .c(n_16339), .d(n_17649), .o(n_17752) );
oa22f02 FE_RC_3006_0 ( .a(n_28336), .b(n_32358), .c(n_32287), .d(n_32384), .o(n_32431) );
ao22s04 FE_RC_3008_0 ( .a(n_32057), .b(n_32324), .c(n_32058), .d(n_32343), .o(n_32427) );
oa22f02 FE_RC_3010_0 ( .a(n_28336), .b(n_32394), .c(n_32566), .d(n_32463), .o(n_32511) );
na02m01 TIMEBOOST_cell_1459 ( .a(n_33785), .b(n_33733), .o(TIMEBOOST_net_344) );
in01s02 FE_RC_3012_0 ( .a(n_27438), .o(FE_RN_1282_0) );
na02m02 TIMEBOOST_cell_1460 ( .a(TIMEBOOST_net_344), .b(n_33833), .o(n_33906) );
oa22m02 FE_RC_3015_0 ( .a(FE_OFN1183_n_24059), .b(n_27727), .c(n_27796), .d(n_27705), .o(n_27749) );
in01s01 FE_RC_3017_0 ( .a(n_27146), .o(FE_RN_1284_0) );
in01s03 FE_RC_3018_0 ( .a(n_27568), .o(FE_RN_1285_0) );
no02m02 TIMEBOOST_cell_1463 ( .a(n_33717), .b(FE_OCP_RBN2570_n_33735), .o(TIMEBOOST_net_346) );
in01m01 FE_RC_301_0 ( .a(n_25479), .o(FE_RN_93_0) );
no02s04 TIMEBOOST_cell_1464 ( .a(TIMEBOOST_net_346), .b(FE_OCP_RBN4913_n_33833), .o(n_33882) );
no02m06 TIMEBOOST_cell_1569 ( .a(FE_OCP_RBN4137_n_7743), .b(n_8258), .o(TIMEBOOST_net_399) );
in01s01 FE_RC_3025_0 ( .a(FE_RN_469_0), .o(FE_RN_1287_0) );
in01f02 FE_RC_3026_0 ( .a(n_29034), .o(FE_RN_1288_0) );
no02f06 FE_RC_3027_0 ( .a(FE_RN_1288_0), .b(FE_RN_1287_0), .o(FE_RN_1289_0) );
in01s01 TIMEBOOST_cell_8892 ( .a(n_1206), .o(TIMEBOOST_net_2936) );
in01s02 FE_RC_3029_0 ( .a(FE_RN_456_0), .o(FE_RN_1290_0) );
in01s06 FE_RC_302_0 ( .a(n_25813), .o(FE_RN_94_0) );
in01m02 FE_RC_3030_0 ( .a(n_24139), .o(FE_RN_1291_0) );
no02m06 FE_RC_3031_0 ( .a(FE_RN_1290_0), .b(FE_RN_1291_0), .o(FE_RN_1292_0) );
no02m08 FE_RC_3032_0 ( .a(FE_RN_1292_0), .b(FE_RN_457_0), .o(n_24222) );
in01s02 FE_RC_3037_0 ( .a(n_45489), .o(FE_RN_1294_0) );
in01m02 FE_RC_3038_0 ( .a(FE_RN_1294_0), .o(FE_RN_1293_0) );
no02f06 TIMEBOOST_cell_4408 ( .a(TIMEBOOST_net_1294), .b(n_1222), .o(n_1230) );
oa22m04 FE_RC_3043_0 ( .a(n_20568), .b(n_21037), .c(FE_OCP_RBN4348_n_20568), .d(n_21002), .o(n_21203) );
ao22m04 FE_RC_3045_0 ( .a(n_26465), .b(n_26500), .c(n_26501), .d(n_26466), .o(n_26657) );
oa22s06 FE_RC_3047_0 ( .a(n_17377), .b(n_17660), .c(n_17376), .d(n_17695), .o(n_17835) );
ao22s04 FE_RC_3048_0 ( .a(n_27468), .b(n_27645), .c(n_27467), .d(n_27634), .o(n_27743) );
no02s01 TIMEBOOST_cell_6913 ( .a(n_23809), .b(n_23743), .o(TIMEBOOST_net_2215) );
in01s01 FE_RC_3050_0 ( .a(n_22501), .o(FE_RN_1296_0) );
in01s01 FE_RC_3051_0 ( .a(FE_RN_1296_0), .o(FE_RN_1295_0) );
no03s02 TIMEBOOST_cell_2158 ( .a(n_17104), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_11_), .c(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17210) );
na02m04 TIMEBOOST_cell_4054 ( .a(TIMEBOOST_net_1117), .b(n_25455), .o(FE_RN_1171_0) );
oa22f04 FE_RC_3058_0 ( .a(n_25426), .b(n_25702), .c(n_25396), .d(FE_OCP_RBN5995_n_25702), .o(n_25826) );
ao22f08 FE_RC_3059_0 ( .a(n_44441), .b(n_25785), .c(n_25507), .d(n_25818), .o(n_25915) );
no02m10 FE_RC_3062_0 ( .a(n_32554), .b(FE_OCP_RBN6532_n_32791), .o(FE_RN_1299_0) );
in01s08 FE_RC_3064_0 ( .a(FE_RN_47_0), .o(FE_RN_1300_0) );
in01s10 FE_RC_3065_0 ( .a(n_23388), .o(FE_RN_1301_0) );
na02s10 FE_RC_3066_0 ( .a(FE_RN_1300_0), .b(FE_RN_1301_0), .o(FE_RN_1302_0) );
no02m10 FE_RC_3067_0 ( .a(FE_OCP_RBN2462_n_23345), .b(FE_RN_1302_0), .o(n_47245) );
oa22s06 FE_RC_3068_0 ( .a(FE_RN_881_0), .b(FE_RN_880_0), .c(n_12038), .d(n_12039), .o(n_12232) );
ao22f06 FE_RC_306_0 ( .a(n_25903), .b(n_25534), .c(n_25533), .d(n_25902), .o(n_25999) );
in01m02 FE_RC_3071_0 ( .a(FE_OCPN1073_n_12638), .o(FE_RN_1303_0) );
in01m02 FE_RC_3072_0 ( .a(n_12983), .o(FE_RN_1304_0) );
no02m06 FE_RC_3073_0 ( .a(FE_RN_1303_0), .b(FE_RN_1304_0), .o(FE_RN_1305_0) );
no02f08 FE_RC_3074_0 ( .a(FE_RN_995_0), .b(FE_RN_1305_0), .o(n_13141) );
ao22f02 FE_RC_3077_0 ( .a(n_33267), .b(n_33687), .c(n_33268), .d(n_33688), .o(n_33771) );
in01s01 FE_RC_3079_0 ( .a(n_23759), .o(FE_RN_1307_0) );
ao22f06 FE_RC_307_0 ( .a(n_25824), .b(n_25893), .c(FE_OFN747_n_22641), .d(FE_OCP_RBN5196_n_25893), .o(n_25982) );
in01s01 FE_RC_3080_0 ( .a(FE_RN_1307_0), .o(FE_RN_1306_0) );
oa22m06 FE_RC_3081_0 ( .a(FE_RN_1308_0), .b(n_33773), .c(n_33322), .d(n_33807), .o(n_33872) );
in01s01 FE_RC_3082_0 ( .a(n_33321), .o(FE_RN_1309_0) );
in01s01 FE_RC_3083_0 ( .a(FE_RN_1309_0), .o(FE_RN_1308_0) );
in01s01 FE_RC_3089_0 ( .a(n_15635), .o(FE_RN_1310_0) );
oa22f04 FE_RC_308_0 ( .a(n_25478), .b(FE_OCP_RBN3106_n_25849), .c(n_25477), .d(n_25849), .o(n_25938) );
in01s02 FE_RC_3090_0 ( .a(n_15907), .o(FE_RN_1311_0) );
no02f06 TIMEBOOST_cell_8508 ( .a(n_29630), .b(n_29507), .o(TIMEBOOST_net_2741) );
no02f01 TIMEBOOST_cell_8666 ( .a(n_31079), .b(n_30987), .o(TIMEBOOST_net_2820) );
in01s01 FE_RC_3097_0 ( .a(n_30790), .o(FE_RN_1314_0) );
in01s01 FE_RC_3098_0 ( .a(FE_RN_1314_0), .o(FE_RN_1313_0) );
oa22f04 FE_RC_3099_0 ( .a(n_26493), .b(n_26849), .c(n_26848), .d(n_26494), .o(n_27010) );
oa22m02 FE_RC_3103_0 ( .a(n_17349), .b(n_17333), .c(n_17392), .d(n_17350), .o(n_17594) );
oa22f02 FE_RC_3105_0 ( .a(n_32287), .b(n_32428), .c(n_28336), .d(n_32380), .o(n_32467) );
oa22f02 FE_RC_3108_0 ( .a(FE_OFN1183_n_24059), .b(n_27714), .c(n_27845), .d(n_27683), .o(n_27737) );
oa22f02 FE_RC_3109_0 ( .a(FE_OFN1183_n_24059), .b(n_27726), .c(n_27796), .d(FE_OCP_RBN6259_n_27726), .o(n_27748) );
oa22m02 FE_RC_3110_0 ( .a(n_22907), .b(n_22829), .c(n_22580), .d(n_22800), .o(n_22908) );
na02f04 TIMEBOOST_cell_4508 ( .a(TIMEBOOST_net_1344), .b(n_6190), .o(n_6297) );
in01m01 FE_RC_3116_0 ( .a(n_23461), .o(FE_RN_1315_0) );
in01s06 FE_RC_3117_0 ( .a(n_23165), .o(FE_RN_1316_0) );
na02s06 FE_RC_3118_0 ( .a(FE_RN_1315_0), .b(FE_RN_1316_0), .o(FE_RN_1317_0) );
na02s02 TIMEBOOST_cell_4219 ( .a(n_12531), .b(n_12387), .o(TIMEBOOST_net_1200) );
no02f04 TIMEBOOST_cell_8780 ( .a(FE_OCP_RBN2981_n_14814), .b(FE_OCP_RBN2834_n_13962), .o(TIMEBOOST_net_2877) );
in01s01 FE_RC_3125_0 ( .a(n_12393), .o(FE_RN_1322_0) );
in01s02 FE_RC_3126_0 ( .a(FE_RN_1322_0), .o(FE_RN_1319_0) );
ao22m04 FE_RC_312_0 ( .a(n_26143), .b(n_25695), .c(n_26142), .d(n_25696), .o(n_26276) );
ao22m06 FE_RC_3136_0 ( .a(FE_RN_1323_0), .b(FE_OCP_RBN2667_n_24408), .c(n_23920), .d(n_24408), .o(n_24510) );
in01s01 FE_RC_3137_0 ( .a(n_23919), .o(FE_RN_1324_0) );
in01s01 FE_RC_3138_0 ( .a(FE_RN_1324_0), .o(FE_RN_1323_0) );
na03f06 TIMEBOOST_cell_8429 ( .a(n_6463), .b(n_6393), .c(n_6404), .o(n_6535) );
no02s01 TIMEBOOST_cell_1537 ( .a(n_45808), .b(n_754), .o(TIMEBOOST_net_383) );
in01m04 FE_RC_3147_0 ( .a(FE_RN_1327_0), .o(n_22556) );
no02s01 TIMEBOOST_cell_1538 ( .a(TIMEBOOST_net_383), .b(n_970), .o(n_45817) );
oa22f02 FE_RC_3149_0 ( .a(n_22961), .b(n_22903), .c(n_22833), .d(FE_OCP_RBN5351_n_22903), .o(n_22963) );
oa22m02 FE_RC_3153_0 ( .a(n_17584), .b(n_17594), .c(n_16339), .d(n_17565), .o(n_17654) );
oa22f10 FE_RC_3154_0 ( .a(n_27893), .b(FE_OCP_RBN5324_n_27885), .c(n_27859), .d(FE_OCP_RBN5323_n_27893), .o(n_28035) );
in01s01 FE_RC_3165_0 ( .a(FE_RN_1328_0), .o(n_23691) );
na02s01 FE_RC_3166_0 ( .a(FE_OCPN1610_n_23503), .b(FE_RN_1329_0), .o(n_23827) );
in01s01 FE_RC_3167_0 ( .a(n_23556), .o(FE_RN_1330_0) );
in01s01 FE_RC_3168_0 ( .a(n_23481), .o(FE_RN_1331_0) );
in01s01 FE_RC_3169_0 ( .a(n_23443), .o(FE_RN_1332_0) );
in01s01 FE_RC_3170_0 ( .a(n_23640), .o(FE_RN_1333_0) );
na02s01 FE_RC_3171_0 ( .a(FE_RN_1332_0), .b(FE_RN_1333_0), .o(FE_RN_1328_0) );
na02s01 FE_RC_3172_0 ( .a(FE_RN_1331_0), .b(FE_RN_1328_0), .o(FE_RN_1329_0) );
no02s02 TIMEBOOST_cell_1776 ( .a(TIMEBOOST_net_502), .b(n_43316), .o(n_43407) );
na02s01 FE_RC_3174_0 ( .a(n_23517), .b(FE_RN_1334_0), .o(n_23930) );
oa22s02 FE_RC_317_0 ( .a(n_27459), .b(n_45619), .c(n_27460), .d(n_27715), .o(n_27804) );
na02s02 FE_RC_3187_0 ( .a(n_37956), .b(n_37955), .o(FE_RN_1346_0) );
no02s06 FE_RC_3188_0 ( .a(FE_RN_1346_0), .b(n_38016), .o(FE_RN_1347_0) );
na02f08 FE_RC_3189_0 ( .a(n_38338), .b(FE_RN_1347_0), .o(n_38205) );
na02s01 FE_RC_3190_0 ( .a(n_41949), .b(n_41947), .o(FE_RN_1348_0) );
na02s01 FE_RC_3191_0 ( .a(FE_RN_1348_0), .b(n_42201), .o(FE_RN_1349_0) );
na02f08 FE_RC_3192_0 ( .a(n_42639), .b(FE_RN_1349_0), .o(n_42654) );
no02f08 FE_RC_3194_0 ( .a(n_42811), .b(FE_RN_1350_0), .o(n_42833) );
na03f40 FE_RC_3196_0 ( .a(n_40647), .b(n_40653), .c(n_40654), .o(n_40664) );
no02s01 TIMEBOOST_cell_1614 ( .a(TIMEBOOST_net_421), .b(n_2892), .o(n_4587) );
no02m08 TIMEBOOST_cell_5972 ( .a(TIMEBOOST_net_1837), .b(n_44775), .o(n_40881) );
in01s02 FE_RC_31_0 ( .a(n_17780), .o(FE_RN_10_0) );
na03s04 FE_RC_3205_0 ( .a(n_41730), .b(n_41748), .c(n_41749), .o(FE_RN_1355_0) );
no02f08 FE_RC_3206_0 ( .a(n_41939), .b(FE_RN_1355_0), .o(n_41962) );
oa22f04 FE_RC_3207_0 ( .a(n_41764), .b(FE_OCP_RBN5744_n_42043), .c(n_41765), .d(n_42043), .o(n_42122) );
in01s06 FE_RC_3208_0 ( .a(FE_RN_1356_0), .o(n_17656) );
no02s06 FE_RC_3209_0 ( .a(n_17683), .b(FE_OCPN937_n_17684), .o(FE_RN_1356_0) );
na02s01 FE_RC_3210_0 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_1_), .b(FE_OCP_RBN6440_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_RN_1357_0) );
na02s02 FE_RC_3211_0 ( .a(FE_RN_1357_0), .b(n_6607), .o(n_6649) );
oa22m02 FE_RC_3212_0 ( .a(FE_OCP_RBN2629_n_2737), .b(n_3591), .c(n_3615), .d(n_47017), .o(n_3761) );
in01s01 FE_RC_3213_0 ( .a(n_30145), .o(FE_RN_1358_0) );
no02f06 FE_RC_3214_0 ( .a(n_45630), .b(FE_RN_1358_0), .o(FE_RN_1359_0) );
ao12f06 FE_RC_3215_0 ( .a(FE_RN_1359_0), .b(FE_RN_525_0), .c(n_45630), .o(n_30428) );
na03f10 TIMEBOOST_cell_8202 ( .a(n_28008), .b(n_27941), .c(n_27896), .o(n_28086) );
na02s06 FE_RC_3218_0 ( .a(n_27175), .b(n_27227), .o(FE_RN_1360_0) );
no02s06 FE_RC_3219_0 ( .a(n_27476), .b(FE_RN_1360_0), .o(n_27535) );
na02m40 FE_RC_3226_0 ( .a(FE_OCP_RBN6471_delay_xor_ln21_unr15_stage6_stallmux_q_3_), .b(n_44061), .o(FE_RN_1364_0) );
na02s02 TIMEBOOST_cell_6990 ( .a(TIMEBOOST_net_2253), .b(FE_OCP_RBN3017_n_20404), .o(n_20499) );
na02s01 TIMEBOOST_cell_6601 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_12_), .b(n_40493), .o(TIMEBOOST_net_2058) );
in01s01 FE_RC_3236_0 ( .a(FE_RN_1371_0), .o(FE_RN_1370_0) );
no02s02 FE_RC_3237_0 ( .a(n_33270), .b(FE_RN_1370_0), .o(FE_RN_1372_0) );
na02m04 FE_RC_3238_0 ( .a(n_33635), .b(FE_RN_1372_0), .o(n_33655) );
in01s01 FE_RC_3239_0 ( .a(n_33199), .o(FE_RN_1373_0) );
in01s01 FE_RC_3240_0 ( .a(FE_RN_1373_0), .o(FE_RN_1371_0) );
in01s02 FE_RC_3241_0 ( .a(n_11997), .o(FE_RN_1374_0) );
in01s02 FE_RC_3242_0 ( .a(n_11998), .o(FE_RN_1375_0) );
na02s02 TIMEBOOST_cell_8114 ( .a(n_11465), .b(n_11464), .o(TIMEBOOST_net_2688) );
na02s02 TIMEBOOST_cell_7066 ( .a(TIMEBOOST_net_2291), .b(n_11557), .o(n_11745) );
in01s01 FE_RC_3245_0 ( .a(n_12393), .o(FE_RN_1377_0) );
in01s06 FE_RC_3246_0 ( .a(n_12394), .o(FE_RN_1378_0) );
in01s02 FE_RC_3249_0 ( .a(n_31058), .o(FE_RN_1380_0) );
no02s01 TIMEBOOST_cell_8498 ( .a(n_37730), .b(n_37632), .o(TIMEBOOST_net_2736) );
no03f20 TIMEBOOST_cell_3468 ( .a(n_27938), .b(FE_OCP_RBN2039_n_44722), .c(n_28058), .o(n_28083) );
no02s01 TIMEBOOST_cell_1599 ( .a(n_34852), .b(n_34372), .o(TIMEBOOST_net_414) );
in01s01 FE_RC_3259_0 ( .a(n_29561), .o(FE_RN_1386_0) );
in01s02 FE_RC_3260_0 ( .a(FE_RN_1386_0), .o(FE_RN_1384_0) );
in01s06 FE_RC_3261_0 ( .a(n_12396), .o(FE_RN_1387_0) );
in01s04 FE_RC_3262_0 ( .a(FE_RN_1389_0), .o(FE_RN_1388_0) );
in01m08 FE_RC_3263_0 ( .a(FE_RN_1390_0), .o(n_12571) );
no02f06 TIMEBOOST_cell_7533 ( .a(TIMEBOOST_net_2397), .b(FE_RN_1672_0), .o(TIMEBOOST_net_1040) );
in01s02 FE_RC_3265_0 ( .a(FE_OCPN1657_n_12368), .o(FE_RN_1391_0) );
in01s02 FE_RC_3266_0 ( .a(FE_RN_1391_0), .o(FE_RN_1389_0) );
no02s01 TIMEBOOST_cell_7047 ( .a(n_4556), .b(n_4316), .o(TIMEBOOST_net_2282) );
in01s02 FE_RC_3273_0 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_13_), .o(FE_RN_1396_0) );
in01s01 FE_RC_3274_0 ( .a(FE_OCP_RBN2414_n_44722), .o(FE_RN_1397_0) );
no03f04 TIMEBOOST_cell_5176 ( .a(n_25037), .b(n_25038), .c(n_25036), .o(TIMEBOOST_net_1536) );
no02m06 TIMEBOOST_cell_3931 ( .a(n_29345), .b(n_28847), .o(TIMEBOOST_net_1056) );
na02m10 FE_RC_3277_0 ( .a(n_28385), .b(FE_RN_1399_0), .o(FE_RN_1401_0) );
oa12f08 FE_RC_3278_0 ( .a(FE_RN_1401_0), .b(FE_RN_1402_0), .c(n_28385), .o(n_28453) );
no03m20 TIMEBOOST_cell_3442 ( .a(n_32602), .b(n_32599), .c(n_32522), .o(TIMEBOOST_net_25) );
in01f06 FE_RC_3280_0 ( .a(FE_OCPN3549_n_28381), .o(FE_RN_1402_0) );
in01s01 FE_RC_3281_0 ( .a(n_28005), .o(FE_RN_1404_0) );
in01s01 FE_RC_3282_0 ( .a(FE_RN_1404_0), .o(FE_RN_1400_0) );
in01s01 FE_RC_3283_0 ( .a(n_33604), .o(FE_RN_1405_0) );
na02f10 FE_RC_3284_0 ( .a(FE_OCP_RBN5713_n_44102), .b(FE_RN_1405_0), .o(n_34203) );
in01s06 FE_RC_3285_0 ( .a(FE_RN_1406_0), .o(n_12270) );
no02s06 FE_RC_3286_0 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_6_), .b(n_12100), .o(FE_RN_1406_0) );
in01s01 FE_RC_3290_0 ( .a(n_12438), .o(FE_RN_1409_0) );
na02s02 FE_RC_3291_0 ( .a(n_12491), .b(FE_RN_1409_0), .o(n_12500) );
no02s01 TIMEBOOST_cell_5319 ( .a(TIMEBOOST_net_1607), .b(n_35882), .o(n_35959) );
na02s10 FE_RC_3293_0 ( .a(n_16936), .b(n_16900), .o(FE_RN_1410_0) );
no02s06 TIMEBOOST_cell_5017 ( .a(TIMEBOOST_net_1456), .b(n_18990), .o(n_19077) );
na02m04 TIMEBOOST_cell_6821 ( .a(n_16404), .b(n_16369), .o(TIMEBOOST_net_2168) );
no02m08 TIMEBOOST_cell_6678 ( .a(TIMEBOOST_net_2096), .b(n_24782), .o(n_24894) );
na02m10 FE_RC_3298_0 ( .a(FE_RN_1414_0), .b(FE_RN_1410_0), .o(n_17194) );
na02s02 TIMEBOOST_cell_8716 ( .a(FE_RN_273_0), .b(FE_OCP_RBN5559_n_1853), .o(TIMEBOOST_net_2845) );
no02m04 TIMEBOOST_cell_1818 ( .a(TIMEBOOST_net_523), .b(n_16234), .o(n_16325) );
in01s02 FE_RC_3300_0 ( .a(n_12667), .o(FE_RN_1416_0) );
in01s02 FE_RC_3301_0 ( .a(FE_RN_1417_0), .o(n_12728) );
no03s02 TIMEBOOST_cell_8242 ( .a(n_24162), .b(n_23763), .c(n_23764), .o(TIMEBOOST_net_2403) );
in01s01 FE_RC_3305_0 ( .a(n_12955), .o(FE_RN_1420_0) );
in01s02 FE_RC_3307_0 ( .a(FE_RN_1421_0), .o(n_12620) );
na02s02 FE_RC_3308_0 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_17_), .b(n_12565), .o(FE_RN_1421_0) );
ao22s10 FE_RC_3312_0 ( .a(n_44365), .b(FE_OCP_RBN1121_delay_xor_ln22_unr12_stage5_stallmux_q_2_), .c(delay_xor_ln22_unr12_stage5_stallmux_q_2_), .d(FE_OCP_RBN7107_n_44365), .o(n_16970) );
in01m02 FE_RC_3313_0 ( .a(n_18343), .o(FE_RN_1424_0) );
na02f04 FE_RC_3315_0 ( .a(n_18650), .b(FE_RN_1424_0), .o(FE_RN_1425_0) );
na02s10 FE_RC_3316_0 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_1_), .b(FE_OCP_RBN7008_n_44962), .o(FE_RN_1426_0) );
in01m01 FE_RC_3323_0 ( .a(FE_OCP_RBN4100_n_12880), .o(FE_RN_1431_0) );
in01s03 FE_RC_3324_0 ( .a(FE_RN_1431_0), .o(n_13195) );
ao22s06 FE_RC_3329_0 ( .a(n_33368), .b(n_33805), .c(n_33326), .d(n_33870), .o(n_33871) );
na02m02 FE_RC_3330_0 ( .a(n_18678), .b(FE_OFN737_n_17093), .o(FE_RN_1434_0) );
na02m04 FE_RC_3331_0 ( .a(FE_RN_1434_0), .b(n_18646), .o(n_18824) );
in01s10 FE_RC_3332_0 ( .a(n_27962), .o(FE_RN_1435_0) );
in01s10 FE_RC_3333_0 ( .a(n_27966), .o(FE_RN_1436_0) );
no02m02 FE_RC_3337_0 ( .a(n_18713), .b(n_17732), .o(FE_RN_1438_0) );
no02m04 FE_RC_3338_0 ( .a(n_18824), .b(FE_RN_1438_0), .o(n_18858) );
in01s02 FE_RC_3339_0 ( .a(n_12547), .o(FE_RN_1439_0) );
no02m02 FE_RC_3340_0 ( .a(FE_OCP_RBN3703_n_12904), .b(FE_RN_1439_0), .o(FE_RN_1440_0) );
no02s04 FE_RC_3342_0 ( .a(FE_OCP_RBN4037_n_12904), .b(n_12547), .o(FE_RN_1442_0) );
no02m06 FE_RC_3343_0 ( .a(FE_RN_1442_0), .b(FE_RN_1440_0), .o(n_13098) );
in01s01 FE_RC_3350_0 ( .a(n_18357), .o(FE_RN_1446_0) );
no02m08 FE_RC_3351_0 ( .a(FE_RN_1446_0), .b(n_19088), .o(n_19116) );
ao22f06 FE_RC_3352_0 ( .a(n_14225), .b(n_14887), .c(n_14265), .d(n_14886), .o(n_14982) );
oa22f06 FE_RC_3353_0 ( .a(n_28675), .b(n_28965), .c(n_28674), .d(n_28966), .o(n_29055) );
na02s01 FE_RC_3355_0 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_24_), .b(FE_RN_1447_0), .o(FE_RN_1448_0) );
na02s04 FE_RC_3356_0 ( .a(n_13866), .b(FE_RN_1450_0), .o(FE_RN_1449_0) );
na02m06 FE_RC_3357_0 ( .a(FE_RN_1449_0), .b(FE_RN_1448_0), .o(n_13955) );
in01s01 FE_RC_3358_0 ( .a(n_12929), .o(FE_RN_1451_0) );
in01s02 FE_RC_3359_0 ( .a(FE_RN_1451_0), .o(FE_RN_1447_0) );
na02s02 TIMEBOOST_cell_4279 ( .a(n_13277), .b(n_13424), .o(TIMEBOOST_net_1230) );
in01s01 FE_RC_3360_0 ( .a(n_47250), .o(FE_RN_1452_0) );
in01s01 FE_RC_3361_0 ( .a(FE_RN_1452_0), .o(FE_RN_1450_0) );
na02m06 FE_RC_3362_0 ( .a(FE_OFN773_n_25834), .b(n_29167), .o(FE_RN_1453_0) );
na02m10 FE_RC_3363_0 ( .a(n_29316), .b(FE_RN_1453_0), .o(n_29339) );
no02m04 FE_RC_3364_0 ( .a(FE_OCP_RBN2539_n_12880), .b(n_13335), .o(FE_RN_1454_0) );
no02m08 FE_RC_3365_0 ( .a(FE_RN_1454_0), .b(n_13390), .o(n_13436) );
in01s01 FE_RC_3366_0 ( .a(FE_OCPN1926_n_34516), .o(FE_RN_1455_0) );
no02s10 FE_RC_3367_0 ( .a(FE_OCP_RBN6044_n_35487), .b(FE_RN_1455_0), .o(n_35575) );
in01s01 FE_RC_3368_0 ( .a(FE_OFN4795_n_13195), .o(FE_RN_1456_0) );
in01f02 FE_RC_3369_0 ( .a(FE_RN_1457_0), .o(n_14605) );
ao22s04 FE_RC_336_0 ( .a(n_1462), .b(n_1558), .c(n_792), .d(n_1780), .o(n_1590) );
no02f02 FE_RC_3370_0 ( .a(FE_RN_1456_0), .b(n_14462), .o(FE_RN_1457_0) );
in01s01 FE_RC_3373_0 ( .a(FE_RN_1458_0), .o(FE_RN_1460_0) );
in01s01 FE_RC_3374_0 ( .a(FE_RN_1460_0), .o(n_19218) );
in01s01 FE_RC_3375_0 ( .a(n_27014), .o(FE_RN_1461_0) );
na02f04 FE_RC_3377_0 ( .a(n_30580), .b(FE_RN_1461_0), .o(FE_RN_1462_0) );
no02s01 FE_RC_3378_0 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_23_), .b(n_23599), .o(FE_RN_1463_0) );
no02m08 FE_RC_3379_0 ( .a(FE_RN_1463_0), .b(n_24285), .o(n_24340) );
ao22s03 FE_RC_337_0 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_6_), .b(n_1528), .c(n_1549), .d(n_1590), .o(n_1591) );
na02m02 TIMEBOOST_cell_7983 ( .a(TIMEBOOST_net_2622), .b(n_5176), .o(n_5321) );
in01s02 FE_RC_3383_0 ( .a(n_14466), .o(FE_RN_1467_0) );
na02m02 FE_RC_3384_0 ( .a(n_14478), .b(FE_RN_1467_0), .o(FE_RN_1468_0) );
in01s01 FE_RC_3385_0 ( .a(FE_OCP_RBN2078_n_14149), .o(FE_RN_1469_0) );
na02m04 FE_RC_3386_0 ( .a(FE_RN_1468_0), .b(FE_RN_1469_0), .o(FE_RN_1470_0) );
na02m06 FE_RC_3387_0 ( .a(FE_RN_1466_0), .b(FE_RN_1470_0), .o(n_14672) );
no02s01 TIMEBOOST_cell_5267 ( .a(TIMEBOOST_net_1581), .b(n_39149), .o(n_39173) );
na02s06 TIMEBOOST_cell_8671 ( .a(TIMEBOOST_net_2822), .b(n_35687), .o(n_35822) );
na02s06 FE_RC_3390_0 ( .a(n_33964), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(FE_RN_1472_0) );
na02f08 FE_RC_3391_0 ( .a(n_33962), .b(FE_RN_1472_0), .o(n_33983) );
in01s01 FE_RC_3394_0 ( .a(FE_OCPN1234_n_33341), .o(FE_RN_1474_0) );
na02m01 FE_RC_3395_0 ( .a(n_44100), .b(FE_RN_1474_0), .o(n_34117) );
na02m08 FE_RC_3397_0 ( .a(FE_OFN743_delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n_24612), .o(FE_RN_1475_0) );
na02m08 FE_RC_3398_0 ( .a(n_24800), .b(FE_RN_1475_0), .o(n_24870) );
na02s01 TIMEBOOST_cell_6867 ( .a(n_32556), .b(n_32555), .o(TIMEBOOST_net_2192) );
in01m01 FE_RC_3401_0 ( .a(n_19213), .o(n_19207) );
no02s02 FE_RC_3402_0 ( .a(n_19181), .b(n_19213), .o(n_19271) );
na02f06 FE_RC_3403_0 ( .a(n_33925), .b(n_33880), .o(FE_RN_1477_0) );
na02f08 FE_RC_3404_0 ( .a(FE_RN_1477_0), .b(n_33881), .o(n_34017) );
in01s01 FE_RC_3405_0 ( .a(FE_OCP_RBN2757_n_13796), .o(FE_RN_1478_0) );
in01f02 FE_RC_3406_0 ( .a(FE_RN_1479_0), .o(n_14612) );
no02f02 FE_RC_3407_0 ( .a(n_14554), .b(FE_RN_1478_0), .o(FE_RN_1479_0) );
ao22m06 FE_RC_3408_0 ( .a(n_15450), .b(n_15989), .c(FE_RN_1480_0), .d(n_15990), .o(n_16146) );
in01s01 FE_RC_3409_0 ( .a(n_15449), .o(FE_RN_1481_0) );
in01s01 FE_RC_3410_0 ( .a(FE_RN_1481_0), .o(FE_RN_1480_0) );
oa22m04 FE_RC_3411_0 ( .a(n_34745), .b(FE_OCP_RBN6753_n_35049), .c(n_34746), .d(n_35049), .o(n_35130) );
na03f04 TIMEBOOST_cell_7303 ( .a(n_39822), .b(n_39816), .c(n_39802), .o(n_39876) );
na03f08 TIMEBOOST_cell_7304 ( .a(TIMEBOOST_net_1351), .b(n_39846), .c(FE_RN_1093_0), .o(FE_RN_1094_0) );
na02s02 FE_RC_3421_0 ( .a(n_14419), .b(FE_OCP_RBN3070_n_15275), .o(FE_RN_1487_0) );
na02f04 FE_RC_3422_0 ( .a(FE_RN_1487_0), .b(n_15504), .o(n_15547) );
in01s01 FE_RC_3423_0 ( .a(FE_RN_1486_0), .o(FE_RN_1488_0) );
in01s03 FE_RC_3424_0 ( .a(FE_RN_1488_0), .o(n_14419) );
in01s02 FE_RC_3428_0 ( .a(n_35294), .o(FE_RN_1491_0) );
na02m02 FE_RC_3429_0 ( .a(n_35275), .b(FE_RN_1491_0), .o(FE_RN_1492_0) );
na02m04 FE_RC_3431_0 ( .a(FE_RN_1492_0), .b(n_35180), .o(FE_RN_1493_0) );
no02s01 FE_RC_3432_0 ( .a(n_30577), .b(n_30173), .o(FE_RN_1494_0) );
na02m08 FE_RC_3433_0 ( .a(FE_RN_1494_0), .b(n_30558), .o(n_30603) );
ao22f02 FE_RC_3437_0 ( .a(n_45013), .b(n_20733), .c(n_45050), .d(n_20734), .o(n_20857) );
no02m02 FE_RC_3439_0 ( .a(FE_RN_1185_0), .b(n_26442), .o(FE_RN_1496_0) );
in01s01 FE_RC_3440_0 ( .a(n_45024), .o(FE_RN_1497_0) );
in01s06 FE_RC_3441_0 ( .a(FE_RN_1498_0), .o(n_21316) );
no02m04 FE_RC_3442_0 ( .a(FE_RN_1497_0), .b(n_21157), .o(FE_RN_1498_0) );
oa22f04 FE_RC_344_0 ( .a(FE_OCP_RBN5663_n_2438), .b(FE_OCP_RBN6642_n_3502), .c(FE_OCP_RBN5653_n_2438), .d(n_3502), .o(n_3018) );
no02s02 FE_RC_3451_0 ( .a(n_25359), .b(n_25358), .o(FE_RN_1505_0) );
no02m02 FE_RC_3452_0 ( .a(n_25656), .b(FE_RN_1505_0), .o(n_25678) );
na02f06 FE_RC_3454_0 ( .a(FE_OCP_RBN3149_n_15553), .b(n_15648), .o(n_15688) );
no02s01 FE_RC_3455_0 ( .a(FE_OCPN1336_n_25673), .b(FE_RN_1508_0), .o(FE_RN_1507_0) );
na02m08 FE_RC_3456_0 ( .a(FE_RN_1507_0), .b(n_26263), .o(n_26376) );
in01s01 FE_RC_3457_0 ( .a(n_25648), .o(FE_RN_1509_0) );
in01s01 FE_RC_3458_0 ( .a(FE_RN_1509_0), .o(FE_RN_1508_0) );
oa22s01 FE_RC_345_0 ( .a(n_1124), .b(n_44652), .c(n_1100), .d(n_44637), .o(n_1303) );
na02s01 FE_RC_3461_0 ( .a(FE_OCP_RBN2064_n_19353), .b(n_19461), .o(FE_RN_1511_0) );
in01s01 FE_RC_3462_0 ( .a(n_20429), .o(FE_RN_1512_0) );
na02s06 FE_RC_3463_0 ( .a(FE_RN_1511_0), .b(FE_RN_1512_0), .o(FE_RN_1513_0) );
na02m10 FE_RC_3464_0 ( .a(FE_RN_1513_0), .b(n_20926), .o(n_20947) );
in01s02 FE_RC_3465_0 ( .a(n_21192), .o(FE_RN_1514_0) );
no02f04 FE_RC_3466_0 ( .a(FE_RN_1514_0), .b(n_21202), .o(n_21240) );
oa22f02 FE_RC_3467_0 ( .a(n_46973), .b(n_17336), .c(n_17753), .d(n_17187), .o(n_17337) );
oa22s01 FE_RC_346_0 ( .a(n_1152), .b(n_44652), .c(n_1138), .d(n_44623), .o(n_1311) );
in01s01 FE_RC_3473_0 ( .a(n_22043), .o(FE_RN_1518_0) );
na02s01 FE_RC_3474_0 ( .a(FE_RN_1518_0), .b(FE_OCP_RBN1161_n_20763), .o(FE_RN_1519_0) );
na02s03 FE_RC_3475_0 ( .a(n_44275), .b(FE_RN_1519_0), .o(n_22170) );
in01s01 FE_RC_3476_0 ( .a(n_20867), .o(FE_RN_1520_0) );
no02s10 FE_RC_3477_0 ( .a(n_22288), .b(FE_RN_1520_0), .o(n_22554) );
oa22s01 FE_RC_347_0 ( .a(n_1211), .b(n_44652), .c(n_1204), .d(n_44623), .o(n_1317) );
in01s01 FE_RC_3480_0 ( .a(n_20867), .o(FE_RN_1523_0) );
na02m06 FE_RC_3482_0 ( .a(n_21708), .b(n_21849), .o(FE_RN_1524_0) );
na02m06 FE_RC_3483_0 ( .a(FE_OCP_RBN3328_n_21616), .b(FE_RN_1524_0), .o(n_21923) );
in01m02 FE_RC_3484_0 ( .a(FE_RN_1525_0), .o(n_16461) );
na02s02 FE_RC_3485_0 ( .a(FE_OCP_RBN2905_n_14590), .b(n_16319), .o(FE_RN_1525_0) );
in01m04 FE_RC_3489_0 ( .a(FE_RN_1528_0), .o(n_26532) );
no02f02 FE_RC_3490_0 ( .a(FE_OCP_DRV_N1488_n_24848), .b(n_26440), .o(FE_RN_1528_0) );
in01m02 FE_RC_3491_0 ( .a(n_21363), .o(FE_RN_1529_0) );
in01f02 FE_RC_3492_0 ( .a(n_21289), .o(FE_RN_1530_0) );
in01f02 FE_RC_3494_0 ( .a(n_21224), .o(FE_RN_1531_0) );
in01f02 FE_RC_3495_0 ( .a(n_21227), .o(FE_RN_1532_0) );
no02f04 TIMEBOOST_cell_1632 ( .a(TIMEBOOST_net_430), .b(n_8881), .o(FE_RN_2025_0) );
no02m06 FE_RC_3500_0 ( .a(FE_RN_1784_0), .b(n_15463), .o(n_15496) );
in01s01 FE_RC_3506_0 ( .a(n_27117), .o(FE_RN_1540_0) );
in01s01 FE_RC_3507_0 ( .a(FE_RN_1540_0), .o(FE_RN_1535_0) );
in01s02 FE_RC_3508_0 ( .a(n_22063), .o(FE_RN_1541_0) );
oa22f04 FE_RC_350_0 ( .a(n_42086), .b(n_41766), .c(n_41767), .d(n_42085), .o(n_42144) );
no02f06 FE_RC_3510_0 ( .a(n_22237), .b(FE_RN_1542_0), .o(n_22446) );
no02f04 FE_RC_3511_0 ( .a(n_15225), .b(n_15137), .o(FE_RN_1543_0) );
no02f06 FE_RC_3512_0 ( .a(FE_RN_1543_0), .b(n_45523), .o(n_15415) );
in01s01 FE_RC_3513_0 ( .a(FE_OCPN1281_n_21007), .o(FE_RN_1544_0) );
na02f04 FE_RC_3514_0 ( .a(FE_RN_1544_0), .b(n_46969), .o(n_21044) );
na02s06 FE_RC_3516_0 ( .a(n_17417), .b(FE_RN_1545_0), .o(n_17523) );
in01s01 FE_RC_3517_0 ( .a(n_28447), .o(FE_RN_1546_0) );
no02f08 TIMEBOOST_cell_4953 ( .a(TIMEBOOST_net_1424), .b(n_28310), .o(n_28368) );
in01s02 FE_RC_3519_0 ( .a(FE_RN_1548_0), .o(n_28607) );
na02m04 TIMEBOOST_cell_8641 ( .a(TIMEBOOST_net_2807), .b(n_30825), .o(n_30930) );
na04m20 TIMEBOOST_cell_5696 ( .a(n_36943), .b(FE_RN_163_0), .c(n_36944), .d(FE_RN_162_0), .o(n_37144) );
in01s01 FE_RC_3522_0 ( .a(n_28646), .o(FE_RN_1550_0) );
na02f06 TIMEBOOST_cell_6751 ( .a(FE_OCP_RBN3073_n_15706), .b(FE_RN_1486_0), .o(TIMEBOOST_net_2133) );
no02f08 TIMEBOOST_cell_7915 ( .a(TIMEBOOST_net_2588), .b(TIMEBOOST_net_893), .o(n_39628) );
in01s06 FE_RC_3526_0 ( .a(n_28647), .o(FE_RN_1553_0) );
no02s02 TIMEBOOST_cell_1691 ( .a(n_3477), .b(n_3364), .o(TIMEBOOST_net_460) );
in01m04 FE_RC_3529_0 ( .a(FE_OCPN1608_n_18176), .o(FE_RN_1554_0) );
in01s03 FE_RC_3530_0 ( .a(n_18177), .o(FE_RN_1555_0) );
na02s01 TIMEBOOST_cell_6037 ( .a(n_37574), .b(n_37556), .o(TIMEBOOST_net_1870) );
na02s02 TIMEBOOST_cell_5117 ( .a(TIMEBOOST_net_1506), .b(n_29749), .o(n_29779) );
na02s02 TIMEBOOST_cell_8769 ( .a(TIMEBOOST_net_2871), .b(n_14586), .o(TIMEBOOST_net_2464) );
no02m08 TIMEBOOST_cell_1950 ( .a(TIMEBOOST_net_589), .b(n_22998), .o(n_23175) );
no02s04 TIMEBOOST_cell_1597 ( .a(n_35130), .b(n_30633), .o(TIMEBOOST_net_413) );
in01s02 FE_RC_3537_0 ( .a(n_10458), .o(FE_RN_1558_0) );
no02f04 TIMEBOOST_cell_3066 ( .a(n_19114), .b(FE_OCPN1709_FE_OFN739_n_17093), .o(TIMEBOOST_net_824) );
na02f08 TIMEBOOST_cell_6684 ( .a(TIMEBOOST_net_2099), .b(FE_RN_978_0), .o(n_38616) );
no02s02 TIMEBOOST_cell_1643 ( .a(n_19565), .b(n_19064), .o(TIMEBOOST_net_436) );
oa22s02 FE_RC_3541_0 ( .a(n_6398), .b(n_6489), .c(n_6399), .d(n_6499), .o(n_6643) );
oa22f04 FE_RC_3542_0 ( .a(n_6447), .b(n_6574), .c(n_6448), .d(n_6558), .o(n_6720) );
ao22f08 FE_RC_3544_0 ( .a(n_40696), .b(FE_OCP_RBN5545_n_45145), .c(n_40339), .d(FE_OCP_RBN5545_n_45145), .o(n_40743) );
na02s01 TIMEBOOST_cell_3922 ( .a(TIMEBOOST_net_1051), .b(FE_OCP_RBN4133_n_38028), .o(n_38214) );
in01m10 FE_RC_3546_0 ( .a(n_27968), .o(FE_RN_1561_0) );
in01m08 FE_RC_3547_0 ( .a(FE_RN_1562_0), .o(n_28002) );
no02s03 TIMEBOOST_cell_5165 ( .a(TIMEBOOST_net_1530), .b(n_34128), .o(FE_RN_2247_0) );
ao22s02 FE_RC_3550_0 ( .a(n_1421), .b(FE_OCP_RBN5515_n_1472), .c(n_1467), .d(n_1472), .o(n_1588) );
oa22s02 FE_RC_3551_0 ( .a(FE_RN_1563_0), .b(FE_OCP_RBN6537_n_1614), .c(FE_RN_1564_0), .d(n_1614), .o(n_1701) );
in01s01 FE_RC_3552_0 ( .a(n_1438), .o(FE_RN_1564_0) );
in01s01 FE_RC_3553_0 ( .a(FE_RN_1564_0), .o(FE_RN_1563_0) );
oa22s02 FE_RC_3554_0 ( .a(n_36604), .b(n_36719), .c(n_36579), .d(n_36718), .o(n_36766) );
na02m08 TIMEBOOST_cell_7064 ( .a(TIMEBOOST_net_2290), .b(n_11227), .o(n_11327) );
no02s01 TIMEBOOST_cell_3950 ( .a(TIMEBOOST_net_1065), .b(n_20037), .o(n_20068) );
in01m20 FE_RC_3558_0 ( .a(n_23022), .o(FE_RN_1566_0) );
in01m10 FE_RC_3559_0 ( .a(FE_RN_1567_0), .o(n_23045) );
in01s20 FE_RC_355_0 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_3_), .o(FE_RN_105_0) );
na02m04 TIMEBOOST_cell_3951 ( .a(n_24421), .b(FE_OFN743_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(TIMEBOOST_net_1066) );
oa22m04 FE_RC_3561_0 ( .a(n_12659), .b(n_13062), .c(n_12660), .d(n_13008), .o(n_13228) );
ao22f06 FE_RC_3562_0 ( .a(n_39202), .b(n_39517), .c(n_39201), .d(n_39516), .o(n_39586) );
ao22f08 FE_RC_3563_0 ( .a(FE_RN_1568_0), .b(FE_OCP_RBN3081_n_39514), .c(FE_RN_1569_0), .d(n_39514), .o(n_39584) );
in01s02 FE_RC_3564_0 ( .a(n_39173), .o(FE_RN_1569_0) );
in01s02 FE_RC_3565_0 ( .a(FE_RN_1569_0), .o(FE_RN_1568_0) );
in01s06 FE_RC_3566_0 ( .a(FE_RN_1570_0), .o(FE_RN_1571_0) );
in01m04 FE_RC_3567_0 ( .a(FE_RN_53_0), .o(FE_RN_1572_0) );
na02m08 FE_RC_3568_0 ( .a(FE_RN_1571_0), .b(FE_RN_1572_0), .o(FE_RN_1573_0) );
no02m08 FE_RC_3569_0 ( .a(FE_OCP_RBN2479_n_47245), .b(FE_RN_1573_0), .o(n_23504) );
no02s02 TIMEBOOST_cell_1547 ( .a(n_38622), .b(FE_OFN5092_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(TIMEBOOST_net_388) );
in01s06 FE_RC_3570_0 ( .a(n_23131), .o(FE_RN_1574_0) );
in01m01 FE_RC_3571_0 ( .a(FE_RN_1574_0), .o(FE_RN_1570_0) );
in01m01 FE_RC_3573_0 ( .a(n_32621), .o(FE_RN_1577_0) );
no02m10 FE_RC_3574_0 ( .a(FE_RN_1579_0), .b(FE_RN_1577_0), .o(FE_RN_1578_0) );
in01m20 FE_RC_3576_0 ( .a(n_32855), .o(FE_RN_1579_0) );
in01s01 FE_RC_3578_0 ( .a(n_1850), .o(FE_RN_1580_0) );
no02f08 TIMEBOOST_cell_5085 ( .a(TIMEBOOST_net_1490), .b(n_18987), .o(n_19058) );
no03s02 TIMEBOOST_cell_8363 ( .a(n_3809), .b(n_3891), .c(n_3850), .o(n_4152) );
oa22f02 FE_RC_3582_0 ( .a(n_32287), .b(n_32255), .c(FE_OFN621_n_28336), .d(n_32240), .o(n_32289) );
oa22s02 FE_RC_3583_0 ( .a(n_3615), .b(n_3616), .c(FE_OFN4763_n_3029), .d(n_3610), .o(n_3776) );
no02s01 TIMEBOOST_cell_1723 ( .a(n_19268), .b(FE_OCP_RBN1139_n_19270), .o(TIMEBOOST_net_476) );
no02m06 TIMEBOOST_cell_7599 ( .a(TIMEBOOST_net_2430), .b(FE_OCP_RBN2765_n_38530), .o(n_38591) );
in01s02 FE_RC_3586_0 ( .a(n_12543), .o(FE_RN_1585_0) );
in01m02 FE_RC_3587_0 ( .a(FE_RN_1586_0), .o(n_12579) );
na03m08 TIMEBOOST_cell_8400 ( .a(n_15896), .b(n_15737), .c(n_15943), .o(n_16144) );
in01s04 FE_RC_3589_0 ( .a(n_12541), .o(FE_RN_1587_0) );
no02m02 TIMEBOOST_cell_6706 ( .a(TIMEBOOST_net_2110), .b(n_3261), .o(n_3379) );
in01s02 FE_RC_3590_0 ( .a(FE_RN_1587_0), .o(FE_RN_1584_0) );
in01s01 FE_RC_3592_0 ( .a(n_43083), .o(FE_RN_1588_0) );
in01s01 FE_RC_3593_0 ( .a(n_43121), .o(FE_RN_1589_0) );
no02s02 FE_RC_3594_0 ( .a(FE_RN_1588_0), .b(FE_RN_1589_0), .o(FE_RN_1590_0) );
no02s10 FE_RC_3595_0 ( .a(FE_OCP_RBN4456_n_43103), .b(FE_RN_1590_0), .o(n_43162) );
ao22s02 FE_RC_3596_0 ( .a(FE_OFN4765_n_3029), .b(FE_OCP_RBN5876_n_3848), .c(n_3082), .d(n_3848), .o(n_4011) );
in01s20 FE_RC_3597_0 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_5_), .o(FE_RN_1591_0) );
in01s06 FE_RC_3598_0 ( .a(FE_OCP_RBN3871_n_44061), .o(FE_RN_1592_0) );
no02f06 TIMEBOOST_cell_3902 ( .a(FE_RN_2725_0), .b(TIMEBOOST_net_1041), .o(n_19025) );
na03s08 TIMEBOOST_cell_8334 ( .a(FE_RN_672_0), .b(FE_RN_673_0), .c(FE_RN_674_0), .o(FE_RN_676_0) );
ao22s02 FE_RC_35_0 ( .a(n_1454), .b(n_1602), .c(n_1453), .d(FE_OCP_RBN6536_n_1602), .o(n_1658) );
na02s06 TIMEBOOST_cell_6869 ( .a(n_32578), .b(n_32582), .o(TIMEBOOST_net_2193) );
ao22s02 FE_RC_3601_0 ( .a(n_43580), .b(n_43780), .c(n_43579), .d(n_43779), .o(n_43835) );
oa22f06 FE_RC_3602_0 ( .a(FE_OCP_RBN6567_n_12714), .b(FE_OCP_RBN2530_n_13151), .c(n_12714), .d(n_13151), .o(n_13334) );
ao22f02 FE_RC_3603_0 ( .a(n_37579), .b(n_37575), .c(n_37581), .d(n_37644), .o(n_37657) );
in01s10 FE_RC_3604_0 ( .a(n_45200), .o(FE_RN_1594_0) );
in01s01 TIMEBOOST_cell_8893 ( .a(TIMEBOOST_net_2936), .o(TIMEBOOST_net_2937) );
no02s02 TIMEBOOST_cell_6832 ( .a(TIMEBOOST_net_2173), .b(n_31730), .o(TIMEBOOST_net_1749) );
oa22m02 FE_RC_3608_0 ( .a(n_7606), .b(n_8819), .c(n_7605), .d(n_8863), .o(n_8923) );
in01s01 FE_RC_3609_0 ( .a(n_33402), .o(FE_RN_1597_0) );
in01m04 FE_RC_360_0 ( .a(n_20309), .o(FE_RN_109_0) );
in01s02 FE_RC_3610_0 ( .a(n_33898), .o(FE_RN_1598_0) );
no02s06 FE_RC_3611_0 ( .a(FE_RN_1597_0), .b(FE_RN_1598_0), .o(FE_RN_1599_0) );
no02s08 FE_RC_3612_0 ( .a(FE_RN_1599_0), .b(n_33922), .o(n_34427) );
in01s01 FE_RC_3615_0 ( .a(FE_OCP_RBN2574_n_2558), .o(FE_RN_1600_0) );
in01s01 FE_RC_3616_0 ( .a(n_2763), .o(FE_RN_1601_0) );
na02s01 TIMEBOOST_cell_4244 ( .a(TIMEBOOST_net_1212), .b(n_18850), .o(TIMEBOOST_net_626) );
na02s02 TIMEBOOST_cell_4245 ( .a(FE_OCPN1908_n_17921), .b(n_17922), .o(TIMEBOOST_net_1213) );
no02s04 TIMEBOOST_cell_1802 ( .a(TIMEBOOST_net_515), .b(n_30471), .o(n_30512) );
in01f08 FE_RC_361_0 ( .a(FE_RN_110_0), .o(n_20616) );
ao22f04 FE_RC_3620_0 ( .a(n_38784), .b(n_38735), .c(n_38734), .d(n_38769), .o(n_38818) );
oa22m04 FE_RC_3621_0 ( .a(FE_OCP_RBN3089_n_4872), .b(FE_OCP_RBN3124_n_5121), .c(n_4900), .d(n_5121), .o(n_5300) );
ao22f04 FE_RC_3622_0 ( .a(n_38705), .b(n_38694), .c(n_38706), .d(n_38693), .o(n_38753) );
oa22f02 FE_RC_3623_0 ( .a(n_38653), .b(n_38678), .c(n_38666), .d(FE_OCP_RBN5816_n_38678), .o(n_38739) );
oa22m02 FE_RC_3624_0 ( .a(n_5389), .b(n_5250), .c(n_5249), .d(n_5361), .o(n_5531) );
oa22s02 FE_RC_3626_0 ( .a(FE_OCP_RBN5807_n_47018), .b(n_3781), .c(FE_OCP_RBN5806_n_47018), .d(n_3780), .o(n_3968) );
oa22s02 FE_RC_3628_0 ( .a(FE_OCP_RBN2627_n_2737), .b(n_47020), .c(FE_OCP_RBN5660_n_2438), .d(n_3231), .o(n_3259) );
no02s02 TIMEBOOST_cell_3086 ( .a(n_2682), .b(n_2681), .o(TIMEBOOST_net_834) );
oa22s02 FE_RC_3630_0 ( .a(n_4714), .b(n_4850), .c(n_4715), .d(n_4849), .o(n_5003) );
in01s01 FE_RC_3632_0 ( .a(FE_OFN321_n_2929), .o(FE_RN_1603_0) );
in01s01 FE_RC_3633_0 ( .a(n_2538), .o(FE_RN_1604_0) );
no02m06 TIMEBOOST_cell_6807 ( .a(TIMEBOOST_net_1138), .b(n_39575), .o(TIMEBOOST_net_2161) );
no02f08 TIMEBOOST_cell_6808 ( .a(TIMEBOOST_net_2161), .b(FE_OCP_RBN3224_n_39575), .o(n_39629) );
ao22f04 FE_RC_3636_0 ( .a(n_10320), .b(n_10317), .c(n_10318), .d(n_10321), .o(n_10480) );
oa22m02 FE_RC_3638_0 ( .a(n_40144), .b(n_40503), .c(n_40143), .d(n_40504), .o(n_40544) );
no03m06 FE_RC_3639_0 ( .a(n_5797), .b(n_5672), .c(n_5601), .o(n_5905) );
ao22m06 FE_RC_3641_0 ( .a(n_25692), .b(FE_OCP_RBN3205_n_26042), .c(n_25691), .d(n_26042), .o(n_26171) );
ao22m04 FE_RC_3642_0 ( .a(n_5904), .b(n_6068), .c(n_5921), .d(n_6067), .o(n_6165) );
oa22m02 FE_RC_3643_0 ( .a(n_44570), .b(FE_OCP_RBN5817_n_8687), .c(FE_OCP_RBN5780_n_44570), .d(n_8687), .o(n_9001) );
oa22s02 FE_RC_3644_0 ( .a(FE_OCP_RBN2744_n_14114), .b(FE_OCP_RBN6801_n_15156), .c(FE_RN_1606_0), .d(FE_OCP_RBN6802_n_15156), .o(n_15523) );
in01s01 FE_RC_3645_0 ( .a(n_14274), .o(FE_RN_1607_0) );
in01s01 FE_RC_3646_0 ( .a(FE_RN_1607_0), .o(FE_RN_1606_0) );
oa22m04 FE_RC_3648_0 ( .a(n_6456), .b(n_6503), .c(n_6493), .d(FE_OCP_RBN6239_n_6456), .o(n_6627) );
oa22s02 FE_RC_3649_0 ( .a(FE_OFN4787_n_46137), .b(n_6567), .c(FE_OFN770_n_46196), .d(FE_OCP_RBN6249_n_6567), .o(n_46186) );
oa22f06 FE_RC_364_0 ( .a(n_42897), .b(n_42585), .c(n_42586), .d(n_42896), .o(n_42959) );
oa22m04 FE_RC_3650_0 ( .a(n_6554), .b(n_6443), .c(n_6442), .d(n_6572), .o(n_6739) );
ao22f04 FE_RC_3655_0 ( .a(n_16865), .b(n_17083), .c(n_16864), .d(n_17123), .o(n_17334) );
oa22f02 FE_RC_3656_0 ( .a(n_17336), .b(n_17440), .c(n_17753), .d(n_17334), .o(n_17476) );
no03m08 TIMEBOOST_cell_7496 ( .a(n_37609), .b(n_37117), .c(n_37608), .o(TIMEBOOST_net_2379) );
oa22f04 FE_RC_3662_0 ( .a(FE_OCP_RBN6170_n_6059), .b(n_6130), .c(n_6059), .d(n_6115), .o(n_6214) );
oa22m02 FE_RC_3663_0 ( .a(n_36748), .b(FE_OCP_RBN6235_n_36780), .c(n_36780), .d(n_36749), .o(n_36829) );
in01s01 FE_RC_3664_0 ( .a(n_23680), .o(FE_RN_1611_0) );
in01m01 FE_RC_3665_0 ( .a(n_24067), .o(FE_RN_1612_0) );
na02m02 FE_RC_3666_0 ( .a(FE_RN_1611_0), .b(FE_RN_1612_0), .o(FE_RN_1613_0) );
no02m04 FE_RC_3667_0 ( .a(n_24068), .b(FE_RN_1613_0), .o(n_24081) );
no02f02 TIMEBOOST_cell_1729 ( .a(n_15552), .b(n_14452), .o(TIMEBOOST_net_479) );
ao22f08 FE_RC_3669_0 ( .a(n_44028), .b(n_40629), .c(n_40639), .d(n_40630), .o(n_40668) );
ao22s06 FE_RC_3670_0 ( .a(n_6579), .b(n_6638), .c(n_6656), .d(n_6637), .o(n_6835) );
in01s01 FE_RC_3672_0 ( .a(n_41406), .o(FE_RN_1614_0) );
in01s01 FE_RC_3673_0 ( .a(n_41407), .o(FE_RN_1615_0) );
no02s02 FE_RC_3674_0 ( .a(FE_RN_1614_0), .b(FE_RN_1615_0), .o(FE_RN_1616_0) );
no02m04 FE_RC_3675_0 ( .a(FE_OCP_RBN6620_n_41381), .b(FE_RN_1616_0), .o(n_41453) );
in01s01 FE_RC_3676_0 ( .a(n_2394), .o(FE_RN_1617_0) );
in01s01 FE_RC_3677_0 ( .a(n_2419), .o(FE_RN_1618_0) );
no03m06 TIMEBOOST_cell_8289 ( .a(FE_OCP_RBN5741_n_4336), .b(n_4336), .c(FE_OCP_RBN5821_n_3437), .o(TIMEBOOST_net_1574) );
na02m08 TIMEBOOST_cell_7805 ( .a(TIMEBOOST_net_2533), .b(n_10939), .o(n_11089) );
ao22s02 FE_RC_3680_0 ( .a(FE_OCP_RBN2492_FE_RN_1367_0), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_23_), .c(n_28606), .d(FE_OCP_RBN6556_n_28458), .o(n_28699) );
oa22s02 FE_RC_3681_0 ( .a(n_1491), .b(FE_RN_398_0), .c(n_1494), .d(FE_RN_399_0), .o(n_1585) );
ao22m04 FE_RC_3682_0 ( .a(n_7732), .b(n_8943), .c(n_7733), .d(n_8944), .o(n_9091) );
ao22s01 FE_RC_3683_0 ( .a(n_17409), .b(FE_OCP_RBN7103_n_44365), .c(delay_xor_ln21_unr12_stage5_stallmux_q_6_), .d(FE_OCP_RBN7104_n_44365), .o(n_17485) );
oa22m02 FE_RC_3684_0 ( .a(FE_OCP_RBN4138_n_7743), .b(FE_OCP_RBN2785_n_8767), .c(FE_OCPN935_n_7802), .d(n_8767), .o(n_8870) );
in01s01 FE_RC_3689_0 ( .a(n_43526), .o(FE_RN_1620_0) );
na02s01 TIMEBOOST_cell_3359 ( .a(TIMEBOOST_net_970), .b(n_26974), .o(n_27031) );
no02s02 TIMEBOOST_cell_3360 ( .a(n_31991), .b(n_47273), .o(TIMEBOOST_net_971) );
oa22f02 FE_RC_3693_0 ( .a(n_24207), .b(FE_OCP_RBN1023_n_24125), .c(n_24125), .d(n_24269), .o(n_24291) );
ao22f02 FE_RC_3694_0 ( .a(n_43539), .b(n_43894), .c(n_43540), .d(n_43895), .o(n_43912) );
oa22f04 FE_RC_3696_0 ( .a(n_23486), .b(n_26464), .c(n_23590), .d(FE_OCP_RBN3274_n_26464), .o(n_26583) );
oa22m02 FE_RC_3698_0 ( .a(n_40598), .b(n_40576), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .d(n_40568), .o(n_40580) );
ao22s04 FE_RC_3699_0 ( .a(n_10416), .b(n_10808), .c(n_10798), .d(n_10415), .o(n_10944) );
ao22s02 FE_RC_369_0 ( .a(n_12185), .b(n_11877), .c(n_11878), .d(n_47211), .o(n_12316) );
oa22s06 FE_RC_36_0 ( .a(n_17792), .b(n_17884), .c(n_17793), .d(n_17842), .o(n_17942) );
oa22m02 FE_RC_3700_0 ( .a(FE_OFN787_n_46285), .b(n_12117), .c(FE_OCP_RBN3352_FE_OFN760_n_46337), .d(FE_OCP_RBN6253_n_12117), .o(n_46352) );
oa22m02 FE_RC_3702_0 ( .a(FE_OFN787_n_46285), .b(n_12162), .c(FE_OCP_RBN3352_FE_OFN760_n_46337), .d(n_12132), .o(n_46349) );
oa22s04 FE_RC_3704_0 ( .a(n_11701), .b(n_11954), .c(n_11700), .d(n_11982), .o(n_12158) );
oa22s02 FE_RC_3705_0 ( .a(FE_OCP_RBN6865_n_46285), .b(n_12158), .c(FE_OFN765_n_46337), .d(n_12133), .o(n_46348) );
oa22s02 FE_RC_3706_0 ( .a(n_24059), .b(n_27693), .c(n_27845), .d(n_27666), .o(n_27731) );
in01s01 FE_RC_3709_0 ( .a(FE_OCP_RBN4087_n_12880), .o(FE_RN_1623_0) );
in01f02 FE_RC_3710_0 ( .a(n_13693), .o(FE_RN_1624_0) );
na03s02 TIMEBOOST_cell_4770 ( .a(n_9639), .b(n_9447), .c(n_9464), .o(n_9883) );
na02m01 TIMEBOOST_cell_6029 ( .a(n_1891), .b(n_1892), .o(TIMEBOOST_net_1866) );
oa22m06 FE_RC_3713_0 ( .a(n_13172), .b(n_13711), .c(n_13180), .d(n_13665), .o(n_13751) );
in01s02 FE_RC_3714_0 ( .a(FE_OCP_RBN2056_n_13784), .o(FE_RN_1626_0) );
na02f06 FE_RC_3716_0 ( .a(FE_OCP_RBN2065_n_13913), .b(FE_RN_1626_0), .o(FE_RN_1628_0) );
na02f08 FE_RC_3717_0 ( .a(FE_RN_1628_0), .b(FE_RN_471_0), .o(n_14092) );
oa22f06 FE_RC_3719_0 ( .a(n_15610), .b(n_15613), .c(n_15609), .d(n_15615), .o(n_15889) );
na02s01 TIMEBOOST_cell_8822 ( .a(FE_OCP_RBN4254_n_3705), .b(n_3258), .o(TIMEBOOST_net_2898) );
na03m08 FE_RC_3723_0 ( .a(n_41577), .b(n_41479), .c(n_41488), .o(n_41578) );
ao22f04 FE_RC_3724_0 ( .a(FE_RN_1629_0), .b(n_33656), .c(n_33251), .d(n_33655), .o(n_33728) );
in01s01 FE_RC_3725_0 ( .a(n_33250), .o(FE_RN_1630_0) );
in01s02 FE_RC_3726_0 ( .a(FE_RN_1630_0), .o(FE_RN_1629_0) );
no02s02 TIMEBOOST_cell_1652 ( .a(TIMEBOOST_net_440), .b(n_4385), .o(n_4386) );
ao22m02 FE_RC_3728_0 ( .a(FE_OCPN935_n_7802), .b(n_8764), .c(FE_OCP_RBN4146_n_7743), .d(n_8765), .o(n_8879) );
oa22f04 FE_RC_3729_0 ( .a(FE_OCP_RBN4146_n_7743), .b(n_8828), .c(FE_OCP_DRV_N3506_n_8189), .d(n_8842), .o(n_8974) );
in01s01 FE_RC_3730_0 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_5_), .o(FE_RN_1631_0) );
na02s02 TIMEBOOST_cell_3994 ( .a(TIMEBOOST_net_1087), .b(n_2469), .o(n_2623) );
no02m02 TIMEBOOST_cell_5293 ( .a(TIMEBOOST_net_1594), .b(n_9682), .o(TIMEBOOST_net_1292) );
no02f06 TIMEBOOST_cell_7685 ( .a(TIMEBOOST_net_2473), .b(TIMEBOOST_net_314), .o(n_42150) );
oa22m04 FE_RC_3737_0 ( .a(FE_OCP_RBN6162_FE_RN_1136_0), .b(n_11324), .c(n_11323), .d(FE_RN_1136_0), .o(n_11403) );
ao22f06 FE_RC_3739_0 ( .a(n_14403), .b(n_14474), .c(n_14404), .d(n_14448), .o(n_14641) );
no02s04 TIMEBOOST_cell_1602 ( .a(TIMEBOOST_net_415), .b(FE_RN_2437_0), .o(FE_RN_2438_0) );
ao22f04 FE_RC_3745_0 ( .a(n_13709), .b(n_13211), .c(n_13212), .d(n_13695), .o(n_13818) );
ao22m04 FE_RC_374_0 ( .a(n_28643), .b(n_28978), .c(n_28644), .d(n_28977), .o(n_29062) );
oa22m04 FE_RC_3751_0 ( .a(n_45747), .b(n_11638), .c(n_11639), .d(n_45748), .o(n_12117) );
no03f10 FE_RC_3752_0 ( .a(n_40649), .b(n_40637), .c(n_40655), .o(n_40659) );
oa22f04 FE_RC_3759_0 ( .a(n_37060), .b(n_37509), .c(n_37059), .d(FE_OCP_RBN2482_n_37509), .o(n_37606) );
in01s06 FE_RC_3761_0 ( .a(n_32572), .o(FE_RN_1639_0) );
na02m08 FE_RC_3762_0 ( .a(FE_OCP_RBN6519_n_32706), .b(FE_RN_1639_0), .o(FE_RN_1640_0) );
no02s01 TIMEBOOST_cell_1619 ( .a(n_47254), .b(n_34256), .o(TIMEBOOST_net_424) );
oa22m04 FE_RC_3764_0 ( .a(FE_OCP_RBN6752_n_30273), .b(n_30501), .c(n_30273), .d(n_30512), .o(n_30608) );
na02s01 TIMEBOOST_cell_2940 ( .a(n_18140), .b(n_18230), .o(TIMEBOOST_net_761) );
oa22m06 FE_RC_3766_0 ( .a(n_12681), .b(n_13410), .c(n_12682), .d(n_13411), .o(n_13497) );
oa22m02 FE_RC_3767_0 ( .a(n_23414), .b(n_26171), .c(FE_OCPN1334_n_23467), .d(n_26200), .o(n_26320) );
in01s01 FE_RC_3768_0 ( .a(FE_RN_1641_0), .o(FE_RN_1642_0) );
in01s01 FE_RC_3769_0 ( .a(FE_RN_1642_0), .o(FE_OCPN1334_n_23467) );
oa22m02 FE_RC_3772_0 ( .a(n_17336), .b(n_17459), .c(n_17753), .d(n_17441), .o(n_17552) );
na02m40 FE_RC_3776_0 ( .a(n_45224), .b(FE_OCP_RBN3818_n_45622), .o(n_11774) );
na02m40 FE_RC_3777_0 ( .a(n_22597), .b(n_44061), .o(n_22708) );
in01s03 FE_RC_3778_0 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_2_), .o(FE_RN_1644_0) );
no02s06 FE_RC_3779_0 ( .a(n_45224), .b(FE_RN_1644_0), .o(FE_RN_1645_0) );
ao22s04 FE_RC_377_0 ( .a(n_6613), .b(n_6679), .c(n_6734), .d(n_6612), .o(n_6804) );
no02s10 FE_RC_3780_0 ( .a(n_11844), .b(FE_RN_1645_0), .o(n_11829) );
na02f04 TIMEBOOST_cell_1549 ( .a(n_8439), .b(n_8506), .o(TIMEBOOST_net_389) );
in01s20 FE_RC_3782_0 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_3_), .o(FE_RN_1646_0) );
no02m06 TIMEBOOST_cell_5652 ( .a(n_11257), .b(n_11244), .o(TIMEBOOST_net_1774) );
no03m08 TIMEBOOST_cell_2276 ( .a(n_33135), .b(n_33186), .c(n_33181), .o(FE_RN_1994_0) );
na02s20 FE_RC_3785_0 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_3_), .b(FE_OCP_RBN7008_n_44962), .o(FE_RN_1648_0) );
na02m20 FE_RC_3786_0 ( .a(n_32433), .b(FE_RN_1648_0), .o(n_32472) );
in01s03 FE_RC_3791_0 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_4_), .o(FE_RN_1651_0) );
no02m08 TIMEBOOST_cell_1620 ( .a(n_34727), .b(TIMEBOOST_net_424), .o(n_34829) );
no02s02 TIMEBOOST_cell_6930 ( .a(TIMEBOOST_net_2223), .b(n_2392), .o(TIMEBOOST_net_1493) );
in01m06 FE_RC_3796_0 ( .a(n_23000), .o(FE_RN_1654_0) );
ao22f08 FE_RC_3797_0 ( .a(FE_RN_1654_0), .b(FE_OCP_RBN5543_n_23044), .c(n_23000), .d(n_45311), .o(n_23193) );
in01s01 FE_RC_3798_0 ( .a(FE_RN_1656_0), .o(FE_RN_1655_0) );
no02s01 FE_RC_3799_0 ( .a(FE_RN_1655_0), .b(n_23170), .o(n_23334) );
in01s04 FE_RC_3800_0 ( .a(n_23170), .o(FE_RN_1657_0) );
no02f08 TIMEBOOST_cell_2927 ( .a(n_29232), .b(TIMEBOOST_net_754), .o(n_29349) );
in01s02 FE_RC_3805_0 ( .a(n_12017), .o(FE_RN_1659_0) );
na02s10 FE_RC_3806_0 ( .a(n_12352), .b(FE_RN_1659_0), .o(FE_RN_1660_0) );
in01s02 FE_RC_3807_0 ( .a(n_12017), .o(FE_RN_1661_0) );
oa12s10 FE_RC_3808_0 ( .a(FE_RN_1660_0), .b(FE_RN_1661_0), .c(n_12352), .o(n_12428) );
in01s01 FE_RC_3809_0 ( .a(n_11863), .o(FE_RN_1662_0) );
in01s01 FE_RC_380_0 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_3_), .o(FE_RN_114_0) );
na02s01 FE_RC_3810_0 ( .a(FE_RN_1662_0), .b(FE_RN_1664_0), .o(FE_RN_1663_0) );
no02f08 FE_RC_3811_0 ( .a(FE_RN_1663_0), .b(n_12449), .o(n_12459) );
in01s01 FE_RC_3812_0 ( .a(n_11960), .o(FE_RN_1665_0) );
in01s01 FE_RC_3813_0 ( .a(FE_RN_1665_0), .o(FE_RN_1664_0) );
in01s01 FE_RC_3814_0 ( .a(n_23571), .o(FE_RN_1666_0) );
in01s01 FE_RC_3815_0 ( .a(n_23826), .o(FE_RN_1667_0) );
na02s02 TIMEBOOST_cell_7844 ( .a(n_35343), .b(n_35340), .o(TIMEBOOST_net_2553) );
no02s01 TIMEBOOST_cell_1898 ( .a(TIMEBOOST_net_563), .b(n_17081), .o(n_17134) );
in01f04 FE_RC_3818_0 ( .a(n_23637), .o(FE_RN_1669_0) );
no02f04 FE_RC_3819_0 ( .a(n_23542), .b(n_23571), .o(FE_RN_1670_0) );
in01s01 FE_RC_381_0 ( .a(FE_OCP_RBN6439_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_RN_115_0) );
na02f04 FE_RC_3820_0 ( .a(FE_RN_1670_0), .b(n_23626), .o(FE_RN_1671_0) );
na02f06 FE_RC_3821_0 ( .a(FE_RN_1669_0), .b(FE_RN_1671_0), .o(FE_RN_1672_0) );
in01m04 FE_RC_3822_0 ( .a(n_23626), .o(FE_RN_1673_0) );
na03s20 TIMEBOOST_cell_8694 ( .a(n_32688), .b(n_32623), .c(FE_OCP_RBN4633_n_44962), .o(TIMEBOOST_net_2834) );
no02s01 TIMEBOOST_cell_1907 ( .a(FE_OCP_RBN1845_n_30492), .b(n_31599), .o(TIMEBOOST_net_568) );
no02s06 FE_RC_382_0 ( .a(FE_RN_114_0), .b(FE_RN_115_0), .o(FE_RN_116_0) );
in01s01 FE_RC_3833_0 ( .a(FE_RN_1070_0), .o(FE_RN_1680_0) );
in01m02 FE_RC_3834_0 ( .a(n_24323), .o(FE_RN_1681_0) );
na02s01 TIMEBOOST_cell_2024 ( .a(n_19274), .b(TIMEBOOST_net_626), .o(n_19416) );
no04s03 TIMEBOOST_cell_7367 ( .a(n_25032), .b(n_25090), .c(n_25033), .d(n_25083), .o(TIMEBOOST_net_2085) );
no02s06 FE_RC_383_0 ( .a(n_6716), .b(FE_RN_116_0), .o(n_6598) );
in01s01 FE_RC_3840_0 ( .a(n_19637), .o(n_19621) );
na02s02 FE_RC_3841_0 ( .a(n_19637), .b(n_19617), .o(n_19690) );
in01f04 FE_RC_3846_0 ( .a(FE_RN_959_0), .o(n_20186) );
in01f02 FE_RC_3848_0 ( .a(n_20186), .o(n_20188) );
na02f02 FE_RC_3849_0 ( .a(FE_OCP_RBN6380_n_20125), .b(FE_RN_959_0), .o(n_20189) );
in01s01 FE_RC_384_0 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_3_), .o(FE_RN_117_0) );
in01f01 FE_RC_3850_0 ( .a(n_20222), .o(FE_RN_1688_0) );
no02f02 FE_RC_3851_0 ( .a(FE_RN_1688_0), .b(n_20261), .o(n_20279) );
in01m01 FE_RC_3852_0 ( .a(n_20261), .o(FE_RN_1689_0) );
na02f02 FE_RC_3853_0 ( .a(FE_RN_1689_0), .b(n_20222), .o(n_20280) );
in01s01 FE_RC_385_0 ( .a(FE_OCP_RBN6439_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_RN_118_0) );
in01m02 FE_RC_3865_0 ( .a(FE_RN_1697_0), .o(n_21092) );
in01s01 FE_RC_3869_0 ( .a(n_22705), .o(n_44364) );
na02m08 TIMEBOOST_cell_3854 ( .a(TIMEBOOST_net_1017), .b(n_23504), .o(n_23581) );
in01s01 FE_RC_3870_0 ( .a(n_22463), .o(FE_RN_1699_0) );
no02s02 FE_RC_3871_0 ( .a(n_22705), .b(FE_RN_1699_0), .o(FE_RN_1700_0) );
no02s02 FE_RC_3872_0 ( .a(FE_RN_1700_0), .b(n_22370), .o(n_22744) );
oa22f08 FE_RC_3880_0 ( .a(n_16745), .b(n_16801), .c(FE_OCP_RBN5322_n_16745), .d(n_16802), .o(n_16987) );
oa22f04 FE_RC_3882_0 ( .a(FE_OCP_RBN2820_n_13962), .b(n_14763), .c(FE_OCP_RBN5777_n_13796), .d(FE_OCP_RBN1597_n_14763), .o(n_14872) );
oa22f04 FE_RC_3884_0 ( .a(n_28677), .b(FE_RN_1738_0), .c(n_28676), .d(FE_OCP_RBN7024_FE_RN_1738_0), .o(n_29054) );
ao22m06 FE_RC_3885_0 ( .a(n_23689), .b(n_24072), .c(n_23690), .d(n_24043), .o(n_24102) );
oa22f04 FE_RC_3887_0 ( .a(n_24469), .b(n_44621), .c(FE_OCP_RBN2693_n_24436), .d(n_24862), .o(n_24945) );
ao22f04 FE_RC_3891_0 ( .a(n_20690), .b(n_20730), .c(n_20647), .d(n_20731), .o(n_20886) );
oa22f04 FE_RC_3892_0 ( .a(FE_OCPN1677_n_27062), .b(FE_OCP_RBN1856_n_30731), .c(FE_OFN1196_n_27014), .d(n_30731), .o(n_30847) );
oa22f02 FE_RC_3893_0 ( .a(FE_OCPN5294_n_30584), .b(n_30747), .c(FE_OCP_RBN2107_n_30747), .d(n_27014), .o(n_30769) );
ao22f02 FE_RC_3894_0 ( .a(n_45070), .b(FE_OCP_RBN6382_n_21087), .c(n_45023), .d(n_21087), .o(n_21233) );
na03s10 FE_RC_389_0 ( .a(n_30021), .b(n_29952), .c(n_29956), .o(n_30022) );
oa22s04 FE_RC_3900_0 ( .a(n_31827), .b(n_32220), .c(n_31828), .d(n_32219), .o(n_32310) );
oa22s02 FE_RC_3901_0 ( .a(n_32122), .b(n_32360), .c(n_32123), .d(n_44213), .o(n_32516) );
oa22m10 FE_RC_3903_0 ( .a(n_17072), .b(n_17192), .c(n_17020), .d(n_17073), .o(n_17340) );
oa22f08 FE_RC_3905_0 ( .a(n_27868), .b(n_27825), .c(n_27751), .d(FE_OCP_RBN1804_n_27825), .o(n_28009) );
oa22m02 FE_RC_3906_0 ( .a(n_12500), .b(n_12690), .c(n_12501), .d(n_12691), .o(n_12771) );
ao22m04 FE_RC_3907_0 ( .a(n_18219), .b(FE_OCP_RBN2043_n_18269), .c(n_18218), .d(FE_OCP_RBN2042_n_18269), .o(n_18375) );
ao22f04 FE_RC_3909_0 ( .a(n_19222), .b(FE_OCP_RBN4082_n_18899), .c(FE_OFN739_n_17093), .d(n_18899), .o(n_19005) );
oa22m04 FE_RC_3912_0 ( .a(n_18538), .b(n_19281), .c(n_18537), .d(n_19280), .o(n_19390) );
ao22f02 FE_RC_3913_0 ( .a(FE_OCP_RBN1019_n_24165), .b(n_24312), .c(n_25265), .d(n_24311), .o(n_24503) );
oa22m02 FE_RC_3918_0 ( .a(FE_OFN748_n_22641), .b(n_25933), .c(FE_RN_1793_0), .d(n_25934), .o(n_26097) );
oa22f02 FE_RC_3919_0 ( .a(n_25971), .b(FE_OCP_RBN1862_n_26049), .c(n_26004), .d(n_26049), .o(n_26267) );
oa22m04 FE_RC_391_0 ( .a(n_32128), .b(FE_OCP_RBN1877_n_32382), .c(n_32129), .d(n_32382), .o(n_32546) );
oa22f02 FE_RC_3925_0 ( .a(FE_OCP_RBN7057_n_36677), .b(n_36738), .c(n_36677), .d(n_36737), .o(n_36782) );
ao22m04 FE_RC_3926_0 ( .a(n_32134), .b(n_45754), .c(n_32135), .d(n_45755), .o(n_32395) );
oa22f02 FE_RC_3927_0 ( .a(n_36797), .b(n_36842), .c(n_36796), .d(n_36831), .o(n_36885) );
no02s01 TIMEBOOST_cell_6675 ( .a(FE_OCP_RBN5394_cordic_combinational_sub_ln23_0_unr12_z_0_), .b(FE_OCP_RBN5392_cordic_combinational_sub_ln23_0_unr12_z_0_), .o(TIMEBOOST_net_2095) );
na03s01 TIMEBOOST_cell_8287 ( .a(n_44102), .b(FE_OCP_RBN5629_n_33976), .c(n_34303), .o(n_34452) );
in01s02 FE_RC_392_0 ( .a(n_15187), .o(FE_RN_120_0) );
na02s80 FE_RC_3930_0 ( .a(n_32564), .b(n_44962), .o(n_32632) );
na02m20 FE_RC_3931_0 ( .a(n_32564), .b(n_44962), .o(FE_RN_1702_0) );
na02m10 FE_RC_3932_0 ( .a(FE_RN_1702_0), .b(FE_RN_1426_0), .o(n_32647) );
oa22m08 FE_RC_3936_0 ( .a(n_22820), .b(n_22746), .c(FE_OCP_RBN2385_n_22820), .d(n_22747), .o(n_22899) );
in01m02 FE_RC_393_0 ( .a(n_15434), .o(FE_RN_121_0) );
na02m04 FE_RC_394_0 ( .a(FE_RN_121_0), .b(FE_RN_120_0), .o(FE_RN_122_0) );
in01s01 FE_RC_3950_0 ( .a(FE_RN_1715_0), .o(FE_RN_1714_0) );
no02s01 FE_RC_3951_0 ( .a(n_32835), .b(FE_RN_1714_0), .o(n_33168) );
in01s04 FE_RC_3952_0 ( .a(n_32835), .o(FE_RN_1716_0) );
na02s01 FE_RC_3956_0 ( .a(FE_RN_1717_0), .b(FE_RN_650_0), .o(n_33484) );
na02s01 FE_RC_3957_0 ( .a(FE_RN_1717_0), .b(FE_RN_650_0), .o(FE_RN_1718_0) );
no02s01 FE_RC_3958_0 ( .a(n_33135), .b(FE_RN_1718_0), .o(n_33501) );
na02f06 FE_RC_395_0 ( .a(FE_RN_122_0), .b(n_15475), .o(n_46982) );
na02s08 TIMEBOOST_cell_4897 ( .a(n_12234), .b(TIMEBOOST_net_1396), .o(n_12298) );
na03s02 TIMEBOOST_cell_4912 ( .a(n_40934), .b(n_40878), .c(n_40928), .o(TIMEBOOST_net_1404) );
in01m03 FE_RC_3966_0 ( .a(FE_RN_1722_0), .o(n_18339) );
no02m02 FE_RC_3967_0 ( .a(n_47248), .b(n_19014), .o(FE_RN_1722_0) );
in01s01 FE_RC_3979_0 ( .a(n_28548), .o(FE_RN_1733_0) );
in01s01 FE_RC_3980_0 ( .a(n_28632), .o(FE_RN_1734_0) );
no02s02 FE_RC_3981_0 ( .a(FE_RN_1733_0), .b(FE_RN_1734_0), .o(FE_RN_1735_0) );
in01s01 FE_RC_3982_0 ( .a(n_28609), .o(FE_RN_1736_0) );
na02f04 FE_RC_3983_0 ( .a(n_28894), .b(FE_RN_1736_0), .o(FE_RN_1737_0) );
na02f06 FE_RC_3985_0 ( .a(FE_RN_1737_0), .b(FE_RN_1735_0), .o(FE_RN_1738_0) );
in01s01 FE_RC_3990_0 ( .a(n_33196), .o(FE_RN_1741_0) );
in01f04 FE_RC_3991_0 ( .a(n_33648), .o(FE_RN_1742_0) );
na02f08 FE_RC_3992_0 ( .a(FE_RN_1741_0), .b(FE_RN_1742_0), .o(FE_RN_1743_0) );
na02f08 FE_RC_3993_0 ( .a(FE_RN_1743_0), .b(FE_RN_1045_0), .o(n_33735) );
in01s02 FE_RC_3994_0 ( .a(n_13010), .o(FE_RN_1744_0) );
oa22f06 FE_RC_3996_0 ( .a(n_18509), .b(n_18956), .c(n_18510), .d(n_18955), .o(n_19064) );
ao22m04 FE_RC_3997_0 ( .a(n_13154), .b(FE_OCP_RBN2554_n_13141), .c(n_13141), .d(FE_OCP_RBN2579_n_13154), .o(n_13331) );
ao22f04 FE_RC_4003_0 ( .a(n_17815), .b(FE_OCP_RBN7031_n_18981), .c(n_17783), .d(n_18981), .o(n_19075) );
in01s02 FE_RC_4004_0 ( .a(FE_OCPN1253_n_23815), .o(FE_RN_1748_0) );
no02m08 FE_RC_4005_0 ( .a(n_24274), .b(FE_RN_1748_0), .o(n_24325) );
na02f06 FE_RC_4007_0 ( .a(n_29318), .b(FE_RN_1750_0), .o(n_29389) );
in01s01 FE_RC_4008_0 ( .a(FE_OCP_DRV_N1889_n_29317), .o(FE_RN_1750_0) );
no02m04 FE_RC_4009_0 ( .a(n_29318), .b(FE_RN_1750_0), .o(n_29340) );
in01s03 FE_RC_400_0 ( .a(n_28001), .o(FE_RN_123_0) );
oa22f04 FE_RC_4010_0 ( .a(FE_OFN773_n_25834), .b(FE_OCP_RBN2610_n_29298), .c(n_29379), .d(n_29298), .o(n_29399) );
na02m06 FE_RC_4011_0 ( .a(FE_OCP_RBN4112_n_12880), .b(n_13497), .o(FE_RN_1751_0) );
na02f08 FE_RC_4012_0 ( .a(FE_RN_1751_0), .b(n_13529), .o(n_13599) );
in01s01 FE_RC_4015_0 ( .a(FE_OCPN1728_n_34096), .o(FE_RN_1753_0) );
no02s06 FE_RC_4016_0 ( .a(FE_RN_1753_0), .b(n_34097), .o(n_34114) );
na02f08 FE_RC_4017_0 ( .a(n_41924), .b(n_41941), .o(FE_RN_1754_0) );
na02f08 FE_RC_4018_0 ( .a(FE_RN_1754_0), .b(n_41789), .o(n_41995) );
in01s03 FE_RC_401_0 ( .a(n_28226), .o(FE_RN_124_0) );
no02s02 TIMEBOOST_cell_1911 ( .a(FE_OCPN6931_n_22156), .b(FE_OCP_RBN4462_n_44267), .o(TIMEBOOST_net_570) );
na02s01 TIMEBOOST_cell_5284 ( .a(FE_OCP_RBN4351_n_20456), .b(FE_OCP_RBN2711_n_19599), .o(TIMEBOOST_net_1590) );
in01s01 FE_RC_4023_0 ( .a(FE_OCPN1696_n_13721), .o(FE_RN_1757_0) );
na02m06 FE_RC_4024_0 ( .a(FE_RN_1757_0), .b(n_13722), .o(n_13753) );
in01s01 FE_RC_4025_0 ( .a(n_23874), .o(FE_RN_1758_0) );
na02f08 FE_RC_4026_0 ( .a(FE_RN_1758_0), .b(n_24566), .o(n_24598) );
na02f04 FE_RC_4027_0 ( .a(n_13625), .b(n_13538), .o(FE_RN_1760_0) );
no02f04 FE_RC_4028_0 ( .a(FE_RN_1760_0), .b(n_13606), .o(FE_RN_1761_0) );
no02f04 FE_RC_4029_0 ( .a(n_13608), .b(n_13606), .o(FE_RN_1762_0) );
na02s06 FE_RC_402_0 ( .a(FE_RN_123_0), .b(FE_RN_124_0), .o(FE_RN_125_0) );
in01s01 FE_RC_4031_0 ( .a(n_13625), .o(FE_RN_1763_0) );
in01s01 FE_RC_4032_0 ( .a(FE_RN_1763_0), .o(FE_RN_1759_0) );
in01s01 FE_RC_4034_0 ( .a(n_19537), .o(FE_RN_1764_0) );
na02s02 FE_RC_4035_0 ( .a(FE_RN_1764_0), .b(n_19528), .o(n_19597) );
in01m02 FE_RC_4036_0 ( .a(n_24719), .o(FE_RN_1765_0) );
in01f04 FE_RC_4039_0 ( .a(FE_RN_1766_0), .o(n_20029) );
no02f04 TIMEBOOST_cell_1668 ( .a(TIMEBOOST_net_448), .b(n_26128), .o(n_26083) );
na02f02 FE_RC_4040_0 ( .a(FE_OCP_RBN5029_n_18678), .b(n_19922), .o(FE_RN_1766_0) );
na02f04 TIMEBOOST_cell_7825 ( .a(TIMEBOOST_net_2543), .b(n_26100), .o(n_26140) );
ao22f06 FE_RC_4043_0 ( .a(FE_OCP_RBN1833_n_14197), .b(n_14246), .c(n_14153), .d(n_14248), .o(n_14450) );
in01s01 FE_RC_4055_0 ( .a(n_8799), .o(FE_RN_1774_0) );
no02s04 TIMEBOOST_cell_1984 ( .a(n_33411), .b(TIMEBOOST_net_606), .o(n_33494) );
no02s01 TIMEBOOST_cell_8628 ( .a(FE_OCP_RBN3307_n_43022), .b(n_42953), .o(TIMEBOOST_net_2801) );
no02f04 FE_RC_4060_0 ( .a(FE_RN_1775_0), .b(FE_RN_1778_0), .o(n_9125) );
in01s01 FE_RC_4061_0 ( .a(FE_OCP_RBN1134_n_19077), .o(FE_RN_1779_0) );
na02s02 FE_RC_4062_0 ( .a(n_20372), .b(FE_RN_1779_0), .o(n_20469) );
in01s02 FE_RC_4063_0 ( .a(n_35012), .o(FE_RN_1780_0) );
in01f02 FE_RC_4064_0 ( .a(n_35078), .o(FE_RN_1781_0) );
in01s01 FE_RC_4069_0 ( .a(FE_OCPN1391_n_15462), .o(FE_RN_1784_0) );
na02f06 FE_RC_4070_0 ( .a(FE_RN_1784_0), .b(n_15463), .o(n_15497) );
ao22f06 FE_RC_4079_0 ( .a(n_42481), .b(n_42887), .c(n_42480), .d(n_42886), .o(n_42947) );
no03s10 TIMEBOOST_cell_7113 ( .a(TIMEBOOST_net_1828), .b(n_17189), .c(n_17126), .o(n_17479) );
in01s01 FE_RC_4080_0 ( .a(n_34870), .o(FE_RN_1789_0) );
no02s08 FE_RC_4081_0 ( .a(FE_OCP_RBN6048_n_35487), .b(FE_RN_1789_0), .o(n_35690) );
na02s01 FE_RC_4083_0 ( .a(n_34894), .b(FE_RN_1790_0), .o(FE_RN_1791_0) );
na02s06 FE_RC_4084_0 ( .a(FE_OCP_RBN3168_n_44211), .b(FE_RN_1791_0), .o(n_35683) );
in01s01 FE_RC_4085_0 ( .a(n_34947), .o(FE_RN_1792_0) );
in01s01 FE_RC_4086_0 ( .a(FE_RN_1792_0), .o(FE_RN_1790_0) );
in01s01 FE_RC_4087_0 ( .a(FE_OFN748_n_22641), .o(FE_RN_1793_0) );
in01m04 FE_RC_408_0 ( .a(n_28292), .o(FE_RN_127_0) );
na02f04 TIMEBOOST_cell_5659 ( .a(TIMEBOOST_net_1777), .b(n_11326), .o(n_11411) );
no02s01 TIMEBOOST_cell_3382 ( .a(FE_OCP_RBN6872_n_31520), .b(n_31017), .o(TIMEBOOST_net_982) );
in01s01 FE_RC_4092_0 ( .a(FE_OCPUNCON3485_n_31012), .o(FE_RN_1796_0) );
no02f04 FE_RC_4093_0 ( .a(n_31013), .b(FE_RN_1796_0), .o(n_31086) );
in01s01 FE_RC_4094_0 ( .a(FE_OCPUNCON3485_n_31012), .o(FE_RN_1797_0) );
na02f04 FE_RC_4095_0 ( .a(n_31013), .b(FE_RN_1797_0), .o(n_31035) );
no03f08 FE_RC_4096_0 ( .a(n_26306), .b(n_26225), .c(n_26217), .o(n_26378) );
na02m02 FE_RC_4097_0 ( .a(n_26292), .b(n_26218), .o(FE_RN_1798_0) );
no02f04 FE_RC_4098_0 ( .a(n_26378), .b(FE_RN_1798_0), .o(n_26445) );
in01f06 FE_RC_409_0 ( .a(FE_RN_128_0), .o(n_28348) );
in01s01 FE_RC_4102_0 ( .a(FE_RN_1184_0), .o(n_21794) );
na02m02 TIMEBOOST_cell_7973 ( .a(TIMEBOOST_net_2617), .b(n_4143), .o(n_4720) );
na02f06 FE_RC_4111_0 ( .a(n_39689), .b(n_39717), .o(FE_RN_1805_0) );
na02f08 FE_RC_4112_0 ( .a(FE_RN_1805_0), .b(n_39724), .o(n_39750) );
in01s01 FE_RC_4128_0 ( .a(FE_OCPN1671_n_39371), .o(FE_RN_1818_0) );
na02s10 FE_RC_4129_0 ( .a(n_39812), .b(FE_RN_1818_0), .o(n_39866) );
in01s01 FE_RC_4130_0 ( .a(n_43256), .o(FE_RN_1819_0) );
in01s01 FE_RC_4131_0 ( .a(n_43692), .o(FE_RN_1820_0) );
na02s06 FE_RC_4132_0 ( .a(FE_RN_1820_0), .b(FE_RN_1819_0), .o(FE_RN_1821_0) );
no02f08 FE_RC_4133_0 ( .a(n_43664), .b(FE_RN_1821_0), .o(n_43721) );
ao22m04 FE_RC_4135_0 ( .a(FE_RN_1270_0), .b(n_36481), .c(FE_RN_1271_0), .d(n_36514), .o(n_36545) );
na02s02 TIMEBOOST_cell_3836 ( .a(TIMEBOOST_net_1008), .b(FE_RN_783_0), .o(FE_RN_785_0) );
no02s01 FE_RC_4138_0 ( .a(n_40042), .b(n_40001), .o(FE_RN_1822_0) );
na02f08 FE_RC_4139_0 ( .a(FE_RN_1822_0), .b(n_40422), .o(n_40466) );
oa22s01 FE_RC_4140_0 ( .a(n_36720), .b(n_36734), .c(n_36721), .d(n_36733), .o(n_36776) );
na02s02 FE_RC_4141_0 ( .a(n_40069), .b(n_40073), .o(FE_RN_1823_0) );
no02s06 FE_RC_4142_0 ( .a(FE_RN_1823_0), .b(n_40113), .o(FE_RN_1824_0) );
na02f10 FE_RC_4143_0 ( .a(FE_RN_1824_0), .b(n_40472), .o(n_40524) );
oa22m02 FE_RC_4144_0 ( .a(n_36763), .b(n_36894), .c(n_36764), .d(n_36867), .o(n_36895) );
oa22m02 FE_RC_4145_0 ( .a(n_40598), .b(n_40579), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .d(n_44958), .o(n_40587) );
in01s01 FE_RC_4147_0 ( .a(n_18356), .o(FE_RN_1825_0) );
in01s04 FE_RC_4148_0 ( .a(n_18339), .o(FE_RN_1826_0) );
na02m08 FE_RC_4149_0 ( .a(FE_RN_1826_0), .b(FE_RN_1825_0), .o(FE_RN_1827_0) );
no02m10 FE_RC_4150_0 ( .a(FE_OCP_RBN5032_n_18951), .b(FE_RN_1827_0), .o(n_19088) );
oa22f02 FE_RC_4153_0 ( .a(FE_OCPN869_n_45003), .b(FE_OCP_RBN5208_n_20412), .c(n_45065), .d(n_20412), .o(n_20542) );
oa22f04 FE_RC_4154_0 ( .a(FE_OCPN869_n_45003), .b(FE_OCP_RBN4644_n_20420), .c(n_45065), .d(n_20420), .o(n_20549) );
ao22m04 FE_RC_4157_0 ( .a(n_22038), .b(FE_OCP_RBN5212_n_21987), .c(n_22039), .d(n_21987), .o(n_22068) );
no02f04 TIMEBOOST_cell_4370 ( .a(TIMEBOOST_net_1275), .b(n_8739), .o(n_8786) );
oa22f04 FE_RC_415_0 ( .a(FE_OCP_RBN6649_n_13818), .b(n_14052), .c(FE_OCP_RBN6646_n_13818), .d(n_14088), .o(n_14278) );
ao22f04 FE_RC_4161_0 ( .a(n_19264), .b(n_19748), .c(n_19301), .d(n_19749), .o(n_19894) );
oa22f04 FE_RC_4162_0 ( .a(n_20226), .b(FE_OCP_RBN1836_n_20209), .c(n_20241), .d(n_20209), .o(n_20336) );
oa22m04 FE_RC_4164_0 ( .a(n_35307), .b(n_35532), .c(n_35323), .d(n_35499), .o(n_35595) );
oa22f04 FE_RC_4169_0 ( .a(n_22492), .b(n_22573), .c(n_22493), .d(n_22593), .o(n_22750) );
na02m08 TIMEBOOST_cell_1800 ( .a(TIMEBOOST_net_514), .b(n_30355), .o(n_30452) );
ao22f02 FE_RC_4177_0 ( .a(n_20540), .b(FE_OCP_RBN5330_n_20678), .c(n_20500), .d(n_20678), .o(n_20877) );
na02s10 FE_RC_4183_0 ( .a(n_44365), .b(FE_OCP_RBN7118_delay_xor_ln22_unr12_stage5_stallmux_q_0_), .o(n_16745) );
in01s04 FE_RC_4184_0 ( .a(FE_RN_1828_0), .o(n_12097) );
na02s04 FE_RC_4185_0 ( .a(n_11941), .b(delay_add_ln22_unr8_stage4_stallmux_q_2_), .o(FE_RN_1828_0) );
in01s02 FE_RC_4186_0 ( .a(n_11991), .o(FE_RN_1829_0) );
in01s02 FE_RC_4187_0 ( .a(n_11908), .o(FE_RN_1830_0) );
no02f08 TIMEBOOST_cell_1760 ( .a(TIMEBOOST_net_494), .b(n_39526), .o(n_39577) );
no02s02 TIMEBOOST_cell_1701 ( .a(n_3758), .b(n_3529), .o(TIMEBOOST_net_465) );
no02m06 TIMEBOOST_cell_1670 ( .a(TIMEBOOST_net_449), .b(n_31158), .o(n_31239) );
in01m04 FE_RC_4195_0 ( .a(FE_RN_1834_0), .o(n_12420) );
no02m04 FE_RC_4196_0 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_10_), .b(n_12350), .o(FE_RN_1834_0) );
ao22s02 FE_RC_419_0 ( .a(FE_OCP_RBN6524_n_6649), .b(n_6571), .c(n_6642), .d(n_6649), .o(n_6759) );
in01s01 FE_RC_4202_0 ( .a(n_6887), .o(FE_RN_1838_0) );
no02s01 FE_RC_4203_0 ( .a(n_6826), .b(FE_RN_1838_0), .o(FE_RN_1839_0) );
na02s02 FE_RC_4204_0 ( .a(FE_RN_1839_0), .b(FE_RN_816_0), .o(FE_RN_1840_0) );
oa22s02 FE_RC_420_0 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(FE_OCP_RBN5435_delay_xor_ln22_unr6_stage3_stallmux_q_0_), .d(FE_OCP_RBN5434_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6654) );
in01s01 FE_RC_4210_0 ( .a(n_18595), .o(FE_RN_1844_0) );
in01s01 FE_RC_4211_0 ( .a(FE_RN_1844_0), .o(FE_RN_1842_0) );
in01s02 FE_RC_4212_0 ( .a(n_23881), .o(FE_RN_1845_0) );
no02s06 FE_RC_4213_0 ( .a(FE_RN_1845_0), .b(n_24208), .o(FE_RN_1846_0) );
ao12s06 FE_RC_4215_0 ( .a(FE_RN_1846_0), .b(FE_RN_1845_0), .c(n_24208), .o(n_24293) );
in01s01 FE_RC_4218_0 ( .a(FE_OCPN1377_n_17836), .o(FE_RN_1849_0) );
na02f04 FE_RC_4219_0 ( .a(FE_RN_1849_0), .b(n_19243), .o(n_19318) );
in01m06 FE_RC_421_0 ( .a(n_28229), .o(FE_RN_129_0) );
oa22f04 FE_RC_4228_0 ( .a(n_13626), .b(FE_RN_1761_0), .c(FE_RN_1759_0), .d(FE_RN_1762_0), .o(n_13683) );
in01s02 FE_RC_422_0 ( .a(n_28230), .o(FE_RN_130_0) );
oa22m06 FE_RC_4230_0 ( .a(n_7514), .b(n_8476), .c(n_7513), .d(n_8461), .o(n_8599) );
in01s01 FE_RC_4231_0 ( .a(n_13148), .o(FE_RN_1855_0) );
in01s04 FE_RC_4232_0 ( .a(FE_RN_1856_0), .o(n_14511) );
no02m04 FE_RC_4233_0 ( .a(FE_RN_1855_0), .b(n_14372), .o(FE_RN_1856_0) );
ao22f06 FE_RC_4234_0 ( .a(n_14821), .b(n_14747), .c(n_14439), .d(n_14746), .o(n_14865) );
ao22f06 FE_RC_4235_0 ( .a(FE_OCP_RBN6701_n_14444), .b(n_14913), .c(n_14912), .d(FE_OCP_RBN6703_n_14444), .o(n_15021) );
in01s01 FE_RC_4236_0 ( .a(n_20321), .o(n_20349) );
na02m10 TIMEBOOST_cell_975 ( .a(FE_RN_1299_0), .b(FE_OCP_RBN6527_n_44962), .o(TIMEBOOST_net_102) );
in01s01 FE_RC_4238_0 ( .a(n_38930), .o(FE_RN_1857_0) );
na02s04 FE_RC_4239_0 ( .a(FE_RN_1857_0), .b(n_38847), .o(n_38951) );
no02s01 TIMEBOOST_cell_8663 ( .a(TIMEBOOST_net_2818), .b(n_31706), .o(n_31743) );
no02s01 FE_RC_4240_0 ( .a(FE_RN_1858_0), .b(FE_RN_1859_0), .o(FE_RN_1860_0) );
no02s06 FE_RC_4241_0 ( .a(FE_RN_1860_0), .b(FE_OCP_RBN4328_n_38878), .o(n_39026) );
in01s01 FE_RC_4242_0 ( .a(n_38564), .o(FE_RN_1861_0) );
in01s01 FE_RC_4243_0 ( .a(FE_RN_1861_0), .o(FE_RN_1859_0) );
in01s01 FE_RC_4244_0 ( .a(n_38562), .o(FE_RN_1862_0) );
in01s01 FE_RC_4245_0 ( .a(FE_RN_1862_0), .o(FE_RN_1858_0) );
in01m03 FE_RC_4247_0 ( .a(FE_RN_1863_0), .o(n_9928) );
na02m02 FE_RC_4248_0 ( .a(FE_OCP_RBN6678_n_8288), .b(n_9704), .o(FE_RN_1863_0) );
na03s02 TIMEBOOST_cell_6027 ( .a(n_18841), .b(n_18840), .c(n_18839), .o(TIMEBOOST_net_1865) );
na02m02 FE_RC_4251_0 ( .a(n_8750), .b(n_9724), .o(FE_RN_1865_0) );
na02f06 FE_RC_4254_0 ( .a(n_35377), .b(n_35360), .o(FE_RN_1867_0) );
na02f08 FE_RC_4255_0 ( .a(FE_RN_1867_0), .b(n_35375), .o(n_35467) );
no02m02 FE_RC_4257_0 ( .a(n_20721), .b(n_20638), .o(n_20759) );
no02m02 TIMEBOOST_cell_1679 ( .a(FE_OCP_RBN4240_n_44594), .b(n_9169), .o(TIMEBOOST_net_454) );
in01s01 FE_RC_4265_0 ( .a(FE_OCP_RBN2892_n_14460), .o(FE_RN_1872_0) );
no02f04 FE_RC_4266_0 ( .a(FE_RN_1872_0), .b(n_16218), .o(n_16272) );
in01s03 FE_RC_4267_0 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(FE_RN_1873_0) );
in01f08 FE_RC_4268_0 ( .a(FE_RN_1874_0), .o(n_39656) );
na02m04 TIMEBOOST_cell_2043 ( .a(n_41941), .b(n_41785), .o(TIMEBOOST_net_636) );
in01m02 FE_RC_4270_0 ( .a(n_26196), .o(FE_RN_1875_0) );
no02f01 FE_RC_4271_0 ( .a(n_23414), .b(FE_RN_1875_0), .o(FE_RN_1876_0) );
no02f02 FE_RC_4272_0 ( .a(n_26359), .b(FE_RN_1876_0), .o(n_26390) );
in01m02 FE_RC_4273_0 ( .a(n_26202), .o(FE_RN_1877_0) );
na02f04 FE_RC_4274_0 ( .a(n_26445), .b(FE_RN_1877_0), .o(FE_RN_1878_0) );
oa12f04 FE_RC_4276_0 ( .a(FE_RN_1878_0), .b(FE_RN_1877_0), .c(n_26445), .o(n_26627) );
in01s01 FE_RC_4285_0 ( .a(n_30572), .o(FE_RN_1885_0) );
in01s01 FE_RC_4286_0 ( .a(FE_RN_1885_0), .o(FE_RN_1883_0) );
na02s06 FE_RC_4288_0 ( .a(n_22553), .b(FE_RN_1886_0), .o(n_22591) );
in01m20 FE_RC_4294_0 ( .a(FE_OCPN1400_n_28095), .o(FE_RN_1888_0) );
in01s10 FE_RC_4295_0 ( .a(n_28092), .o(FE_RN_1889_0) );
na02m20 FE_RC_4296_0 ( .a(FE_RN_1888_0), .b(FE_RN_1889_0), .o(FE_RN_1890_0) );
na02s04 TIMEBOOST_cell_2817 ( .a(TIMEBOOST_net_699), .b(n_1648), .o(n_1742) );
no03s02 TIMEBOOST_cell_8262 ( .a(n_9089), .b(n_9112), .c(n_9113), .o(n_9314) );
ao22m04 FE_RC_4299_0 ( .a(FE_OCPN1709_FE_OFN739_n_17093), .b(n_19008), .c(n_17783), .d(n_19033), .o(n_19110) );
oa22s06 FE_RC_429_0 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_0_), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(FE_OCP_RBN6435_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .d(n_6510), .o(n_6590) );
in01s02 FE_RC_42_0 ( .a(n_17741), .o(FE_RN_12_0) );
ao22s04 FE_RC_4305_0 ( .a(n_23844), .b(n_24308), .c(n_23845), .d(n_24307), .o(n_24421) );
ao22s06 FE_RC_430_0 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n_6542), .c(delay_xor_ln21_unr6_stage3_stallmux_q_2_), .d(FE_OCP_RBN5434_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6616) );
in01s02 FE_RC_4312_0 ( .a(n_17669), .o(FE_RN_1894_0) );
in01s06 FE_RC_4313_0 ( .a(n_17642), .o(FE_RN_1895_0) );
no02m08 FE_RC_4314_0 ( .a(FE_RN_1894_0), .b(FE_RN_1895_0), .o(FE_RN_1896_0) );
na02m08 FE_RC_4315_0 ( .a(FE_RN_1896_0), .b(n_17579), .o(n_17797) );
oa22f08 FE_RC_4316_0 ( .a(FE_OCPN906_n_21956), .b(n_21904), .c(FE_OCPN904_n_21955), .d(n_21903), .o(n_21973) );
in01s01 FE_RC_4317_0 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_8_), .o(FE_RN_1897_0) );
in01s01 FE_RC_4318_0 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_7_), .o(FE_RN_1898_0) );
na02s01 FE_RC_4319_0 ( .a(FE_RN_1897_0), .b(FE_RN_1898_0), .o(FE_RN_1899_0) );
in01s02 FE_RC_431_0 ( .a(n_12581), .o(FE_RN_132_0) );
na02s01 FE_RC_4320_0 ( .a(FE_RN_1899_0), .b(n_1416), .o(n_1601) );
ao22f02 FE_RC_4326_0 ( .a(n_19372), .b(n_19818), .c(n_19342), .d(n_19819), .o(n_19922) );
ao22s02 FE_RC_4327_0 ( .a(n_1539), .b(FE_OCP_RBN5547_n_1733), .c(n_1540), .d(n_1733), .o(n_1822) );
oa22m02 FE_RC_4328_0 ( .a(n_18238), .b(n_18475), .c(n_18239), .d(n_18476), .o(n_18678) );
in01s01 FE_RC_4329_0 ( .a(n_1711), .o(FE_RN_1903_0) );
in01s01 FE_RC_432_0 ( .a(n_12590), .o(FE_RN_133_0) );
in01s01 FE_RC_4330_0 ( .a(n_1712), .o(FE_RN_1904_0) );
no02s02 TIMEBOOST_cell_1711 ( .a(n_15771), .b(n_15336), .o(TIMEBOOST_net_470) );
na03f04 TIMEBOOST_cell_4656 ( .a(FE_OCP_RBN1832_n_14197), .b(n_14153), .c(n_14247), .o(n_14412) );
ao22s02 FE_RC_4333_0 ( .a(n_1474), .b(FE_OCP_RBN2445_n_1675), .c(n_1475), .d(n_1675), .o(n_1727) );
oa22s02 FE_RC_4334_0 ( .a(FE_OCPN3544_n_1448), .b(FE_OCP_RBN6534_n_1577), .c(FE_OCPN3543_n_1448), .d(n_1577), .o(n_1660) );
no02f08 TIMEBOOST_cell_8757 ( .a(TIMEBOOST_net_2865), .b(n_14032), .o(n_14201) );
in01s01 FE_RC_4336_0 ( .a(n_2673), .o(FE_RN_1907_0) );
in01s02 FE_RC_4337_0 ( .a(FE_RN_1908_0), .o(n_2774) );
no02s01 TIMEBOOST_cell_2013 ( .a(n_24645), .b(n_23996), .o(TIMEBOOST_net_621) );
in01s01 FE_RC_4339_0 ( .a(FE_OCP_RBN5648_n_2438), .o(FE_RN_1909_0) );
no02s06 TIMEBOOST_cell_6846 ( .a(TIMEBOOST_net_2180), .b(FE_OCP_RBN6849_n_26358), .o(n_26596) );
in01s01 FE_RC_4340_0 ( .a(n_2746), .o(FE_RN_1910_0) );
no02s02 FE_RC_4341_0 ( .a(FE_RN_1909_0), .b(FE_RN_1910_0), .o(FE_RN_1911_0) );
no02s06 FE_RC_4342_0 ( .a(FE_RN_1911_0), .b(n_2821), .o(n_2840) );
oa22s01 FE_RC_4343_0 ( .a(n_928), .b(FE_OCPN839_n_44672), .c(n_875), .d(n_44637), .o(n_1316) );
oa22s02 FE_RC_4344_0 ( .a(n_1167), .b(FE_OCPN839_n_44672), .c(n_1154), .d(n_44637), .o(n_1314) );
oa22s01 FE_RC_4345_0 ( .a(n_1205), .b(n_44659), .c(n_1200), .d(n_44637), .o(n_1354) );
oa22s01 FE_RC_4346_0 ( .a(n_938), .b(n_44659), .c(FE_OFN1178_n_916), .d(n_44637), .o(n_1337) );
oa22s01 FE_RC_4347_0 ( .a(n_1217), .b(n_44659), .c(n_1216), .d(n_44637), .o(n_1336) );
oa22s02 FE_RC_4348_0 ( .a(n_966), .b(n_44659), .c(n_897), .d(n_44637), .o(n_1327) );
oa22s02 FE_RC_4349_0 ( .a(n_958), .b(n_44659), .c(n_918), .d(n_44637), .o(n_1307) );
no02s02 TIMEBOOST_cell_6907 ( .a(n_23681), .b(n_24067), .o(TIMEBOOST_net_2212) );
oa22s01 FE_RC_4350_0 ( .a(n_1132), .b(n_44652), .c(n_1106), .d(n_44637), .o(n_1350) );
oa22s01 FE_RC_4351_0 ( .a(n_1127), .b(n_44652), .c(n_1088), .d(n_44637), .o(n_1338) );
oa22s01 FE_RC_4352_0 ( .a(n_1189), .b(n_44652), .c(n_1179), .d(n_44637), .o(n_1334) );
oa22s01 FE_RC_4353_0 ( .a(n_1168), .b(n_44652), .c(n_1150), .d(n_44637), .o(n_1333) );
oa22s01 FE_RC_4354_0 ( .a(n_1004), .b(n_44652), .c(n_967), .d(n_44637), .o(n_1328) );
oa22s01 FE_RC_4355_0 ( .a(n_1206), .b(n_44652), .c(n_1201), .d(n_44637), .o(n_1312) );
oa22s01 FE_RC_4356_0 ( .a(n_1048), .b(n_44652), .c(n_998), .d(n_44637), .o(n_1309) );
oa22s02 FE_RC_4357_0 ( .a(n_1010), .b(n_44652), .c(n_993), .d(n_44637), .o(n_1301) );
oa22s01 FE_RC_4358_0 ( .a(n_1164), .b(n_44652), .c(n_1157), .d(n_44637), .o(n_1298) );
oa22m10 FE_RC_4359_0 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_1_), .b(FE_OCP_RBN7114_n_44365), .c(n_44365), .d(FE_OCP_RBN4593_delay_xor_ln22_unr12_stage5_stallmux_q_1_), .o(n_16801) );
in01m06 FE_RC_435_0 ( .a(n_28189), .o(FE_RN_135_0) );
ao22f04 FE_RC_4360_0 ( .a(n_18408), .b(FE_OCP_RBN7025_n_18873), .c(n_18407), .d(n_18873), .o(n_18986) );
oa22s02 FE_RC_4361_0 ( .a(n_2973), .b(n_4132), .c(n_2974), .d(n_4184), .o(n_4396) );
in01s01 FE_RC_4363_0 ( .a(n_4026), .o(FE_RN_1912_0) );
in01s01 FE_RC_4364_0 ( .a(n_4000), .o(FE_RN_1913_0) );
na02s01 TIMEBOOST_cell_4354 ( .a(TIMEBOOST_net_1267), .b(n_20657), .o(n_20703) );
na03f04 TIMEBOOST_cell_8305 ( .a(n_3109), .b(FE_RN_16_0), .c(n_3232), .o(FE_RN_2208_0) );
oa22s02 FE_RC_4367_0 ( .a(n_47019), .b(n_3704), .c(n_3439), .d(FE_OCP_RBN6718_n_3604), .o(n_3824) );
oa22s02 FE_RC_4368_0 ( .a(n_3717), .b(n_3705), .c(n_3715), .d(n_3698), .o(n_3803) );
oa22s02 FE_RC_4369_0 ( .a(n_47341), .b(n_3705), .c(n_3240), .d(n_3604), .o(n_3751) );
in01s03 FE_RC_436_0 ( .a(n_28191), .o(FE_RN_136_0) );
oa22s02 FE_RC_4370_0 ( .a(n_5273), .b(FE_OCP_RBN6201_FE_OFN789_n_46195), .c(n_5196), .d(FE_OFN4789_n_46137), .o(n_46165) );
in01s02 FE_RC_4371_0 ( .a(n_4609), .o(FE_RN_1915_0) );
in01s01 FE_RC_4372_0 ( .a(n_4743), .o(FE_RN_1916_0) );
na02s02 TIMEBOOST_cell_6237 ( .a(n_35539), .b(n_35559), .o(TIMEBOOST_net_1970) );
no02s01 TIMEBOOST_cell_5251 ( .a(TIMEBOOST_net_1573), .b(n_25750), .o(n_25751) );
ao22s02 FE_RC_4375_0 ( .a(n_3217), .b(n_2756), .c(FE_OCP_RBN4147_n_3217), .d(n_2792), .o(n_2899) );
ao22f04 FE_RC_4376_0 ( .a(FE_OCP_RBN3715_n_19241), .b(FE_OCP_RBN2791_FE_RN_368_0), .c(FE_OCPN3570_n_19303), .d(FE_RN_368_0), .o(n_19891) );
oa22f02 FE_RC_4377_0 ( .a(FE_OCPN1394_n_22801), .b(n_22640), .c(n_22617), .d(n_22833), .o(n_22716) );
in01s01 FE_RC_4379_0 ( .a(FE_OCP_RBN1134_n_19077), .o(FE_RN_1918_0) );
na02m08 FE_RC_437_0 ( .a(FE_RN_135_0), .b(FE_RN_136_0), .o(FE_RN_137_0) );
in01s01 FE_RC_4380_0 ( .a(n_20343), .o(FE_RN_1919_0) );
no02s01 FE_RC_4381_0 ( .a(FE_RN_1918_0), .b(FE_RN_1919_0), .o(FE_RN_1920_0) );
no02s06 FE_RC_4382_0 ( .a(FE_RN_1920_0), .b(n_20404), .o(n_20654) );
in01s02 FE_RC_4383_0 ( .a(FE_OCP_RBN1134_n_19077), .o(FE_RN_1921_0) );
in01m01 FE_RC_4384_0 ( .a(n_19325), .o(FE_RN_1922_0) );
no02m02 TIMEBOOST_cell_7741 ( .a(TIMEBOOST_net_2501), .b(n_9390), .o(n_9643) );
na03s06 TIMEBOOST_cell_7742 ( .a(FE_OCP_RBN2851_n_4905), .b(n_3750), .c(FE_OCP_RBN2853_n_4905), .o(TIMEBOOST_net_2502) );
ao22m02 FE_RC_4387_0 ( .a(FE_OCP_RBN2921_n_3878), .b(FE_OCP_RBN3023_n_47011), .c(FE_OCP_RBN6774_n_4046), .d(n_47011), .o(n_4429) );
ao22m02 FE_RC_4388_0 ( .a(FE_OCP_RBN6765_n_3704), .b(n_3971), .c(FE_OCP_RBN6774_n_4046), .d(n_5603), .o(n_4265) );
in01s01 FE_RC_4389_0 ( .a(n_3835), .o(FE_RN_1924_0) );
na02m08 FE_RC_438_0 ( .a(FE_RN_137_0), .b(n_28190), .o(n_28273) );
in01s01 FE_RC_4390_0 ( .a(n_3905), .o(FE_RN_1925_0) );
no02s02 FE_RC_4391_0 ( .a(FE_RN_1924_0), .b(FE_RN_1925_0), .o(FE_RN_1926_0) );
no02m04 TIMEBOOST_cell_8720 ( .a(FE_RN_252_0), .b(FE_RN_253_0), .o(TIMEBOOST_net_2847) );
oa22m02 FE_RC_4393_0 ( .a(FE_OCP_RBN6767_n_3704), .b(n_4376), .c(FE_OCP_RBN2921_n_3878), .d(FE_OCP_RBN5992_n_4376), .o(n_4554) );
oa22s04 FE_RC_4394_0 ( .a(FE_OCP_RBN6774_n_4046), .b(n_4294), .c(FE_OCP_RBN6776_n_4046), .d(FE_OCP_RBN3067_n_4294), .o(n_4552) );
ao22f02 FE_RC_4395_0 ( .a(n_4875), .b(FE_OCP_RBN6842_n_5397), .c(n_4759), .d(n_5397), .o(n_5543) );
in01s02 FE_RC_4396_0 ( .a(n_5310), .o(FE_RN_1927_0) );
in01s01 FE_RC_4397_0 ( .a(n_5426), .o(FE_RN_1928_0) );
no02s04 FE_RC_4398_0 ( .a(FE_RN_1927_0), .b(FE_RN_1928_0), .o(FE_RN_1929_0) );
no02s01 TIMEBOOST_cell_1136 ( .a(TIMEBOOST_net_182), .b(n_41109), .o(n_41178) );
in01s02 FE_RC_43_0 ( .a(n_17742), .o(FE_RN_13_0) );
ao22f02 FE_RC_4400_0 ( .a(FE_OCP_RBN3254_n_5478), .b(n_5503), .c(n_5478), .d(n_5487), .o(n_5656) );
ao22f02 FE_RC_4401_0 ( .a(n_5695), .b(FE_OCP_RBN6124_n_5465), .c(n_5465), .d(n_5696), .o(n_5820) );
oa22m04 FE_RC_4402_0 ( .a(FE_OCP_RBN4360_n_20632), .b(n_20926), .c(n_20632), .d(n_20861), .o(n_20984) );
ao22m08 FE_RC_4403_0 ( .a(n_20658), .b(n_21149), .c(n_20659), .d(n_21150), .o(n_21312) );
in01s02 FE_RC_4404_0 ( .a(n_5677), .o(FE_RN_1930_0) );
in01s02 FE_RC_4405_0 ( .a(n_5911), .o(FE_RN_1931_0) );
no02m04 FE_RC_4406_0 ( .a(FE_RN_1930_0), .b(FE_RN_1931_0), .o(FE_RN_1932_0) );
na02s01 TIMEBOOST_cell_1124 ( .a(TIMEBOOST_net_176), .b(n_33291), .o(n_33351) );
ao22f04 FE_RC_4408_0 ( .a(FE_OCP_RBN6136_n_5816), .b(n_5832), .c(n_5816), .d(n_5833), .o(n_5989) );
in01s03 FE_RC_440_0 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_3_), .o(FE_RN_138_0) );
oa22s02 FE_RC_4410_0 ( .a(n_5066), .b(FE_OCP_RBN6080_n_5346), .c(n_5065), .d(n_5346), .o(n_5490) );
in01s02 FE_RC_4411_0 ( .a(n_4908), .o(FE_RN_1933_0) );
in01m02 FE_RC_4412_0 ( .a(n_5452), .o(FE_RN_1934_0) );
no02s01 TIMEBOOST_cell_1107 ( .a(n_22845), .b(n_22853), .o(TIMEBOOST_net_168) );
no02s01 TIMEBOOST_cell_1108 ( .a(TIMEBOOST_net_168), .b(n_23469), .o(n_23523) );
in01s01 FE_RC_4415_0 ( .a(n_4647), .o(FE_RN_1936_0) );
in01s01 FE_RC_4416_0 ( .a(n_5218), .o(FE_RN_1937_0) );
na02s01 TIMEBOOST_cell_8493 ( .a(TIMEBOOST_net_2733), .b(n_7373), .o(n_7440) );
na02f04 TIMEBOOST_cell_7692 ( .a(n_14786), .b(n_14215), .o(TIMEBOOST_net_2477) );
in01s01 FE_RC_4419_0 ( .a(n_4140), .o(FE_RN_1939_0) );
in01s02 FE_RC_4420_0 ( .a(n_4407), .o(FE_RN_1940_0) );
no02m06 TIMEBOOST_cell_8863 ( .a(TIMEBOOST_net_2918), .b(n_11429), .o(n_11568) );
na02f06 TIMEBOOST_cell_8868 ( .a(n_26084), .b(n_26104), .o(TIMEBOOST_net_2921) );
oa22s04 FE_RC_4423_0 ( .a(n_22167), .b(n_22564), .c(n_22165), .d(FE_OCP_RBN3416_n_22564), .o(n_22718) );
oa22s02 FE_RC_4424_0 ( .a(n_4190), .b(n_4097), .c(n_4096), .d(n_4191), .o(n_4438) );
oa22s03 FE_RC_4425_0 ( .a(n_22385), .b(n_22682), .c(n_22386), .d(n_47207), .o(n_22835) );
oa22f06 FE_RC_4426_0 ( .a(n_22661), .b(n_22490), .c(n_22491), .d(n_22624), .o(n_22818) );
oa22f02 FE_RC_4427_0 ( .a(FE_OCPN1394_n_22801), .b(n_22715), .c(n_22793), .d(n_22670), .o(n_22770) );
oa22s02 FE_RC_4428_0 ( .a(n_22337), .b(n_22685), .c(n_22719), .d(n_22336), .o(n_22874) );
oa22f04 FE_RC_4429_0 ( .a(n_22460), .b(n_22743), .c(FE_RN_1295_0), .d(n_22703), .o(n_22903) );
no02s01 TIMEBOOST_cell_8538 ( .a(FE_RN_889_0), .b(FE_RN_891_0), .o(TIMEBOOST_net_2756) );
in01s01 FE_RC_4430_0 ( .a(n_6215), .o(FE_RN_1942_0) );
in01s02 FE_RC_4431_0 ( .a(n_6332), .o(FE_RN_1943_0) );
na02s04 FE_RC_4432_0 ( .a(FE_RN_1942_0), .b(FE_RN_1943_0), .o(FE_RN_1944_0) );
no02s01 TIMEBOOST_cell_1494 ( .a(TIMEBOOST_net_361), .b(n_8656), .o(n_8707) );
oa22s02 FE_RC_4434_0 ( .a(n_6408), .b(FE_OCP_RBN3445_n_6513), .c(n_6409), .d(n_6513), .o(n_6670) );
no02s02 TIMEBOOST_cell_3861 ( .a(n_37125), .b(n_37272), .o(TIMEBOOST_net_1021) );
oa22s01 FE_RC_4449_0 ( .a(n_1165), .b(n_44652), .c(n_1143), .d(n_44661), .o(n_1295) );
oa22s02 FE_RC_444_0 ( .a(FE_OCP_RBN2631_n_9003), .b(FE_OCPN849_n_7712), .c(FE_OCP_RBN6601_n_7708), .d(n_9003), .o(n_8077) );
oa22s01 FE_RC_4450_0 ( .a(n_1065), .b(n_44652), .c(n_1049), .d(n_44623), .o(n_1304) );
oa22s01 FE_RC_4451_0 ( .a(n_1102), .b(FE_OCPN838_n_44672), .c(n_1064), .d(n_44637), .o(n_1343) );
no02s02 TIMEBOOST_cell_1567 ( .a(n_8342), .b(FE_OCP_RBN6601_n_7708), .o(TIMEBOOST_net_398) );
na02s02 TIMEBOOST_cell_4285 ( .a(FE_OFN738_n_17093), .b(n_18032), .o(TIMEBOOST_net_1233) );
oa22m04 FE_RC_4456_0 ( .a(n_22039), .b(n_21985), .c(n_22038), .d(n_44296), .o(n_22066) );
oa22m04 FE_RC_4457_0 ( .a(n_30147), .b(n_30424), .c(n_30425), .d(n_30148), .o(n_30492) );
ao22f02 FE_RC_4459_0 ( .a(n_30466), .b(n_44439), .c(n_27014), .d(n_30451), .o(n_30542) );
no02s02 TIMEBOOST_cell_1903 ( .a(n_27117), .b(n_27086), .o(TIMEBOOST_net_566) );
ao22m04 FE_RC_4461_0 ( .a(n_45065), .b(n_20325), .c(n_45066), .d(FE_OCP_RBN2095_n_20325), .o(n_20435) );
oa22m08 FE_RC_4462_0 ( .a(n_11763), .b(FE_OCP_RBN2427_n_11907), .c(n_11907), .d(n_11764), .o(n_12062) );
oa22m08 FE_RC_4464_0 ( .a(FE_OCP_RBN3989_n_32772), .b(n_32678), .c(n_32679), .d(n_32772), .o(n_32827) );
in01s06 FE_RC_4466_0 ( .a(n_32634), .o(FE_RN_1954_0) );
in01m06 FE_RC_4467_0 ( .a(n_32818), .o(FE_RN_1955_0) );
na02s20 FE_RC_4468_0 ( .a(FE_RN_1955_0), .b(FE_RN_1954_0), .o(FE_RN_1956_0) );
oa22s04 FE_RC_4471_0 ( .a(n_36236), .b(n_36517), .c(n_36237), .d(n_36516), .o(n_36615) );
oa22s02 FE_RC_4472_0 ( .a(n_36832), .b(n_36770), .c(n_36769), .d(n_36833), .o(n_36874) );
oa22s02 FE_RC_4476_0 ( .a(n_6960), .b(n_6690), .c(n_6689), .d(n_6961), .o(n_7050) );
ao22m04 FE_RC_4477_0 ( .a(n_33287), .b(n_33730), .c(n_33729), .d(n_33288), .o(n_33825) );
in01m02 FE_RC_4478_0 ( .a(n_28332), .o(FE_RN_1957_0) );
in01s02 FE_RC_4479_0 ( .a(n_28334), .o(FE_RN_1958_0) );
oa22m02 FE_RC_447_0 ( .a(FE_OCP_RBN6601_n_7708), .b(FE_OCP_RBN6628_n_8269), .c(FE_OCPN849_n_7712), .d(n_8269), .o(n_8107) );
na02m04 FE_RC_4480_0 ( .a(FE_RN_1957_0), .b(FE_RN_1958_0), .o(FE_RN_1959_0) );
na02m06 FE_RC_4481_0 ( .a(FE_RN_1959_0), .b(n_28333), .o(n_28405) );
in01f06 FE_RC_4484_0 ( .a(n_28308), .o(FE_RN_1960_0) );
in01s02 FE_RC_4485_0 ( .a(n_28309), .o(FE_RN_1961_0) );
no02m10 TIMEBOOST_cell_8470 ( .a(FE_RN_1259_0), .b(FE_RN_1258_0), .o(TIMEBOOST_net_2722) );
no03m08 TIMEBOOST_cell_8458 ( .a(TIMEBOOST_net_1320), .b(n_21351), .c(n_21574), .o(n_21764) );
oa22m04 FE_RC_4489_0 ( .a(n_7486), .b(FE_OCP_RBN6631_n_8111), .c(n_8111), .d(n_7487), .o(n_8221) );
oa22f04 FE_RC_4490_0 ( .a(FE_OCP_RBN2608_FE_OCPN855_n_7721), .b(FE_OCP_RBN4185_n_8288), .c(FE_OCP_RBN2616_FE_OCPN857_n_7802), .d(n_8288), .o(n_8410) );
ao22f04 FE_RC_4493_0 ( .a(n_7661), .b(n_8704), .c(n_7660), .d(n_8703), .o(n_8842) );
oa22f04 FE_RC_4494_0 ( .a(n_28602), .b(n_28948), .c(n_28601), .d(n_28949), .o(n_29030) );
ao22m04 FE_RC_4495_0 ( .a(n_13045), .b(n_13956), .c(n_13046), .d(n_13955), .o(n_14099) );
ao22m04 FE_RC_4496_0 ( .a(n_44352), .b(n_7520), .c(n_7519), .d(FE_OCP_RBN6658_n_44352), .o(n_8380) );
oa22f04 FE_RC_4498_0 ( .a(FE_OFN4796_n_13195), .b(FE_OCP_RBN2076_n_14149), .c(n_14149), .d(n_13418), .o(n_14321) );
oa22m02 FE_RC_4499_0 ( .a(n_8681), .b(n_8554), .c(n_8499), .d(n_8680), .o(n_8838) );
in01s06 FE_RC_449_0 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_3_), .o(FE_RN_141_0) );
na02s04 FE_RC_44_0 ( .a(FE_RN_12_0), .b(FE_RN_13_0), .o(FE_RN_14_0) );
ao22f04 FE_RC_4500_0 ( .a(n_13515), .b(n_14328), .c(FE_OFN4795_n_13195), .d(n_14327), .o(n_14462) );
oa22f02 FE_RC_4501_0 ( .a(n_9173), .b(n_9754), .c(n_9111), .d(n_9855), .o(n_9941) );
ao22m06 FE_RC_4502_0 ( .a(FE_OCP_RBN2535_n_33568), .b(n_33183), .c(n_33568), .d(n_33182), .o(n_33697) );
oa22f04 FE_RC_4503_0 ( .a(n_34558), .b(n_34876), .c(n_34559), .d(n_34877), .o(n_34980) );
oa22f04 FE_RC_4505_0 ( .a(FE_OCPN1083_n_8388), .b(n_8667), .c(n_8750), .d(n_8666), .o(n_8782) );
oa22f02 FE_RC_4507_0 ( .a(FE_OCP_RBN4186_n_8288), .b(n_8602), .c(FE_OCP_RBN6675_n_8288), .d(n_8601), .o(n_8753) );
oa22m02 FE_RC_4508_0 ( .a(n_45091), .b(n_20941), .c(n_45013), .d(FE_OCP_RBN7047_n_20941), .o(n_21072) );
oa22f04 FE_RC_4509_0 ( .a(n_45066), .b(n_20462), .c(n_20461), .d(n_45012), .o(n_20636) );
oa22f04 FE_RC_4512_0 ( .a(n_10366), .b(FE_OCP_RBN6027_n_10445), .c(n_10445), .d(n_10365), .o(n_10568) );
oa22f04 FE_RC_4515_0 ( .a(n_29501), .b(n_29730), .c(n_29530), .d(n_29749), .o(n_29773) );
na02f04 TIMEBOOST_cell_5159 ( .a(TIMEBOOST_net_1527), .b(n_14557), .o(n_14638) );
in01s01 FE_RC_4518_0 ( .a(FE_OCPN1402_FE_OFN1196_n_27014), .o(FE_RN_1963_0) );
in01f02 FE_RC_4519_0 ( .a(n_30619), .o(FE_RN_1964_0) );
no02f04 TIMEBOOST_cell_3862 ( .a(TIMEBOOST_net_1021), .b(n_37447), .o(n_37512) );
no02f08 TIMEBOOST_cell_7010 ( .a(TIMEBOOST_net_2263), .b(n_34827), .o(n_34955) );
na02f08 TIMEBOOST_cell_5438 ( .a(FE_OCP_RBN2108_n_15911), .b(n_14452), .o(TIMEBOOST_net_1667) );
oa22f04 FE_RC_4522_0 ( .a(n_34394), .b(n_34880), .c(n_34395), .d(n_34881), .o(n_34982) );
oa22s04 FE_RC_4524_0 ( .a(n_11745), .b(n_11964), .c(n_11746), .d(n_11987), .o(n_12197) );
oa22m04 FE_RC_4525_0 ( .a(n_11742), .b(n_12022), .c(n_11741), .d(n_11986), .o(n_12217) );
ao22f04 FE_RC_4526_0 ( .a(n_35139), .b(n_35332), .c(n_35140), .d(FE_RN_1493_0), .o(n_35416) );
ao22m04 FE_RC_4527_0 ( .a(n_27062), .b(n_30534), .c(FE_OFN1198_n_27014), .d(FE_OCP_RBN6000_n_30534), .o(n_30625) );
oa22m02 FE_RC_4528_0 ( .a(FE_OCPN1681_n_30614), .b(FE_OCP_RBN5943_n_35207), .c(n_30633), .d(n_35207), .o(n_35231) );
no02m08 TIMEBOOST_cell_5093 ( .a(TIMEBOOST_net_1494), .b(n_19331), .o(n_19467) );
in01s01 FE_RC_4530_0 ( .a(n_30403), .o(FE_RN_1966_0) );
in01s02 FE_RC_4531_0 ( .a(n_30678), .o(FE_RN_1967_0) );
no02s02 FE_RC_4532_0 ( .a(FE_RN_1966_0), .b(FE_RN_1967_0), .o(FE_RN_1968_0) );
na02m04 TIMEBOOST_cell_1096 ( .a(n_23438), .b(TIMEBOOST_net_162), .o(n_23494) );
in01s01 FE_RC_4534_0 ( .a(FE_RN_1132_0), .o(FE_RN_1969_0) );
in01s02 FE_RC_4535_0 ( .a(n_30885), .o(FE_RN_1970_0) );
na02m04 FE_RC_4536_0 ( .a(FE_RN_1969_0), .b(FE_RN_1970_0), .o(FE_RN_1971_0) );
na02m06 FE_RC_4537_0 ( .a(FE_RN_1133_0), .b(FE_RN_1971_0), .o(n_31010) );
oa22f04 FE_RC_4538_0 ( .a(FE_RN_1780_0), .b(n_35078), .c(n_35012), .d(FE_RN_1781_0), .o(n_35198) );
ao22m02 FE_RC_4539_0 ( .a(n_30545), .b(n_34983), .c(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q), .d(n_34960), .o(n_35107) );
no03s03 FE_RC_4540_0 ( .a(n_31947), .b(n_31993), .c(n_31992), .o(n_32021) );
oa22m02 FE_RC_4541_0 ( .a(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n_36709), .c(TIMEBOOST_net_2317), .d(n_36654), .o(n_36722) );
oa22f04 FE_RC_4543_0 ( .a(n_35971), .b(n_36447), .c(n_35972), .d(n_45617), .o(n_36520) );
oa22s02 FE_RC_4551_0 ( .a(n_17136), .b(n_17626), .c(n_17191), .d(n_17600), .o(n_17782) );
ao22f02 FE_RC_4552_0 ( .a(FE_OCP_RBN6035_n_30769), .b(FE_OCP_RBN3722_n_30776), .c(n_30776), .d(n_30769), .o(n_30918) );
oa22f06 FE_RC_4553_0 ( .a(n_31831), .b(n_32196), .c(n_31832), .d(n_32218), .o(n_32311) );
oa22f04 FE_RC_4554_0 ( .a(n_32143), .b(n_31834), .c(n_31833), .d(FE_OCP_RBN3406_n_32143), .o(n_32255) );
na02s02 TIMEBOOST_cell_1687 ( .a(FE_RN_530_0), .b(FE_RN_529_0), .o(TIMEBOOST_net_458) );
no02s02 TIMEBOOST_cell_1795 ( .a(FE_OFN4800_n_44498), .b(n_10883), .o(TIMEBOOST_net_512) );
ao22f04 FE_RC_4561_0 ( .a(n_7495), .b(n_8207), .c(n_7494), .d(n_8206), .o(n_8288) );
in01s01 FE_RC_4563_0 ( .a(n_32704), .o(FE_RN_1975_0) );
in01m04 FE_RC_4564_0 ( .a(FE_RN_257_0), .o(FE_RN_1976_0) );
na02m08 FE_RC_4565_0 ( .a(FE_RN_1975_0), .b(FE_RN_1976_0), .o(FE_RN_1977_0) );
no02s01 TIMEBOOST_cell_8479 ( .a(TIMEBOOST_net_2726), .b(n_37166), .o(n_37201) );
oa22m04 FE_RC_4568_0 ( .a(n_11296), .b(FE_OCP_RBN3359_n_11275), .c(n_11275), .d(n_11274), .o(n_11377) );
ao22f10 FE_RC_4570_0 ( .a(FE_OCP_RBN2028_n_44722), .b(n_44422), .c(FE_OCP_RBN7128_n_44722), .d(n_44420), .o(n_27859) );
oa22s03 FE_RC_4571_0 ( .a(n_22498), .b(FE_OCP_RBN5348_FE_RN_627_0), .c(n_22499), .d(FE_RN_627_0), .o(n_22897) );
in01f20 FE_RC_4572_0 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_3_), .o(FE_RN_1978_0) );
in01s06 FE_RC_4573_0 ( .a(n_44723), .o(FE_RN_1979_0) );
no02s02 TIMEBOOST_cell_4112 ( .a(TIMEBOOST_net_1146), .b(n_36098), .o(n_36268) );
no02s06 TIMEBOOST_cell_8675 ( .a(TIMEBOOST_net_2824), .b(TIMEBOOST_net_2678), .o(n_36612) );
no02s02 TIMEBOOST_cell_6997 ( .a(n_15441), .b(n_15482), .o(TIMEBOOST_net_2257) );
na03f06 FE_RC_4580_0 ( .a(n_16172), .b(n_16205), .c(n_16170), .o(n_16290) );
oa22f04 FE_RC_4581_0 ( .a(n_12961), .b(n_13816), .c(n_12962), .d(n_13815), .o(n_13927) );
ao22m04 FE_RC_4582_0 ( .a(FE_OCP_RBN4106_n_12880), .b(n_14069), .c(n_13195), .d(FE_OCP_RBN2066_n_14069), .o(n_14249) );
ao22f08 FE_RC_4584_0 ( .a(FE_OCP_RBN2068_n_14069), .b(FE_OCP_RBN6378_n_14380), .c(FE_OCP_RBN2070_n_14069), .d(FE_OCP_RBN6379_n_14380), .o(n_14585) );
no02m04 TIMEBOOST_cell_8793 ( .a(TIMEBOOST_net_2883), .b(n_24650), .o(n_24750) );
na02s01 TIMEBOOST_cell_3358 ( .a(n_26865), .b(n_26864), .o(TIMEBOOST_net_970) );
no03s08 TIMEBOOST_cell_8331 ( .a(n_10485), .b(n_10276), .c(n_10484), .o(TIMEBOOST_net_1942) );
oa22f04 FE_RC_4595_0 ( .a(n_23718), .b(n_24018), .c(n_23685), .d(n_24019), .o(n_24079) );
oa22f04 FE_RC_4597_0 ( .a(n_25824), .b(n_25729), .c(FE_OFN747_n_22641), .d(FE_OCP_RBN5200_n_25729), .o(n_25847) );
oa22f02 FE_RC_4598_0 ( .a(n_45091), .b(n_20847), .c(n_45013), .d(n_20848), .o(n_21006) );
oa22f02 FE_RC_4599_0 ( .a(n_26331), .b(n_26400), .c(n_26399), .d(n_26364), .o(n_26522) );
na02m06 FE_RC_45_0 ( .a(FE_RN_14_0), .b(n_17743), .o(n_17841) );
ao22m04 FE_RC_4602_0 ( .a(FE_OCPN1693_n_33140), .b(n_33596), .c(n_33141), .d(n_33595), .o(n_33675) );
ao22s04 FE_RC_4604_0 ( .a(n_45024), .b(FE_OCP_RBN2112_n_20935), .c(n_45010), .d(n_20935), .o(n_21064) );
ao22f02 FE_RC_4607_0 ( .a(FE_OCP_RBN5911_n_44563), .b(n_10225), .c(FE_OFN4775_n_44463), .d(FE_OCP_RBN6015_n_10225), .o(n_10401) );
oa22m04 FE_RC_4609_0 ( .a(n_22419), .b(n_22625), .c(n_22416), .d(FE_OCP_RBN4648_n_22625), .o(n_22819) );
ao22f20 FE_RC_460_0 ( .a(n_27776), .b(FE_OCP_RBN7127_n_44722), .c(n_44759), .d(delay_xor_ln22_unr18_stage7_stallmux_q_2_), .o(n_27827) );
oa22f02 FE_RC_4610_0 ( .a(n_22801), .b(n_22819), .c(n_22793), .d(n_22792), .o(n_22893) );
ao22s02 FE_RC_4611_0 ( .a(n_27246), .b(FE_OCP_RBN6064_n_30908), .c(n_27366), .d(n_30908), .o(n_31023) );
ao22m04 FE_RC_4612_0 ( .a(FE_OFN1196_n_27014), .b(FE_OCP_RBN1846_n_30492), .c(n_30466), .d(n_30492), .o(n_30575) );
in01s01 FE_RC_4613_0 ( .a(FE_RN_1982_0), .o(FE_RN_1981_0) );
no02s01 FE_RC_4614_0 ( .a(n_32800), .b(FE_RN_1981_0), .o(n_33113) );
na02f08 FE_RC_4616_0 ( .a(n_33039), .b(n_32833), .o(FE_RN_1982_0) );
oa22m04 FE_RC_461_0 ( .a(n_12997), .b(n_13533), .c(n_12998), .d(n_13532), .o(n_13616) );
na02s02 TIMEBOOST_cell_1587 ( .a(n_3184), .b(n_3216), .o(TIMEBOOST_net_408) );
na02m04 TIMEBOOST_cell_6822 ( .a(TIMEBOOST_net_2168), .b(n_16472), .o(n_16569) );
no02s02 TIMEBOOST_cell_8837 ( .a(TIMEBOOST_net_2905), .b(n_4681), .o(TIMEBOOST_net_2157) );
na03m08 TIMEBOOST_cell_6517 ( .a(n_24345), .b(FE_OFN743_delay_sub_ln23_0_unr15_stage6_stallmux_q), .c(n_24369), .o(TIMEBOOST_net_1953) );
no02s02 TIMEBOOST_cell_8558 ( .a(n_2913), .b(n_3259), .o(TIMEBOOST_net_2766) );
no02s02 TIMEBOOST_cell_1751 ( .a(FE_OCPN4539_n_20332), .b(FE_OCP_RBN4325_n_20333), .o(TIMEBOOST_net_490) );
na02s02 FE_RC_4635_0 ( .a(n_35780), .b(n_35732), .o(FE_RN_1995_0) );
no02f08 FE_RC_4636_0 ( .a(n_36352), .b(FE_RN_1995_0), .o(n_36381) );
no02m20 FE_RC_4639_0 ( .a(FE_OCP_RBN6320_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_0_), .o(FE_RN_1997_0) );
na02s06 FE_RC_4643_0 ( .a(FE_OCPN1902_n_32712), .b(n_32709), .o(FE_RN_2000_0) );
na02s06 FE_RC_4644_0 ( .a(n_46413), .b(n_32711), .o(FE_RN_2001_0) );
na02s02 TIMEBOOST_cell_1605 ( .a(n_30255), .b(n_30267), .o(TIMEBOOST_net_417) );
in01m01 FE_RC_4647_0 ( .a(n_36011), .o(FE_RN_2003_0) );
na02m04 FE_RC_4648_0 ( .a(n_36416), .b(FE_RN_2003_0), .o(n_36445) );
in01s01 FE_RC_4649_0 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_5_), .o(FE_RN_2004_0) );
ao22m02 FE_RC_464_0 ( .a(n_12600), .b(n_13175), .c(n_12599), .d(n_13176), .o(n_13335) );
na02s01 FE_RC_4650_0 ( .a(FE_RN_2004_0), .b(n_6874), .o(n_6992) );
na02s01 FE_RC_4652_0 ( .a(n_34328), .b(n_34570), .o(n_34415) );
in01s01 FE_RC_4660_0 ( .a(n_19533), .o(FE_RN_2009_0) );
in01s02 FE_RC_4661_0 ( .a(FE_RN_2010_0), .o(n_19617) );
na02s02 FE_RC_4662_0 ( .a(n_19528), .b(FE_RN_2009_0), .o(FE_RN_2010_0) );
in01s02 FE_RC_4665_0 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_13_), .o(FE_RN_2012_0) );
na02s10 FE_RC_4666_0 ( .a(FE_OCP_RBN2414_n_44722), .b(n_28044), .o(FE_RN_2013_0) );
in01s01 FE_RC_4667_0 ( .a(FE_OCP_RBN2039_n_44722), .o(FE_RN_2014_0) );
na02f02 TIMEBOOST_cell_7845 ( .a(TIMEBOOST_net_2553), .b(n_35444), .o(n_35472) );
na02f04 FE_RC_4669_0 ( .a(FE_RN_2015_0), .b(n_27972), .o(FE_RN_2016_0) );
ao22f08 FE_RC_4670_0 ( .a(FE_RN_2012_0), .b(FE_RN_2013_0), .c(FE_RN_2014_0), .d(FE_RN_2016_0), .o(FE_RN_2017_0) );
na02f10 FE_RC_4671_0 ( .a(FE_RN_2017_0), .b(n_28359), .o(n_28383) );
no02s01 FE_RC_4672_0 ( .a(n_27710), .b(n_27712), .o(FE_RN_2018_0) );
no02s06 FE_RC_4673_0 ( .a(FE_RN_2018_0), .b(n_28467), .o(n_28510) );
in01s01 TIMEBOOST_cell_8899 ( .a(TIMEBOOST_net_2942), .o(TIMEBOOST_net_2943) );
na03s02 TIMEBOOST_cell_7560 ( .a(FE_RN_697_0), .b(n_25135), .c(FE_RN_699_0), .o(TIMEBOOST_net_2411) );
in01s01 FE_RC_4677_0 ( .a(FE_OCP_RBN2599_n_7743), .o(FE_RN_2021_0) );
no02m04 TIMEBOOST_cell_4148 ( .a(TIMEBOOST_net_1164), .b(n_36669), .o(TIMEBOOST_net_974) );
no02s02 TIMEBOOST_cell_4149 ( .a(n_16118), .b(n_16843), .o(TIMEBOOST_net_1165) );
ao22m04 FE_RC_467_0 ( .a(n_12794), .b(n_13575), .c(n_12793), .d(n_13576), .o(n_13661) );
na02s02 TIMEBOOST_cell_4181 ( .a(n_22230), .b(n_22474), .o(TIMEBOOST_net_1181) );
na02f06 TIMEBOOST_cell_8568 ( .a(FE_OCP_RBN2085_n_14911), .b(FE_OCP_RBN2834_n_13962), .o(TIMEBOOST_net_2771) );
no02f06 FE_RC_4682_0 ( .a(FE_RN_2023_0), .b(FE_RN_2025_0), .o(n_9113) );
in01m06 FE_RC_4685_0 ( .a(FE_RN_2027_0), .o(n_32845) );
no02m08 FE_RC_4686_0 ( .a(n_32784), .b(delay_add_ln22_unr20_stage8_stallmux_q_3_), .o(FE_RN_2027_0) );
ao22m04 FE_RC_468_0 ( .a(n_12647), .b(n_13299), .c(n_12648), .d(n_13298), .o(n_13388) );
na02s06 FE_RC_4692_0 ( .a(FE_OCP_RBN6556_n_28458), .b(n_28606), .o(FE_RN_2031_0) );
na02m08 FE_RC_4693_0 ( .a(FE_RN_2031_0), .b(n_28979), .o(n_29039) );
in01s01 FE_RC_4694_0 ( .a(FE_OCP_RBN6685_FE_OCPN4529_FE_OCP_RBN2748_n_8474), .o(FE_RN_2032_0) );
na02m02 FE_RC_4696_0 ( .a(FE_RN_2032_0), .b(n_9809), .o(FE_RN_2033_0) );
na02s10 FE_RC_4698_0 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_1_), .b(FE_OCP_RBN7129_n_44722), .o(n_27738) );
oa22m02 FE_RC_469_0 ( .a(n_28732), .b(n_29117), .c(n_28733), .d(n_29116), .o(n_29217) );
na02f02 FE_RC_4700_0 ( .a(n_19915), .b(FE_OCP_DRV_N1898_n_18287), .o(FE_RN_2034_0) );
na02s20 FE_RC_4703_0 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_1_), .b(FE_OCP_RBN7015_n_44962), .o(FE_RN_2036_0) );
na02f20 FE_RC_4704_0 ( .a(n_32578), .b(FE_RN_2036_0), .o(n_32520) );
in01s01 FE_RC_4705_0 ( .a(n_12956), .o(FE_RN_2037_0) );
in01s01 FE_RC_4706_0 ( .a(n_46415), .o(FE_RN_2038_0) );
no02s01 FE_RC_4707_0 ( .a(FE_RN_2037_0), .b(FE_RN_2038_0), .o(FE_RN_2039_0) );
in01m06 FE_RC_4708_0 ( .a(FE_RN_2040_0), .o(n_13957) );
na02m08 FE_RC_4709_0 ( .a(n_13866), .b(FE_RN_2039_0), .o(FE_RN_2040_0) );
ao22f04 FE_RC_470_0 ( .a(n_28997), .b(n_28625), .c(n_28998), .d(n_28624), .o(n_29091) );
in01m02 FE_RC_4710_0 ( .a(n_14321), .o(FE_RN_2041_0) );
na02m02 TIMEBOOST_cell_1988 ( .a(TIMEBOOST_net_608), .b(n_29039), .o(n_29065) );
na02s06 TIMEBOOST_cell_4922 ( .a(n_7063), .b(n_7062), .o(TIMEBOOST_net_1409) );
in01s01 FE_RC_4713_0 ( .a(n_33017), .o(FE_RN_2043_0) );
in01m01 FE_RC_4714_0 ( .a(n_33386), .o(FE_RN_2044_0) );
no02m02 FE_RC_4715_0 ( .a(FE_RN_2043_0), .b(FE_RN_2044_0), .o(FE_RN_2045_0) );
na02m02 FE_RC_4716_0 ( .a(n_33388), .b(FE_RN_2045_0), .o(n_33412) );
in01s01 FE_RC_4722_0 ( .a(FE_OCPN1291_n_29439), .o(FE_RN_2049_0) );
no02f06 FE_RC_4723_0 ( .a(n_29440), .b(FE_RN_2049_0), .o(n_29466) );
in01m03 FE_RC_4725_0 ( .a(n_29258), .o(FE_RN_2051_0) );
in01s01 FE_RC_4733_0 ( .a(FE_OCP_DRV_N4503_n_28888), .o(FE_RN_2056_0) );
no02s04 FE_RC_4734_0 ( .a(FE_RN_2056_0), .b(n_29841), .o(n_29893) );
no02s10 FE_RC_4739_0 ( .a(n_31605), .b(n_31664), .o(FE_RN_2059_0) );
na02f20 FE_RC_4740_0 ( .a(n_31959), .b(FE_RN_2059_0), .o(n_32000) );
in01s01 FE_RC_4741_0 ( .a(n_27062), .o(FE_RN_2060_0) );
no02m04 FE_RC_4742_0 ( .a(FE_RN_2060_0), .b(n_30818), .o(FE_RN_1144_0) );
in01s01 FE_RC_4746_0 ( .a(n_45024), .o(FE_RN_2063_0) );
no02m02 FE_RC_4748_0 ( .a(FE_RN_2063_0), .b(n_21072), .o(FE_RN_2064_0) );
in01s02 FE_RC_474_0 ( .a(n_13829), .o(FE_RN_145_0) );
no02f06 FE_RC_4750_0 ( .a(n_33715), .b(FE_RN_2288_0), .o(n_33731) );
na02f06 FE_RC_4753_0 ( .a(n_20903), .b(n_20930), .o(FE_RN_2067_0) );
na02f08 FE_RC_4754_0 ( .a(FE_RN_2067_0), .b(n_20957), .o(n_21054) );
ao22m04 FE_RC_4755_0 ( .a(FE_OCPN1679_n_27315), .b(FE_OCP_RBN6085_n_31010), .c(n_27366), .d(n_31010), .o(n_31111) );
in01s01 FE_RC_4756_0 ( .a(n_31740), .o(FE_RN_2068_0) );
na02s04 FE_RC_4757_0 ( .a(FE_RN_2068_0), .b(n_31765), .o(n_31805) );
in01s02 FE_RC_4758_0 ( .a(n_31048), .o(FE_RN_2069_0) );
in01m02 FE_RC_4759_0 ( .a(n_30930), .o(FE_RN_2070_0) );
na02m01 TIMEBOOST_cell_5287 ( .a(TIMEBOOST_net_1591), .b(n_3547), .o(n_3758) );
in01s01 FE_RC_4766_0 ( .a(FE_OCPUNCON3491_n_30322), .o(FE_RN_2074_0) );
na02f06 FE_RC_4767_0 ( .a(n_31449), .b(FE_RN_2074_0), .o(n_31477) );
in01m02 FE_RC_4768_0 ( .a(FE_RN_2075_0), .o(n_45523) );
na02s02 FE_RC_4769_0 ( .a(n_15001), .b(n_13476), .o(FE_RN_2075_0) );
no02f02 TIMEBOOST_cell_5288 ( .a(FE_OCP_RBN5331_n_20843), .b(n_20790), .o(TIMEBOOST_net_1592) );
in01s01 FE_RC_4770_0 ( .a(n_1669), .o(FE_RN_2076_0) );
in01s01 FE_RC_4771_0 ( .a(n_1645), .o(FE_RN_2077_0) );
in01s01 TIMEBOOST_cell_8901 ( .a(TIMEBOOST_net_2944), .o(TIMEBOOST_net_2945) );
na02s01 FE_RC_4773_0 ( .a(n_1682), .b(n_1681), .o(FE_RN_2079_0) );
na02s01 FE_RC_4774_0 ( .a(n_1646), .b(n_1645), .o(FE_RN_2080_0) );
na03m02 TIMEBOOST_cell_3525 ( .a(FE_OCP_RBN4032_n_37690), .b(n_37755), .c(TIMEBOOST_net_729), .o(n_37772) );
no02s02 TIMEBOOST_cell_1832 ( .a(TIMEBOOST_net_530), .b(n_31765), .o(n_31850) );
na02m04 TIMEBOOST_cell_5617 ( .a(TIMEBOOST_net_1756), .b(n_11363), .o(n_11494) );
no02s02 TIMEBOOST_cell_1921 ( .a(n_22554), .b(n_22411), .o(TIMEBOOST_net_575) );
in01s02 FE_RC_4779_0 ( .a(n_1748), .o(FE_RN_2084_0) );
na02s01 FE_RC_4780_0 ( .a(n_1741), .b(FE_RN_2084_0), .o(FE_RN_2085_0) );
no02s01 FE_RC_4781_0 ( .a(n_1749), .b(FE_RN_2085_0), .o(FE_RN_2086_0) );
oa22s04 FE_RC_4782_0 ( .a(n_1742), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_22_), .c(n_1686), .d(n_1787), .o(FE_RN_2087_0) );
na02s01 FE_RC_4783_0 ( .a(n_1596), .b(n_1597), .o(FE_RN_2088_0) );
oa12f06 FE_RC_4784_0 ( .a(FE_RN_2087_0), .b(FE_RN_2088_0), .c(n_45718), .o(FE_RN_2089_0) );
na02f08 FE_RC_4785_0 ( .a(FE_RN_2089_0), .b(FE_RN_2086_0), .o(n_2148) );
no02s02 FE_RC_4786_0 ( .a(n_37017), .b(n_37004), .o(FE_RN_2090_0) );
na02m06 FE_RC_4787_0 ( .a(FE_RN_2090_0), .b(n_37133), .o(FE_RN_2091_0) );
no02f08 FE_RC_4788_0 ( .a(FE_RN_2091_0), .b(n_37299), .o(n_37380) );
ao22m04 FE_RC_478_0 ( .a(n_13022), .b(n_13929), .c(n_13023), .d(n_13928), .o(n_14069) );
na03s08 FE_RC_4791_0 ( .a(n_39061), .b(n_39060), .c(n_38951), .o(n_39062) );
ao22f08 FE_RC_4792_0 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_4_), .b(n_6957), .c(n_6763), .d(n_6585), .o(n_6900) );
na02s01 TIMEBOOST_cell_5249 ( .a(TIMEBOOST_net_1572), .b(n_26606), .o(n_26687) );
na02s01 FE_RC_4794_0 ( .a(n_34440), .b(n_34186), .o(n_34493) );
na02s01 FE_RC_4795_0 ( .a(n_34186), .b(n_34440), .o(FE_RN_2092_0) );
no02s01 FE_RC_4796_0 ( .a(n_34204), .b(FE_RN_2092_0), .o(n_34574) );
in01m06 FE_RC_4797_0 ( .a(n_34192), .o(FE_RN_2093_0) );
no02f08 FE_RC_4798_0 ( .a(n_34204), .b(FE_RN_2093_0), .o(FE_RN_2094_0) );
ao22s06 FE_RC_47_0 ( .a(n_17394), .b(FE_OCP_RBN7103_n_44365), .c(delay_xor_ln22_unr12_stage5_stallmux_q_6_), .d(FE_OCP_RBN5511_n_44365), .o(n_17581) );
in01s01 FE_RC_4800_0 ( .a(FE_OCP_RBN4096_n_12880), .o(FE_RN_2095_0) );
no02f04 FE_RC_4802_0 ( .a(FE_RN_2095_0), .b(FE_RN_2154_0), .o(FE_RN_2097_0) );
no02f08 FE_RC_4803_0 ( .a(n_13788), .b(FE_RN_2097_0), .o(n_13886) );
in01s02 FE_RC_4804_0 ( .a(FE_OCP_DRV_N1407_n_28550), .o(FE_RN_2098_0) );
no02f08 FE_RC_4805_0 ( .a(n_28935), .b(FE_RN_2098_0), .o(n_28976) );
in01s01 FE_RC_4808_0 ( .a(n_11769), .o(FE_RN_2100_0) );
no02s06 FE_RC_4809_0 ( .a(n_11694), .b(FE_RN_2100_0), .o(FE_RN_2101_0) );
in01m20 FE_RC_4813_0 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_2_), .o(FE_RN_2103_0) );
na03s02 TIMEBOOST_cell_2251 ( .a(n_1911), .b(n_1758), .c(n_1933), .o(TIMEBOOST_net_343) );
no02f08 TIMEBOOST_cell_1558 ( .a(TIMEBOOST_net_393), .b(n_30518), .o(n_30663) );
oa22f06 FE_RC_4816_0 ( .a(n_36268), .b(FE_OCP_RBN3381_n_36547), .c(n_36269), .d(n_36547), .o(n_36651) );
na02s02 FE_RC_4817_0 ( .a(n_12106), .b(n_12105), .o(FE_RN_2105_0) );
oa12s02 FE_RC_4818_0 ( .a(FE_RN_2105_0), .b(n_12106), .c(n_12105), .o(n_12230) );
in01s01 FE_RC_481_0 ( .a(n_28701), .o(FE_RN_147_0) );
na02s01 FE_RC_4821_0 ( .a(n_7891), .b(n_7857), .o(FE_RN_2107_0) );
no02f08 FE_RC_4822_0 ( .a(n_8337), .b(FE_RN_2107_0), .o(n_8369) );
in01s01 FE_RC_4823_0 ( .a(n_7963), .o(FE_RN_2108_0) );
in01s01 FE_RC_4824_0 ( .a(n_7999), .o(FE_RN_2109_0) );
no02s02 FE_RC_4825_0 ( .a(n_8058), .b(FE_RN_2109_0), .o(FE_RN_2110_0) );
no02s01 FE_RC_4826_0 ( .a(n_8012), .b(n_7980), .o(FE_RN_2111_0) );
na02s01 FE_RC_4827_0 ( .a(FE_RN_2111_0), .b(n_8014), .o(FE_RN_2112_0) );
oa22f06 FE_RC_4828_0 ( .a(FE_RN_2110_0), .b(FE_RN_2108_0), .c(FE_RN_2112_0), .d(n_8613), .o(n_8684) );
na03m08 FE_RC_4829_0 ( .a(n_9465), .b(FE_OCP_RBN5881_FE_RN_314_0), .c(n_9504), .o(n_9627) );
in01f02 FE_RC_482_0 ( .a(n_29092), .o(FE_RN_148_0) );
no03m04 TIMEBOOST_cell_8250 ( .a(n_7724), .b(n_7458), .c(n_7753), .o(n_7884) );
no02f06 TIMEBOOST_cell_8756 ( .a(n_13858), .b(n_14001), .o(TIMEBOOST_net_2865) );
no02s06 TIMEBOOST_cell_5137 ( .a(TIMEBOOST_net_1516), .b(n_8973), .o(n_9190) );
in01s40 FE_RC_4833_0 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_0_), .o(FE_RN_2115_0) );
na02s40 FE_RC_4834_0 ( .a(FE_RN_2115_0), .b(n_44061), .o(n_22769) );
in01s06 FE_RC_4835_0 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_1_), .o(FE_RN_2116_0) );
na02s08 FE_RC_4836_0 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(FE_RN_2116_0), .o(n_6607) );
in01m40 FE_RC_4837_0 ( .a(n_45204), .o(FE_RN_2117_0) );
na02m20 FE_RC_4838_0 ( .a(FE_RN_2117_0), .b(n_44061), .o(n_22634) );
ao22f04 FE_RC_4839_0 ( .a(n_37065), .b(n_37492), .c(n_37066), .d(n_46952), .o(n_37577) );
na02f06 FE_RC_483_0 ( .a(FE_RN_148_0), .b(FE_RN_147_0), .o(FE_RN_149_0) );
na02s04 TIMEBOOST_cell_2139 ( .a(n_11604), .b(n_11664), .o(TIMEBOOST_net_684) );
oa22s02 FE_RC_4846_0 ( .a(n_6745), .b(n_6598), .c(FE_OCP_RBN6529_n_6745), .d(n_6599), .o(n_6780) );
no02s06 TIMEBOOST_cell_6150 ( .a(TIMEBOOST_net_1926), .b(n_35113), .o(n_35219) );
no02f06 TIMEBOOST_cell_8759 ( .a(TIMEBOOST_net_2866), .b(n_29481), .o(n_29529) );
na02f08 FE_RC_484_0 ( .a(FE_RN_149_0), .b(n_29122), .o(n_46960) );
ao22s02 FE_RC_4850_0 ( .a(n_2218), .b(n_2293), .c(n_2245), .d(n_2622), .o(n_2342) );
in01s10 FE_RC_4851_0 ( .a(n_23229), .o(FE_RN_2124_0) );
in01m06 FE_RC_4852_0 ( .a(FE_RN_62_0), .o(FE_RN_2125_0) );
na02f10 FE_RC_4853_0 ( .a(FE_RN_2124_0), .b(FE_RN_2125_0), .o(FE_RN_2126_0) );
no02f10 FE_RC_4854_0 ( .a(FE_RN_2126_0), .b(n_23126), .o(n_23246) );
in01m02 FE_RC_4855_0 ( .a(FE_RN_2127_0), .o(n_20239) );
na02m02 FE_RC_4856_0 ( .a(FE_OCPN5101_n_18918), .b(n_20184), .o(FE_RN_2127_0) );
no02f06 TIMEBOOST_cell_4040 ( .a(TIMEBOOST_net_1110), .b(n_39584), .o(TIMEBOOST_net_892) );
no02s01 TIMEBOOST_cell_4041 ( .a(n_15970), .b(n_16210), .o(TIMEBOOST_net_1111) );
oa22m08 FE_RC_4859_0 ( .a(n_39247), .b(n_39477), .c(n_39248), .d(n_39478), .o(n_39559) );
in01s01 FE_RC_4860_0 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_1_), .o(FE_RN_2129_0) );
no02m01 FE_RC_4861_0 ( .a(FE_RN_2129_0), .b(n_6948), .o(FE_RN_2130_0) );
na04m08 TIMEBOOST_cell_7313 ( .a(n_6102), .b(n_6065), .c(FE_OCP_RBN4454_n_6102), .d(n_6064), .o(n_6196) );
no03s08 TIMEBOOST_cell_8197 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_11_), .b(n_45180), .c(n_40674), .o(TIMEBOOST_net_113) );
no02s06 FE_RC_4864_0 ( .a(FE_RN_2132_0), .b(FE_RN_2130_0), .o(n_6973) );
oa22m04 FE_RC_4867_0 ( .a(n_4671), .b(n_4736), .c(FE_OCPN4545_FE_OCP_RBN2850_n_3645), .d(n_4730), .o(n_4916) );
no02s02 FE_RC_4868_0 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_29_), .b(FE_OCP_RBN3938_n_46254), .o(FE_RN_2134_0) );
no02s10 FE_RC_4869_0 ( .a(n_37563), .b(FE_RN_2134_0), .o(n_37609) );
ao22m06 FE_RC_4870_0 ( .a(n_23012), .b(n_23101), .c(n_23011), .d(n_23126), .o(n_23225) );
in01s01 FE_RC_4871_0 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_0_), .o(FE_RN_2135_0) );
no02s06 FE_RC_4872_0 ( .a(FE_RN_2135_0), .b(n_6654), .o(n_6669) );
ao22m02 FE_RC_4873_0 ( .a(n_18240), .b(n_18563), .c(n_18241), .d(n_18562), .o(n_18713) );
in01s01 FE_RC_4874_0 ( .a(n_25418), .o(FE_RN_2136_0) );
na02m08 FE_RC_4875_0 ( .a(n_25786), .b(n_24438), .o(FE_RN_2137_0) );
na02f08 FE_RC_4876_0 ( .a(FE_RN_2136_0), .b(FE_RN_2137_0), .o(FE_RN_2138_0) );
na02s01 FE_RC_4877_0 ( .a(n_24458), .b(n_25486), .o(FE_RN_2139_0) );
no02s02 TIMEBOOST_cell_4557 ( .a(FE_OCPN919_n_17042), .b(n_17070), .o(TIMEBOOST_net_1369) );
na02s04 TIMEBOOST_cell_5687 ( .a(TIMEBOOST_net_1791), .b(n_11575), .o(n_11856) );
na02m08 TIMEBOOST_cell_5475 ( .a(TIMEBOOST_net_1685), .b(n_21786), .o(n_21873) );
in01s01 FE_RC_4881_0 ( .a(n_7321), .o(FE_RN_2142_0) );
in01s02 FE_RC_4882_0 ( .a(FE_RN_2143_0), .o(n_7654) );
no02s01 FE_RC_4883_0 ( .a(FE_RN_2142_0), .b(n_7612), .o(FE_RN_2143_0) );
in01s02 FE_RC_4884_0 ( .a(n_2261), .o(FE_RN_2144_0) );
no02m06 FE_RC_4885_0 ( .a(n_2332), .b(FE_RN_2144_0), .o(FE_RN_2145_0) );
no02m08 FE_RC_4886_0 ( .a(n_2258), .b(FE_RN_2145_0), .o(n_2508) );
ao22f04 FE_RC_4889_0 ( .a(n_34536), .b(n_34872), .c(n_34507), .d(n_34822), .o(n_34921) );
in01m02 FE_RC_4892_0 ( .a(n_46991), .o(FE_RN_2149_0) );
oa22m04 FE_RC_4893_0 ( .a(FE_OCP_RBN5613_n_7730), .b(n_46991), .c(FE_OCP_RBN5606_n_7730), .d(FE_RN_2149_0), .o(n_8154) );
in01s01 FE_RC_4894_0 ( .a(FE_OCPN3557_n_7673), .o(FE_RN_2150_0) );
no02s06 FE_RC_4895_0 ( .a(FE_RN_2150_0), .b(n_7674), .o(n_7727) );
in01s01 FE_RC_4896_0 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_8_), .o(FE_RN_2151_0) );
na02s02 FE_RC_4897_0 ( .a(FE_RN_2151_0), .b(n_7050), .o(n_7107) );
in01f02 FE_RC_4902_0 ( .a(n_13836), .o(FE_RN_2154_0) );
no02f10 FE_RC_4905_0 ( .a(n_23067), .b(n_23066), .o(FE_RN_2156_0) );
ao12f10 FE_RC_4906_0 ( .a(FE_RN_2156_0), .b(n_23066), .c(n_23067), .o(n_23189) );
ao22f04 FE_RC_4908_0 ( .a(n_9982), .b(n_10062), .c(n_10095), .d(n_9983), .o(n_10274) );
oa22f06 FE_RC_4909_0 ( .a(FE_OCP_RBN2936_n_8981), .b(n_10865), .c(n_10712), .d(n_10863), .o(n_11008) );
na02s02 TIMEBOOST_cell_1689 ( .a(n_19615), .b(FE_RN_527_0), .o(TIMEBOOST_net_459) );
oa22s04 FE_RC_4911_0 ( .a(n_7361), .b(n_8074), .c(n_7362), .d(n_8075), .o(n_8187) );
in01s04 FE_RC_4912_0 ( .a(FE_RN_2157_0), .o(n_17791) );
no02s04 FE_RC_4913_0 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_6_), .b(n_17667), .o(FE_RN_2157_0) );
ao22m06 FE_RC_4914_0 ( .a(n_44155), .b(n_22772), .c(n_22677), .d(n_22771), .o(n_22942) );
in01s02 FE_RC_4917_0 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_15_), .o(FE_RN_2159_0) );
na02s02 TIMEBOOST_cell_6028 ( .a(TIMEBOOST_net_1865), .b(n_18813), .o(n_18931) );
no02m04 TIMEBOOST_cell_8721 ( .a(TIMEBOOST_net_2847), .b(n_12478), .o(n_12523) );
na02f08 FE_RC_4920_0 ( .a(n_33382), .b(FE_RN_2161_0), .o(FE_RN_1717_0) );
in01s01 FE_RC_4921_0 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_18_), .o(FE_RN_2162_0) );
no02s06 FE_RC_4922_0 ( .a(FE_RN_2162_0), .b(n_32860), .o(n_32897) );
in01m06 FE_RC_4924_0 ( .a(FE_RN_2164_0), .o(n_39668) );
na02s01 TIMEBOOST_cell_5940 ( .a(TIMEBOOST_net_1821), .b(n_1479), .o(FE_RN_2559_0) );
in01s01 FE_RC_4926_0 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(FE_RN_2165_0) );
no02f06 FE_RC_4927_0 ( .a(FE_RN_2165_0), .b(n_39523), .o(FE_RN_2166_0) );
ao12f04 FE_RC_4928_0 ( .a(FE_RN_2166_0), .b(n_45840), .c(n_39523), .o(n_39592) );
in01m04 FE_RC_4929_0 ( .a(n_32800), .o(FE_RN_2167_0) );
ao22s02 FE_RC_4931_0 ( .a(n_3113), .b(n_3639), .c(n_4719), .d(n_3638), .o(n_3661) );
in01s01 FE_RC_4932_0 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_14_), .o(FE_RN_2168_0) );
na02s06 FE_RC_4933_0 ( .a(FE_RN_2168_0), .b(n_28447), .o(n_28491) );
in01s01 FE_RC_4934_0 ( .a(n_38512), .o(FE_RN_2169_0) );
no02s06 FE_RC_4935_0 ( .a(FE_RN_2169_0), .b(FE_OCP_RBN5897_n_38806), .o(n_38987) );
ao22m02 FE_RC_4937_0 ( .a(n_5907), .b(n_6017), .c(n_5996), .d(n_5910), .o(n_6108) );
in01m04 FE_RC_4938_0 ( .a(FE_RN_2170_0), .o(FE_OCPN895_n_28506) );
na02f06 FE_RC_4939_0 ( .a(n_28452), .b(n_28453), .o(FE_RN_2170_0) );
in01s01 FE_RC_4940_0 ( .a(n_37912), .o(FE_RN_2171_0) );
na02s06 FE_RC_4941_0 ( .a(n_37945), .b(FE_RN_2171_0), .o(n_37975) );
oa22s06 FE_RC_4942_0 ( .a(n_17247), .b(n_17085), .c(n_17245), .d(n_17086), .o(n_17348) );
na02s03 TIMEBOOST_cell_5116 ( .a(n_29550), .b(n_29523), .o(TIMEBOOST_net_1506) );
in01s02 FE_RC_4944_0 ( .a(n_11694), .o(FE_RN_2173_0) );
in01s06 FE_RC_4945_0 ( .a(FE_RN_2174_0), .o(n_12038) );
no02s01 TIMEBOOST_cell_3893 ( .a(n_28679), .b(n_28680), .o(TIMEBOOST_net_1037) );
in01s06 FE_RC_4947_0 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_4_), .o(FE_RN_2175_0) );
na02m08 TIMEBOOST_cell_5037 ( .a(TIMEBOOST_net_1466), .b(n_19708), .o(n_19806) );
no02f04 TIMEBOOST_cell_5038 ( .a(n_44871), .b(n_37889), .o(TIMEBOOST_net_1467) );
in01s02 FE_RC_4950_0 ( .a(n_9425), .o(FE_RN_2177_0) );
no02m02 FE_RC_4951_0 ( .a(n_9611), .b(FE_RN_2177_0), .o(FE_RN_2178_0) );
ao12f02 FE_RC_4953_0 ( .a(FE_RN_2178_0), .b(n_9611), .c(FE_RN_2177_0), .o(n_9788) );
no02m01 FE_RC_4954_0 ( .a(n_7730), .b(n_7832), .o(FE_RN_2180_0) );
no02m08 FE_RC_4955_0 ( .a(n_7948), .b(FE_RN_2180_0), .o(n_7985) );
oa22s02 FE_RC_4956_0 ( .a(n_3743), .b(n_3875), .c(n_3799), .d(FE_OCP_RBN5916_n_3875), .o(n_4099) );
na02s01 FE_RC_4957_0 ( .a(n_37392), .b(n_37393), .o(FE_RN_2181_0) );
na02s02 FE_RC_4958_0 ( .a(FE_RN_2181_0), .b(n_37893), .o(n_37956) );
ao22m04 FE_RC_4959_0 ( .a(n_12593), .b(FE_OCP_RBN5582_n_12802), .c(n_12592), .d(FE_OCP_RBN5584_n_12802), .o(n_13005) );
in01s01 FE_RC_495_0 ( .a(n_13257), .o(FE_RN_150_0) );
oa22f02 FE_RC_4961_0 ( .a(FE_OCP_RBN4139_n_7743), .b(n_8402), .c(FE_OCP_RBN5635_n_7708), .d(FE_OCP_RBN2734_n_8402), .o(n_8525) );
in01s01 FE_RC_4962_0 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_16_), .o(FE_RN_2182_0) );
in01s01 FE_RC_4963_0 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_17_), .o(FE_RN_2183_0) );
no02s01 FE_RC_4964_0 ( .a(FE_RN_2182_0), .b(FE_RN_2183_0), .o(FE_RN_2184_0) );
no02m06 FE_RC_4965_0 ( .a(FE_RN_2184_0), .b(FE_OCP_RBN2469_n_33034), .o(n_33135) );
ao22m04 FE_RC_4968_0 ( .a(n_7541), .b(n_8547), .c(n_7540), .d(n_8546), .o(n_8664) );
ao22m04 FE_RC_4969_0 ( .a(FE_OCP_RBN4040_n_37707), .b(n_37775), .c(n_37734), .d(n_37776), .o(n_37848) );
in01s04 FE_RC_496_0 ( .a(n_14194), .o(FE_RN_151_0) );
in01s01 FE_RC_4970_0 ( .a(n_8069), .o(FE_RN_2186_0) );
na02m02 FE_RC_4972_0 ( .a(FE_RN_2186_0), .b(n_8776), .o(FE_RN_2187_0) );
in01s01 FE_RC_4978_0 ( .a(FE_OCP_RBN2540_n_12880), .o(FE_RN_2191_0) );
in01m04 FE_RC_4979_0 ( .a(FE_RN_2192_0), .o(n_47253) );
no02s06 FE_RC_497_0 ( .a(FE_RN_151_0), .b(FE_RN_150_0), .o(FE_RN_152_0) );
no02m04 FE_RC_4980_0 ( .a(FE_RN_2191_0), .b(n_13483), .o(FE_RN_2192_0) );
in01s01 FE_RC_4981_0 ( .a(n_18366), .o(FE_RN_2193_0) );
in01s02 FE_RC_4982_0 ( .a(n_18718), .o(FE_RN_2194_0) );
no02m04 FE_RC_4983_0 ( .a(FE_RN_2193_0), .b(FE_RN_2194_0), .o(FE_RN_2195_0) );
na02m04 FE_RC_4984_0 ( .a(FE_OCP_RBN7023_n_18650), .b(FE_RN_2195_0), .o(n_18799) );
in01s01 FE_RC_4985_0 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_7_), .o(FE_RN_2196_0) );
in01s04 FE_RC_4986_0 ( .a(FE_RN_2197_0), .o(n_32821) );
no02s02 TIMEBOOST_cell_1629 ( .a(n_3705), .b(FE_RN_2301_0), .o(TIMEBOOST_net_429) );
na02f06 TIMEBOOST_cell_7993 ( .a(TIMEBOOST_net_2627), .b(n_26180), .o(n_26361) );
in01s01 FE_RC_4991_0 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_6_), .o(FE_RN_2200_0) );
no04f06 TIMEBOOST_cell_5743 ( .a(n_33567), .b(n_34037), .c(n_47249), .d(n_33642), .o(n_33693) );
na02m02 TIMEBOOST_cell_8677 ( .a(TIMEBOOST_net_2825), .b(n_36692), .o(n_36706) );
na02f02 FE_RC_4996_0 ( .a(n_9655), .b(n_9603), .o(FE_RN_2202_0) );
na02f04 FE_RC_4997_0 ( .a(n_9633), .b(FE_RN_2202_0), .o(n_9921) );
in01s02 FE_RC_4998_0 ( .a(n_9396), .o(FE_RN_2203_0) );
in01s02 FE_RC_4999_0 ( .a(n_9387), .o(FE_RN_2204_0) );
na02s06 TIMEBOOST_cell_4209 ( .a(n_12253), .b(n_12252), .o(TIMEBOOST_net_1195) );
oa22m02 FE_RC_5000_0 ( .a(FE_RN_2203_0), .b(n_9387), .c(n_9396), .d(FE_RN_2204_0), .o(n_9641) );
in01s01 FE_RC_5001_0 ( .a(n_7925), .o(FE_RN_2205_0) );
in01f02 FE_RC_5002_0 ( .a(FE_RN_2206_0), .o(n_8651) );
na02f02 FE_RC_5003_0 ( .a(FE_RN_2205_0), .b(n_8580), .o(FE_RN_2206_0) );
no02s02 TIMEBOOST_cell_4139 ( .a(n_11439), .b(n_10613), .o(TIMEBOOST_net_1160) );
in01f04 FE_RC_5005_0 ( .a(FE_RN_2208_0), .o(n_3303) );
no02m06 TIMEBOOST_cell_4146 ( .a(TIMEBOOST_net_1163), .b(n_36630), .o(n_36751) );
na02m02 FE_RC_5009_0 ( .a(FE_OCP_RBN6724_n_44055), .b(n_9284), .o(FE_RN_2210_0) );
in01s01 FE_RC_5010_0 ( .a(n_44055), .o(FE_RN_2211_0) );
oa12m02 FE_RC_5011_0 ( .a(FE_RN_2210_0), .b(FE_RN_2211_0), .c(n_9284), .o(n_9519) );
na02m02 FE_RC_5012_0 ( .a(n_9605), .b(n_9781), .o(FE_RN_2212_0) );
no02m02 FE_RC_5013_0 ( .a(n_9605), .b(n_9781), .o(FE_RN_2213_0) );
oa12f02 FE_RC_5014_0 ( .a(FE_RN_2212_0), .b(FE_RN_2213_0), .c(n_9506), .o(n_9655) );
in01s01 FE_RC_5015_0 ( .a(n_18335), .o(FE_RN_2214_0) );
in01s02 FE_RC_5016_0 ( .a(FE_RN_2215_0), .o(FE_RN_519_0) );
no02s02 FE_RC_5017_0 ( .a(n_18864), .b(FE_RN_2214_0), .o(FE_RN_2215_0) );
oa22m08 FE_RC_5020_0 ( .a(n_24224), .b(n_23760), .c(FE_RN_1306_0), .d(n_24225), .o(n_24305) );
oa22s02 FE_RC_5022_0 ( .a(n_3274), .b(FE_OCP_RBN6659_n_2829), .c(n_2664), .d(n_2829), .o(n_2930) );
in01s01 FE_RC_5024_0 ( .a(n_8232), .o(FE_RN_2217_0) );
in01m04 FE_RC_5025_0 ( .a(FE_RN_2218_0), .o(n_9570) );
no02s04 FE_RC_5026_0 ( .a(FE_RN_2217_0), .b(n_9450), .o(FE_RN_2218_0) );
in01s01 FE_RC_5027_0 ( .a(n_8232), .o(FE_RN_2219_0) );
no02s06 FE_RC_5029_0 ( .a(n_9342), .b(FE_RN_2219_0), .o(FE_RN_2220_0) );
in01f02 FE_RC_5031_0 ( .a(FE_RN_2222_0), .o(n_9077) );
ao22f04 FE_RC_5033_0 ( .a(FE_OCP_RBN4150_n_13616), .b(n_13713), .c(n_13616), .d(n_13746), .o(n_13849) );
oa22m10 FE_RC_5034_0 ( .a(n_32752), .b(n_45741), .c(n_32680), .d(FE_OCP_RBN5524_n_32752), .o(n_32829) );
ao22f04 FE_RC_5035_0 ( .a(n_5998), .b(n_6021), .c(n_5997), .d(FE_OCP_RBN6169_n_6021), .o(n_6135) );
oa22m04 FE_RC_5036_0 ( .a(n_18032), .b(n_19353), .c(n_19218), .d(FE_OCP_RBN2063_n_19353), .o(n_19462) );
ao22s20 FE_RC_5039_0 ( .a(n_32622), .b(FE_OCP_RBN7013_n_44962), .c(delay_xor_ln22_unr21_stage8_stallmux_q_4_), .d(FE_OCP_RBN4633_n_44962), .o(n_32680) );
oa22s02 FE_RC_5040_0 ( .a(FE_OFN770_n_46196), .b(FE_OCP_RBN3454_n_6557), .c(FE_OFN4787_n_46137), .d(n_6557), .o(n_46185) );
no02m02 FE_RC_5042_0 ( .a(n_13272), .b(n_14519), .o(FE_RN_2224_0) );
in01s03 FE_RC_5043_0 ( .a(n_24810), .o(FE_RN_2225_0) );
no02s08 FE_RC_5044_0 ( .a(n_24975), .b(FE_RN_2225_0), .o(n_24992) );
ao22m02 FE_RC_5045_0 ( .a(FE_OCPN931_n_7817), .b(n_8637), .c(FE_OCP_RBN2598_n_7743), .d(FE_OCP_RBN5746_n_8637), .o(n_8790) );
oa22f04 FE_RC_5046_0 ( .a(FE_OCP_RBN2714_n_24501), .b(n_44423), .c(n_24555), .d(n_24990), .o(n_25102) );
na02s03 FE_RC_5047_0 ( .a(n_13757), .b(n_12935), .o(FE_RN_2226_0) );
in01s01 FE_RC_5049_0 ( .a(FE_OFN4808_n_28820), .o(FE_RN_2227_0) );
na02m08 FE_RC_5050_0 ( .a(FE_RN_2227_0), .b(n_29347), .o(FE_RN_2228_0) );
in01s01 FE_RC_5051_0 ( .a(FE_OFN4808_n_28820), .o(FE_RN_2229_0) );
oa12m08 FE_RC_5052_0 ( .a(FE_RN_2228_0), .b(FE_RN_2229_0), .c(n_29347), .o(n_29448) );
oa22m04 FE_RC_5053_0 ( .a(n_28845), .b(FE_OCP_RBN5672_n_29425), .c(n_29425), .d(n_28846), .o(n_29553) );
in01s01 FE_RC_5054_0 ( .a(FE_OCPN1722_n_29060), .o(FE_RN_2230_0) );
na02s10 FE_RC_5055_0 ( .a(n_29922), .b(FE_RN_2230_0), .o(n_29952) );
ao22s04 FE_RC_5056_0 ( .a(n_7736), .b(n_8914), .c(n_7735), .d(n_8921), .o(n_9057) );
ao22m20 FE_RC_5058_0 ( .a(n_44962), .b(n_32615), .c(delay_xor_ln22_unr21_stage8_stallmux_q_2_), .d(FE_OCP_RBN7015_n_44962), .o(n_32663) );
na02m02 FE_RC_5059_0 ( .a(FE_RN_1065_0), .b(n_19470), .o(FE_RN_2231_0) );
oa12f02 FE_RC_5060_0 ( .a(FE_RN_2231_0), .b(n_19470), .c(FE_RN_1065_0), .o(n_19601) );
in01s01 FE_RC_5061_0 ( .a(FE_OCPN1327_n_16192), .o(FE_RN_2232_0) );
no02s06 FE_RC_5062_0 ( .a(FE_OCP_RBN6175_n_16923), .b(FE_RN_2232_0), .o(n_17120) );
in01s01 FE_RC_5063_0 ( .a(FE_OCP_RBN3084_n_15314), .o(FE_RN_2233_0) );
no02m10 FE_RC_5064_0 ( .a(n_16912), .b(FE_RN_2233_0), .o(n_17045) );
no02s02 FE_RC_5065_0 ( .a(n_4400), .b(n_4277), .o(FE_RN_2234_0) );
no02s04 FE_RC_5066_0 ( .a(n_4304), .b(FE_RN_2234_0), .o(n_4572) );
in01m02 FE_RC_5067_0 ( .a(n_29624), .o(FE_RN_2235_0) );
in01s01 FE_RC_5068_0 ( .a(n_29615), .o(FE_RN_2236_0) );
no02f02 FE_RC_5069_0 ( .a(FE_RN_2235_0), .b(FE_RN_2236_0), .o(FE_RN_2237_0) );
no02f02 FE_RC_5070_0 ( .a(FE_RN_2237_0), .b(n_29808), .o(FE_RN_2238_0) );
in01s01 FE_RC_5071_0 ( .a(n_29615), .o(FE_RN_2239_0) );
no02s02 FE_RC_5072_0 ( .a(FE_OCP_RBN5719_n_29624), .b(FE_RN_2239_0), .o(FE_RN_2240_0) );
ao12f02 FE_RC_5073_0 ( .a(FE_RN_2238_0), .b(FE_RN_2240_0), .c(n_29808), .o(n_29839) );
ao22m04 FE_RC_5074_0 ( .a(FE_OCPN1741_n_18591), .b(n_19393), .c(n_18592), .d(FE_OCP_RBN2663_n_19393), .o(n_19538) );
in01s02 FE_RC_5075_0 ( .a(FE_RN_2241_0), .o(FE_OCPN1913_n_2669) );
no02s02 FE_RC_5076_0 ( .a(n_2622), .b(n_2623), .o(FE_RN_2241_0) );
ao22m06 FE_RC_5077_0 ( .a(n_15369), .b(n_15906), .c(n_15370), .d(n_15820), .o(n_16084) );
in01m03 FE_RC_5078_0 ( .a(FE_RN_2242_0), .o(n_29984) );
no02m02 FE_RC_5079_0 ( .a(FE_OCP_DRV_N1468_n_28775), .b(n_29839), .o(FE_RN_2242_0) );
oa22f04 FE_RC_5080_0 ( .a(n_38722), .b(FE_OCP_RBN2897_n_38750), .c(n_38720), .d(n_38750), .o(n_38800) );
oa22s02 FE_RC_5081_0 ( .a(n_6418), .b(n_6351), .c(n_6350), .d(n_6388), .o(n_6529) );
ao22m06 FE_RC_5082_0 ( .a(n_24624), .b(FE_OCP_RBN5717_n_24718), .c(n_24718), .d(FE_OFN5074_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24875) );
na02m04 FE_RC_5083_0 ( .a(n_13338), .b(n_13400), .o(FE_RN_2243_0) );
na02m06 FE_RC_5084_0 ( .a(FE_RN_2243_0), .b(n_13360), .o(n_13397) );
in01m04 FE_RC_5085_0 ( .a(FE_RN_2244_0), .o(n_9355) );
no02m04 FE_RC_5086_0 ( .a(FE_OCP_RBN6630_n_8269), .b(n_9125), .o(FE_RN_2244_0) );
ao22f08 FE_RC_5087_0 ( .a(n_24620), .b(n_24798), .c(n_22280), .d(n_24799), .o(n_24891) );
na02f06 FE_RC_5088_0 ( .a(n_19877), .b(n_19739), .o(FE_RN_2245_0) );
na02f08 FE_RC_5089_0 ( .a(FE_RN_2245_0), .b(n_19770), .o(n_19854) );
ao22m02 FE_RC_5090_0 ( .a(n_2249), .b(n_2702), .c(n_2230), .d(n_1978), .o(n_2344) );
in01s01 TIMEBOOST_cell_5918 ( .a(TIMEBOOST_net_1806), .o(TIMEBOOST_net_1807) );
no02s01 TIMEBOOST_cell_2902 ( .a(n_33063), .b(n_33104), .o(TIMEBOOST_net_742) );
no02s06 FE_RC_5093_0 ( .a(FE_RN_2247_0), .b(n_34135), .o(FE_RN_2248_0) );
na02s04 FE_RC_5094_0 ( .a(n_34144), .b(n_34146), .o(FE_RN_2249_0) );
in01s02 FE_RC_5095_0 ( .a(n_34187), .o(FE_RN_2250_0) );
no02m04 FE_RC_5096_0 ( .a(FE_RN_2249_0), .b(FE_RN_2250_0), .o(FE_RN_2251_0) );
no02f08 TIMEBOOST_cell_8817 ( .a(TIMEBOOST_net_2895), .b(n_15357), .o(TIMEBOOST_net_1539) );
no02s01 TIMEBOOST_cell_5302 ( .a(n_19967), .b(n_19945), .o(TIMEBOOST_net_1599) );
in01s01 FE_RC_5100_0 ( .a(FE_OCPN4542_FE_OCP_RBN2812_n_8835), .o(FE_RN_2253_0) );
na02s02 FE_RC_5101_0 ( .a(FE_RN_2253_0), .b(n_10148), .o(n_10324) );
in01s01 FE_RC_5102_0 ( .a(FE_OCP_RBN2717_n_8242), .o(FE_RN_2254_0) );
in01s02 FE_RC_5103_0 ( .a(FE_RN_2255_0), .o(n_9366) );
na02s02 FE_RC_5104_0 ( .a(FE_RN_2254_0), .b(n_9087), .o(FE_RN_2255_0) );
in01s01 FE_RC_5107_0 ( .a(FE_OCPN3589_n_21419), .o(FE_RN_2257_0) );
no02m01 FE_RC_5108_0 ( .a(FE_RN_2257_0), .b(FE_OCP_RBN4468_n_44267), .o(n_22194) );
in01s01 FE_RC_5109_0 ( .a(FE_OCPN1312_FE_OCP_RBN1024_n_24125), .o(FE_RN_2258_0) );
oa22f02 FE_RC_510_0 ( .a(n_14714), .b(n_14658), .c(n_14657), .d(n_14715), .o(n_14814) );
na02m06 FE_RC_5111_0 ( .a(FE_RN_2258_0), .b(FE_OCP_RBN2910_n_25178), .o(FE_RN_2259_0) );
in01s02 FE_RC_5112_0 ( .a(n_14190), .o(FE_RN_2260_0) );
na02s01 TIMEBOOST_cell_6388 ( .a(TIMEBOOST_net_2045), .b(n_27393), .o(n_27523) );
no02m04 TIMEBOOST_cell_4969 ( .a(TIMEBOOST_net_1432), .b(n_37515), .o(TIMEBOOST_net_1203) );
ao22f04 FE_RC_5118_0 ( .a(FE_OCP_RBN2676_n_8163), .b(n_8370), .c(FE_OCP_RBN2677_n_8163), .d(n_8439), .o(n_8489) );
ao22m04 FE_RC_5119_0 ( .a(n_5093), .b(n_5429), .c(n_5094), .d(n_5428), .o(n_5555) );
oa22f04 FE_RC_5120_0 ( .a(n_23963), .b(n_24721), .c(n_23962), .d(n_24720), .o(n_24857) );
no02m06 FE_RC_5121_0 ( .a(n_21429), .b(n_21509), .o(FE_RN_2264_0) );
na02m08 FE_RC_5122_0 ( .a(FE_RN_2264_0), .b(n_21558), .o(n_21658) );
no02f06 TIMEBOOST_cell_2865 ( .a(TIMEBOOST_net_723), .b(FE_RN_2082_0), .o(n_45718) );
na02f06 TIMEBOOST_cell_6735 ( .a(FE_OCP_RBN1601_n_14638), .b(FE_OCP_RBN4202_n_13796), .o(TIMEBOOST_net_2125) );
na02s08 FE_RC_5125_0 ( .a(FE_RN_2266_0), .b(n_34463), .o(n_34514) );
no02s01 FE_RC_5126_0 ( .a(n_33541), .b(n_33583), .o(FE_RN_2267_0) );
no02s06 FE_RC_5127_0 ( .a(FE_RN_2267_0), .b(FE_OCP_RBN6665_n_34297), .o(n_34490) );
oa22f08 FE_RC_5128_0 ( .a(n_20266), .b(n_20208), .c(FE_OCPN1316_n_20265), .d(n_20207), .o(n_20299) );
in01s01 FE_RC_5129_0 ( .a(n_45073), .o(FE_RN_2268_0) );
in01m06 FE_RC_5130_0 ( .a(FE_RN_2269_0), .o(n_21507) );
na02m04 FE_RC_5131_0 ( .a(FE_RN_2268_0), .b(n_21361), .o(FE_RN_2269_0) );
oa22m04 FE_RC_5133_0 ( .a(n_5095), .b(n_5561), .c(n_5096), .d(n_5562), .o(n_5693) );
no02m04 FE_RC_5134_0 ( .a(FE_OCP_RBN4441_n_5891), .b(n_5812), .o(FE_RN_2270_0) );
na02m04 FE_RC_5135_0 ( .a(FE_RN_2270_0), .b(n_6015), .o(FE_RN_2271_0) );
na03m20 TIMEBOOST_cell_4586 ( .a(FE_RN_1594_0), .b(FE_OCP_RBN2030_n_44722), .c(n_27911), .o(n_28036) );
no03f08 TIMEBOOST_cell_5866 ( .a(n_16682), .b(n_16600), .c(FE_OCP_RBN4458_FE_RN_1190_0), .o(n_16749) );
na02f04 FE_RC_5138_0 ( .a(n_5879), .b(FE_RN_2273_0), .o(FE_RN_2274_0) );
na02s06 FE_RC_5139_0 ( .a(FE_RN_2271_0), .b(FE_RN_2274_0), .o(n_6077) );
ao22f04 FE_RC_513_0 ( .a(FE_OCP_RBN7131_n_29262), .b(n_45186), .c(FE_OCP_RBN7130_n_29262), .d(n_29451), .o(n_29577) );
in01s01 FE_RC_5140_0 ( .a(n_7725), .o(FE_RN_2275_0) );
in01m02 FE_RC_5141_0 ( .a(FE_RN_2276_0), .o(n_8392) );
na02m02 FE_RC_5142_0 ( .a(FE_RN_2275_0), .b(n_8271), .o(FE_RN_2276_0) );
in01m02 FE_RC_5143_0 ( .a(FE_RN_2277_0), .o(FE_OCP_RBN4440_n_5891) );
no02m01 FE_RC_5144_0 ( .a(n_5746), .b(FE_OCP_RBN3066_n_4294), .o(FE_RN_2277_0) );
oa22f02 FE_RC_5145_0 ( .a(n_14809), .b(n_14884), .c(n_14810), .d(n_14885), .o(n_14985) );
oa22m04 FE_RC_5146_0 ( .a(n_24461), .b(n_24719), .c(FE_RN_1765_0), .d(n_24486), .o(n_24826) );
in01s01 FE_RC_5148_0 ( .a(n_8676), .o(FE_RN_2278_0) );
na02m02 FE_RC_5149_0 ( .a(n_7929), .b(FE_RN_2278_0), .o(FE_RN_2279_0) );
oa12m02 FE_RC_5150_0 ( .a(FE_RN_2279_0), .b(FE_OCP_RBN6579_n_8676), .c(n_7929), .o(n_8115) );
ao22f02 FE_RC_5151_0 ( .a(n_5136), .b(n_5532), .c(n_5137), .d(FE_OCP_RBN4400_n_5532), .o(n_5627) );
oa22m04 FE_RC_5152_0 ( .a(n_25562), .b(n_25845), .c(FE_OCP_RBN2978_n_25562), .d(n_25846), .o(n_25934) );
in01s01 FE_RC_5154_0 ( .a(FE_OCP_RBN2833_n_13962), .o(FE_RN_2280_0) );
na02f02 FE_RC_5155_0 ( .a(FE_RN_2280_0), .b(n_14768), .o(FE_RN_2281_0) );
oa12f02 FE_RC_5156_0 ( .a(FE_RN_2281_0), .b(n_14768), .c(FE_OCP_RBN5799_n_13962), .o(n_14873) );
no02m04 TIMEBOOST_cell_5592 ( .a(n_31850), .b(n_31835), .o(TIMEBOOST_net_1744) );
in01s02 FE_RC_5158_0 ( .a(FE_RN_2283_0), .o(FE_OCP_RBN4444_n_5849) );
na02s03 TIMEBOOST_cell_8600 ( .a(n_39130), .b(n_39068), .o(TIMEBOOST_net_2787) );
oa22f02 FE_RC_5162_0 ( .a(n_10068), .b(n_9987), .c(n_10047), .d(FE_OCP_RBN6004_n_10068), .o(n_10326) );
in01s01 FE_RC_5163_0 ( .a(FE_OCP_DRV_N1417_n_32985), .o(FE_RN_2284_0) );
na02f04 FE_RC_5164_0 ( .a(n_33780), .b(FE_RN_2284_0), .o(n_33880) );
oa22m02 FE_RC_5165_0 ( .a(n_9856), .b(n_9801), .c(FE_OCP_RBN5981_n_9856), .d(n_9800), .o(n_10015) );
ao22f04 FE_RC_5166_0 ( .a(n_15295), .b(n_15655), .c(n_15294), .d(n_15698), .o(n_15861) );
in01s01 FE_RC_5167_0 ( .a(n_7788), .o(FE_RN_2285_0) );
in01s01 FE_RC_5168_0 ( .a(n_7311), .o(FE_RN_2286_0) );
na02s01 FE_RC_5169_0 ( .a(n_7788), .b(n_7311), .o(FE_RN_2287_0) );
oa22f02 FE_RC_516_0 ( .a(n_15071), .b(FE_OCP_RBN5982_n_15160), .c(FE_OCP_RBN4343_n_15071), .d(n_15160), .o(n_15314) );
ao22s04 FE_RC_5170_0 ( .a(FE_RN_2286_0), .b(FE_RN_2285_0), .c(FE_RN_2287_0), .d(n_7745), .o(n_7810) );
oa22f04 FE_RC_5171_0 ( .a(n_24262), .b(FE_OCP_RBN4158_n_24222), .c(n_24222), .d(FE_OCP_RBN983_n_24262), .o(n_24426) );
in01s01 FE_RC_5172_0 ( .a(FE_OCPN1321_n_33714), .o(FE_RN_2288_0) );
na02f06 FE_RC_5173_0 ( .a(FE_RN_2288_0), .b(n_33715), .o(n_33777) );
ao22m04 FE_RC_5174_0 ( .a(n_26265), .b(n_25725), .c(n_25724), .d(n_26266), .o(n_26398) );
no02m06 FE_RC_5176_0 ( .a(FE_RN_1185_0), .b(n_26553), .o(FE_RN_2289_0) );
oa22f04 FE_RC_5177_0 ( .a(n_9030), .b(n_9042), .c(FE_OCP_RBN5883_n_9042), .d(FE_OCP_RBN2922_n_9030), .o(n_9247) );
oa22m02 FE_RC_5178_0 ( .a(n_33752), .b(n_33750), .c(n_33769), .d(FE_OCP_RBN1811_n_33750), .o(n_33868) );
ao22s04 FE_RC_5179_0 ( .a(n_24137), .b(FE_OCP_RBN4148_n_24173), .c(n_24121), .d(n_24173), .o(n_24306) );
oa22f06 FE_RC_5180_0 ( .a(FE_OCPN1338_n_25775), .b(n_26502), .c(n_25776), .d(n_26503), .o(n_26622) );
oa22m04 FE_RC_5183_0 ( .a(n_11181), .b(FE_OCP_RBN6134_n_11221), .c(n_11221), .d(n_11217), .o(n_11308) );
oa22f02 FE_RC_5184_0 ( .a(n_10757), .b(n_10790), .c(n_10758), .d(n_10789), .o(n_10906) );
in01s01 FE_RC_5185_0 ( .a(n_45066), .o(FE_RN_2291_0) );
no02f04 FE_RC_5186_0 ( .a(n_20719), .b(FE_RN_2291_0), .o(FE_RN_1490_0) );
no02m10 TIMEBOOST_cell_1039 ( .a(FE_RN_236_0), .b(n_18026), .o(TIMEBOOST_net_134) );
no02f06 TIMEBOOST_cell_5405 ( .a(TIMEBOOST_net_1650), .b(n_26795), .o(n_26911) );
no02m10 TIMEBOOST_cell_1040 ( .a(TIMEBOOST_net_134), .b(n_18115), .o(n_18177) );
na02s04 FE_RC_5190_0 ( .a(n_3977), .b(n_4275), .o(FE_RN_2294_0) );
na02s04 FE_RC_5191_0 ( .a(FE_RN_2294_0), .b(n_4329), .o(n_4553) );
oa22f08 FE_RC_5192_0 ( .a(n_16440), .b(n_16596), .c(n_16463), .d(FE_OCP_RBN3360_n_16596), .o(n_16702) );
ao22m06 FE_RC_5193_0 ( .a(FE_OCP_RBN3103_n_20710), .b(n_21014), .c(FE_OCP_RBN4364_n_20710), .d(n_21015), .o(n_21163) );
na02s02 FE_RC_5196_0 ( .a(n_35824), .b(n_35784), .o(FE_RN_2296_0) );
na02s06 FE_RC_5197_0 ( .a(FE_OCP_RBN4910_n_44222), .b(FE_RN_2296_0), .o(FE_RN_2297_0) );
na02m10 FE_RC_5198_0 ( .a(n_36013), .b(FE_RN_2297_0), .o(n_36071) );
oa22f04 FE_RC_5202_0 ( .a(n_16489), .b(FE_OCP_RBN6135_n_16553), .c(n_16553), .d(n_16514), .o(n_16638) );
in01s01 FE_RC_5205_0 ( .a(n_3666), .o(FE_RN_2301_0) );
na02f06 TIMEBOOST_cell_7786 ( .a(n_42223), .b(n_42208), .o(TIMEBOOST_net_2524) );
na02s01 TIMEBOOST_cell_6639 ( .a(n_18568), .b(n_18664), .o(TIMEBOOST_net_2077) );
ao22m02 FE_RC_5208_0 ( .a(n_45070), .b(n_20950), .c(n_45032), .d(n_20949), .o(n_21084) );
in01s01 FE_RC_5211_0 ( .a(FE_OCP_RBN2892_n_14460), .o(FE_RN_2304_0) );
na02m06 FE_RC_5212_0 ( .a(FE_RN_2304_0), .b(n_16218), .o(n_16436) );
in01s01 FE_RC_5213_0 ( .a(n_45073), .o(FE_RN_2305_0) );
in01m04 FE_RC_5214_0 ( .a(FE_RN_2306_0), .o(n_21397) );
na02m02 FE_RC_5215_0 ( .a(FE_RN_2305_0), .b(n_21233), .o(FE_RN_2306_0) );
in01s02 FE_RC_5219_0 ( .a(n_26666), .o(FE_RN_2309_0) );
na02s06 FE_RC_5220_0 ( .a(FE_OCP_RBN6871_FE_RN_2289_0), .b(FE_RN_2309_0), .o(FE_RN_2310_0) );
no02f08 FE_RC_5221_0 ( .a(n_26785), .b(FE_RN_2310_0), .o(n_26920) );
na02s01 FE_RC_5222_0 ( .a(FE_OCP_RBN3181_n_10477), .b(FE_OCP_RBN4385_n_10570), .o(FE_RN_2311_0) );
na02s06 FE_RC_5223_0 ( .a(FE_OCP_RBN4482_n_11439), .b(FE_RN_2311_0), .o(n_11664) );
no02f06 FE_RC_5224_0 ( .a(n_21707), .b(n_21659), .o(FE_RN_2312_0) );
no02f08 FE_RC_5225_0 ( .a(FE_RN_2312_0), .b(n_21660), .o(n_21811) );
oa22s02 FE_RC_5226_0 ( .a(FE_OFN4787_n_46137), .b(n_6646), .c(FE_OFN770_n_46196), .d(n_6670), .o(n_46190) );
oa22m02 FE_RC_5230_0 ( .a(n_11501), .b(n_11553), .c(n_11500), .d(n_11523), .o(n_11778) );
oa22m02 FE_RC_5231_0 ( .a(n_11750), .b(n_11947), .c(n_11749), .d(n_11913), .o(n_12144) );
oa22f02 FE_RC_5232_0 ( .a(FE_OCPN5280_n_30614), .b(n_35262), .c(n_30633), .d(n_35281), .o(n_35340) );
in01s02 FE_RC_5233_0 ( .a(n_35326), .o(FE_RN_2314_0) );
na02m06 FE_RC_5234_0 ( .a(n_35342), .b(FE_RN_2314_0), .o(n_35358) );
oa22m02 FE_RC_5235_0 ( .a(FE_OCP_RBN6865_n_46285), .b(n_11731), .c(FE_OCP_RBN4448_FE_OFN760_n_46337), .d(n_11682), .o(n_46363) );
oa22s02 FE_RC_5236_0 ( .a(FE_OCP_RBN6865_n_46285), .b(n_11778), .c(FE_OCP_RBN4448_FE_OFN760_n_46337), .d(n_11725), .o(n_46361) );
no02m04 FE_RC_5239_0 ( .a(n_25963), .b(n_27121), .o(FE_RN_2316_0) );
no02m06 FE_RC_5240_0 ( .a(n_27086), .b(FE_RN_2316_0), .o(n_27276) );
oa22f04 FE_RC_5242_0 ( .a(n_35225), .b(n_35347), .c(n_35346), .d(n_35226), .o(n_35421) );
oa22m02 FE_RC_5243_0 ( .a(FE_OCP_RBN6865_n_46285), .b(n_12145), .c(FE_OFN765_n_46337), .d(n_12102), .o(n_46353) );
oa22m04 FE_RC_5244_0 ( .a(n_11743), .b(n_11980), .c(n_11744), .d(FE_OCP_RBN3437_n_11980), .o(n_12162) );
in01s01 FE_RC_5245_0 ( .a(FE_OCP_RBN5206_n_20504), .o(FE_RN_2317_0) );
no02m06 FE_RC_5246_0 ( .a(FE_RN_2317_0), .b(n_22005), .o(n_22027) );
in01s06 FE_RC_5249_0 ( .a(FE_RN_2318_0), .o(n_17515) );
na02s02 FE_RC_5250_0 ( .a(n_17233), .b(n_17250), .o(FE_RN_2318_0) );
in01m04 FE_RC_5251_0 ( .a(FE_OCP_RBN6839_FE_RN_2660_0), .o(FE_RN_2319_0) );
no02f08 FE_RC_5252_0 ( .a(FE_RN_2319_0), .b(n_31443), .o(n_31492) );
in01s04 FE_RC_5253_0 ( .a(FE_RN_2320_0), .o(n_27192) );
na02m04 FE_RC_5254_0 ( .a(n_25363), .b(n_26844), .o(FE_RN_2320_0) );
in01f02 FE_RC_5255_0 ( .a(FE_RN_2321_0), .o(n_21792) );
no02m02 FE_RC_5256_0 ( .a(n_20059), .b(n_21656), .o(FE_RN_2321_0) );
na02f06 FE_RC_5257_0 ( .a(n_21353), .b(n_21159), .o(FE_RN_2322_0) );
na02f08 FE_RC_5258_0 ( .a(FE_RN_2322_0), .b(n_21186), .o(n_21470) );
in01s01 FE_RC_5260_0 ( .a(n_27416), .o(FE_RN_2323_0) );
na02s01 FE_RC_5261_0 ( .a(n_25810), .b(FE_RN_2323_0), .o(FE_RN_2324_0) );
na02m08 FE_RC_5262_0 ( .a(FE_RN_2324_0), .b(n_27167), .o(n_27206) );
oa22m04 FE_RC_5264_0 ( .a(n_27582), .b(n_27489), .c(n_27488), .d(n_45745), .o(n_27655) );
oa22s02 FE_RC_5265_0 ( .a(n_17315), .b(FE_OCP_RBN3427_n_17510), .c(n_17316), .d(n_17510), .o(n_17687) );
oa22s02 FE_RC_5266_0 ( .a(n_17313), .b(n_17557), .c(n_17314), .d(n_17558), .o(n_17725) );
in01s01 FE_RC_5267_0 ( .a(FE_OCP_RBN1032_n_25844), .o(FE_RN_2325_0) );
no02s06 FE_RC_5268_0 ( .a(FE_RN_2325_0), .b(FE_OCP_RBN6218_n_27110), .o(n_27464) );
in01s01 FE_RC_5269_0 ( .a(FE_OCPUNCON3481_n_21058), .o(FE_RN_2326_0) );
ao22f06 FE_RC_526_0 ( .a(n_30219), .b(n_30453), .c(n_30218), .d(n_30454), .o(n_30541) );
no02f04 FE_RC_5270_0 ( .a(n_21059), .b(FE_RN_2326_0), .o(n_21174) );
no02s01 FE_RC_5271_0 ( .a(FE_RN_1883_0), .b(n_30573), .o(FE_RN_2327_0) );
no02s08 FE_RC_5272_0 ( .a(FE_RN_2327_0), .b(n_31835), .o(n_31953) );
in01s01 FE_RC_5273_0 ( .a(n_25598), .o(FE_RN_2328_0) );
no02s06 FE_RC_5274_0 ( .a(FE_RN_2328_0), .b(n_27098), .o(n_27183) );
in01f02 FE_RC_5275_0 ( .a(n_26401), .o(FE_RN_2329_0) );
in01f02 FE_RC_5276_0 ( .a(n_26390), .o(FE_RN_2330_0) );
ao22f02 FE_RC_5277_0 ( .a(n_26390), .b(FE_RN_2329_0), .c(FE_RN_2330_0), .d(n_26401), .o(n_26588) );
na02s01 FE_RC_5281_0 ( .a(n_30326), .b(n_30327), .o(FE_RN_2333_0) );
na02m08 FE_RC_5282_0 ( .a(FE_RN_2333_0), .b(n_31783), .o(n_31836) );
oa22m02 FE_RC_5283_0 ( .a(n_36787), .b(n_36789), .c(n_36788), .d(n_36798), .o(n_36866) );
in01m04 FE_RC_5284_0 ( .a(FE_RN_2334_0), .o(n_26586) );
na02f02 FE_RC_5285_0 ( .a(FE_OCP_DRV_N1488_n_24848), .b(n_26440), .o(FE_RN_2334_0) );
no02f04 FE_RC_5286_0 ( .a(n_26337), .b(n_26412), .o(FE_RN_2335_0) );
no02f08 FE_RC_5287_0 ( .a(FE_RN_2335_0), .b(n_26338), .o(n_26506) );
oa22m01 FE_RC_5288_0 ( .a(FE_OCPN5262_n_27536), .b(n_31239), .c(n_27366), .d(FE_OCP_RBN3272_n_31239), .o(n_31360) );
oa22f02 FE_RC_5289_0 ( .a(n_31081), .b(FE_OCPN5286_n_30708), .c(n_27131), .d(n_31026), .o(n_31099) );
oa22f04 FE_RC_5290_0 ( .a(n_27306), .b(n_27614), .c(n_27305), .d(n_27615), .o(n_27714) );
oa22m04 FE_RC_5291_0 ( .a(n_27267), .b(FE_OCP_RBN6255_FE_RN_1283_0), .c(n_27268), .d(FE_RN_1283_0), .o(n_27727) );
in01s01 FE_RC_5292_0 ( .a(n_27494), .o(FE_RN_2336_0) );
oa22f04 FE_RC_5294_0 ( .a(FE_RN_2336_0), .b(FE_OCP_RBN6256_FE_RN_2452_0), .c(FE_RN_2452_0), .d(n_27494), .o(n_27726) );
oa22s04 FE_RC_5296_0 ( .a(n_27399), .b(n_27681), .c(n_27398), .d(n_27682), .o(n_27772) );
oa22s02 FE_RC_5298_0 ( .a(n_27490), .b(n_27701), .c(n_27491), .d(n_27702), .o(n_27799) );
oa22f04 FE_RC_5299_0 ( .a(n_27493), .b(n_27723), .c(n_27492), .d(FE_OCP_RBN1876_n_27723), .o(n_27835) );
oa22s02 FE_RC_5302_0 ( .a(n_27484), .b(n_27688), .c(n_27485), .d(n_44360), .o(n_27781) );
ao22f04 FE_RC_5313_0 ( .a(n_19964), .b(n_19686), .c(n_19687), .d(n_19963), .o(n_20072) );
in01s02 FE_RC_5315_0 ( .a(n_17888), .o(FE_RN_2344_0) );
in01s02 FE_RC_5316_0 ( .a(n_17889), .o(FE_RN_2345_0) );
na02s02 TIMEBOOST_cell_5668 ( .a(n_17201), .b(n_17043), .o(TIMEBOOST_net_1782) );
no04f10 TIMEBOOST_cell_6417 ( .a(n_28029), .b(n_28028), .c(n_28117), .d(n_28118), .o(n_28248) );
in01s06 FE_RC_5319_0 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_3_), .o(FE_RN_2347_0) );
no02s04 TIMEBOOST_cell_6117 ( .a(TIMEBOOST_net_436), .b(n_19566), .o(TIMEBOOST_net_1910) );
na03m04 TIMEBOOST_cell_7359 ( .a(FE_OCP_RBN6133_n_11169), .b(n_11114), .c(n_11202), .o(n_11301) );
oa22m04 FE_RC_5323_0 ( .a(n_18262), .b(n_18412), .c(n_18261), .d(n_18438), .o(n_18600) );
oa22s01 FE_RC_5324_0 ( .a(n_1099), .b(n_44652), .c(n_1098), .d(n_44661), .o(n_1294) );
oa22f04 FE_RC_5325_0 ( .a(n_19419), .b(n_19421), .c(FE_OCPN1290_n_19384), .d(n_19423), .o(n_19555) );
oa22m02 FE_RC_5326_0 ( .a(FE_OCP_RBN5027_n_18515), .b(n_18433), .c(n_18468), .d(FE_OCP_RBN5028_n_18515), .o(n_18789) );
ao22s04 FE_RC_5327_0 ( .a(FE_RN_1123_0), .b(n_30601), .c(n_30369), .d(FE_RN_1124_0), .o(n_30733) );
oa22m04 FE_RC_5328_0 ( .a(n_20434), .b(n_20799), .c(n_20460), .d(n_20819), .o(n_20941) );
ao22f04 FE_RC_5329_0 ( .a(n_30997), .b(n_31161), .c(n_30998), .d(n_31160), .o(n_31304) );
oa22m04 FE_RC_5330_0 ( .a(n_27366), .b(n_30888), .c(FE_OCPN1763_n_30708), .d(n_30943), .o(n_30965) );
oa22m04 FE_RC_5332_0 ( .a(n_22459), .b(n_22612), .c(n_22500), .d(n_22598), .o(n_22774) );
in01s01 FE_RC_5335_0 ( .a(n_23848), .o(FE_RN_2350_0) );
in01s02 FE_RC_5336_0 ( .a(n_24251), .o(FE_RN_2351_0) );
no02s06 FE_RC_5337_0 ( .a(FE_RN_2350_0), .b(FE_RN_2351_0), .o(FE_RN_2352_0) );
no02s08 FE_RC_5338_0 ( .a(FE_RN_2352_0), .b(FE_RN_510_0), .o(n_24366) );
oa22m08 FE_RC_5339_0 ( .a(n_23880), .b(n_24489), .c(n_23879), .d(n_24490), .o(n_24612) );
ao22f04 FE_RC_5340_0 ( .a(n_22207), .b(n_24797), .c(n_24828), .d(n_24918), .o(n_24967) );
na02s02 TIMEBOOST_cell_2078 ( .a(TIMEBOOST_net_653), .b(n_42362), .o(n_42387) );
ao22m04 FE_RC_5342_0 ( .a(n_26785), .b(n_26747), .c(n_26758), .d(n_46934), .o(n_26844) );
oa22s06 FE_RC_5343_0 ( .a(n_27482), .b(n_27684), .c(n_27483), .d(n_27703), .o(n_27800) );
oa22s02 FE_RC_5344_0 ( .a(FE_OFN1183_n_24059), .b(FE_OCP_RBN6258_n_27743), .c(n_27796), .d(n_27743), .o(n_27815) );
no02s01 TIMEBOOST_cell_1621 ( .a(n_3135), .b(n_3026), .o(TIMEBOOST_net_425) );
ao22m04 FE_RC_5346_0 ( .a(n_12578), .b(FE_OCP_RBN5576_n_12727), .c(n_12577), .d(FE_OCP_RBN5574_n_12727), .o(n_12902) );
ao22f04 FE_RC_5347_0 ( .a(FE_OCP_RBN5019_n_13726), .b(n_13840), .c(n_13814), .d(FE_OCP_RBN6638_n_13726), .o(n_14004) );
ao22m08 FE_RC_5349_0 ( .a(FE_RN_1026_0), .b(FE_OCP_RBN2560_n_13084), .c(FE_RN_1027_0), .d(n_13711), .o(n_13732) );
oa22f10 FE_RC_5350_0 ( .a(n_27827), .b(n_27831), .c(FE_OCP_RBN5040_n_27827), .d(n_27832), .o(n_27939) );
ao22s06 FE_RC_5352_0 ( .a(n_44696), .b(n_44723), .c(n_44695), .d(FE_OCP_RBN7128_n_44722), .o(n_27888) );
oa22m08 FE_RC_5353_0 ( .a(n_11833), .b(n_11773), .c(n_11772), .d(n_11927), .o(n_12021) );
oa22m02 FE_RC_5356_0 ( .a(n_12574), .b(n_13059), .c(n_12575), .d(n_13060), .o(n_13232) );
ao22f02 FE_RC_5358_0 ( .a(FE_OCP_RBN5710_n_13984), .b(n_14287), .c(n_14336), .d(n_13984), .o(n_14519) );
in01s01 FE_RC_5359_0 ( .a(n_12935), .o(FE_RN_2353_0) );
na02m06 FE_RC_5361_0 ( .a(FE_RN_2353_0), .b(FE_OCP_RBN5664_n_13757), .o(FE_RN_2355_0) );
na02f08 FE_RC_5362_0 ( .a(FE_RN_2226_0), .b(FE_RN_2355_0), .o(n_13858) );
ao22f04 FE_RC_5363_0 ( .a(n_13630), .b(FE_OCP_RBN1593_n_13557), .c(FE_OCP_RBN1592_n_13557), .d(n_13629), .o(n_13722) );
oa22f04 FE_RC_5364_0 ( .a(FE_OCP_RBN2061_n_13813), .b(n_13659), .c(n_13673), .d(n_13813), .o(n_13890) );
oa22m06 FE_RC_5366_0 ( .a(FE_OCP_RBN2772_n_45521), .b(n_13514), .c(n_13515), .d(n_45521), .o(n_14539) );
oa22f02 FE_RC_5368_0 ( .a(n_14824), .b(FE_OCP_RBN5759_n_14444), .c(FE_OCP_RBN6702_n_14444), .d(n_14891), .o(n_14962) );
oa22f04 FE_RC_5369_0 ( .a(n_14755), .b(n_14803), .c(n_14802), .d(n_14773), .o(n_14911) );
oa22f04 FE_RC_5371_0 ( .a(n_15059), .b(n_14976), .c(n_14975), .d(n_15060), .o(n_15206) );
ao22m04 FE_RC_5372_0 ( .a(n_14618), .b(n_16088), .c(n_14588), .d(FE_OCP_RBN3178_n_16088), .o(FE_RN_1151_0) );
oa22m04 FE_RC_5373_0 ( .a(n_17320), .b(n_17522), .c(n_17319), .d(n_17566), .o(n_17697) );
oa22s03 FE_RC_5374_0 ( .a(n_17318), .b(n_17516), .c(n_17317), .d(n_17559), .o(n_17723) );
ao22m04 FE_RC_5376_0 ( .a(n_17268), .b(n_17446), .c(n_17452), .d(n_17269), .o(n_17587) );
oa22f04 FE_RC_5379_0 ( .a(n_14560), .b(n_14659), .c(n_14485), .d(n_14660), .o(n_14763) );
oa22f02 FE_RC_537_0 ( .a(n_16396), .b(n_16609), .c(n_16626), .d(n_16397), .o(n_16719) );
oa22f02 FE_RC_5380_0 ( .a(n_14889), .b(n_14852), .c(n_14874), .d(n_14890), .o(n_14991) );
oa22f08 FE_RC_5383_0 ( .a(FE_RN_444_0), .b(FE_RN_443_0), .c(FE_RN_445_0), .d(n_32638), .o(n_32653) );
ao22s06 FE_RC_5385_0 ( .a(FE_RN_1377_0), .b(FE_RN_1378_0), .c(FE_RN_1319_0), .d(n_12394), .o(n_12463) );
no02s02 TIMEBOOST_cell_1671 ( .a(n_3279), .b(n_3173), .o(TIMEBOOST_net_450) );
oa22f02 FE_RC_5389_0 ( .a(n_22709), .b(n_22801), .c(n_22793), .d(FE_OCP_RBN3456_n_22709), .o(n_22766) );
oa22s02 FE_RC_5390_0 ( .a(n_20231), .b(n_22897), .c(n_22793), .d(n_22856), .o(n_22957) );
oa22s02 FE_RC_5391_0 ( .a(n_22801), .b(n_22857), .c(n_22793), .d(n_22790), .o(n_22892) );
oa22s02 FE_RC_5392_0 ( .a(n_22961), .b(n_22902), .c(n_20252), .d(n_22862), .o(n_22962) );
ao22m04 FE_RC_5393_0 ( .a(n_31156), .b(FE_RN_538_0), .c(FE_RN_539_0), .d(n_31305), .o(n_31446) );
ao22m02 FE_RC_5396_0 ( .a(n_17213), .b(n_17275), .c(n_17214), .d(n_17287), .o(n_17475) );
no03s02 FE_RC_5397_0 ( .a(n_17036), .b(n_17137), .c(n_17027), .o(FE_RN_1545_0) );
oa22f04 FE_RC_5398_0 ( .a(FE_OCP_DRV_N3526_n_17031), .b(n_17513), .c(FE_OCP_DRV_N3528_n_17071), .d(n_17492), .o(n_17685) );
ao22f04 FE_RC_5400_0 ( .a(n_15377), .b(n_15660), .c(n_15629), .d(n_15376), .o(n_15817) );
in01s02 FE_RC_5402_0 ( .a(FE_OCP_DRV_N1410_n_12416), .o(FE_RN_2356_0) );
in01s01 FE_RC_5403_0 ( .a(n_12362), .o(FE_RN_2357_0) );
no02s01 TIMEBOOST_cell_1774 ( .a(TIMEBOOST_net_501), .b(n_21748), .o(n_21718) );
no02s10 TIMEBOOST_cell_1808 ( .a(FE_RN_329_0), .b(TIMEBOOST_net_518), .o(n_16086) );
oa22m02 FE_RC_5406_0 ( .a(FE_OFN1181_n_13195), .b(n_14114), .c(n_13515), .d(FE_OCP_RBN2741_n_14114), .o(n_14271) );
oa22f04 FE_RC_5407_0 ( .a(n_25633), .b(n_25355), .c(n_25356), .d(n_25602), .o(n_25729) );
in01s01 FE_RC_5408_0 ( .a(n_23995), .o(FE_RN_2359_0) );
in01s01 FE_RC_5409_0 ( .a(n_24645), .o(FE_RN_2360_0) );
na02s02 FE_RC_5410_0 ( .a(FE_RN_2359_0), .b(FE_RN_2360_0), .o(FE_RN_2361_0) );
na02s02 TIMEBOOST_cell_8128 ( .a(n_22288), .b(n_20859), .o(TIMEBOOST_net_2695) );
ao22f04 FE_RC_5413_0 ( .a(FE_OCP_RBN2652_n_29448), .b(n_29690), .c(n_30310), .d(n_29689), .o(n_29753) );
oa22s06 FE_RC_5414_0 ( .a(n_15671), .b(n_15818), .c(n_15672), .d(n_15819), .o(n_16011) );
oa22f04 FE_RC_5415_0 ( .a(FE_OCP_RBN3419_n_32130), .b(n_32346), .c(n_32130), .d(n_32330), .o(n_32471) );
oa22m08 FE_RC_5418_0 ( .a(n_11786), .b(n_11817), .c(n_11704), .d(n_11818), .o(n_12005) );
oa22f04 FE_RC_5419_0 ( .a(n_14412), .b(n_14244), .c(n_14285), .d(n_14413), .o(n_14554) );
in01f02 FE_RC_541_0 ( .a(n_16536), .o(FE_RN_153_0) );
na03m20 TIMEBOOST_cell_5692 ( .a(n_11774), .b(n_45622), .c(FE_OCP_RBN6318_n_45224), .o(n_11817) );
na02s06 TIMEBOOST_cell_4910 ( .a(n_47210), .b(n_6903), .o(TIMEBOOST_net_1403) );
na03s10 TIMEBOOST_cell_7112 ( .a(n_32598), .b(TIMEBOOST_net_588), .c(n_32641), .o(n_32699) );
no02m04 FE_RC_5428_0 ( .a(n_23371), .b(n_23361), .o(FE_RN_2367_0) );
na02f06 FE_RC_5429_0 ( .a(n_23456), .b(FE_RN_2367_0), .o(FE_RN_2368_0) );
in01f04 FE_RC_542_0 ( .a(n_16566), .o(FE_RN_154_0) );
na02f08 FE_RC_5430_0 ( .a(FE_RN_2368_0), .b(FE_RN_2366_0), .o(n_23579) );
na02f04 TIMEBOOST_cell_5109 ( .a(TIMEBOOST_net_1502), .b(n_8880), .o(FE_RN_2023_0) );
no02f06 TIMEBOOST_cell_5110 ( .a(FE_RN_762_0), .b(FE_RN_760_0), .o(TIMEBOOST_net_1503) );
na02s01 TIMEBOOST_cell_1409 ( .a(n_23838), .b(n_23722), .o(TIMEBOOST_net_319) );
in01s02 FE_RC_5440_0 ( .a(n_23481), .o(FE_RN_2376_0) );
no02s04 TIMEBOOST_cell_8594 ( .a(n_19725), .b(FE_OCP_RBN5681_n_19177), .o(TIMEBOOST_net_2784) );
na03s08 TIMEBOOST_cell_8180 ( .a(FE_RN_2173_0), .b(delay_xor_ln22_unr9_stage4_stallmux_q_7_), .c(n_45697), .o(FE_RN_2174_0) );
no03s08 TIMEBOOST_cell_8474 ( .a(FE_OCP_RBN2426_n_11907), .b(FE_RN_918_0), .c(FE_RN_1829_0), .o(TIMEBOOST_net_2724) );
in01m04 FE_RC_5444_0 ( .a(n_23481), .o(FE_RN_2380_0) );
no02m06 TIMEBOOST_cell_8864 ( .a(FE_OCP_RBN3396_n_11486), .b(n_11530), .o(TIMEBOOST_net_2919) );
na03m04 TIMEBOOST_cell_7268 ( .a(FE_OCP_RBN2951_n_3867), .b(FE_OCPN4828_FE_OCP_RBN4275_n_3700), .c(TIMEBOOST_net_1652), .o(n_4081) );
na02f04 TIMEBOOST_cell_8802 ( .a(FE_OCP_RBN3071_n_15433), .b(n_14452), .o(TIMEBOOST_net_2888) );
na02s01 TIMEBOOST_cell_1410 ( .a(TIMEBOOST_net_319), .b(n_24610), .o(n_24770) );
na02m02 FE_RC_5455_0 ( .a(n_18866), .b(FE_OFN737_n_17093), .o(FE_RN_2388_0) );
na02f04 FE_RC_5456_0 ( .a(n_18858), .b(FE_RN_2388_0), .o(n_18945) );
na02m04 FE_RC_5457_0 ( .a(n_24860), .b(n_24919), .o(FE_RN_2390_0) );
no02f06 FE_RC_5458_0 ( .a(n_24924), .b(FE_RN_2390_0), .o(FE_RN_2391_0) );
no02m08 FE_RC_5459_0 ( .a(n_24924), .b(n_24923), .o(FE_RN_2392_0) );
no03s08 TIMEBOOST_cell_6405 ( .a(FE_RN_1651_0), .b(FE_OCP_RBN6310_n_45224), .c(n_11737), .o(n_11991) );
oa22f08 FE_RC_5460_0 ( .a(FE_RN_2391_0), .b(n_24920), .c(FE_RN_2389_0), .d(FE_RN_2392_0), .o(n_25074) );
in01s01 FE_RC_5461_0 ( .a(n_24919), .o(FE_RN_2393_0) );
in01s01 FE_RC_5462_0 ( .a(FE_RN_2393_0), .o(FE_RN_2389_0) );
ao22f02 FE_RC_5463_0 ( .a(n_30140), .b(n_30388), .c(n_30139), .d(n_30379), .o(n_30451) );
in01s01 FE_RC_5465_0 ( .a(n_19170), .o(FE_RN_2394_0) );
in01m04 FE_RC_5466_0 ( .a(FE_RN_2395_0), .o(n_19323) );
no02m04 FE_RC_5467_0 ( .a(FE_RN_2394_0), .b(n_19206), .o(FE_RN_2395_0) );
na02s04 FE_RC_5468_0 ( .a(n_17900), .b(n_19206), .o(FE_RN_2396_0) );
na02m08 FE_RC_5469_0 ( .a(FE_RN_2396_0), .b(n_19323), .o(n_19380) );
no02s01 TIMEBOOST_cell_1959 ( .a(n_12086), .b(n_12079), .o(TIMEBOOST_net_594) );
no02s02 TIMEBOOST_cell_2910 ( .a(n_12975), .b(n_12947), .o(TIMEBOOST_net_746) );
no02s06 FE_RC_5472_0 ( .a(n_28649), .b(n_28705), .o(FE_RN_2398_0) );
na02f10 FE_RC_5473_0 ( .a(n_29218), .b(FE_RN_2398_0), .o(n_29232) );
in01s02 FE_RC_5474_0 ( .a(FE_RN_1420_0), .o(FE_RN_2399_0) );
na02m06 TIMEBOOST_cell_7003 ( .a(n_44492), .b(FE_OCP_RBN3212_n_10568), .o(TIMEBOOST_net_2260) );
in01s01 FE_RC_5477_0 ( .a(FE_RN_1384_0), .o(FE_RN_2401_0) );
in01f04 FE_RC_5478_0 ( .a(FE_RN_2402_0), .o(n_29585) );
no02f04 FE_RC_5479_0 ( .a(n_29518), .b(FE_RN_2401_0), .o(FE_RN_2402_0) );
in01s01 FE_RC_5481_0 ( .a(FE_OCP_RBN3707_n_18716), .o(FE_RN_2403_0) );
no02f06 FE_RC_5482_0 ( .a(n_20070), .b(FE_RN_2403_0), .o(n_20125) );
in01m06 FE_RC_5483_0 ( .a(n_45209), .o(FE_RN_2404_0) );
na02s20 FE_RC_5484_0 ( .a(n_45224), .b(FE_RN_2404_0), .o(n_11786) );
no02s01 FE_RC_5488_0 ( .a(n_23851), .b(n_23850), .o(FE_RN_2407_0) );
na02m08 FE_RC_5489_0 ( .a(FE_RN_2407_0), .b(n_24445), .o(n_24500) );
na03m10 TIMEBOOST_cell_7115 ( .a(FE_RN_1578_0), .b(n_32689), .c(n_32851), .o(n_32889) );
in01s02 FE_RC_5490_0 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_0_), .o(FE_RN_2408_0) );
na02s06 FE_RC_5491_0 ( .a(n_27888), .b(FE_RN_2408_0), .o(n_27910) );
in01s01 FE_RC_5494_0 ( .a(n_45008), .o(FE_RN_2410_0) );
in01f02 FE_RC_5495_0 ( .a(FE_RN_2411_0), .o(n_20760) );
na02f02 FE_RC_5496_0 ( .a(n_20542), .b(FE_RN_2410_0), .o(FE_RN_2411_0) );
in01f01 FE_RC_5497_0 ( .a(n_29566), .o(FE_RN_2412_0) );
no03f08 TIMEBOOST_cell_8232 ( .a(n_18285), .b(n_18263), .c(n_18300), .o(n_18343) );
na03m04 TIMEBOOST_cell_4742 ( .a(n_4920), .b(n_4741), .c(n_4856), .o(n_5101) );
no02s04 FE_RC_5500_0 ( .a(n_24624), .b(n_24518), .o(FE_RN_2414_0) );
no02m08 FE_RC_5501_0 ( .a(FE_RN_2414_0), .b(n_24778), .o(n_24800) );
in01s01 FE_RC_5505_0 ( .a(FE_RN_462_0), .o(FE_RN_2417_0) );
in01s02 FE_RC_5506_0 ( .a(FE_OCP_RBN1016_n_13601), .o(FE_RN_2418_0) );
na02s04 FE_RC_5507_0 ( .a(FE_RN_2417_0), .b(FE_RN_2418_0), .o(FE_RN_2419_0) );
na02m06 TIMEBOOST_cell_8511 ( .a(TIMEBOOST_net_2742), .b(n_13408), .o(n_13511) );
in01s01 FE_RC_5509_0 ( .a(n_13262), .o(FE_RN_2420_0) );
in01m04 FE_RC_5510_0 ( .a(FE_RN_2421_0), .o(n_14093) );
na02m04 FE_RC_5511_0 ( .a(FE_RN_2420_0), .b(n_13997), .o(FE_RN_2421_0) );
in01m04 FE_RC_5512_0 ( .a(FE_RN_2422_0), .o(FE_RN_1099_0) );
no02m04 FE_RC_5513_0 ( .a(n_47251), .b(n_29407), .o(FE_RN_2422_0) );
in01f04 FE_RC_5514_0 ( .a(FE_RN_2423_0), .o(n_26220) );
no02f03 FE_RC_5515_0 ( .a(n_26087), .b(FE_RN_1793_0), .o(FE_RN_2423_0) );
na02s01 FE_RC_5518_0 ( .a(n_31795), .b(n_30350), .o(FE_RN_2425_0) );
na02m08 FE_RC_5519_0 ( .a(n_31518), .b(FE_RN_2425_0), .o(n_31549) );
in01s01 FE_RC_5520_0 ( .a(FE_OCPN3531_n_26468), .o(FE_RN_2426_0) );
no02f04 FE_RC_5521_0 ( .a(n_26469), .b(FE_RN_2426_0), .o(n_26559) );
in01s01 FE_RC_5524_0 ( .a(FE_OCPN1291_n_29439), .o(FE_RN_2428_0) );
na02f06 FE_RC_5525_0 ( .a(n_29440), .b(FE_RN_2428_0), .o(n_29516) );
no02f06 FE_RC_5526_0 ( .a(n_31141), .b(n_31163), .o(FE_RN_2429_0) );
no02f08 FE_RC_5527_0 ( .a(FE_RN_2429_0), .b(n_31162), .o(n_31308) );
in01s06 FE_RC_5528_0 ( .a(FE_RN_2430_0), .o(n_27620) );
no02s06 FE_RC_5529_0 ( .a(n_27598), .b(n_27549), .o(FE_RN_2430_0) );
in01f06 FE_RC_5530_0 ( .a(FE_RN_2431_0), .o(n_30843) );
na02f06 FE_RC_5531_0 ( .a(n_30727), .b(FE_OCPN1676_n_27062), .o(FE_RN_2431_0) );
in01s01 FE_RC_5532_0 ( .a(n_46419), .o(FE_RN_2432_0) );
in01s01 FE_RC_5533_0 ( .a(n_15144), .o(FE_RN_2433_0) );
na02s02 FE_RC_5534_0 ( .a(FE_RN_2432_0), .b(FE_RN_2433_0), .o(FE_RN_2434_0) );
no02s10 TIMEBOOST_cell_1017 ( .a(FE_RN_2522_0), .b(n_28226), .o(TIMEBOOST_net_123) );
no03m04 TIMEBOOST_cell_2219 ( .a(FE_RN_2196_0), .b(n_32740), .c(n_32741), .o(FE_RN_2197_0) );
in01s02 FE_RC_5537_0 ( .a(n_15219), .o(FE_RN_2437_0) );
na02f02 TIMEBOOST_cell_4537 ( .a(n_11238), .b(n_11044), .o(TIMEBOOST_net_1359) );
no02f04 FE_RC_5539_0 ( .a(FE_RN_2438_0), .b(FE_OCP_RBN3099_n_15561), .o(FE_RN_2439_0) );
no02s10 TIMEBOOST_cell_1018 ( .a(TIMEBOOST_net_123), .b(FE_OCP_RBN5375_n_28123), .o(n_28271) );
no02s06 FE_RC_5541_0 ( .a(FE_OCP_RBN5329_n_15047), .b(n_14340), .o(FE_RN_2440_0) );
na02s06 FE_RC_5542_0 ( .a(n_14340), .b(FE_OCP_RBN5329_n_15047), .o(FE_RN_2441_0) );
ao12m08 FE_RC_5543_0 ( .a(FE_RN_2440_0), .b(FE_RN_2441_0), .c(n_15151), .o(n_15276) );
in01f02 FE_RC_5544_0 ( .a(FE_RN_2442_0), .o(n_15392) );
no02f02 FE_RC_5545_0 ( .a(FE_RN_1141_0), .b(FE_OCP_RBN2103_n_15286), .o(FE_RN_2442_0) );
in01s01 FE_RC_5546_0 ( .a(n_14452), .o(FE_RN_2443_0) );
in01m04 FE_RC_5547_0 ( .a(FE_RN_2444_0), .o(n_16233) );
na02m04 FE_RC_5548_0 ( .a(FE_RN_2443_0), .b(n_16095), .o(FE_RN_2444_0) );
in01s01 FE_RC_5549_0 ( .a(FE_OCP_RBN2087_n_14911), .o(FE_RN_2445_0) );
no02s04 FE_RC_5550_0 ( .a(FE_RN_2445_0), .b(n_16622), .o(n_16682) );
in01s02 FE_RC_5551_0 ( .a(n_16665), .o(FE_RN_2446_0) );
ao22m04 FE_RC_5552_0 ( .a(n_16716), .b(n_16665), .c(FE_RN_2446_0), .d(n_16735), .o(n_16791) );
no02s01 TIMEBOOST_cell_1545 ( .a(n_42443), .b(n_42444), .o(TIMEBOOST_net_387) );
na02m06 TIMEBOOST_cell_4268 ( .a(TIMEBOOST_net_1224), .b(n_8101), .o(FE_RN_188_0) );
ao22f04 FE_RC_5557_0 ( .a(n_23029), .b(FE_OCP_RBN2450_n_23246), .c(n_23030), .d(n_23246), .o(n_23347) );
na02s01 TIMEBOOST_cell_6387 ( .a(FE_OCPN945_n_27287), .b(FE_OCP_RBN3275_n_26464), .o(TIMEBOOST_net_2045) );
na04s08 TIMEBOOST_cell_8213 ( .a(n_22562), .b(FE_OCPN1049_n_23581), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_), .d(n_23574), .o(n_23680) );
in01s02 FE_RC_555_0 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_5_), .o(FE_RN_162_0) );
ao22f04 FE_RC_5560_0 ( .a(FE_OCP_RBN4144_n_7743), .b(n_8465), .c(FE_OCPN931_n_7817), .d(n_8498), .o(n_8608) );
ao22m04 FE_RC_5561_0 ( .a(n_13912), .b(n_14286), .c(FE_OCPN1250_n_13882), .d(n_14186), .o(n_14372) );
na02s02 TIMEBOOST_cell_7980 ( .a(n_5025), .b(n_4441), .o(TIMEBOOST_net_2621) );
ao22m08 FE_RC_5563_0 ( .a(FE_OCP_RBN2653_n_29448), .b(FE_OFN775_n_25834), .c(FE_RN_1384_0), .d(n_29448), .o(n_29545) );
in01s01 FE_RC_5564_0 ( .a(FE_RN_2448_0), .o(FE_RN_2449_0) );
in01s02 FE_RC_5565_0 ( .a(FE_RN_2449_0), .o(FE_OFN775_n_25834) );
oa22m04 FE_RC_5566_0 ( .a(n_18032), .b(FE_OCP_RBN1824_n_19434), .c(FE_OFN738_n_17093), .d(n_19434), .o(n_19561) );
oa22f04 FE_RC_5568_0 ( .a(FE_OCP_RBN1820_n_13858), .b(n_14034), .c(FE_OCP_RBN1819_n_13858), .d(n_14071), .o(n_14197) );
ao22m06 FE_RC_5569_0 ( .a(n_10468), .b(n_10731), .c(n_10467), .d(n_10764), .o(n_10878) );
in01s20 FE_RC_556_0 ( .a(n_36918), .o(FE_RN_163_0) );
oa22f02 FE_RC_5570_0 ( .a(n_29704), .b(n_29788), .c(n_29763), .d(n_29717), .o(n_29845) );
ao22f04 FE_RC_5571_0 ( .a(n_19889), .b(n_19998), .c(n_19997), .d(n_19863), .o(n_20070) );
no02s02 TIMEBOOST_cell_1889 ( .a(n_11087), .b(FE_OCP_RBN5955_FE_OFN4772_n_44463), .o(TIMEBOOST_net_559) );
oa22f02 FE_RC_5574_0 ( .a(n_23447), .b(n_26290), .c(FE_RN_1641_0), .d(n_26291), .o(n_26442) );
ao22f06 FE_RC_5575_0 ( .a(n_34335), .b(n_34829), .c(n_34334), .d(n_34793), .o(n_34934) );
oa22f06 FE_RC_5576_0 ( .a(n_16423), .b(n_16419), .c(FE_OCPN1324_n_14577), .d(n_16426), .o(n_16526) );
ao22m08 FE_RC_5578_0 ( .a(n_20784), .b(n_21165), .c(n_20785), .d(n_21196), .o(n_21358) );
no02s02 FE_RC_5579_0 ( .a(n_27568), .b(n_27277), .o(FE_RN_2450_0) );
no02s06 TIMEBOOST_cell_6019 ( .a(FE_OCP_RBN2483_FE_RN_657_0), .b(n_33019), .o(TIMEBOOST_net_1861) );
no02m06 FE_RC_5582_0 ( .a(FE_RN_2450_0), .b(FE_OCP_RBN6242_n_27436), .o(FE_RN_2452_0) );
oa22f04 FE_RC_5583_0 ( .a(n_21645), .b(n_21927), .c(n_21678), .d(n_21895), .o(n_21983) );
oa22m02 FE_RC_5584_0 ( .a(n_36739), .b(n_36760), .c(n_36740), .d(n_36759), .o(n_36792) );
oa22s04 FE_RC_5585_0 ( .a(n_31796), .b(n_32243), .c(n_31797), .d(n_32225), .o(n_32339) );
oa22f10 FE_RC_5587_0 ( .a(n_32575), .b(n_32523), .c(n_32601), .d(FE_OCP_RBN4919_n_32575), .o(n_32655) );
na02m08 TIMEBOOST_cell_4911 ( .a(TIMEBOOST_net_1403), .b(n_7000), .o(n_7060) );
na02s01 TIMEBOOST_cell_1581 ( .a(n_25169), .b(n_24999), .o(TIMEBOOST_net_405) );
na02s01 TIMEBOOST_cell_6109 ( .a(n_42392), .b(n_42125), .o(TIMEBOOST_net_1906) );
no02m08 TIMEBOOST_cell_4945 ( .a(TIMEBOOST_net_1420), .b(n_28231), .o(n_28306) );
na02s02 TIMEBOOST_cell_5265 ( .a(TIMEBOOST_net_1580), .b(n_24653), .o(n_24766) );
no02f04 TIMEBOOST_cell_1608 ( .a(TIMEBOOST_net_418), .b(n_38863), .o(n_39086) );
oa22m08 FE_RC_5595_0 ( .a(n_22992), .b(n_22985), .c(n_22993), .d(n_23040), .o(n_23136) );
na03s03 TIMEBOOST_cell_8275 ( .a(FE_OCP_RBN5723_n_47022), .b(n_2913), .c(n_3132), .o(n_3214) );
oa22s04 FE_RC_5597_0 ( .a(n_7597), .b(FE_OCP_RBN2817_n_8939), .c(n_7596), .d(n_8939), .o(n_9082) );
ao22f08 FE_RC_5598_0 ( .a(n_28083), .b(FE_OCP_RBN5376_n_28123), .c(n_28084), .d(n_28123), .o(n_28207) );
ao22m08 FE_RC_5599_0 ( .a(FE_OCP_RBN6162_FE_RN_1136_0), .b(n_11370), .c(FE_OCP_RBN3377_n_44342), .d(n_11371), .o(n_11475) );
ao22m06 FE_RC_5600_0 ( .a(n_34005), .b(n_34084), .c(FE_OCP_RBN5627_n_33976), .d(n_34083), .o(n_34183) );
ao22f04 FE_RC_5601_0 ( .a(n_25623), .b(n_26000), .c(n_25622), .d(n_26022), .o(n_26152) );
ao22f06 FE_RC_5602_0 ( .a(n_25594), .b(n_25940), .c(n_25593), .d(n_25918), .o(n_26020) );
ao22f04 FE_RC_5604_0 ( .a(FE_OCPN904_n_21955), .b(n_21924), .c(FE_OCPN906_n_21956), .d(n_21923), .o(n_22005) );
ao22f06 FE_RC_5605_0 ( .a(n_16291), .b(n_16324), .c(n_16325), .d(n_16287), .o(n_16474) );
oa22m04 FE_RC_5607_0 ( .a(n_17457), .b(n_17381), .c(n_17380), .d(n_17495), .o(n_17630) );
ao22s02 FE_RC_5608_0 ( .a(n_22462), .b(n_44364), .c(n_22464), .d(n_22705), .o(n_22790) );
oa22f04 FE_RC_5609_0 ( .a(n_19033), .b(n_19518), .c(n_20307), .d(n_19475), .o(n_19666) );
oa22f02 FE_RC_5610_0 ( .a(n_38654), .b(n_38778), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .d(n_38628), .o(n_38673) );
oa22m04 FE_RC_5611_0 ( .a(FE_OCP_RBN2460_n_12365), .b(n_12110), .c(n_12111), .d(n_12365), .o(n_12453) );
oa22s06 FE_RC_5613_0 ( .a(n_17869), .b(n_17907), .c(n_17868), .d(n_17908), .o(n_18038) );
ao22m06 FE_RC_5614_0 ( .a(FE_RN_2453_0), .b(n_36501), .c(n_36197), .d(FE_OCP_RBN6150_n_36501), .o(n_36559) );
in01s01 FE_RC_5615_0 ( .a(n_36196), .o(FE_RN_2454_0) );
in01s02 FE_RC_5616_0 ( .a(FE_RN_2454_0), .o(FE_RN_2453_0) );
no02m04 TIMEBOOST_cell_1675 ( .a(n_26037), .b(n_23353), .o(TIMEBOOST_net_452) );
oa22m08 FE_RC_5618_0 ( .a(FE_OCP_RBN7017_n_32687), .b(n_32647), .c(FE_OCP_RBN7016_n_32687), .d(FE_OCP_RBN1803_n_32647), .o(n_32770) );
oa22m04 FE_RC_5619_0 ( .a(n_20499), .b(n_20620), .c(n_20465), .d(n_20653), .o(n_20804) );
na02f08 TIMEBOOST_cell_2957 ( .a(TIMEBOOST_net_769), .b(n_2240), .o(n_2318) );
in01s01 FE_RC_5621_0 ( .a(n_20703), .o(FE_RN_2456_0) );
in01s01 FE_RC_5622_0 ( .a(FE_RN_2456_0), .o(FE_RN_2455_0) );
oa22s02 FE_RC_5624_0 ( .a(n_27481), .b(n_27692), .c(n_27480), .d(n_27717), .o(n_27805) );
oa22s02 FE_RC_5625_0 ( .a(n_27523), .b(n_27695), .c(n_27524), .d(n_27673), .o(n_27783) );
oa22f02 FE_RC_5628_0 ( .a(n_30706), .b(n_30658), .c(n_30657), .d(FE_OCP_RBN6032_n_30706), .o(n_30860) );
na02s04 TIMEBOOST_cell_1688 ( .a(TIMEBOOST_net_458), .b(n_20024), .o(FE_RN_532_0) );
no02s02 TIMEBOOST_cell_2916 ( .a(n_18932), .b(n_18882), .o(TIMEBOOST_net_749) );
oa22m06 FE_RC_5631_0 ( .a(n_36301), .b(n_36560), .c(n_36302), .d(n_36546), .o(n_36669) );
oa22f02 FE_RC_5632_0 ( .a(FE_OCPN1394_n_22801), .b(n_22596), .c(n_22580), .d(n_22570), .o(n_22629) );
oa22s02 FE_RC_5634_0 ( .a(n_27487), .b(n_27610), .c(n_27486), .d(n_27624), .o(n_27720) );
no02m10 TIMEBOOST_cell_2967 ( .a(n_41294), .b(TIMEBOOST_net_774), .o(n_41327) );
oa22s01 FE_RC_5640_0 ( .a(n_17336), .b(n_17782), .c(n_16339), .d(n_17756), .o(n_17829) );
no02s06 TIMEBOOST_cell_6749 ( .a(n_24601), .b(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(TIMEBOOST_net_2132) );
no02s08 TIMEBOOST_cell_6750 ( .a(TIMEBOOST_net_2132), .b(n_24602), .o(n_24788) );
no02m08 FE_RC_5643_0 ( .a(n_32684), .b(n_32810), .o(FE_RN_2458_0) );
na02m08 FE_RC_5644_0 ( .a(n_32684), .b(n_32810), .o(FE_RN_2459_0) );
ao12m08 FE_RC_5645_0 ( .a(FE_RN_2458_0), .b(FE_RN_2459_0), .c(n_32770), .o(n_32848) );
no02f08 FE_RC_5646_0 ( .a(n_28098), .b(n_27865), .o(FE_RN_2460_0) );
na02f08 FE_RC_5647_0 ( .a(n_28098), .b(n_27865), .o(FE_RN_2461_0) );
ao12f08 FE_RC_5648_0 ( .a(FE_RN_2460_0), .b(FE_RN_2461_0), .c(n_28009), .o(n_28120) );
na02f08 FE_RC_5649_0 ( .a(n_28234), .b(n_28182), .o(FE_RN_2462_0) );
na02f08 FE_RC_5650_0 ( .a(FE_RN_2462_0), .b(n_28183), .o(n_28322) );
in01s06 FE_RC_5651_0 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_5_), .o(FE_RN_2463_0) );
in01s02 FE_RC_5652_0 ( .a(n_23137), .o(FE_RN_2464_0) );
no02m02 TIMEBOOST_cell_2928 ( .a(n_29193), .b(n_28767), .o(TIMEBOOST_net_755) );
in01f04 FE_RC_5654_0 ( .a(n_23197), .o(FE_RN_2466_0) );
no02s04 TIMEBOOST_cell_1719 ( .a(n_20336), .b(n_45066), .o(TIMEBOOST_net_474) );
na02f06 FE_RC_5656_0 ( .a(n_23270), .b(FE_RN_2467_0), .o(FE_RN_1656_0) );
na02s01 FE_RC_5657_0 ( .a(FE_OCPN5228_n_33917), .b(n_33820), .o(FE_RN_2468_0) );
no02s02 FE_RC_5658_0 ( .a(n_33917), .b(n_33820), .o(FE_RN_2469_0) );
oa12m04 FE_RC_5659_0 ( .a(FE_RN_2468_0), .b(FE_RN_2469_0), .c(n_33868), .o(n_33940) );
in01f02 FE_RC_5660_0 ( .a(FE_RN_2470_0), .o(n_19348) );
no02s01 TIMEBOOST_cell_1997 ( .a(n_37875), .b(n_37910), .o(TIMEBOOST_net_613) );
in01s01 FE_RC_5663_0 ( .a(FE_OCPN5277_n_13329), .o(FE_RN_2471_0) );
no02m08 FE_RC_5664_0 ( .a(FE_RN_2471_0), .b(n_14585), .o(n_14611) );
in01s02 FE_RC_5666_0 ( .a(n_20477), .o(FE_RN_2472_0) );
no02f04 TIMEBOOST_cell_2134 ( .a(TIMEBOOST_net_681), .b(n_5858), .o(n_5955) );
in01s02 FE_RC_5674_0 ( .a(n_20828), .o(FE_RN_2477_0) );
in01f02 FE_RC_5675_0 ( .a(FE_RN_2478_0), .o(n_20944) );
na02m02 FE_RC_5676_0 ( .a(FE_RN_2477_0), .b(n_20825), .o(FE_RN_2478_0) );
in01s01 FE_RC_5677_0 ( .a(n_14588), .o(FE_RN_2479_0) );
in01f02 FE_RC_5678_0 ( .a(FE_RN_2480_0), .o(n_16206) );
no02m02 FE_RC_5679_0 ( .a(FE_RN_2479_0), .b(n_16095), .o(FE_RN_2480_0) );
no02s02 TIMEBOOST_cell_6962 ( .a(TIMEBOOST_net_2239), .b(n_3299), .o(TIMEBOOST_net_1904) );
na02s02 TIMEBOOST_cell_3110 ( .a(FE_RN_899_0), .b(FE_RN_897_0), .o(TIMEBOOST_net_846) );
in01s02 FE_RC_5687_0 ( .a(n_44040), .o(FE_RN_2485_0) );
na02s02 TIMEBOOST_cell_8848 ( .a(n_16453), .b(n_16454), .o(TIMEBOOST_net_2911) );
no02s01 TIMEBOOST_cell_5442 ( .a(n_4875), .b(FE_OCPN3584_n_4556), .o(TIMEBOOST_net_1669) );
no02s02 FE_RC_5690_0 ( .a(n_30592), .b(n_30593), .o(FE_RN_2487_0) );
in01s06 FE_RC_5691_0 ( .a(n_31819), .o(FE_RN_2488_0) );
no02s10 FE_RC_5692_0 ( .a(FE_RN_2488_0), .b(FE_RN_2487_0), .o(FE_RN_2489_0) );
no02f20 FE_RC_5693_0 ( .a(n_32081), .b(FE_RN_2489_0), .o(n_32142) );
na02s01 FE_RC_5694_0 ( .a(FE_OCP_RBN2106_n_30619), .b(n_30729), .o(FE_RN_2490_0) );
in01s01 FE_RC_5695_0 ( .a(n_31518), .o(FE_RN_2491_0) );
na02s06 FE_RC_5696_0 ( .a(FE_RN_2490_0), .b(FE_RN_2491_0), .o(FE_RN_2492_0) );
na02s10 FE_RC_5697_0 ( .a(n_31685), .b(FE_RN_2492_0), .o(FE_RN_2493_0) );
no02m20 FE_RC_5698_0 ( .a(FE_RN_2493_0), .b(n_32000), .o(n_32088) );
no02s02 FE_RC_5699_0 ( .a(n_22591), .b(FE_RN_625_0), .o(FE_RN_2494_0) );
oa22f08 FE_RC_569_0 ( .a(n_45511), .b(n_40631), .c(n_40601), .d(FE_OCP_RBN2410_n_40631), .o(n_40663) );
no02s06 FE_RC_5700_0 ( .a(FE_RN_2494_0), .b(FE_RN_622_0), .o(FE_RN_627_0) );
oa22m02 FE_RC_5701_0 ( .a(n_18259), .b(FE_OCP_RBN5325_n_18653), .c(n_18260), .d(n_18653), .o(n_18866) );
na03m06 TIMEBOOST_cell_7200 ( .a(n_14437), .b(n_14399), .c(n_14461), .o(n_14590) );
oa22f06 FE_RC_5704_0 ( .a(n_36194), .b(n_36535), .c(n_36195), .d(n_44168), .o(n_36632) );
oa22s04 FE_RC_5705_0 ( .a(n_31858), .b(n_32224), .c(n_31859), .d(n_32242), .o(n_32338) );
ao22m10 FE_RC_5707_0 ( .a(FE_OCP_RBN2392_n_16970), .b(n_16972), .c(n_16970), .d(FE_OCP_RBN5018_n_16972), .o(n_17230) );
ao22f04 FE_RC_5709_0 ( .a(n_13418), .b(n_14252), .c(FE_OFN4795_n_13195), .d(n_14273), .o(n_14468) );
oa22f04 FE_RC_5710_0 ( .a(FE_OCP_RBN2089_n_14964), .b(n_14907), .c(n_14924), .d(n_14964), .o(n_15083) );
ao22f04 FE_RC_5711_0 ( .a(n_21289), .b(FE_RN_1529_0), .c(n_21363), .d(FE_RN_1530_0), .o(n_21503) );
na03m08 FE_RC_5712_0 ( .a(n_22185), .b(FE_RN_1541_0), .c(FE_OCP_RBN5049_FE_RN_606_0), .o(FE_RN_1542_0) );
ao22m10 FE_RC_5714_0 ( .a(n_17129), .b(FE_RN_485_0), .c(FE_RN_486_0), .d(n_16984), .o(n_17243) );
oa22m08 FE_RC_5715_0 ( .a(n_11734), .b(n_11788), .c(FE_OCP_RBN3702_n_11788), .d(n_11735), .o(n_11941) );
ao22f10 FE_RC_5716_0 ( .a(n_27970), .b(FE_OCP_RBN1805_n_27934), .c(n_27912), .d(n_27934), .o(n_28085) );
in01f01 FE_RC_5717_0 ( .a(n_18343), .o(FE_RN_2495_0) );
in01s02 FE_RC_5718_0 ( .a(n_18319), .o(FE_RN_2496_0) );
na02m04 FE_RC_5719_0 ( .a(FE_RN_2495_0), .b(FE_RN_2496_0), .o(FE_RN_2497_0) );
no02f04 FE_RC_5720_0 ( .a(FE_RN_2497_0), .b(FE_OCP_RBN7023_n_18650), .o(n_18760) );
ao22m02 FE_RC_5721_0 ( .a(n_12888), .b(FE_OCP_RBN2044_n_12907), .c(n_12907), .d(n_12889), .o(n_13096) );
oa22f04 FE_RC_5722_0 ( .a(n_33060), .b(n_33492), .c(n_33059), .d(n_45627), .o(n_33567) );
oa22f04 FE_RC_5723_0 ( .a(n_28604), .b(FE_OCP_RBN1808_n_28968), .c(n_28603), .d(n_28968), .o(n_29056) );
oa22m02 FE_RC_5724_0 ( .a(n_13010), .b(n_13144), .c(n_13146), .d(FE_RN_1744_0), .o(n_13225) );
oa22m04 FE_RC_5725_0 ( .a(n_25738), .b(n_29163), .c(FE_OFN773_n_25834), .d(FE_OCP_RBN2566_n_29163), .o(n_29271) );
oa22f02 FE_RC_5726_0 ( .a(n_18950), .b(n_18826), .c(n_18949), .d(n_18859), .o(n_19011) );
oa22f02 FE_RC_5727_0 ( .a(n_19170), .b(n_19241), .c(FE_OCP_RBN3713_n_19241), .d(n_18010), .o(n_19377) );
oa22s04 FE_RC_5729_0 ( .a(FE_OCP_RBN6651_n_13818), .b(n_15156), .c(FE_OCPN1077_n_13831), .d(n_15194), .o(n_15266) );
in01s01 FE_RC_572_0 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_3_), .o(FE_RN_168_0) );
ao22f04 FE_RC_5730_0 ( .a(n_35135), .b(n_35289), .c(n_35288), .d(n_35137), .o(n_35383) );
ao22f04 FE_RC_5731_0 ( .a(n_30466), .b(FE_OCP_RBN1847_n_30428), .c(n_27014), .d(n_30428), .o(n_30500) );
ao22m04 FE_RC_5732_0 ( .a(n_30276), .b(n_30736), .c(n_30275), .d(n_30735), .o(n_30849) );
oa22m04 FE_RC_5733_0 ( .a(n_45091), .b(n_21003), .c(n_45024), .d(n_21004), .o(n_21157) );
oa22m02 FE_RC_5734_0 ( .a(n_45010), .b(n_20984), .c(n_45070), .d(n_20985), .o(n_21127) );
oa22m04 FE_RC_5735_0 ( .a(n_30930), .b(FE_RN_2069_0), .c(n_31048), .d(FE_RN_2070_0), .o(n_31198) );
ao22f04 FE_RC_5738_0 ( .a(n_21709), .b(n_21745), .c(n_21685), .d(n_21768), .o(n_21874) );
oa22m04 FE_RC_5739_0 ( .a(n_21726), .b(n_21945), .c(n_21701), .d(n_21944), .o(n_22037) );
in01s02 FE_RC_573_0 ( .a(n_22738), .o(FE_RN_169_0) );
oa22f06 FE_RC_5740_0 ( .a(n_36005), .b(n_36492), .c(n_36004), .d(n_36493), .o(n_36569) );
oa22s06 FE_RC_5741_0 ( .a(n_36094), .b(n_36506), .c(n_36093), .d(n_36507), .o(n_36594) );
oa22s01 FE_RC_5742_0 ( .a(n_17584), .b(n_17811), .c(n_16339), .d(n_17781), .o(n_17855) );
in01s40 FE_RC_5743_0 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_3_), .o(FE_RN_2498_0) );
na02s40 FE_RC_5744_0 ( .a(FE_OCP_RBN7106_n_44365), .b(FE_RN_2498_0), .o(n_17040) );
in01s03 FE_RC_5745_0 ( .a(n_45209), .o(FE_RN_2499_0) );
no02m08 TIMEBOOST_cell_5021 ( .a(n_24081), .b(TIMEBOOST_net_1458), .o(n_24157) );
na02s01 TIMEBOOST_cell_5022 ( .a(n_37929), .b(n_37969), .o(TIMEBOOST_net_1459) );
in01s20 FE_RC_5748_0 ( .a(FE_RN_1364_0), .o(FE_RN_2501_0) );
no02m40 FE_RC_5749_0 ( .a(FE_RN_2501_0), .b(n_22990), .o(n_23040) );
no02s06 FE_RC_574_0 ( .a(FE_RN_169_0), .b(FE_RN_168_0), .o(FE_RN_170_0) );
in01s01 FE_RC_5750_0 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_), .o(FE_RN_2502_0) );
na02m03 FE_RC_5751_0 ( .a(n_6517), .b(FE_RN_2502_0), .o(FE_RN_2503_0) );
na02f10 FE_RC_5752_0 ( .a(n_6966), .b(FE_RN_2503_0), .o(n_6762) );
ao22s10 FE_RC_5753_0 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_5_), .b(FE_OCP_RBN6466_n_44061), .c(FE_OCP_RBN2272_delay_xor_ln22_unr15_stage6_stallmux_q_5_), .d(FE_OCP_RBN5507_n_44061), .o(n_22937) );
oa22f08 FE_RC_5754_0 ( .a(n_32582), .b(n_32520), .c(n_32522), .d(n_32521), .o(n_32638) );
in01s01 FE_RC_5756_0 ( .a(n_11882), .o(FE_RN_2504_0) );
na02s02 FE_RC_5757_0 ( .a(n_11907), .b(FE_RN_2504_0), .o(n_11908) );
in01m10 FE_RC_5758_0 ( .a(n_36878), .o(FE_RN_2505_0) );
na02m10 FE_RC_5759_0 ( .a(n_36921), .b(FE_RN_2505_0), .o(FE_RN_2506_0) );
no02s06 FE_RC_575_0 ( .a(n_22855), .b(FE_RN_170_0), .o(n_22983) );
na02m10 FE_RC_5760_0 ( .a(FE_RN_2506_0), .b(n_36897), .o(n_37058) );
no02s06 FE_RC_5763_0 ( .a(n_6698), .b(n_6896), .o(FE_RN_2508_0) );
na02s06 FE_RC_5764_0 ( .a(n_6698), .b(n_6896), .o(FE_RN_2509_0) );
ao12s06 FE_RC_5765_0 ( .a(FE_RN_2508_0), .b(FE_RN_2509_0), .c(n_6835), .o(n_6945) );
in01s02 FE_RC_5769_0 ( .a(FE_RN_2512_0), .o(n_6891) );
in01m08 FE_RC_576_0 ( .a(n_37032), .o(FE_RN_171_0) );
no02s02 FE_RC_5770_0 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_3_), .b(n_6804), .o(FE_RN_2512_0) );
no02s01 TIMEBOOST_cell_3920 ( .a(TIMEBOOST_net_1050), .b(n_38112), .o(n_38183) );
in01f10 FE_RC_5772_0 ( .a(n_27999), .o(FE_RN_2514_0) );
in01m10 FE_RC_5773_0 ( .a(FE_RN_2515_0), .o(n_28028) );
na02s01 TIMEBOOST_cell_6108 ( .a(TIMEBOOST_net_1905), .b(n_42201), .o(n_42341) );
no02m06 FE_RC_5775_0 ( .a(n_11767), .b(n_11994), .o(FE_RN_2516_0) );
ao12m06 FE_RC_5776_0 ( .a(FE_RN_2516_0), .b(FE_RN_2517_0), .c(n_11994), .o(n_12195) );
in01s02 FE_RC_5777_0 ( .a(n_11767), .o(FE_RN_2518_0) );
in01s02 FE_RC_5778_0 ( .a(FE_RN_2518_0), .o(FE_RN_2517_0) );
no02m08 FE_RC_5779_0 ( .a(n_12176), .b(n_12069), .o(FE_RN_2519_0) );
in01m08 FE_RC_577_0 ( .a(n_37031), .o(FE_RN_172_0) );
no02m08 FE_RC_5780_0 ( .a(FE_RN_2519_0), .b(n_12097), .o(n_12292) );
in01s06 FE_RC_5781_0 ( .a(n_28058), .o(FE_RN_2520_0) );
in01s10 FE_RC_5782_0 ( .a(n_28219), .o(FE_RN_2521_0) );
na02s10 FE_RC_5783_0 ( .a(FE_RN_2521_0), .b(FE_RN_2520_0), .o(FE_RN_2522_0) );
na03m04 TIMEBOOST_cell_8181 ( .a(n_28399), .b(FE_RN_731_0), .c(FE_RN_732_0), .o(FE_RN_734_0) );
in01f04 FE_RC_5785_0 ( .a(FE_RN_2523_0), .o(n_28182) );
no02f06 FE_RC_5786_0 ( .a(n_28086), .b(delay_add_ln22_unr17_stage7_stallmux_q_4_), .o(FE_RN_2523_0) );
in01s01 FE_RC_5787_0 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_6_), .o(FE_RN_2524_0) );
na02s02 FE_RC_5788_0 ( .a(FE_RN_2524_0), .b(n_6990), .o(n_7063) );
no02f08 FE_RC_578_0 ( .a(FE_RN_172_0), .b(FE_RN_171_0), .o(FE_RN_173_0) );
in01s02 FE_RC_5791_0 ( .a(FE_RN_2527_0), .o(FE_RN_2526_0) );
na02f08 FE_RC_5792_0 ( .a(n_7031), .b(FE_RN_2526_0), .o(n_7083) );
in01s01 FE_RC_5793_0 ( .a(n_6683), .o(FE_RN_2528_0) );
in01s01 FE_RC_5794_0 ( .a(FE_RN_2528_0), .o(FE_RN_2527_0) );
in01s06 FE_RC_5795_0 ( .a(FE_RN_969_0), .o(FE_RN_2529_0) );
in01s06 FE_RC_5796_0 ( .a(n_17579), .o(FE_RN_2530_0) );
na02s06 TIMEBOOST_cell_8543 ( .a(TIMEBOOST_net_2758), .b(n_34320), .o(n_34433) );
no03f08 TIMEBOOST_cell_2364 ( .a(n_41374), .b(n_41322), .c(n_41370), .o(n_41405) );
in01s02 FE_RC_5799_0 ( .a(FE_RN_2532_0), .o(n_12424) );
ao22s04 FE_RC_57_0 ( .a(FE_OCP_RBN5653_n_2438), .b(n_3080), .c(FE_OCP_RBN5663_n_2438), .d(n_3597), .o(n_3116) );
no02s02 FE_RC_5800_0 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_9_), .b(n_12342), .o(FE_RN_2532_0) );
in01s01 FE_RC_5803_0 ( .a(n_6767), .o(FE_RN_2535_0) );
no02s02 FE_RC_5804_0 ( .a(FE_RN_2535_0), .b(n_6836), .o(FE_RN_2536_0) );
in01s01 FE_RC_5805_0 ( .a(n_6737), .o(FE_RN_2537_0) );
no03s04 TIMEBOOST_cell_8238 ( .a(n_37795), .b(n_37823), .c(TIMEBOOST_net_298), .o(n_37861) );
in01s01 FE_RC_5807_0 ( .a(FE_RN_2534_0), .o(FE_RN_2539_0) );
no02m04 TIMEBOOST_cell_1702 ( .a(TIMEBOOST_net_465), .b(n_3821), .o(n_5629) );
in01s01 FE_RC_5809_0 ( .a(n_6717), .o(FE_RN_2541_0) );
no02m02 TIMEBOOST_cell_1704 ( .a(TIMEBOOST_net_466), .b(n_3722), .o(n_4041) );
no03f04 TIMEBOOST_cell_2433 ( .a(FE_OCP_RBN1816_n_33873), .b(FE_OCP_RBN1814_n_33846), .c(n_33901), .o(n_34010) );
na02m04 TIMEBOOST_cell_8642 ( .a(FE_RN_1933_0), .b(FE_RN_1934_0), .o(TIMEBOOST_net_2808) );
in01s02 FE_RC_5813_0 ( .a(n_6676), .o(FE_RN_2544_0) );
in01s02 FE_RC_5814_0 ( .a(FE_RN_2544_0), .o(FE_RN_2534_0) );
in01s01 FE_RC_5818_0 ( .a(n_1722), .o(FE_RN_2548_0) );
in01s01 FE_RC_5819_0 ( .a(FE_RN_2548_0), .o(FE_RN_2546_0) );
no02s01 TIMEBOOST_cell_6587 ( .a(n_28176), .b(n_28175), .o(TIMEBOOST_net_2051) );
no02m04 TIMEBOOST_cell_6056 ( .a(TIMEBOOST_net_1879), .b(n_2266), .o(n_2332) );
in01s01 FE_RC_5822_0 ( .a(n_1387), .o(FE_RN_2550_0) );
in01s01 FE_RC_5823_0 ( .a(n_1480), .o(FE_RN_2551_0) );
no02s01 FE_RC_5824_0 ( .a(FE_RN_2551_0), .b(FE_RN_2550_0), .o(FE_RN_2552_0) );
in01s01 FE_RC_5825_0 ( .a(FE_RN_2554_0), .o(FE_RN_2553_0) );
na02s01 FE_RC_5826_0 ( .a(FE_RN_2552_0), .b(FE_RN_2553_0), .o(FE_RN_2555_0) );
in01s01 FE_RC_5827_0 ( .a(n_1780), .o(FE_RN_2556_0) );
in01s01 FE_RC_5828_0 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_28_), .o(FE_RN_2557_0) );
na02s01 TIMEBOOST_cell_2818 ( .a(n_46107), .b(n_32422), .o(TIMEBOOST_net_700) );
no02s01 TIMEBOOST_cell_5562 ( .a(n_22134), .b(n_44277), .o(TIMEBOOST_net_1729) );
na02s02 FE_RC_5831_0 ( .a(n_1840), .b(FE_RN_2559_0), .o(FE_RN_2560_0) );
na02s06 TIMEBOOST_cell_8542 ( .a(FE_RN_2734_0), .b(n_34297), .o(TIMEBOOST_net_2758) );
na02s20 TIMEBOOST_cell_7426 ( .a(FE_OCPN1649_n_44734), .b(delay_xor_ln22_unr18_stage7_stallmux_q_6_), .o(TIMEBOOST_net_2344) );
in01s01 FE_RC_5834_0 ( .a(n_1431), .o(FE_RN_2562_0) );
in01s01 FE_RC_5835_0 ( .a(FE_RN_2562_0), .o(FE_RN_2554_0) );
in01s01 FE_RC_5836_0 ( .a(n_32957), .o(FE_RN_2563_0) );
na02m10 FE_RC_5837_0 ( .a(n_33411), .b(FE_RN_2563_0), .o(n_33475) );
in01s01 FE_RC_5838_0 ( .a(n_33231), .o(FE_RN_2564_0) );
na02m08 FE_RC_5839_0 ( .a(n_33674), .b(FE_RN_2564_0), .o(n_33707) );
na02m10 FE_RC_583_0 ( .a(FE_OCP_RBN6518_n_32706), .b(FE_OCP_RBN5517_n_32436), .o(FE_RN_176_0) );
ao22f01 FE_RC_5840_0 ( .a(n_18198), .b(n_18360), .c(n_18199), .d(n_18318), .o(n_18515) );
no02m06 TIMEBOOST_cell_6677 ( .a(n_24746), .b(n_24546), .o(TIMEBOOST_net_2096) );
in01s01 FE_RC_5843_0 ( .a(n_7092), .o(FE_RN_2567_0) );
in01s01 FE_RC_5844_0 ( .a(FE_RN_2567_0), .o(FE_RN_2566_0) );
in01s01 FE_RC_5845_0 ( .a(n_12865), .o(FE_RN_2568_0) );
ao22m02 FE_RC_5846_0 ( .a(n_12800), .b(n_12865), .c(FE_RN_2568_0), .d(FE_OCP_RBN2510_n_12800), .o(n_12949) );
na02m08 TIMEBOOST_cell_6694 ( .a(TIMEBOOST_net_2104), .b(n_34514), .o(n_34591) );
no03s02 TIMEBOOST_cell_5811 ( .a(TIMEBOOST_net_1599), .b(n_20151), .c(TIMEBOOST_net_1112), .o(n_20245) );
in01s02 FE_RC_5849_0 ( .a(FE_RN_2569_0), .o(FE_RN_2571_0) );
in01s04 FE_RC_5850_0 ( .a(FE_RN_2571_0), .o(n_7702) );
in01f02 FE_RC_5854_0 ( .a(n_29141), .o(FE_RN_2574_0) );
oa22f04 FE_RC_5855_0 ( .a(FE_RN_2574_0), .b(n_29057), .c(n_29141), .d(n_29058), .o(n_29299) );
in01s01 FE_RC_5856_0 ( .a(FE_OCPN1307_n_23677), .o(FE_RN_2575_0) );
no02m08 FE_RC_5857_0 ( .a(FE_RN_2575_0), .b(n_24200), .o(n_24248) );
in01s01 FE_RC_5858_0 ( .a(n_28764), .o(FE_RN_2576_0) );
na02m06 FE_RC_5859_0 ( .a(FE_RN_2576_0), .b(n_29273), .o(FE_RN_2577_0) );
in01s01 FE_RC_5860_0 ( .a(n_28764), .o(FE_RN_2578_0) );
oa12f06 FE_RC_5861_0 ( .a(FE_RN_2577_0), .b(FE_RN_2578_0), .c(n_29273), .o(n_29378) );
no02s01 FE_RC_5862_0 ( .a(FE_RN_1842_0), .b(n_18594), .o(FE_RN_2579_0) );
na02m08 FE_RC_5863_0 ( .a(FE_RN_2579_0), .b(n_19080), .o(n_19105) );
in01m02 FE_RC_5864_0 ( .a(n_19135), .o(FE_RN_2580_0) );
ao22m02 FE_RC_5865_0 ( .a(n_19135), .b(FE_OCP_RBN5035_n_19055), .c(FE_RN_2580_0), .d(FE_OCP_RBN5377_n_19055), .o(n_19315) );
in01s01 FE_RC_5866_0 ( .a(FE_OCP_DRV_N1441_n_17836), .o(FE_RN_2581_0) );
no02f02 FE_RC_5867_0 ( .a(n_19243), .b(FE_RN_2581_0), .o(FE_RN_2470_0) );
in01s01 FE_RC_5868_0 ( .a(FE_OCPN5281_n_24425), .o(FE_RN_2582_0) );
no02f04 FE_RC_5869_0 ( .a(n_24426), .b(FE_RN_2582_0), .o(n_24494) );
ao22m06 FE_RC_5870_0 ( .a(n_25859), .b(FE_OCP_RBN2651_n_29470), .c(n_29630), .d(n_29470), .o(n_29594) );
in01m02 FE_RC_5871_0 ( .a(n_13529), .o(FE_RN_2583_0) );
oa22m02 FE_RC_5872_0 ( .a(n_13497), .b(n_13529), .c(FE_RN_2583_0), .d(n_13562), .o(n_13647) );
in01f02 FE_RC_5873_0 ( .a(n_19110), .o(FE_RN_2584_0) );
na02m08 TIMEBOOST_cell_4987 ( .a(TIMEBOOST_net_1441), .b(n_12450), .o(FE_RN_405_0) );
na02f02 TIMEBOOST_cell_6692 ( .a(TIMEBOOST_net_2103), .b(n_14201), .o(n_14334) );
na02s01 FE_RC_5876_0 ( .a(n_13190), .b(n_13101), .o(FE_RN_2586_0) );
no02f04 FE_RC_5877_0 ( .a(FE_RN_2586_0), .b(n_14100), .o(n_14123) );
no02s01 FE_RC_5878_0 ( .a(n_2660), .b(n_2661), .o(FE_RN_2587_0) );
na02s01 FE_RC_5879_0 ( .a(n_2712), .b(FE_RN_2587_0), .o(FE_RN_2588_0) );
no02f08 FE_RC_5880_0 ( .a(n_3212), .b(FE_RN_2588_0), .o(n_3227) );
ao22f04 FE_RC_5881_0 ( .a(n_38183), .b(n_38499), .c(n_38184), .d(n_38500), .o(n_38569) );
in01s01 FE_RC_5882_0 ( .a(n_2720), .o(FE_RN_2589_0) );
no03s20 TIMEBOOST_cell_2184 ( .a(n_27864), .b(n_27918), .c(n_27919), .o(n_28012) );
na02f08 FE_RC_5884_0 ( .a(n_3227), .b(FE_RN_2590_0), .o(n_3291) );
na02f06 FE_RC_5885_0 ( .a(n_19774), .b(n_19704), .o(FE_RN_2591_0) );
no02f08 FE_RC_5886_0 ( .a(FE_RN_2591_0), .b(n_19736), .o(n_19924) );
in01s02 FE_RC_5887_0 ( .a(n_19799), .o(FE_RN_2592_0) );
no02m02 TIMEBOOST_cell_5211 ( .a(TIMEBOOST_net_1553), .b(n_34788), .o(TIMEBOOST_net_853) );
no02f04 FE_RC_5890_0 ( .a(n_19799), .b(FE_OCP_RBN6374_n_19722), .o(FE_RN_2595_0) );
no03s02 TIMEBOOST_cell_5212 ( .a(n_3138), .b(n_3170), .c(TIMEBOOST_net_1092), .o(TIMEBOOST_net_1554) );
na03s08 FE_RC_5892_0 ( .a(n_34460), .b(n_34401), .c(n_34398), .o(FE_RN_2596_0) );
no02f10 FE_RC_5893_0 ( .a(n_34820), .b(FE_RN_2596_0), .o(n_34767) );
no02s06 FE_RC_5894_0 ( .a(n_34490), .b(n_34514), .o(FE_RN_2597_0) );
in01s01 FE_RC_5895_0 ( .a(n_34406), .o(FE_RN_2598_0) );
na02m08 FE_RC_5896_0 ( .a(n_34767), .b(FE_RN_2598_0), .o(FE_RN_2599_0) );
na02m10 FE_RC_5897_0 ( .a(FE_RN_2599_0), .b(FE_RN_2597_0), .o(n_34873) );
in01f02 FE_RC_5898_0 ( .a(FE_RN_2600_0), .o(n_8800) );
na02f02 FE_RC_5899_0 ( .a(n_8739), .b(n_8678), .o(FE_RN_2600_0) );
oa22f02 FE_RC_58_0 ( .a(n_18457), .b(n_19041), .c(n_18456), .d(n_19059), .o(n_19219) );
in01s01 FE_RC_5900_0 ( .a(FE_OCPN3529_n_28829), .o(FE_RN_2601_0) );
na02s02 FE_RC_5901_0 ( .a(FE_RN_2601_0), .b(n_29831), .o(n_29864) );
in01s01 FE_RC_5904_0 ( .a(n_29031), .o(FE_RN_2603_0) );
na02s10 FE_RC_5905_0 ( .a(n_29922), .b(FE_RN_2603_0), .o(n_30021) );
in01s01 FE_RC_5907_0 ( .a(FE_OCP_RBN4081_n_18899), .o(FE_RN_2604_0) );
na02m08 FE_RC_5908_0 ( .a(FE_RN_2604_0), .b(n_20228), .o(n_20285) );
in01f02 FE_RC_5909_0 ( .a(FE_RN_2605_0), .o(n_25175) );
in01s01 FE_RC_590_0 ( .a(n_17581), .o(FE_RN_177_0) );
na02f02 FE_RC_5910_0 ( .a(n_23892), .b(n_25114), .o(FE_RN_2605_0) );
in01m02 FE_RC_5911_0 ( .a(n_45520), .o(FE_RN_2606_0) );
na02f04 FE_RC_5912_0 ( .a(FE_RN_2606_0), .b(FE_OCP_RBN5776_n_13796), .o(FE_RN_2607_0) );
na02f06 FE_RC_5913_0 ( .a(n_14801), .b(FE_RN_2607_0), .o(n_14856) );
in01s01 FE_RC_5914_0 ( .a(FE_OCP_RBN5622_n_18986), .o(FE_RN_2608_0) );
no02m06 FE_RC_5915_0 ( .a(FE_RN_2608_0), .b(n_20249), .o(n_20309) );
in01s02 FE_RC_5916_0 ( .a(n_35059), .o(FE_RN_2609_0) );
in01m08 FE_RC_5917_0 ( .a(FE_RN_2610_0), .o(n_35123) );
no02m08 FE_RC_5918_0 ( .a(n_35012), .b(FE_RN_2609_0), .o(FE_RN_2610_0) );
in01s01 FE_RC_5919_0 ( .a(n_38859), .o(FE_RN_2611_0) );
in01m02 FE_RC_5920_0 ( .a(FE_RN_2612_0), .o(n_38885) );
na02s02 FE_RC_5921_0 ( .a(FE_RN_2611_0), .b(FE_OCP_RBN6758_n_38806), .o(FE_RN_2612_0) );
in01s01 FE_RC_5922_0 ( .a(FE_OCP_RBN1134_n_19077), .o(FE_RN_2613_0) );
na02m02 FE_RC_5923_0 ( .a(FE_RN_2613_0), .b(n_20372), .o(FE_RN_442_0) );
no02s03 FE_RC_5924_0 ( .a(FE_OCP_RBN6764_FE_RN_2259_0), .b(n_25295), .o(FE_RN_2614_0) );
na02f06 FE_RC_5925_0 ( .a(n_25654), .b(FE_RN_2614_0), .o(n_25676) );
ao22f04 FE_RC_5926_0 ( .a(n_9550), .b(n_9583), .c(n_9551), .d(n_9626), .o(n_9819) );
in01s01 FE_RC_5927_0 ( .a(FE_OCP_DRV_N4505_n_13476), .o(FE_RN_2615_0) );
no02f02 FE_RC_5928_0 ( .a(n_15001), .b(FE_RN_2615_0), .o(n_15137) );
in01s01 FE_RC_5929_0 ( .a(n_45008), .o(FE_RN_2616_0) );
na02s06 FE_RC_592_0 ( .a(FE_RN_177_0), .b(FE_OCP_RBN6370_n_17582), .o(FE_RN_179_0) );
no02f04 FE_RC_5930_0 ( .a(n_20549), .b(FE_RN_2616_0), .o(FE_RN_578_0) );
in01s01 FE_RC_5931_0 ( .a(n_20345), .o(FE_RN_2618_0) );
in01s01 FE_RC_5932_0 ( .a(n_20914), .o(FE_RN_2619_0) );
no02s02 FE_RC_5933_0 ( .a(FE_RN_2617_0), .b(n_20914), .o(FE_RN_2620_0) );
oa22f06 FE_RC_5934_0 ( .a(FE_RN_2619_0), .b(FE_RN_2618_0), .c(FE_RN_2620_0), .d(n_20820), .o(n_20849) );
in01s01 FE_RC_5935_0 ( .a(n_20345), .o(FE_RN_2621_0) );
in01s01 FE_RC_5936_0 ( .a(FE_RN_2621_0), .o(FE_RN_2617_0) );
in01s01 FE_RC_5937_0 ( .a(FE_OCPN1690_n_10105), .o(FE_RN_2622_0) );
no02s03 FE_RC_5938_0 ( .a(FE_RN_2622_0), .b(n_10106), .o(n_10197) );
na02s06 FE_RC_5939_0 ( .a(n_39012), .b(n_39013), .o(FE_RN_2623_0) );
na02s02 TIMEBOOST_cell_3917 ( .a(n_7749), .b(n_7366), .o(TIMEBOOST_net_1049) );
no02s08 FE_RC_5940_0 ( .a(n_39081), .b(FE_RN_2623_0), .o(FE_RN_2624_0) );
na02f10 FE_RC_5941_0 ( .a(n_39220), .b(FE_RN_2624_0), .o(n_39293) );
in01m02 FE_RC_5942_0 ( .a(n_35399), .o(FE_RN_2625_0) );
in01s02 FE_RC_5943_0 ( .a(n_35303), .o(FE_RN_2626_0) );
ao22m04 FE_RC_5944_0 ( .a(FE_RN_2625_0), .b(n_35303), .c(FE_RN_2626_0), .d(n_35399), .o(n_35483) );
ao22m02 FE_RC_5945_0 ( .a(n_10060), .b(FE_OCP_RBN3069_n_9910), .c(n_9910), .d(n_10019), .o(n_10225) );
in01s01 FE_RC_5946_0 ( .a(n_30220), .o(FE_RN_2627_0) );
na02s01 FE_RC_5947_0 ( .a(FE_OCPN6269_n_30599), .b(FE_RN_2627_0), .o(FE_RN_2628_0) );
oa12s01 FE_RC_5948_0 ( .a(FE_RN_2628_0), .b(FE_OCPN6269_n_30599), .c(n_30221), .o(n_30697) );
in01s01 FE_RC_5949_0 ( .a(FE_RN_1313_0), .o(FE_RN_2629_0) );
na02s01 FE_RC_5950_0 ( .a(n_30220), .b(FE_RN_2629_0), .o(FE_RN_2630_0) );
oa12s01 FE_RC_5951_0 ( .a(FE_RN_2630_0), .b(n_30220), .c(FE_OCPN1402_FE_OFN1196_n_27014), .o(FE_RN_2631_0) );
na02s02 FE_RC_5952_0 ( .a(n_30599), .b(FE_RN_2631_0), .o(FE_RN_2632_0) );
no02s01 FE_RC_5953_0 ( .a(n_30221), .b(FE_OCPN1402_FE_OFN1196_n_27014), .o(FE_RN_2633_0) );
in01s01 FE_RC_5954_0 ( .a(FE_RN_1313_0), .o(FE_RN_2634_0) );
ao12s02 FE_RC_5955_0 ( .a(FE_RN_2633_0), .b(n_30221), .c(FE_RN_2634_0), .o(FE_RN_2635_0) );
in01s01 FE_RC_5957_0 ( .a(n_45069), .o(FE_RN_2636_0) );
no02f02 FE_RC_5958_0 ( .a(FE_RN_2636_0), .b(n_20771), .o(FE_RN_1500_0) );
in01s01 FE_RC_5959_0 ( .a(FE_RN_2638_0), .o(FE_RN_2637_0) );
na02m03 FE_RC_5960_0 ( .a(n_10194), .b(FE_RN_2637_0), .o(n_47263) );
in01s01 FE_RC_5961_0 ( .a(FE_OCP_RBN2812_n_8835), .o(FE_RN_2639_0) );
in01s01 FE_RC_5962_0 ( .a(FE_RN_2639_0), .o(FE_RN_2638_0) );
in01s01 FE_RC_5963_0 ( .a(FE_OCPN5265_n_20852), .o(FE_RN_2640_0) );
na02f04 FE_RC_5964_0 ( .a(n_20853), .b(FE_RN_2640_0), .o(n_20883) );
in01s01 FE_RC_5965_0 ( .a(FE_OCPN1639_n_35367), .o(FE_RN_2641_0) );
na02f06 FE_RC_5966_0 ( .a(n_35368), .b(FE_RN_2641_0), .o(n_35410) );
in01s01 FE_RC_5967_0 ( .a(n_45010), .o(FE_RN_2642_0) );
no02m02 FE_RC_5968_0 ( .a(FE_RN_2642_0), .b(n_20951), .o(FE_RN_1697_0) );
in01s01 FE_RC_5969_0 ( .a(FE_OCPN5231_n_35594), .o(FE_RN_2643_0) );
na02m04 FE_RC_5970_0 ( .a(FE_RN_2643_0), .b(n_35595), .o(n_35650) );
in01s01 FE_RC_5971_0 ( .a(n_39189), .o(FE_RN_2644_0) );
na02f04 FE_RC_5972_0 ( .a(n_39450), .b(FE_RN_2644_0), .o(FE_RN_2645_0) );
in01s01 FE_RC_5973_0 ( .a(n_39189), .o(FE_RN_2646_0) );
oa12f04 FE_RC_5974_0 ( .a(FE_RN_2645_0), .b(FE_RN_2646_0), .c(n_39450), .o(n_39523) );
in01s01 FE_RC_5977_0 ( .a(FE_OCPN5223_n_10357), .o(FE_RN_2648_0) );
na02s06 FE_RC_5978_0 ( .a(n_10672), .b(FE_RN_2648_0), .o(n_10732) );
in01f02 FE_RC_5979_0 ( .a(n_15531), .o(FE_RN_2649_0) );
no04f08 TIMEBOOST_cell_7139 ( .a(n_23441), .b(n_23426), .c(n_23142), .d(n_23143), .o(n_23555) );
in01s01 TIMEBOOST_cell_7389 ( .a(TIMEBOOST_net_2324), .o(TIMEBOOST_net_2325) );
ao22f06 FE_RC_5983_0 ( .a(n_15371), .b(n_15805), .c(n_15372), .d(n_15852), .o(n_16041) );
na02s01 FE_RC_5984_0 ( .a(n_9148), .b(FE_OCPN1092_n_9014), .o(FE_RN_2652_0) );
na02s01 FE_RC_5985_0 ( .a(FE_OCP_RBN4356_n_10100), .b(FE_RN_2652_0), .o(FE_RN_2653_0) );
na02s06 FE_RC_5986_0 ( .a(n_10711), .b(FE_RN_2653_0), .o(n_10760) );
in01s01 FE_RC_5987_0 ( .a(n_45024), .o(FE_RN_2654_0) );
in01m02 FE_RC_5988_0 ( .a(FE_RN_2655_0), .o(n_21287) );
no02m02 FE_RC_5989_0 ( .a(FE_RN_2654_0), .b(n_21127), .o(FE_RN_2655_0) );
no02s02 TIMEBOOST_cell_1622 ( .a(TIMEBOOST_net_425), .b(n_3177), .o(n_4953) );
in01m02 FE_RC_5990_0 ( .a(n_30956), .o(FE_RN_2656_0) );
in01m02 FE_RC_5991_0 ( .a(n_30926), .o(FE_RN_2657_0) );
ao22m04 FE_RC_5992_0 ( .a(FE_RN_2656_0), .b(n_30926), .c(FE_RN_2657_0), .d(n_30956), .o(n_31126) );
no02s02 FE_RC_5993_0 ( .a(n_4998), .b(n_5021), .o(FE_RN_2658_0) );
na02m02 FE_RC_5994_0 ( .a(FE_RN_2658_0), .b(n_5272), .o(n_5348) );
in01s01 FE_RC_5995_0 ( .a(FE_OCP_DRV_N6897_FE_OCPN1679_n_27315), .o(FE_RN_2659_0) );
no02s04 FE_RC_5997_0 ( .a(FE_RN_2659_0), .b(n_31101), .o(FE_RN_2660_0) );
no02s01 FE_RC_5998_0 ( .a(FE_OCPUNCON1759_n_35644), .b(FE_RN_2661_0), .o(FE_RN_2662_0) );
no02s06 FE_RC_5999_0 ( .a(FE_RN_2662_0), .b(n_44222), .o(n_35693) );
in01s01 FE_RC_6000_0 ( .a(n_34707), .o(FE_RN_2663_0) );
in01s01 FE_RC_6001_0 ( .a(FE_RN_2663_0), .o(FE_RN_2661_0) );
in01s02 FE_RC_6002_0 ( .a(n_35831), .o(FE_RN_2664_0) );
in01s06 FE_RC_6003_0 ( .a(FE_RN_2665_0), .o(n_35869) );
no03m08 FE_RC_6004_0 ( .a(n_35696), .b(n_35752), .c(FE_RN_2664_0), .o(FE_RN_2665_0) );
ao22f02 FE_RC_6005_0 ( .a(n_26137), .b(FE_OCP_RBN6089_n_26304), .c(n_26304), .d(n_26138), .o(n_26440) );
no02s02 TIMEBOOST_cell_5131 ( .a(TIMEBOOST_net_1513), .b(n_34565), .o(n_34622) );
no02f04 TIMEBOOST_cell_8775 ( .a(TIMEBOOST_net_2874), .b(n_14956), .o(n_15009) );
no02f08 FE_RC_6008_0 ( .a(FE_RN_2668_0), .b(n_35872), .o(FE_RN_2669_0) );
no02s06 FE_RC_6009_0 ( .a(n_35755), .b(n_35754), .o(FE_RN_2670_0) );
no02f06 TIMEBOOST_cell_1676 ( .a(TIMEBOOST_net_452), .b(n_26121), .o(n_26302) );
no02m02 TIMEBOOST_cell_1351 ( .a(n_13453), .b(FE_OCP_RBN2540_n_12880), .o(TIMEBOOST_net_290) );
in01s01 TIMEBOOST_cell_8887 ( .a(TIMEBOOST_net_2930), .o(TIMEBOOST_net_2931) );
in01s01 FE_RC_6012_0 ( .a(n_35667), .o(FE_RN_2672_0) );
in01s02 FE_RC_6013_0 ( .a(FE_RN_2672_0), .o(FE_RN_2666_0) );
in01m04 FE_RC_6014_0 ( .a(FE_RN_2673_0), .o(n_26766) );
na02s02 FE_RC_6015_0 ( .a(n_26522), .b(n_25013), .o(FE_RN_2673_0) );
in01s01 FE_RC_6016_0 ( .a(n_21505), .o(FE_RN_2674_0) );
na02s04 FE_RC_6017_0 ( .a(n_21506), .b(FE_RN_2674_0), .o(FE_OCPN903_n_21955) );
na02s01 TIMEBOOST_cell_1145 ( .a(n_37541), .b(n_37540), .o(TIMEBOOST_net_187) );
no02f04 TIMEBOOST_cell_2069 ( .a(n_42051), .b(n_42196), .o(TIMEBOOST_net_649) );
oa22f04 FE_RC_601_0 ( .a(n_37461), .b(n_37141), .c(n_37140), .d(n_37462), .o(n_37581) );
na02s01 TIMEBOOST_cell_1146 ( .a(TIMEBOOST_net_187), .b(n_37475), .o(n_37543) );
no02m04 FE_RC_6021_0 ( .a(n_31465), .b(FE_RN_2675_0), .o(n_31584) );
no02s06 FE_RC_6022_0 ( .a(n_35911), .b(n_35910), .o(FE_RN_2676_0) );
na02f10 FE_RC_6023_0 ( .a(n_36376), .b(FE_RN_2676_0), .o(n_36410) );
na03m20 FE_RC_6027_0 ( .a(n_39866), .b(n_39924), .c(n_39925), .o(FE_RN_2679_0) );
no02f08 FE_RC_6028_0 ( .a(FE_RN_2679_0), .b(n_40050), .o(n_40124) );
no02s01 FE_RC_6029_0 ( .a(FE_OCP_RBN6038_n_30733), .b(FE_OCP_RBN6055_n_46957), .o(FE_RN_2680_0) );
ao22f04 FE_RC_602_0 ( .a(n_37181), .b(FE_OCP_RBN2463_n_37449), .c(n_37180), .d(n_37449), .o(n_37535) );
no02s03 FE_RC_6030_0 ( .a(FE_OCP_RBN4472_n_31819), .b(FE_RN_2680_0), .o(n_47273) );
in01s01 FE_RC_6031_0 ( .a(FE_OCPN1435_n_21278), .o(FE_RN_2681_0) );
na02s02 FE_RC_6032_0 ( .a(FE_RN_2681_0), .b(n_22249), .o(n_22330) );
in01s01 FE_RC_6033_0 ( .a(n_25595), .o(FE_RN_2682_0) );
na02s06 FE_RC_6034_0 ( .a(FE_RN_2682_0), .b(n_27103), .o(n_27157) );
na02s03 FE_RC_6035_0 ( .a(n_17595), .b(n_17190), .o(FE_RN_2683_0) );
na02m03 FE_RC_6036_0 ( .a(FE_RN_2683_0), .b(n_17445), .o(n_17689) );
na02s04 TIMEBOOST_cell_8707 ( .a(TIMEBOOST_net_2840), .b(FE_OCP_RBN2443_n_44798), .o(FE_RN_904_0) );
no02f10 TIMEBOOST_cell_1446 ( .a(TIMEBOOST_net_337), .b(FE_OCP_RBN7030_n_44259), .o(n_33833) );
na02s06 FE_RC_6039_0 ( .a(FE_RN_2685_0), .b(n_27274), .o(FE_RN_2686_0) );
na02s06 FE_RC_6040_0 ( .a(n_27554), .b(n_27189), .o(FE_RN_2687_0) );
no02s10 FE_RC_6041_0 ( .a(FE_RN_2687_0), .b(FE_RN_2686_0), .o(n_27593) );
na02s06 FE_RC_6042_0 ( .a(n_40037), .b(n_40074), .o(FE_RN_2688_0) );
no02f10 FE_RC_6043_0 ( .a(FE_RN_2688_0), .b(n_40466), .o(n_40472) );
oa22s02 FE_RC_6044_0 ( .a(n_22377), .b(n_22687), .c(n_22378), .d(n_22721), .o(n_22875) );
in01f02 FE_RC_6045_0 ( .a(n_32471), .o(FE_RN_2689_0) );
oa22f01 FE_RC_6046_0 ( .a(n_28336), .b(FE_RN_2689_0), .c(n_32566), .d(n_32471), .o(n_32545) );
oa22m06 FE_RC_6048_0 ( .a(n_22339), .b(n_22722), .c(FE_OCPN5306_n_22338), .d(n_22756), .o(n_22914) );
oa22m04 FE_RC_6049_0 ( .a(n_17321), .b(n_17514), .c(n_17322), .d(n_17493), .o(n_17686) );
in01f08 FE_RC_6050_0 ( .a(n_32279), .o(FE_OCP_RBN5218_n_32279) );
in01s01 FE_RC_6055_0 ( .a(n_17688), .o(FE_RN_2693_0) );
oa22s01 FE_RC_6056_0 ( .a(n_17584), .b(n_17688), .c(FE_RN_2693_0), .d(n_16339), .o(n_17750) );
in01m02 FE_RC_6057_0 ( .a(n_17591), .o(FE_RN_2694_0) );
oa22f02 FE_RC_6058_0 ( .a(FE_OCP_RBN3199_n_15599), .b(n_17591), .c(FE_RN_2694_0), .d(n_17753), .o(n_17647) );
in01s02 FE_RC_6059_0 ( .a(n_32326), .o(FE_RN_2695_0) );
no02s01 TIMEBOOST_cell_1411 ( .a(n_24182), .b(n_23769), .o(TIMEBOOST_net_320) );
in01s01 FE_RC_6061_0 ( .a(FE_RN_375_0), .o(FE_RN_2697_0) );
no02s04 TIMEBOOST_cell_1412 ( .a(TIMEBOOST_net_320), .b(n_24183), .o(n_24251) );
in01s02 FE_RC_6063_0 ( .a(n_32120), .o(FE_RN_2699_0) );
no02m08 FE_RC_6064_0 ( .a(FE_OCP_RBN5218_n_32279), .b(n_32326), .o(FE_RN_2700_0) );
no02m08 FE_RC_6065_0 ( .a(FE_RN_2700_0), .b(n_32020), .o(FE_RN_2701_0) );
in01s01 FE_RC_6067_0 ( .a(n_12212), .o(FE_RN_2702_0) );
oa22s02 FE_RC_6068_0 ( .a(FE_OFN787_n_46285), .b(n_12212), .c(FE_RN_2702_0), .d(FE_OFN765_n_46337), .o(n_46345) );
oa22f04 FE_RC_6069_0 ( .a(n_12705), .b(FE_OCP_RBN1589_n_13460), .c(n_12684), .d(n_13460), .o(n_13557) );
ao22m06 FE_RC_6070_0 ( .a(FE_OCP_RBN5510_FE_RN_1997_0), .b(n_11814), .c(FE_OCP_RBN5509_FE_RN_1997_0), .d(n_11813), .o(n_12036) );
oa22f04 FE_RC_6071_0 ( .a(FE_OCP_RBN5326_n_29292), .b(n_29258), .c(n_29292), .d(FE_RN_2051_0), .o(n_29392) );
ao22f04 FE_RC_6072_0 ( .a(n_30869), .b(FE_OCP_RBN7053_n_30867), .c(n_30867), .d(n_30870), .o(n_30978) );
ao22s02 FE_RC_6073_0 ( .a(n_20704), .b(n_21178), .c(FE_RN_2455_0), .d(n_21177), .o(n_21346) );
in01s02 FE_RC_6074_0 ( .a(n_31234), .o(FE_RN_2703_0) );
in01s02 FE_RC_6075_0 ( .a(n_31463), .o(FE_RN_2704_0) );
na02f06 TIMEBOOST_cell_5537 ( .a(TIMEBOOST_net_1716), .b(n_36550), .o(n_36626) );
no02s01 TIMEBOOST_cell_5538 ( .a(n_43388), .b(FE_OCP_RBN3308_n_43022), .o(TIMEBOOST_net_1717) );
oa22f08 FE_RC_6078_0 ( .a(FE_RN_495_0), .b(FE_RN_496_0), .c(FE_RN_497_0), .d(n_27104), .o(n_27244) );
oa22m04 FE_RC_6079_0 ( .a(n_22270), .b(n_22639), .c(n_22307), .d(FE_OCP_RBN6231_n_22639), .o(n_22829) );
no03f06 FE_RC_6080_0 ( .a(n_16171), .b(n_16236), .c(n_16166), .o(n_16237) );
ao22m10 FE_RC_6082_0 ( .a(FE_OCP_RBN3815_n_45209), .b(FE_OCP_RBN6319_n_45224), .c(n_45209), .d(n_45224), .o(n_11760) );
in01m80 FE_RC_6083_0 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_3_), .o(FE_RN_2706_0) );
na02m80 FE_RC_6084_0 ( .a(FE_RN_2706_0), .b(n_44962), .o(n_32433) );
ao22s06 FE_RC_6086_0 ( .a(FE_OCP_RBN7117_delay_xor_ln22_unr12_stage5_stallmux_q_0_), .b(FE_OCP_RBN7111_n_44365), .c(delay_xor_ln22_unr12_stage5_stallmux_q_0_), .d(FE_OCP_RBN7106_n_44365), .o(n_16799) );
na02m08 FE_RC_6087_0 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_1_), .b(FE_OCP_RBN6307_n_45224), .o(FE_RN_2708_0) );
na02m08 FE_RC_6088_0 ( .a(n_11762), .b(FE_RN_2708_0), .o(n_11813) );
in01s06 FE_RC_6089_0 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_0_), .o(FE_RN_2709_0) );
na02f04 TIMEBOOST_cell_1705 ( .a(FE_OCP_RBN2837_n_13962), .b(n_15353), .o(TIMEBOOST_net_467) );
na02s10 FE_RC_6090_0 ( .a(FE_RN_2709_0), .b(n_16829), .o(n_16857) );
oa22m08 FE_RC_6091_0 ( .a(n_22769), .b(n_22672), .c(n_22575), .d(n_22673), .o(n_22827) );
na02s02 TIMEBOOST_cell_4065 ( .a(n_44579), .b(n_9157), .o(TIMEBOOST_net_1123) );
in01m01 FE_RC_6093_0 ( .a(n_17084), .o(FE_RN_2710_0) );
no02s10 FE_RC_6094_0 ( .a(n_17192), .b(n_17133), .o(FE_RN_2711_0) );
na02s10 FE_RC_6095_0 ( .a(FE_RN_2711_0), .b(FE_RN_2710_0), .o(n_17442) );
oa22m10 FE_RC_6096_0 ( .a(n_32659), .b(n_32754), .c(n_32660), .d(n_32715), .o(n_32784) );
no02s06 FE_RC_6097_0 ( .a(n_17192), .b(n_17084), .o(n_17126) );
no02s02 TIMEBOOST_cell_6865 ( .a(n_36999), .b(n_37070), .o(TIMEBOOST_net_2191) );
in01s10 FE_RC_6099_0 ( .a(n_32704), .o(FE_RN_2712_0) );
in01m08 FE_RC_6100_0 ( .a(FE_RN_176_0), .o(FE_RN_2713_0) );
na02m10 FE_RC_6101_0 ( .a(FE_RN_2712_0), .b(FE_RN_2713_0), .o(FE_RN_2714_0) );
no02m10 FE_RC_6102_0 ( .a(FE_RN_2714_0), .b(n_32643), .o(n_32721) );
oa22m10 FE_RC_6103_0 ( .a(n_27966), .b(FE_RN_1435_0), .c(n_27962), .d(FE_RN_1436_0), .o(n_28116) );
na02f02 TIMEBOOST_cell_8027 ( .a(TIMEBOOST_net_2644), .b(n_16855), .o(TIMEBOOST_net_1761) );
in01s04 FE_RC_6105_0 ( .a(n_28530), .o(FE_RN_2715_0) );
no02m08 FE_RC_6106_0 ( .a(n_28571), .b(FE_RN_2715_0), .o(FE_RN_2716_0) );
na02f08 FE_RC_6107_0 ( .a(n_28871), .b(FE_RN_2716_0), .o(n_28935) );
in01m01 FE_RC_6108_0 ( .a(n_18264), .o(FE_RN_2717_0) );
na02m04 FE_RC_6109_0 ( .a(n_18313), .b(FE_RN_2717_0), .o(FE_RN_2718_0) );
in01s01 FE_RC_610_0 ( .a(n_37471), .o(FE_RN_183_0) );
in01s02 FE_RC_6110_0 ( .a(n_18278), .o(FE_RN_2719_0) );
no02f01 TIMEBOOST_cell_4036 ( .a(n_20081), .b(TIMEBOOST_net_1108), .o(n_20194) );
in01s02 FE_RC_6112_0 ( .a(n_18278), .o(FE_RN_2721_0) );
no03s03 TIMEBOOST_cell_3623 ( .a(FE_RN_1600_0), .b(FE_RN_1601_0), .c(n_2748), .o(n_2859) );
na03m04 TIMEBOOST_cell_3620 ( .a(n_34184), .b(n_34160), .c(n_44102), .o(n_34221) );
no02f04 FE_RC_6118_0 ( .a(n_18892), .b(FE_OFN739_n_17093), .o(FE_RN_2725_0) );
no03s03 TIMEBOOST_cell_5851 ( .a(n_46938), .b(FE_OCP_RBN3307_n_43022), .c(n_43270), .o(n_43327) );
in01s06 FE_RC_611_0 ( .a(n_37078), .o(FE_RN_184_0) );
na02m06 FE_RC_6121_0 ( .a(delay_sub_ln23_0_unr21_stage8_stallmux_q), .b(n_33976), .o(FE_RN_2726_0) );
na02m08 FE_RC_6122_0 ( .a(FE_RN_2726_0), .b(n_34078), .o(n_34124) );
in01s01 FE_RC_6123_0 ( .a(FE_OCPN1373_n_34051), .o(FE_RN_2727_0) );
no02f06 FE_RC_6124_0 ( .a(FE_RN_2727_0), .b(n_34052), .o(n_34095) );
no02s06 FE_RC_6125_0 ( .a(FE_RN_1384_0), .b(n_29477), .o(FE_RN_2728_0) );
no02m08 FE_RC_6126_0 ( .a(FE_RN_2728_0), .b(n_29475), .o(n_29494) );
na02s02 FE_RC_6127_0 ( .a(n_19218), .b(n_19219), .o(FE_RN_2729_0) );
na02m08 FE_RC_6128_0 ( .a(n_19388), .b(FE_RN_2729_0), .o(n_19517) );
na02s01 FE_RC_6129_0 ( .a(n_13000), .b(n_12967), .o(FE_RN_2730_0) );
na02s10 FE_RC_612_0 ( .a(FE_RN_184_0), .b(FE_RN_183_0), .o(FE_RN_185_0) );
no02m04 FE_RC_6130_0 ( .a(FE_RN_2730_0), .b(n_13957), .o(n_13995) );
no02s01 TIMEBOOST_cell_7079 ( .a(FE_OCP_RBN6001_n_30534), .b(FE_OCP_RBN6008_n_30608), .o(TIMEBOOST_net_2298) );
in01s01 FE_RC_6132_0 ( .a(FE_OFN4792_n_13195), .o(FE_RN_2731_0) );
na02f04 FE_RC_6133_0 ( .a(FE_RN_2731_0), .b(FE_RN_2154_0), .o(FE_RN_2732_0) );
na02f08 FE_RC_6134_0 ( .a(FE_RN_2732_0), .b(n_13789), .o(n_13887) );
in01s02 FE_RC_6135_0 ( .a(n_34294), .o(FE_RN_2734_0) );
no02m02 TIMEBOOST_cell_8596 ( .a(n_30737), .b(FE_OCPN1404_n_30823), .o(TIMEBOOST_net_2785) );
na02s02 TIMEBOOST_cell_8750 ( .a(FE_RN_1603_0), .b(FE_RN_1604_0), .o(TIMEBOOST_net_2862) );
in01s01 FE_RC_6138_0 ( .a(FE_RN_2733_0), .o(FE_RN_2736_0) );
in01s02 FE_RC_6139_0 ( .a(FE_RN_2736_0), .o(n_34294) );
na02f04 FE_RC_6141_0 ( .a(n_24661), .b(n_24761), .o(FE_RN_2737_0) );
na02f06 FE_RC_6142_0 ( .a(FE_RN_2737_0), .b(n_24698), .o(n_24760) );
in01s01 FE_RC_6143_0 ( .a(FE_OCPN5102_FE_OCP_RBN5029_n_18678), .o(FE_RN_2738_0) );
no02m03 FE_RC_6144_0 ( .a(FE_RN_2738_0), .b(n_19922), .o(n_20005) );
no02m06 FE_RC_6145_0 ( .a(n_22207), .b(n_24684), .o(FE_RN_2739_0) );
no02f08 FE_RC_6146_0 ( .a(FE_RN_2739_0), .b(n_24870), .o(n_24918) );
na02s06 FE_RC_6147_0 ( .a(n_34241), .b(n_34242), .o(FE_RN_2740_0) );
no02f10 FE_RC_6148_0 ( .a(n_34632), .b(FE_RN_2740_0), .o(n_34661) );
in01s01 FE_RC_6149_0 ( .a(FE_OCP_RBN4084_n_13453), .o(FE_RN_2741_0) );
na02m06 FE_RC_6150_0 ( .a(FE_RN_2741_0), .b(n_14672), .o(n_14754) );
oa22f04 FE_RC_6151_0 ( .a(FE_RN_2742_0), .b(n_20003), .c(n_19838), .d(n_20028), .o(n_20095) );
in01m02 FE_RC_6152_0 ( .a(n_19813), .o(FE_RN_2743_0) );
in01f02 FE_RC_6153_0 ( .a(FE_RN_2743_0), .o(FE_RN_2742_0) );
in01s01 FE_RC_6154_0 ( .a(FE_OCP_RBN4637_n_18600), .o(FE_RN_2744_0) );
no02f04 FE_RC_6155_0 ( .a(n_20095), .b(FE_RN_2744_0), .o(n_20170) );
in01s01 FE_RC_6156_0 ( .a(FE_OCPN4536_n_14543), .o(FE_RN_2745_0) );
na02f06 FE_RC_6157_0 ( .a(FE_RN_2745_0), .b(n_14544), .o(n_14573) );
na02s02 TIMEBOOST_cell_7506 ( .a(n_12652), .b(n_12454), .o(TIMEBOOST_net_2384) );
oa22f02 FE_RC_6159_0 ( .a(n_20194), .b(n_20047), .c(n_20174), .d(n_20046), .o(n_20273) );
in01s04 FE_RC_6160_0 ( .a(n_25182), .o(FE_RN_2746_0) );
in01s04 FE_RC_6161_0 ( .a(n_25154), .o(FE_RN_2747_0) );
in01f02 FE_RC_6162_0 ( .a(n_25155), .o(FE_RN_2748_0) );
na02f08 FE_RC_6163_0 ( .a(FE_RN_2747_0), .b(FE_RN_2748_0), .o(FE_RN_2749_0) );
no02m08 FE_RC_6164_0 ( .a(n_25182), .b(n_25147), .o(FE_RN_2750_0) );
ao22f08 FE_RC_6165_0 ( .a(FE_RN_2746_0), .b(FE_RN_2749_0), .c(FE_RN_2750_0), .d(n_25366), .o(n_25432) );
in01f06 FE_RC_6166_0 ( .a(FE_RN_2751_0), .o(n_35083) );
no02f06 FE_RC_6167_0 ( .a(n_35063), .b(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(FE_RN_2751_0) );
in01s01 FE_RC_6168_0 ( .a(FE_OCP_RBN6639_n_13726), .o(FE_RN_2752_0) );
in01f02 FE_RC_6169_0 ( .a(FE_RN_2753_0), .o(n_15036) );
no02f02 FE_RC_6170_0 ( .a(FE_RN_2752_0), .b(n_14921), .o(FE_RN_2753_0) );
in01s01 FE_RC_6171_0 ( .a(FE_OCPUNCON1750_n_33904), .o(FE_RN_2754_0) );
na02f04 FE_RC_6172_0 ( .a(n_35324), .b(FE_RN_2754_0), .o(n_35360) );
in01s01 FE_RC_6177_0 ( .a(n_25275), .o(FE_RN_2758_0) );
in01s01 FE_RC_6178_0 ( .a(n_25399), .o(FE_RN_2759_0) );
no02s02 FE_RC_6179_0 ( .a(FE_RN_2758_0), .b(FE_RN_2759_0), .o(FE_RN_2760_0) );
in01f02 FE_RC_6180_0 ( .a(FE_RN_2761_0), .o(n_25707) );
na02f02 FE_RC_6181_0 ( .a(n_25656), .b(FE_RN_2760_0), .o(FE_RN_2761_0) );
in01s02 FE_RC_6182_0 ( .a(FE_RN_2635_0), .o(FE_RN_2762_0) );
in01s02 FE_RC_6183_0 ( .a(n_30599), .o(FE_RN_2763_0) );
na02s04 FE_RC_6184_0 ( .a(FE_RN_2762_0), .b(FE_RN_2763_0), .o(FE_RN_2764_0) );
na02m06 FE_RC_6185_0 ( .a(FE_RN_2632_0), .b(FE_RN_2764_0), .o(n_30818) );
na02m04 FE_RC_6186_0 ( .a(n_25458), .b(n_25455), .o(FE_RN_2765_0) );
no02m08 FE_RC_6187_0 ( .a(FE_RN_2765_0), .b(n_25675), .o(n_25726) );
ao22f04 FE_RC_6188_0 ( .a(n_15349), .b(n_15309), .c(n_15308), .d(n_15313), .o(n_15610) );
in01f04 FE_RC_6189_0 ( .a(FE_RN_2766_0), .o(n_25939) );
na03f08 FE_RC_618_0 ( .a(n_37755), .b(n_37756), .c(FE_OCP_RBN4032_n_37690), .o(n_37780) );
no02f04 FE_RC_6190_0 ( .a(n_25847), .b(FE_RN_2767_0), .o(FE_RN_2766_0) );
in01s01 FE_RC_6191_0 ( .a(FE_RN_1106_0), .o(FE_RN_2768_0) );
in01s01 FE_RC_6192_0 ( .a(FE_RN_2768_0), .o(FE_RN_2767_0) );
oa22f04 FE_RC_6193_0 ( .a(n_20877), .b(n_20716), .c(n_20876), .d(n_20960), .o(n_20903) );
oa22f02 FE_RC_6194_0 ( .a(FE_OFN748_n_22641), .b(FE_OCP_RBN1012_n_25826), .c(n_23254), .d(n_25826), .o(n_25920) );
in01m04 FE_RC_6195_0 ( .a(n_35235), .o(FE_RN_2769_0) );
in01f08 FE_RC_6196_0 ( .a(FE_RN_2770_0), .o(n_35365) );
no02f08 FE_RC_6197_0 ( .a(n_35290), .b(FE_RN_2769_0), .o(FE_RN_2770_0) );
in01s01 FE_RC_6198_0 ( .a(FE_OFN747_n_22641), .o(FE_RN_2771_0) );
in01f06 FE_RC_6199_0 ( .a(FE_RN_2772_0), .o(n_26026) );
ao22f04 FE_RC_619_0 ( .a(n_41213), .b(n_40969), .c(FE_OCP_RBN2485_n_41213), .d(n_40970), .o(n_41285) );
in01s02 FE_RC_61_0 ( .a(n_3061), .o(FE_RN_16_0) );
na02f04 FE_RC_6200_0 ( .a(n_25912), .b(FE_RN_2771_0), .o(FE_RN_2772_0) );
na02s03 FE_RC_6201_0 ( .a(n_20489), .b(n_20459), .o(FE_RN_2773_0) );
no02m08 FE_RC_6202_0 ( .a(n_20913), .b(FE_RN_2773_0), .o(n_20932) );
in01s01 FE_RC_6203_0 ( .a(FE_OCP_DRV_N1421_n_35367), .o(FE_RN_2774_0) );
no02f06 FE_RC_6204_0 ( .a(n_35368), .b(FE_RN_2774_0), .o(n_35385) );
no02s06 FE_RC_6205_0 ( .a(n_14239), .b(n_15142), .o(FE_RN_2775_0) );
in01m08 FE_RC_6206_0 ( .a(FE_RN_2776_0), .o(n_15804) );
no02m08 FE_RC_6207_0 ( .a(FE_RN_2775_0), .b(n_15625), .o(FE_RN_2776_0) );
oa22m06 FE_RC_6208_0 ( .a(n_15804), .b(n_15259), .c(FE_OCP_RBN3153_n_15804), .d(n_15298), .o(n_15900) );
in01s01 FE_RC_6209_0 ( .a(n_45024), .o(FE_RN_2777_0) );
no02m04 FE_RC_6210_0 ( .a(FE_RN_2777_0), .b(n_21046), .o(FE_RN_586_0) );
in01s01 TIMEBOOST_cell_5913 ( .a(FE_OFN1_n_43918), .o(TIMEBOOST_net_1802) );
in01m02 FE_RC_6212_0 ( .a(n_21511), .o(FE_RN_2778_0) );
in01m02 FE_RC_6213_0 ( .a(n_21438), .o(FE_RN_2779_0) );
ao22m04 FE_RC_6214_0 ( .a(FE_RN_2778_0), .b(n_21438), .c(FE_RN_2779_0), .d(n_21511), .o(n_21656) );
in01f02 FE_RC_6215_0 ( .a(FE_RN_2780_0), .o(n_21741) );
na02m02 FE_RC_6216_0 ( .a(n_20018), .b(n_21581), .o(FE_RN_2780_0) );
no02s06 TIMEBOOST_cell_1093 ( .a(n_17848), .b(FE_RN_10_0), .o(TIMEBOOST_net_161) );
na02f08 FE_RC_6218_0 ( .a(n_21684), .b(n_21665), .o(FE_RN_2782_0) );
no02s06 TIMEBOOST_cell_1094 ( .a(TIMEBOOST_net_161), .b(n_17923), .o(n_18022) );
oa22m04 FE_RC_621_0 ( .a(FE_OCPN1910_n_40921), .b(n_41256), .c(n_40922), .d(n_41257), .o(n_41312) );
no02f10 FE_RC_6220_0 ( .a(FE_RN_2783_0), .b(n_21617), .o(n_21849) );
in01s04 FE_RC_6221_0 ( .a(n_26580), .o(FE_RN_2784_0) );
no02f08 FE_RC_6222_0 ( .a(n_26781), .b(FE_RN_2784_0), .o(FE_RN_1058_0) );
in01f02 FE_RC_6223_0 ( .a(n_21727), .o(FE_RN_2785_0) );
no02f08 FE_RC_6224_0 ( .a(FE_RN_1184_0), .b(FE_RN_2785_0), .o(FE_RN_2786_0) );
no02f08 FE_RC_6225_0 ( .a(FE_RN_2786_0), .b(n_21676), .o(n_21818) );
in01f02 FE_RC_6226_0 ( .a(n_26564), .o(FE_RN_2787_0) );
in01m02 FE_RC_6227_0 ( .a(n_26516), .o(FE_RN_2788_0) );
in01s01 FE_RC_6229_0 ( .a(FE_OCPN1933_n_26801), .o(FE_RN_2789_0) );
no02m06 TIMEBOOST_cell_1746 ( .a(TIMEBOOST_net_487), .b(n_26355), .o(n_26519) );
na02m06 FE_RC_6230_0 ( .a(FE_RN_2789_0), .b(n_26802), .o(n_26877) );
na02m04 FE_RC_6231_0 ( .a(n_26473), .b(n_26467), .o(FE_RN_2790_0) );
no02m10 FE_RC_6232_0 ( .a(FE_OCP_RBN3356_FE_RN_1058_0), .b(FE_RN_2790_0), .o(n_26987) );
ao22f06 FE_RC_6233_0 ( .a(FE_OCPN1303_n_35945), .b(n_36431), .c(FE_OCPN1304_n_35945), .d(n_36445), .o(n_36489) );
na03s04 FE_RC_6234_0 ( .a(n_22232), .b(n_22231), .c(n_22153), .o(n_22273) );
oa22s02 FE_RC_6235_0 ( .a(n_36490), .b(n_36234), .c(n_36235), .d(FE_OCP_RBN3371_n_36490), .o(n_36567) );
in01s01 FE_RC_6236_0 ( .a(FE_RN_1523_0), .o(FE_RN_2791_0) );
no02s01 FE_RC_6237_0 ( .a(n_20862), .b(FE_RN_2791_0), .o(FE_RN_2792_0) );
no02s06 FE_RC_6238_0 ( .a(FE_RN_2792_0), .b(n_22121), .o(n_22304) );
no02s01 FE_RC_6239_0 ( .a(n_22187), .b(n_20978), .o(n_22213) );
no02s01 FE_RC_6240_0 ( .a(FE_OCP_DRV_N1430_n_22126), .b(n_22187), .o(n_22212) );
in01s01 FE_RC_6241_0 ( .a(FE_OCP_DRV_N1430_n_22126), .o(FE_RN_2793_0) );
in01s01 FE_RC_6242_0 ( .a(n_20978), .o(FE_RN_2794_0) );
no02s01 FE_RC_6243_0 ( .a(FE_RN_2793_0), .b(FE_RN_2794_0), .o(FE_RN_2795_0) );
no02s06 FE_RC_6244_0 ( .a(n_22187), .b(FE_RN_2795_0), .o(FE_RN_2796_0) );
no02m08 FE_RC_6245_0 ( .a(n_22304), .b(FE_RN_2796_0), .o(n_22445) );
no03s02 FE_RC_6246_0 ( .a(n_22383), .b(n_22292), .c(n_22291), .o(FE_RN_1886_0) );
in01s01 FE_RC_6247_0 ( .a(n_16943), .o(FE_RN_2797_0) );
no02s02 FE_RC_6248_0 ( .a(n_17283), .b(FE_RN_2797_0), .o(FE_RN_2798_0) );
na02s06 FE_RC_6249_0 ( .a(FE_RN_2798_0), .b(n_17402), .o(n_17483) );
no02s01 FE_RC_6250_0 ( .a(n_25757), .b(n_25789), .o(FE_RN_2799_0) );
in01s02 FE_RC_6251_0 ( .a(n_27086), .o(FE_RN_2800_0) );
no02s06 FE_RC_6252_0 ( .a(FE_RN_2800_0), .b(FE_RN_2799_0), .o(FE_RN_2801_0) );
no02f10 FE_RC_6253_0 ( .a(n_27514), .b(FE_RN_2801_0), .o(n_27554) );
oa22m04 FE_RC_6254_0 ( .a(n_22544), .b(n_22303), .c(n_22341), .d(n_22566), .o(n_22684) );
oa22f04 FE_RC_6255_0 ( .a(n_22387), .b(n_22603), .c(n_22340), .d(n_22619), .o(n_22778) );
oa22s06 FE_RC_6256_0 ( .a(n_17385), .b(n_17693), .c(n_17384), .d(n_17658), .o(n_17812) );
ao22f02 FE_RC_625_0 ( .a(n_41344), .b(n_41325), .c(n_41353), .d(FE_OCP_RBN4055_n_41325), .o(n_41364) );
in01s01 FE_RC_6266_0 ( .a(n_30955), .o(FE_RN_2811_0) );
oa22f04 FE_RC_6268_0 ( .a(n_22494), .b(n_22574), .c(n_22558), .d(n_22495), .o(n_22715) );
oa22m04 FE_RC_6269_0 ( .a(n_17344), .b(n_17312), .c(n_17311), .d(n_17404), .o(n_17591) );
oa22s01 FE_RC_6270_0 ( .a(n_20231), .b(n_22874), .c(n_20252), .d(n_44327), .o(n_22947) );
oa22s03 FE_RC_6271_0 ( .a(n_22496), .b(n_22744), .c(n_22497), .d(n_22706), .o(n_22902) );
oa22m06 FE_RC_6272_0 ( .a(n_32120), .b(FE_RN_2698_0), .c(FE_RN_2699_0), .d(FE_RN_2701_0), .o(n_32517) );
oa22m02 FE_RC_6273_0 ( .a(n_36758), .b(n_36790), .c(n_36757), .d(n_36791), .o(n_36845) );
no02s01 TIMEBOOST_cell_6673 ( .a(n_2803), .b(FE_RN_2589_0), .o(TIMEBOOST_net_2094) );
no02s02 TIMEBOOST_cell_6674 ( .a(TIMEBOOST_net_2094), .b(n_2729), .o(FE_RN_2590_0) );
in01s06 FE_RC_6276_0 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_4_), .o(FE_RN_2813_0) );
no02s06 TIMEBOOST_cell_5677 ( .a(TIMEBOOST_net_1786), .b(n_27145), .o(FE_RN_2685_0) );
na02m06 TIMEBOOST_cell_5685 ( .a(TIMEBOOST_net_1790), .b(n_36595), .o(n_36675) );
na02m08 TIMEBOOST_cell_3850 ( .a(TIMEBOOST_net_1015), .b(n_7284), .o(n_7346) );
na02s06 TIMEBOOST_cell_3851 ( .a(n_7085), .b(n_7086), .o(TIMEBOOST_net_1016) );
ao22s04 FE_RC_6281_0 ( .a(n_6616), .b(n_6635), .c(n_6617), .d(FE_OCP_RBN2407_n_6635), .o(n_6798) );
in01s02 FE_RC_6282_0 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_0_), .o(FE_RN_2816_0) );
na02m08 FE_RC_6283_0 ( .a(FE_RN_2816_0), .b(n_22632), .o(n_22674) );
oa22m08 FE_RC_6284_0 ( .a(FE_RN_2000_0), .b(FE_RN_2001_0), .c(n_32711), .d(FE_RN_2002_0), .o(n_32794) );
in01s01 FE_RC_6285_0 ( .a(FE_RN_2817_0), .o(n_47210) );
no02s02 FE_RC_6286_0 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_3_), .b(n_6780), .o(FE_RN_2817_0) );
oa22m08 FE_RC_6287_0 ( .a(n_32730), .b(n_32815), .c(n_32729), .d(n_32816), .o(n_32906) );
in01f04 FE_RC_6288_0 ( .a(FE_RN_2818_0), .o(n_32905) );
no02m04 FE_RC_6289_0 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_5_), .b(n_32827), .o(FE_RN_2818_0) );
in01s10 FE_RC_6290_0 ( .a(FE_OCPN1718_n_28065), .o(FE_RN_2819_0) );
no02m20 FE_RC_6291_0 ( .a(FE_RN_2819_0), .b(FE_OCP_RBN5549_n_28319), .o(n_28385) );
no02m06 TIMEBOOST_cell_8649 ( .a(TIMEBOOST_net_2811), .b(n_39594), .o(FE_RN_2164_0) );
no03s01 TIMEBOOST_cell_2442 ( .a(n_2609), .b(FE_OCP_RBN6611_n_2289), .c(FE_OFN798_n_2620), .o(FE_RN_276_0) );
in01f04 FE_RC_6294_0 ( .a(FE_RN_2821_0), .o(FE_OCPN893_n_28471) );
no02f06 FE_RC_6295_0 ( .a(n_28452), .b(n_28453), .o(FE_RN_2821_0) );
no02f01 TIMEBOOST_cell_1703 ( .a(n_3630), .b(n_3624), .o(TIMEBOOST_net_466) );
in01s01 FE_RC_6297_0 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_), .o(FE_RN_2822_0) );
in01s01 FE_RC_6298_0 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_), .o(FE_RN_2823_0) );
na02s01 FE_RC_6299_0 ( .a(FE_RN_2822_0), .b(FE_RN_2823_0), .o(FE_RN_2824_0) );
ao22f04 FE_RC_629_0 ( .a(n_23732), .b(n_24085), .c(n_24084), .d(n_23731), .o(n_24165) );
na02s08 FE_RC_6300_0 ( .a(FE_RN_2824_0), .b(n_28458), .o(n_28632) );
no02s04 TIMEBOOST_cell_1752 ( .a(TIMEBOOST_net_490), .b(n_20767), .o(n_20819) );
in01s01 FE_RC_6302_0 ( .a(n_6749), .o(FE_RN_2826_0) );
in01s01 FE_RC_6303_0 ( .a(FE_RN_2826_0), .o(FE_RN_2825_0) );
no02s02 TIMEBOOST_cell_8836 ( .a(n_4245), .b(FE_OCP_RBN5977_n_4245), .o(TIMEBOOST_net_2905) );
na02m06 TIMEBOOST_cell_4421 ( .a(FE_OCP_RBN3218_n_15992), .b(FE_OCPN1733_n_14524), .o(TIMEBOOST_net_1301) );
in01s01 FE_RC_6306_0 ( .a(FE_RN_2546_0), .o(FE_RN_2828_0) );
na02s02 FE_RC_6307_0 ( .a(n_1746), .b(FE_RN_2828_0), .o(FE_RN_2829_0) );
no02f10 FE_RC_6308_0 ( .a(n_2148), .b(FE_RN_2829_0), .o(n_2151) );
no02s01 FE_RC_6309_0 ( .a(n_6764), .b(n_6765), .o(FE_RN_2830_0) );
no02s01 TIMEBOOST_cell_1877 ( .a(n_35003), .b(FE_OCP_RBN6076_n_44256), .o(TIMEBOOST_net_553) );
na02s01 FE_RC_6310_0 ( .a(FE_RN_2830_0), .b(n_6813), .o(FE_RN_2831_0) );
no02f08 FE_RC_6311_0 ( .a(n_7480), .b(FE_RN_2831_0), .o(n_7516) );
in01s01 FE_RC_6312_0 ( .a(n_1565), .o(FE_RN_2832_0) );
no02s03 FE_RC_6313_0 ( .a(FE_RN_2832_0), .b(FE_OCP_RBN5595_n_45903), .o(n_2266) );
in01s01 FE_RC_6314_0 ( .a(FE_OCP_DRV_N7074_n_7116), .o(FE_RN_2833_0) );
in01s01 TIMEBOOST_cell_5911 ( .a(FE_OFN1_n_43918), .o(TIMEBOOST_net_1800) );
no02s01 TIMEBOOST_cell_4970 ( .a(n_32973), .b(n_32972), .o(TIMEBOOST_net_1433) );
in01s01 FE_RC_6317_0 ( .a(n_23683), .o(FE_RN_2835_0) );
no02s02 FE_RC_6318_0 ( .a(n_23775), .b(FE_RN_2835_0), .o(FE_RN_2836_0) );
na02m04 FE_RC_6319_0 ( .a(FE_RN_2836_0), .b(n_24122), .o(n_24139) );
no02m01 FE_RC_6320_0 ( .a(FE_RN_2838_0), .b(n_24162), .o(FE_RN_2837_0) );
na02m06 FE_RC_6321_0 ( .a(FE_RN_2837_0), .b(n_24200), .o(n_24224) );
in01s01 FE_RC_6322_0 ( .a(n_23740), .o(FE_RN_2839_0) );
in01s01 FE_RC_6323_0 ( .a(FE_RN_2839_0), .o(FE_RN_2838_0) );
ao22f04 FE_RC_6324_0 ( .a(n_33664), .b(FE_OCP_RBN7029_n_44259), .c(n_44259), .d(FE_OCP_RBN2550_n_33664), .o(n_33780) );
in01s01 FE_RC_6325_0 ( .a(n_28826), .o(FE_RN_2840_0) );
na02m06 FE_RC_6326_0 ( .a(n_29279), .b(FE_RN_2840_0), .o(FE_RN_2841_0) );
in01s01 FE_RC_6327_0 ( .a(n_28826), .o(FE_RN_2842_0) );
oa12m06 FE_RC_6328_0 ( .a(FE_RN_2841_0), .b(FE_RN_2842_0), .c(n_29279), .o(n_29371) );
in01s01 FE_RC_6329_0 ( .a(n_18741), .o(FE_RN_2843_0) );
no02s02 FE_RC_6330_0 ( .a(n_18821), .b(FE_RN_2843_0), .o(FE_RN_2844_0) );
na02s08 FE_RC_6331_0 ( .a(FE_RN_2844_0), .b(n_19210), .o(n_19246) );
in01s02 FE_RC_6332_0 ( .a(FE_OCP_RBN2570_n_33735), .o(FE_RN_2845_0) );
in01m02 FE_RC_6333_0 ( .a(n_33834), .o(FE_RN_2846_0) );
no02s02 TIMEBOOST_cell_4172 ( .a(TIMEBOOST_net_1176), .b(n_36467), .o(n_36543) );
na02m08 TIMEBOOST_cell_5010 ( .a(n_18434), .b(n_18372), .o(TIMEBOOST_net_1453) );
in01s01 FE_RC_6336_0 ( .a(FE_OCP_DRV_N6904_n_33945), .o(FE_RN_2848_0) );
na02f06 FE_RC_6337_0 ( .a(FE_RN_2848_0), .b(n_33946), .o(n_33966) );
na02m01 FE_RC_6338_0 ( .a(FE_OCP_RBN2654_FE_OCPN914_n_8091), .b(FE_OCP_RBN5607_n_7730), .o(FE_RN_2849_0) );
na02m08 FE_RC_6339_0 ( .a(FE_RN_2849_0), .b(n_7985), .o(n_8095) );
na02s01 FE_RC_6340_0 ( .a(n_7827), .b(n_7805), .o(FE_RN_2850_0) );
no02f06 FE_RC_6341_0 ( .a(FE_RN_2850_0), .b(n_8215), .o(n_8283) );
na02s03 FE_RC_6342_0 ( .a(n_17900), .b(n_19110), .o(FE_RN_2851_0) );
na02f08 FE_RC_6343_0 ( .a(n_19474), .b(FE_RN_2851_0), .o(n_19516) );
ao22f02 FE_RC_6344_0 ( .a(n_13437), .b(n_13949), .c(n_13195), .d(n_13960), .o(n_14127) );
ao22m04 FE_RC_6345_0 ( .a(FE_RN_1293_0), .b(n_29732), .c(FE_OCP_RBN2650_n_29470), .d(n_29719), .o(n_29813) );
na02s01 FE_RC_6346_0 ( .a(n_33708), .b(n_34200), .o(FE_RN_2853_0) );
na02m08 FE_RC_6347_0 ( .a(FE_RN_2853_0), .b(FE_OCP_RBN5712_n_44102), .o(n_34192) );
in01s01 FE_RC_6348_0 ( .a(FE_RN_2852_0), .o(FE_RN_2854_0) );
in01s01 FE_RC_6349_0 ( .a(FE_RN_2854_0), .o(n_34200) );
no02s03 TIMEBOOST_cell_1882 ( .a(TIMEBOOST_net_555), .b(n_35827), .o(n_35867) );
in01s01 FE_RC_6351_0 ( .a(n_28830), .o(FE_RN_2855_0) );
na02s04 FE_RC_6352_0 ( .a(FE_RN_2855_0), .b(n_29846), .o(n_29968) );
oa22f02 FE_RC_6353_0 ( .a(n_8189), .b(n_8835), .c(FE_OCP_RBN4146_n_7743), .d(FE_OCP_RBN2813_n_8835), .o(n_8953) );
na02s04 FE_RC_6354_0 ( .a(n_18140), .b(n_19580), .o(FE_RN_2856_0) );
na02m08 FE_RC_6355_0 ( .a(FE_RN_2856_0), .b(n_20002), .o(n_20062) );
in01s01 FE_RC_6356_0 ( .a(n_9012), .o(FE_RN_2857_0) );
na02f02 FE_RC_6357_0 ( .a(FE_RN_2857_0), .b(n_8953), .o(FE_RN_2222_0) );
in01m02 FE_RC_6358_0 ( .a(n_14370), .o(FE_RN_2858_0) );
no02f04 FE_RC_6359_0 ( .a(n_14483), .b(FE_RN_2858_0), .o(n_14552) );
in01s01 FE_RC_6360_0 ( .a(FE_OCP_RBN4084_n_13453), .o(FE_RN_2859_0) );
no02m06 FE_RC_6361_0 ( .a(FE_RN_2859_0), .b(n_14672), .o(n_14697) );
oa22m06 FE_RC_6364_0 ( .a(n_34622), .b(n_34875), .c(n_34623), .d(n_34901), .o(n_34999) );
in01s01 FE_RC_6365_0 ( .a(n_8232), .o(FE_RN_2861_0) );
in01m02 FE_RC_6366_0 ( .a(FE_RN_2862_0), .o(n_9503) );
no02m02 FE_RC_6367_0 ( .a(FE_RN_2861_0), .b(n_9360), .o(FE_RN_2862_0) );
in01s01 FE_RC_6368_0 ( .a(FE_OCP_RBN5622_n_18986), .o(FE_RN_2863_0) );
na02s06 FE_RC_6369_0 ( .a(FE_RN_2863_0), .b(n_20249), .o(n_20311) );
in01s01 FE_RC_636_0 ( .a(n_7447), .o(FE_RN_186_0) );
na02f06 FE_RC_6370_0 ( .a(n_30354), .b(n_30176), .o(n_30409) );
oa22m04 FE_RC_6372_0 ( .a(n_9543), .b(n_9638), .c(n_9569), .d(n_9628), .o(n_9864) );
in01s01 FE_RC_6373_0 ( .a(FE_OCPN1672_n_14055), .o(FE_RN_2864_0) );
no02s08 FE_RC_6374_0 ( .a(FE_OCP_RBN4324_n_15156), .b(FE_RN_2864_0), .o(n_15461) );
in01s01 FE_RC_6375_0 ( .a(FE_OCP_DRV_N6266_FE_OCP_RBN1823_n_19434), .o(FE_RN_2865_0) );
na02s06 FE_RC_6376_0 ( .a(n_20456), .b(FE_RN_2865_0), .o(n_20533) );
ao22f06 FE_RC_6377_0 ( .a(n_30259), .b(n_30623), .c(n_30260), .d(n_30605), .o(n_30731) );
in01s01 FE_RC_6378_0 ( .a(n_45010), .o(FE_RN_2866_0) );
in01f02 FE_RC_6379_0 ( .a(FE_RN_2867_0), .o(n_20980) );
no02s02 TIMEBOOST_cell_7920 ( .a(n_5540), .b(n_5500), .o(TIMEBOOST_net_2591) );
no02f02 FE_RC_6380_0 ( .a(FE_RN_2866_0), .b(n_20857), .o(FE_RN_2867_0) );
na02s02 FE_RC_6381_0 ( .a(FE_OCPN5105_n_30371), .b(FE_RN_2869_0), .o(FE_RN_2868_0) );
no02m08 FE_RC_6382_0 ( .a(n_30676), .b(FE_RN_2868_0), .o(n_30739) );
in01s01 FE_RC_6383_0 ( .a(n_30372), .o(FE_RN_2870_0) );
in01s01 FE_RC_6384_0 ( .a(FE_RN_2870_0), .o(FE_RN_2869_0) );
no02s02 FE_RC_6385_0 ( .a(n_15127), .b(n_47261), .o(FE_RN_2871_0) );
na02s06 FE_RC_6386_0 ( .a(n_15625), .b(FE_RN_2871_0), .o(n_15739) );
oa22f04 FE_RC_6387_0 ( .a(n_10032), .b(n_10203), .c(n_10200), .d(n_10033), .o(n_10399) );
in01s01 FE_RC_6388_0 ( .a(FE_OFN757_n_44464), .o(FE_RN_2872_0) );
in01f02 FE_RC_6389_0 ( .a(FE_RN_2873_0), .o(n_10598) );
in01m06 FE_RC_638_0 ( .a(FE_RN_188_0), .o(n_8186) );
no02f02 FE_RC_6390_0 ( .a(FE_RN_2872_0), .b(n_10513), .o(FE_RN_2873_0) );
in01s01 FE_RC_6391_0 ( .a(n_10464), .o(FE_RN_2874_0) );
in01s02 FE_RC_6392_0 ( .a(n_10465), .o(FE_RN_2875_0) );
ao22f06 FE_RC_6393_0 ( .a(FE_RN_2874_0), .b(FE_RN_2875_0), .c(n_46420), .d(n_10740), .o(n_10779) );
in01s01 FE_RC_6394_0 ( .a(FE_OCPN5219_n_10300), .o(FE_RN_2876_0) );
na02s06 FE_RC_6395_0 ( .a(n_10760), .b(FE_RN_2876_0), .o(n_10827) );
in01s01 FE_RC_6396_0 ( .a(n_31079), .o(n_31097) );
no02s06 TIMEBOOST_cell_8466 ( .a(FE_OCP_RBN6466_n_44061), .b(FE_OCP_RBN1118_delay_xor_ln22_unr15_stage6_stallmux_q_0_), .o(TIMEBOOST_net_2720) );
oa22f02 FE_RC_6398_0 ( .a(n_21326), .b(FE_OCP_RBN3723_n_21442), .c(n_21442), .d(n_21327), .o(n_21581) );
ao22f04 FE_RC_6399_0 ( .a(n_26516), .b(FE_RN_2787_0), .c(FE_RN_2788_0), .d(n_26564), .o(n_26721) );
na02s02 TIMEBOOST_cell_8807 ( .a(TIMEBOOST_net_2890), .b(n_42414), .o(FE_RN_1350_0) );
in01s01 FE_RC_6400_0 ( .a(FE_OCPN5235_n_44162), .o(FE_RN_2877_0) );
no02m04 FE_RC_6401_0 ( .a(FE_RN_2877_0), .b(n_21973), .o(n_22028) );
in01s01 FE_RC_6402_0 ( .a(n_30534), .o(FE_RN_2878_0) );
no02s01 FE_RC_6403_0 ( .a(FE_RN_2878_0), .b(FE_OCP_RBN6812_n_30608), .o(FE_RN_2879_0) );
no02s06 FE_RC_6404_0 ( .a(FE_OCP_RBN3391_n_31819), .b(FE_RN_2879_0), .o(n_31993) );
na02s01 TIMEBOOST_cell_1380 ( .a(n_33764), .b(TIMEBOOST_net_304), .o(n_33931) );
in01s01 FE_RC_6406_0 ( .a(FE_RN_2811_0), .o(FE_RN_2880_0) );
no02s01 TIMEBOOST_cell_1171 ( .a(n_37789), .b(n_37731), .o(TIMEBOOST_net_200) );
no02s01 TIMEBOOST_cell_1172 ( .a(TIMEBOOST_net_200), .b(n_37726), .o(n_37790) );
in01s01 FE_RC_6409_0 ( .a(n_32024), .o(FE_RN_2883_0) );
in01s01 FE_RC_640_0 ( .a(n_7318), .o(FE_RN_189_0) );
no02s02 FE_RC_6410_0 ( .a(FE_RN_2883_0), .b(FE_RN_2882_0), .o(FE_RN_2884_0) );
na02s02 FE_RC_6411_0 ( .a(n_47274), .b(n_31990), .o(FE_RN_2885_0) );
in01s02 FE_RC_6412_0 ( .a(n_32021), .o(FE_RN_2886_0) );
no02s06 FE_RC_6413_0 ( .a(FE_RN_2885_0), .b(FE_RN_2886_0), .o(FE_RN_2887_0) );
no02m08 TIMEBOOST_cell_1413 ( .a(FE_RN_1269_0), .b(n_23824), .o(TIMEBOOST_net_321) );
no02m10 TIMEBOOST_cell_1414 ( .a(n_24127), .b(TIMEBOOST_net_321), .o(n_24274) );
oa22s02 FE_RC_6416_0 ( .a(n_32124), .b(n_32365), .c(n_32125), .d(n_32364), .o(n_32519) );
oa22f04 FE_RC_6417_0 ( .a(n_32975), .b(n_33428), .c(n_32974), .d(n_33427), .o(n_33503) );
ao22m04 FE_RC_6418_0 ( .a(n_18638), .b(FE_OCP_RBN5640_n_19060), .c(n_18637), .d(n_19060), .o(n_19177) );
ao22f04 FE_RC_6419_0 ( .a(n_19134), .b(n_19387), .c(n_19164), .d(n_19386), .o(n_19563) );
in01s01 FE_RC_641_0 ( .a(n_45875), .o(FE_RN_190_0) );
ao22m04 FE_RC_6420_0 ( .a(FE_OCP_RBN4202_n_13796), .b(n_14441), .c(FE_OCP_RBN2762_n_13796), .d(FE_OCP_RBN2815_n_14441), .o(n_14571) );
oa22f04 FE_RC_6421_0 ( .a(n_20671), .b(n_21088), .c(n_20670), .d(n_21089), .o(n_21238) );
oa22f04 FE_RC_6422_0 ( .a(n_21227), .b(FE_RN_1531_0), .c(n_21224), .d(FE_RN_1532_0), .o(n_21435) );
oa22m04 FE_RC_6423_0 ( .a(n_36186), .b(n_45625), .c(n_36187), .d(n_36508), .o(n_36592) );
oa22f04 FE_RC_6424_0 ( .a(n_21132), .b(n_44718), .c(n_21133), .d(n_44717), .o(n_21285) );
na02s04 FE_RC_642_0 ( .a(FE_RN_189_0), .b(FE_RN_190_0), .o(FE_RN_191_0) );
na02s06 FE_RC_643_0 ( .a(FE_RN_191_0), .b(n_7868), .o(n_46991) );
ao22f04 FE_RC_644_0 ( .a(n_38160), .b(n_38447), .c(n_38161), .d(n_38446), .o(n_38534) );
ao22m02 FE_RC_646_0 ( .a(n_7438), .b(n_8044), .c(n_7437), .d(n_8043), .o(n_8163) );
oa22f04 FE_RC_655_0 ( .a(n_41997), .b(n_41779), .c(n_41780), .d(n_41996), .o(n_42051) );
oa22f04 FE_RC_656_0 ( .a(n_7546), .b(n_8381), .c(n_7545), .d(n_8382), .o(n_8498) );
ao22m04 FE_RC_657_0 ( .a(n_7587), .b(n_8434), .c(n_7586), .d(n_8435), .o(n_8548) );
oa22m02 FE_RC_658_0 ( .a(n_8295), .b(n_7452), .c(n_8294), .d(n_7453), .o(n_8402) );
ao22s06 FE_RC_65_0 ( .a(n_18545), .b(n_19003), .c(n_18544), .d(n_19002), .o(n_19148) );
oa22m02 FE_RC_660_0 ( .a(n_7640), .b(n_8523), .c(n_7639), .d(FE_OCP_RBN5716_n_8523), .o(n_8637) );
na02m08 TIMEBOOST_cell_6022 ( .a(TIMEBOOST_net_1862), .b(FE_OCP_RBN2508_n_37720), .o(n_37763) );
oa22m02 FE_RC_669_0 ( .a(delay_sub_ln23_0_unr29_stage10_stallmux_q), .b(n_42169), .c(n_42196), .d(FE_OCP_RBN5844_n_42169), .o(n_42187) );
no02s03 FE_RC_672_0 ( .a(FE_OCP_RBN4211_n_8767), .b(FE_OCP_RBN5822_n_8985), .o(FE_RN_197_0) );
no02s04 FE_RC_673_0 ( .a(FE_RN_197_0), .b(n_8986), .o(n_9087) );
ao22f04 FE_RC_678_0 ( .a(n_20279), .b(n_20376), .c(n_20280), .d(n_20344), .o(n_20504) );
ao22f04 FE_RC_680_0 ( .a(n_20303), .b(n_20414), .c(n_20286), .d(n_20415), .o(n_20545) );
na03m04 TIMEBOOST_cell_3680 ( .a(n_3994), .b(FE_OCP_RBN6770_n_3700), .c(n_4024), .o(n_4300) );
oa22f04 FE_RC_686_0 ( .a(n_20874), .b(n_20905), .c(n_20904), .d(n_20875), .o(n_21059) );
oa22f04 FE_RC_68_0 ( .a(n_18639), .b(n_19108), .c(n_19107), .d(n_18640), .o(n_19241) );
oa22s02 FE_RC_700_0 ( .a(n_22907), .b(n_22901), .c(n_22833), .d(n_22861), .o(n_22960) );
in01s01 FE_RC_701_0 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_23_), .o(FE_RN_198_0) );
in01s06 FE_RC_702_0 ( .a(n_36988), .o(FE_RN_199_0) );
na02s02 TIMEBOOST_cell_3880 ( .a(TIMEBOOST_net_1030), .b(n_46252), .o(n_45890) );
no02m04 TIMEBOOST_cell_8553 ( .a(TIMEBOOST_net_2763), .b(TIMEBOOST_net_2234), .o(n_8235) );
no02s06 TIMEBOOST_cell_1732 ( .a(TIMEBOOST_net_480), .b(FE_RN_326_0), .o(n_47008) );
no03s08 TIMEBOOST_cell_2172 ( .a(n_32547), .b(n_32625), .c(TIMEBOOST_net_587), .o(n_32626) );
in01s01 FE_RC_707_0 ( .a(n_28523), .o(FE_RN_201_0) );
in01s01 FE_RC_708_0 ( .a(n_28533), .o(FE_RN_202_0) );
na02s02 TIMEBOOST_cell_8879 ( .a(TIMEBOOST_net_2926), .b(n_32044), .o(n_32122) );
na02m06 TIMEBOOST_cell_4918 ( .a(n_6968), .b(n_6969), .o(TIMEBOOST_net_1407) );
in01s02 FE_RC_711_0 ( .a(n_32863), .o(FE_RN_204_0) );
na02m04 TIMEBOOST_cell_5657 ( .a(TIMEBOOST_net_1776), .b(n_11350), .o(n_11453) );
in01m04 FE_RC_713_0 ( .a(FE_RN_206_0), .o(n_32923) );
no02s03 TIMEBOOST_cell_1793 ( .a(n_10765), .b(n_10470), .o(TIMEBOOST_net_511) );
ao22f02 FE_RC_720_0 ( .a(n_38153), .b(n_38418), .c(n_38154), .d(n_38419), .o(n_38515) );
no02s01 TIMEBOOST_cell_1591 ( .a(FE_OCP_RBN2816_n_34509), .b(n_34564), .o(TIMEBOOST_net_410) );
ao22f02 FE_RC_723_0 ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .b(n_38515), .c(n_38778), .d(FE_OCP_RBN5690_n_38515), .o(n_38579) );
in01s01 FE_RC_724_0 ( .a(n_28460), .o(FE_RN_210_0) );
in01s02 FE_RC_725_0 ( .a(n_28575), .o(FE_RN_211_0) );
na02s04 FE_RC_726_0 ( .a(FE_RN_210_0), .b(FE_RN_211_0), .o(FE_RN_212_0) );
na02m04 FE_RC_727_0 ( .a(n_28682), .b(FE_RN_212_0), .o(n_28705) );
no02s02 TIMEBOOST_cell_1685 ( .a(n_25369), .b(n_25408), .o(TIMEBOOST_net_457) );
no03s02 FE_RC_729_0 ( .a(n_38111), .b(n_38088), .c(n_38112), .o(n_38113) );
ao22f08 FE_RC_730_0 ( .a(n_39177), .b(n_39469), .c(n_39176), .d(n_39441), .o(n_39553) );
in01s02 FE_RC_731_0 ( .a(n_17713), .o(FE_RN_213_0) );
in01s02 FE_RC_732_0 ( .a(n_17355), .o(FE_RN_214_0) );
na02s06 FE_RC_733_0 ( .a(FE_RN_213_0), .b(FE_RN_214_0), .o(FE_RN_215_0) );
no02f08 FE_RC_734_0 ( .a(n_17736), .b(FE_RN_215_0), .o(n_17787) );
na02m06 TIMEBOOST_cell_2122 ( .a(TIMEBOOST_net_675), .b(n_26976), .o(n_27067) );
oa22f08 FE_RC_738_0 ( .a(n_34533), .b(n_34900), .c(n_34534), .d(n_34874), .o(n_35001) );
oa22f08 FE_RC_741_0 ( .a(n_39226), .b(n_39467), .c(n_39227), .d(n_39466), .o(n_39551) );
oa22m04 FE_RC_742_0 ( .a(n_34304), .b(n_34729), .c(n_34305), .d(n_34715), .o(n_34836) );
in01s01 FE_RC_743_0 ( .a(n_23599), .o(FE_RN_216_0) );
na02s03 TIMEBOOST_cell_8129 ( .a(TIMEBOOST_net_2695), .b(n_22374), .o(n_22492) );
in01s02 FE_RC_745_0 ( .a(FE_RN_218_0), .o(n_23741) );
no02m02 TIMEBOOST_cell_6097 ( .a(n_14229), .b(n_14187), .o(TIMEBOOST_net_1900) );
in01s06 FE_RC_749_0 ( .a(n_11643), .o(FE_RN_220_0) );
na02s10 FE_RC_750_0 ( .a(FE_RN_220_0), .b(FE_OCP_RBN6531_n_11780), .o(FE_RN_221_0) );
no02s10 FE_RC_751_0 ( .a(n_11962), .b(FE_RN_221_0), .o(n_47211) );
no02m04 TIMEBOOST_cell_6998 ( .a(TIMEBOOST_net_2257), .b(n_15569), .o(n_15637) );
no02s01 TIMEBOOST_cell_6095 ( .a(n_34003), .b(FE_OCP_RBN5714_n_44102), .o(TIMEBOOST_net_1899) );
in01s01 FE_RC_757_0 ( .a(n_32791), .o(FE_RN_222_0) );
in01m06 FE_RC_758_0 ( .a(n_32549), .o(FE_RN_223_0) );
no02m04 FE_RC_759_0 ( .a(FE_RN_222_0), .b(FE_RN_223_0), .o(FE_RN_224_0) );
na02f04 TIMEBOOST_cell_7693 ( .a(TIMEBOOST_net_2477), .b(n_14880), .o(n_14917) );
oa22f04 FE_RC_766_0 ( .a(n_41233), .b(n_40949), .c(n_40950), .d(n_41222), .o(n_41302) );
in01s01 FE_RC_769_0 ( .a(n_6539), .o(FE_RN_228_0) );
in01s01 FE_RC_770_0 ( .a(n_6876), .o(FE_RN_229_0) );
no02s02 FE_RC_771_0 ( .a(FE_RN_229_0), .b(FE_RN_228_0), .o(FE_RN_230_0) );
in01s02 FE_RC_773_0 ( .a(n_11983), .o(FE_RN_231_0) );
no02s02 TIMEBOOST_cell_7979 ( .a(TIMEBOOST_net_2620), .b(n_4847), .o(n_5015) );
in01s06 FE_RC_777_0 ( .a(n_18137), .o(FE_RN_234_0) );
in01s10 FE_RC_778_0 ( .a(n_17977), .o(FE_RN_235_0) );
na02s10 FE_RC_779_0 ( .a(FE_RN_235_0), .b(FE_RN_234_0), .o(FE_RN_236_0) );
no02s02 TIMEBOOST_cell_1677 ( .a(n_26037), .b(FE_RN_1793_0), .o(TIMEBOOST_net_453) );
na02s06 FE_RC_785_0 ( .a(n_1402), .b(FE_OCPN3545_n_1705), .o(FE_RN_239_0) );
no02s02 TIMEBOOST_cell_1617 ( .a(n_34687), .b(n_34239), .o(TIMEBOOST_net_423) );
in01s03 FE_RC_788_0 ( .a(n_17967), .o(FE_RN_240_0) );
in01s03 FE_RC_789_0 ( .a(n_17891), .o(FE_RN_241_0) );
na02s03 FE_RC_790_0 ( .a(FE_RN_240_0), .b(FE_RN_241_0), .o(FE_RN_242_0) );
no02m02 TIMEBOOST_cell_1680 ( .a(TIMEBOOST_net_454), .b(n_9110), .o(n_9241) );
no02m02 FE_RC_798_0 ( .a(FE_OCP_RBN2513_n_28699), .b(FE_OCP_RBN2523_n_29017), .o(FE_RN_245_0) );
na02m04 FE_RC_799_0 ( .a(FE_RN_245_0), .b(n_29018), .o(n_29038) );
na02m08 TIMEBOOST_cell_6917 ( .a(FE_OFN741_delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n_24222), .o(TIMEBOOST_net_2217) );
no03f10 FE_RC_801_0 ( .a(n_37173), .b(n_36981), .c(n_37090), .o(n_37209) );
na02s06 FE_RC_804_0 ( .a(FE_OCP_RBN5539_n_23307), .b(FE_OCP_RBN2422_n_23023), .o(FE_RN_248_0) );
no02s01 TIMEBOOST_cell_4147 ( .a(FE_OFN5084_n_36750), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_1164) );
in01s01 FE_RC_806_0 ( .a(n_6932), .o(FE_RN_249_0) );
no02s02 TIMEBOOST_cell_8572 ( .a(n_4220), .b(n_4165), .o(TIMEBOOST_net_2773) );
no02s02 TIMEBOOST_cell_8672 ( .a(n_26009), .b(FE_OFN748_n_22641), .o(TIMEBOOST_net_2823) );
na02s01 TIMEBOOST_cell_6395 ( .a(FE_OCP_RBN6031_n_25997), .b(n_27120), .o(TIMEBOOST_net_2049) );
oa22m04 FE_RC_811_0 ( .a(n_23017), .b(n_23195), .c(n_23212), .d(n_23018), .o(n_23266) );
in01m04 FE_RC_812_0 ( .a(n_12477), .o(FE_RN_252_0) );
in01m01 FE_RC_813_0 ( .a(n_12492), .o(FE_RN_253_0) );
no02s02 TIMEBOOST_cell_7729 ( .a(TIMEBOOST_net_2495), .b(n_26611), .o(n_26645) );
no02s02 TIMEBOOST_cell_1811 ( .a(n_30678), .b(n_30403), .o(TIMEBOOST_net_520) );
in01m06 FE_RC_818_0 ( .a(n_32553), .o(FE_RN_255_0) );
in01s06 FE_RC_819_0 ( .a(n_32579), .o(FE_RN_256_0) );
na02m08 FE_RC_820_0 ( .a(FE_RN_255_0), .b(FE_RN_256_0), .o(FE_RN_257_0) );
no02s08 TIMEBOOST_cell_8683 ( .a(TIMEBOOST_net_2828), .b(TIMEBOOST_net_915), .o(n_21466) );
in01s02 FE_RC_823_0 ( .a(n_23327), .o(FE_RN_259_0) );
in01m04 FE_RC_824_0 ( .a(FE_RN_260_0), .o(n_23404) );
no02f08 TIMEBOOST_cell_1768 ( .a(TIMEBOOST_net_498), .b(n_39589), .o(n_39617) );
na02s01 FE_RC_828_0 ( .a(FE_RN_264_0), .b(FE_RN_265_0), .o(FE_RN_263_0) );
na02f08 FE_RC_829_0 ( .a(FE_RN_263_0), .b(FE_OCP_RBN2443_n_44798), .o(n_40893) );
ao22f06 FE_RC_831_0 ( .a(FE_OCPN1689_n_23167), .b(n_23439), .c(FE_OCPN1688_n_23167), .d(n_23453), .o(n_23539) );
in01s01 FE_RC_832_0 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_), .o(FE_RN_264_0) );
in01s01 FE_RC_833_0 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_), .o(FE_RN_265_0) );
no02s02 FE_RC_834_0 ( .a(FE_RN_265_0), .b(FE_RN_264_0), .o(FE_RN_266_0) );
no02m10 FE_RC_835_0 ( .a(FE_RN_266_0), .b(n_44798), .o(n_40826) );
in01s01 FE_RC_837_0 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_13_), .o(FE_RN_267_0) );
in01s01 FE_RC_838_0 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_12_), .o(FE_RN_268_0) );
no02s01 FE_RC_839_0 ( .a(FE_RN_267_0), .b(FE_RN_268_0), .o(FE_RN_269_0) );
in01s04 FE_RC_83_0 ( .a(n_19859), .o(FE_RN_18_0) );
no02s03 FE_RC_840_0 ( .a(FE_RN_269_0), .b(FE_OCP_RBN4003_n_33015), .o(n_33380) );
no02f08 TIMEBOOST_cell_1638 ( .a(TIMEBOOST_net_433), .b(n_14628), .o(n_14801) );
oa22m04 FE_RC_844_0 ( .a(n_45508), .b(n_40627), .c(n_47203), .d(n_40628), .o(n_40676) );
in01f03 FE_RC_845_0 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_7_), .o(FE_RN_270_0) );
in01s06 FE_RC_846_0 ( .a(FE_OCP_RBN5513_n_44365), .o(FE_RN_271_0) );
no02f04 TIMEBOOST_cell_1682 ( .a(n_45631), .b(TIMEBOOST_net_455), .o(n_30388) );
no02s02 TIMEBOOST_cell_5353 ( .a(TIMEBOOST_net_1624), .b(n_3838), .o(n_5603) );
in01s03 FE_RC_84_0 ( .a(n_20079), .o(FE_RN_19_0) );
in01s01 FE_RC_851_0 ( .a(n_1842), .o(FE_RN_273_0) );
no02f04 TIMEBOOST_cell_6852 ( .a(TIMEBOOST_net_2183), .b(n_44158), .o(n_21271) );
no03f10 TIMEBOOST_cell_546 ( .a(FE_RN_2782_0), .b(n_21507), .c(n_21658), .o(FE_RN_2783_0) );
in01m02 FE_RC_857_0 ( .a(n_2735), .o(FE_RN_277_0) );
in01m02 FE_RC_858_0 ( .a(FE_RN_278_0), .o(n_2821) );
no02m02 FE_RC_859_0 ( .a(FE_RN_276_0), .b(FE_RN_277_0), .o(FE_RN_278_0) );
na02s06 TIMEBOOST_cell_6668 ( .a(TIMEBOOST_net_2091), .b(n_19862), .o(n_19973) );
oa22s02 FE_RC_862_0 ( .a(n_1567), .b(n_1808), .c(n_1568), .d(n_1813), .o(n_1865) );
oa22s02 FE_RC_866_0 ( .a(n_32349), .b(n_32126), .c(n_32127), .d(n_32366), .o(n_32518) );
na02f10 TIMEBOOST_cell_2072 ( .a(TIMEBOOST_net_650), .b(n_34440), .o(n_34632) );
oa22f08 FE_RC_873_0 ( .a(n_32551), .b(n_32583), .c(n_32552), .d(n_32641), .o(n_32671) );
oa22s01 FE_RC_874_0 ( .a(n_32566), .b(n_32516), .c(n_28336), .d(FE_OCP_RBN5352_n_32516), .o(n_32567) );
oa22m01 FE_RC_875_0 ( .a(n_32287), .b(n_32546), .c(n_28336), .d(n_32513), .o(n_32594) );
in01s01 FE_RC_876_0 ( .a(n_37426), .o(FE_RN_282_0) );
in01s02 FE_RC_877_0 ( .a(n_37220), .o(FE_RN_283_0) );
na02s06 FE_RC_878_0 ( .a(FE_RN_282_0), .b(FE_RN_283_0), .o(FE_RN_284_0) );
no02s01 TIMEBOOST_cell_2138 ( .a(TIMEBOOST_net_683), .b(n_40110), .o(n_40249) );
oa22f04 FE_RC_883_0 ( .a(n_12755), .b(n_13267), .c(n_12756), .d(n_13266), .o(n_13453) );
in01s06 FE_RC_884_0 ( .a(n_28011), .o(FE_RN_285_0) );
in01s03 FE_RC_885_0 ( .a(n_28012), .o(FE_RN_286_0) );
no02s02 TIMEBOOST_cell_6717 ( .a(FE_OCP_RBN2659_n_2832), .b(n_2867), .o(TIMEBOOST_net_2116) );
no02m04 TIMEBOOST_cell_6040 ( .a(TIMEBOOST_net_1871), .b(n_24566), .o(TIMEBOOST_net_793) );
oa22m04 FE_RC_888_0 ( .a(n_11802), .b(n_12023), .c(n_11801), .d(n_11988), .o(n_12211) );
oa22s02 FE_RC_889_0 ( .a(n_11804), .b(n_11990), .c(n_11803), .d(n_12025), .o(n_12212) );
oa22f02 FE_RC_88_0 ( .a(n_19238), .b(FE_OCP_RBN5380_n_19428), .c(n_19428), .d(n_19203), .o(n_19591) );
ao22m02 FE_RC_890_0 ( .a(n_12024), .b(n_11809), .c(n_11808), .d(n_11989), .o(n_12067) );
oa22f04 FE_RC_891_0 ( .a(n_12819), .b(n_13343), .c(n_12820), .d(n_13344), .o(n_13489) );
in01s01 FE_RC_892_0 ( .a(n_17661), .o(FE_RN_288_0) );
na03m08 TIMEBOOST_cell_6552 ( .a(n_24993), .b(n_24804), .c(n_44445), .o(n_25098) );
na02s01 TIMEBOOST_cell_7504 ( .a(n_549), .b(n_241), .o(TIMEBOOST_net_2383) );
oa22f02 FE_RC_900_0 ( .a(FE_OFN4787_n_46137), .b(n_6725), .c(FE_OFN770_n_46196), .d(n_6774), .o(n_46193) );
oa22s02 FE_RC_901_0 ( .a(FE_OFN770_n_46196), .b(n_6719), .c(FE_OFN4787_n_46137), .d(n_6701), .o(n_46194) );
oa22s02 FE_RC_914_0 ( .a(FE_OFN770_n_46196), .b(n_6643), .c(FE_OFN4787_n_46137), .d(n_6587), .o(n_46189) );
oa22s04 FE_RC_917_0 ( .a(n_6555), .b(n_6453), .c(n_6454), .d(n_6581), .o(n_6719) );
in01s01 TIMEBOOST_cell_8888 ( .a(n_1065), .o(TIMEBOOST_net_2932) );
no02s02 TIMEBOOST_cell_2015 ( .a(n_13323), .b(n_13120), .o(TIMEBOOST_net_622) );
oa22m02 FE_RC_923_0 ( .a(n_7399), .b(FE_OCP_RBN5693_n_8138), .c(n_7400), .d(n_8138), .o(n_8242) );
oa22f04 FE_RC_925_0 ( .a(n_6465), .b(n_6576), .c(n_6466), .d(n_47335), .o(n_6774) );
oa22s04 FE_RC_926_0 ( .a(n_11739), .b(n_11959), .c(n_11740), .d(n_11985), .o(n_12196) );
oa22s02 FE_RC_929_0 ( .a(FE_OFN787_n_46285), .b(n_12114), .c(FE_OCP_RBN3352_FE_OFN760_n_46337), .d(n_12037), .o(n_46357) );
in01s02 FE_RC_930_0 ( .a(n_24933), .o(FE_RN_294_0) );
in01s06 FE_RC_931_0 ( .a(n_25067), .o(FE_RN_295_0) );
no02s06 TIMEBOOST_cell_6866 ( .a(TIMEBOOST_net_2191), .b(n_37076), .o(n_37185) );
na02f04 TIMEBOOST_cell_5244 ( .a(FE_OCP_RBN2830_n_13962), .b(n_14592), .o(TIMEBOOST_net_1570) );
oa22s02 FE_RC_935_0 ( .a(FE_OFN4787_n_46137), .b(n_6479), .c(FE_OFN770_n_46196), .d(n_46993), .o(n_46181) );
ao22f02 FE_RC_936_0 ( .a(FE_OCP_RBN4160_FE_OCPN857_n_7802), .b(FE_OCP_RBN2716_n_8242), .c(FE_OCP_RBN5647_FE_OCPN855_n_7721), .d(n_8242), .o(n_8335) );
ao22s06 FE_RC_940_0 ( .a(n_24375), .b(n_23967), .c(n_24407), .d(n_23968), .o(n_24506) );
oa22s06 FE_RC_942_0 ( .a(n_6328), .b(n_6347), .c(n_6358), .d(FE_OCP_RBN4488_n_6299), .o(n_6487) );
oa22m02 FE_RC_945_0 ( .a(n_7430), .b(n_8211), .c(n_7431), .d(n_8212), .o(n_8321) );
na02s06 TIMEBOOST_cell_3873 ( .a(n_28270), .b(n_28063), .o(TIMEBOOST_net_1027) );
in01s01 FE_RC_947_0 ( .a(n_47240), .o(FE_RN_298_0) );
na02m06 TIMEBOOST_cell_3874 ( .a(TIMEBOOST_net_1027), .b(n_28271), .o(n_28295) );
oa22m02 FE_RC_951_0 ( .a(FE_OFN4787_n_46137), .b(n_6589), .c(n_6627), .d(FE_OFN770_n_46196), .o(n_46187) );
oa22m02 FE_RC_953_0 ( .a(FE_OFN4787_n_46137), .b(n_6618), .c(n_6648), .d(FE_OFN770_n_46196), .o(n_46188) );
na02s01 TIMEBOOST_cell_7898 ( .a(n_35932), .b(n_35931), .o(TIMEBOOST_net_2580) );
oa22f02 FE_RC_956_0 ( .a(n_46418), .b(n_8497), .c(n_8496), .d(n_8367), .o(n_8597) );
oa22f04 FE_RC_966_0 ( .a(n_13321), .b(n_13838), .c(n_13320), .d(n_13812), .o(n_13960) );
ao22s02 FE_RC_970_0 ( .a(n_17389), .b(n_17694), .c(n_17324), .d(n_17659), .o(n_17729) );
ao22m02 FE_RC_971_0 ( .a(n_8567), .b(FE_OCP_RBN2810_n_8542), .c(n_8566), .d(FE_OCP_RBN2811_n_8542), .o(n_8687) );
ao22f02 FE_RC_973_0 ( .a(FE_OCPN935_n_7802), .b(FE_OCP_RBN5749_n_8599), .c(FE_OCP_RBN4139_n_7743), .d(n_8599), .o(n_8727) );
ao22m02 FE_RC_975_0 ( .a(FE_OCP_RBN5653_n_2438), .b(n_3673), .c(FE_OCP_RBN5649_n_2438), .d(n_3155), .o(n_3189) );
oa22s01 FE_RC_977_0 ( .a(n_17584), .b(n_17835), .c(n_16339), .d(n_47195), .o(n_17880) );
oa22s01 FE_RC_978_0 ( .a(n_17336), .b(n_17812), .c(n_16339), .d(n_17809), .o(n_17879) );
oa22m02 FE_RC_97_0 ( .a(FE_OFN4787_n_46137), .b(n_6700), .c(FE_OFN770_n_46196), .d(n_6739), .o(n_46191) );
oa22m04 FE_RC_980_0 ( .a(n_9493), .b(n_9574), .c(n_9476), .d(n_9573), .o(n_9724) );
oa22m04 FE_RC_984_0 ( .a(n_11748), .b(n_11953), .c(n_11952), .d(n_11747), .o(n_12145) );
oa22m02 FE_RC_985_0 ( .a(FE_OCP_RBN6865_n_46285), .b(n_12131), .c(FE_OFN765_n_46337), .d(n_12060), .o(n_46355) );
oa22m02 FE_RC_986_0 ( .a(FE_OCP_RBN6865_n_46285), .b(n_12068), .c(FE_OFN765_n_46337), .d(n_12064), .o(n_46354) );
oa22m04 FE_RC_989_0 ( .a(n_37574), .b(n_37689), .c(n_37556), .d(n_37755), .o(n_37771) );
no02s01 TIMEBOOST_cell_3122 ( .a(FE_OCPN4857_n_14317), .b(n_15250), .o(TIMEBOOST_net_852) );
in01s01 FE_RC_993_0 ( .a(n_3039), .o(FE_RN_303_0) );
in01s01 FE_RC_994_0 ( .a(n_2604), .o(FE_RN_304_0) );
no02s01 TIMEBOOST_cell_4224 ( .a(TIMEBOOST_net_1202), .b(n_33474), .o(n_33059) );
na02f08 TIMEBOOST_cell_5098 ( .a(FE_OCP_RBN4153_n_29378), .b(FE_OFN773_n_25834), .o(TIMEBOOST_net_1497) );
ao22m02 FE_RC_997_0 ( .a(n_2594), .b(FE_OCP_RBN4212_n_3343), .c(n_3343), .d(n_2595), .o(n_3421) );
na02s04 FE_RC_998_0 ( .a(n_33213), .b(n_33787), .o(FE_RN_306_0) );
in01f04 FE_RC_999_0 ( .a(n_33810), .o(FE_RN_307_0) );
in01m03 FE_RC_9_0 ( .a(n_18052), .o(FE_RN_3_0) );
ms00f80 cos_out_reg_0_ ( .ck(ispd_clk), .d(n_43154), .o(cos_out_0) );
ms00f80 cos_out_reg_10_ ( .ck(ispd_clk), .d(n_43766), .o(cos_out_10) );
ms00f80 cos_out_reg_11_ ( .ck(ispd_clk), .d(n_43797), .o(cos_out_11) );
ms00f80 cos_out_reg_12_ ( .ck(ispd_clk), .d(n_43776), .o(cos_out_12) );
ms00f80 cos_out_reg_13_ ( .ck(ispd_clk), .d(n_43796), .o(cos_out_13) );
ms00f80 cos_out_reg_14_ ( .ck(ispd_clk), .d(n_43818), .o(cos_out_14) );
ms00f80 cos_out_reg_15_ ( .ck(ispd_clk), .d(n_43850), .o(cos_out_15) );
ms00f80 cos_out_reg_16_ ( .ck(ispd_clk), .d(n_43817), .o(cos_out_16) );
ms00f80 cos_out_reg_17_ ( .ck(ispd_clk), .d(n_43852), .o(cos_out_17) );
ms00f80 cos_out_reg_18_ ( .ck(ispd_clk), .d(n_43851), .o(cos_out_18) );
ms00f80 cos_out_reg_19_ ( .ck(ispd_clk), .d(n_43844), .o(cos_out_19) );
ms00f80 cos_out_reg_1_ ( .ck(ispd_clk), .d(n_43288), .o(cos_out_1) );
ms00f80 cos_out_reg_20_ ( .ck(ispd_clk), .d(n_43860), .o(cos_out_20) );
ms00f80 cos_out_reg_21_ ( .ck(ispd_clk), .d(n_43865), .o(cos_out_21) );
ms00f80 cos_out_reg_22_ ( .ck(ispd_clk), .d(n_43870), .o(cos_out_22) );
ms00f80 cos_out_reg_23_ ( .ck(ispd_clk), .d(n_43869), .o(cos_out_23) );
ms00f80 cos_out_reg_24_ ( .ck(ispd_clk), .d(n_43884), .o(cos_out_24) );
ms00f80 cos_out_reg_25_ ( .ck(ispd_clk), .d(n_43886), .o(cos_out_25) );
ms00f80 cos_out_reg_26_ ( .ck(ispd_clk), .d(n_43891), .o(cos_out_26) );
ms00f80 cos_out_reg_27_ ( .ck(ispd_clk), .d(n_43909), .o(cos_out_27) );
ms00f80 cos_out_reg_28_ ( .ck(ispd_clk), .d(n_43904), .o(cos_out_28) );
ms00f80 cos_out_reg_29_ ( .ck(ispd_clk), .d(n_43897), .o(cos_out_29) );
ms00f80 cos_out_reg_2_ ( .ck(ispd_clk), .d(n_43381), .o(cos_out_2) );
ms00f80 cos_out_reg_30_ ( .ck(ispd_clk), .d(n_43906), .o(cos_out_30) );
ms00f80 cos_out_reg_31_ ( .ck(ispd_clk), .d(n_43905), .o(cos_out_31) );
ms00f80 cos_out_reg_3_ ( .ck(ispd_clk), .d(n_43693), .o(cos_out_3) );
ms00f80 cos_out_reg_4_ ( .ck(ispd_clk), .d(n_43694), .o(cos_out_4) );
ms00f80 cos_out_reg_5_ ( .ck(ispd_clk), .d(n_43695), .o(cos_out_5) );
ms00f80 cos_out_reg_6_ ( .ck(ispd_clk), .d(n_43688), .o(cos_out_6) );
ms00f80 cos_out_reg_7_ ( .ck(ispd_clk), .d(n_43702), .o(cos_out_7) );
ms00f80 cos_out_reg_8_ ( .ck(ispd_clk), .d(n_43738), .o(cos_out_8) );
ms00f80 cos_out_reg_9_ ( .ck(ispd_clk), .d(n_43767), .o(cos_out_9) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_14740), .o(delay_add_ln22_unr11_stage5_stallmux_q_0_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N1506_n_16183), .o(delay_add_ln22_unr11_stage5_stallmux_q_10_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_16425), .o(delay_add_ln22_unr11_stage5_stallmux_q_11_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_16602), .o(delay_add_ln22_unr11_stage5_stallmux_q_12_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_46979), .o(delay_add_ln22_unr11_stage5_stallmux_q_13_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_16686), .o(delay_add_ln22_unr11_stage5_stallmux_q_14_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_46977), .o(delay_add_ln22_unr11_stage5_stallmux_q_15_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_16810), .o(delay_add_ln22_unr11_stage5_stallmux_q_16_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_16916), .o(delay_add_ln22_unr11_stage5_stallmux_q_17_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_46974), .o(delay_add_ln22_unr11_stage5_stallmux_q_18_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_17199), .o(delay_add_ln22_unr11_stage5_stallmux_q_19_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_15033), .o(delay_add_ln22_unr11_stage5_stallmux_q_1_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_17294), .o(delay_add_ln22_unr11_stage5_stallmux_q_20_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_17460), .o(delay_add_ln22_unr11_stage5_stallmux_q_21_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_17594), .o(delay_add_ln22_unr11_stage5_stallmux_q_22_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_17630), .o(delay_add_ln22_unr11_stage5_stallmux_q_23_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_17728), .o(delay_add_ln22_unr11_stage5_stallmux_q_24_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_17759), .o(delay_add_ln22_unr11_stage5_stallmux_q_25_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_17782), .o(delay_add_ln22_unr11_stage5_stallmux_q_26_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_17811), .o(delay_add_ln22_unr11_stage5_stallmux_q_27_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_44447), .o(delay_add_ln22_unr11_stage5_stallmux_q_28_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_17835), .o(delay_add_ln22_unr11_stage5_stallmux_q_29_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_15221), .o(delay_add_ln22_unr11_stage5_stallmux_q_2_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_17812), .o(delay_add_ln22_unr11_stage5_stallmux_q_30_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_17834), .o(delay_add_ln22_unr11_stage5_stallmux_q_31_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_15303), .o(delay_add_ln22_unr11_stage5_stallmux_q_3_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_15489), .o(delay_add_ln22_unr11_stage5_stallmux_q_4_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N1500_n_15605), .o(delay_add_ln22_unr11_stage5_stallmux_q_5_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_15751), .o(delay_add_ln22_unr11_stage5_stallmux_q_6_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_15757), .o(delay_add_ln22_unr11_stage5_stallmux_q_7_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N1502_n_15979), .o(delay_add_ln22_unr11_stage5_stallmux_q_8_) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N1504_n_16106), .o(delay_add_ln22_unr11_stage5_stallmux_q_9_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_20715), .o(delay_add_ln22_unr14_stage6_stallmux_q_0_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_21915), .o(delay_add_ln22_unr14_stage6_stallmux_q_10_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_21967), .o(delay_add_ln22_unr14_stage6_stallmux_q_11_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_22016), .o(delay_add_ln22_unr14_stage6_stallmux_q_12_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_22107), .o(delay_add_ln22_unr14_stage6_stallmux_q_13_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_22275), .o(delay_add_ln22_unr14_stage6_stallmux_q_14_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_22392), .o(delay_add_ln22_unr14_stage6_stallmux_q_15_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_22479), .o(delay_add_ln22_unr14_stage6_stallmux_q_16_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_22596), .o(delay_add_ln22_unr14_stage6_stallmux_q_17_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_22631), .o(delay_add_ln22_unr14_stage6_stallmux_q_18_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_22715), .o(delay_add_ln22_unr14_stage6_stallmux_q_19_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_21027), .o(delay_add_ln22_unr14_stage6_stallmux_q_1_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(FE_OCP_RBN6241_n_22622), .o(delay_add_ln22_unr14_stage6_stallmux_q_20_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_22750), .o(delay_add_ln22_unr14_stage6_stallmux_q_21_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(FE_OCP_RBN5051_n_22709), .o(delay_add_ln22_unr14_stage6_stallmux_q_22_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_22774), .o(delay_add_ln22_unr14_stage6_stallmux_q_23_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_22789), .o(delay_add_ln22_unr14_stage6_stallmux_q_24_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_22818), .o(delay_add_ln22_unr14_stage6_stallmux_q_25_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_22819), .o(delay_add_ln22_unr14_stage6_stallmux_q_26_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_22903), .o(delay_add_ln22_unr14_stage6_stallmux_q_27_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_22857), .o(delay_add_ln22_unr14_stage6_stallmux_q_28_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_22902), .o(delay_add_ln22_unr14_stage6_stallmux_q_29_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_21173), .o(delay_add_ln22_unr14_stage6_stallmux_q_2_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_22901), .o(delay_add_ln22_unr14_stage6_stallmux_q_30_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_22897), .o(delay_add_ln22_unr14_stage6_stallmux_q_31_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_21302), .o(delay_add_ln22_unr14_stage6_stallmux_q_3_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_21341), .o(delay_add_ln22_unr14_stage6_stallmux_q_4_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_21486), .o(delay_add_ln22_unr14_stage6_stallmux_q_5_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_21602), .o(delay_add_ln22_unr14_stage6_stallmux_q_6_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_21702), .o(delay_add_ln22_unr14_stage6_stallmux_q_7_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N5362_n_21732), .o(delay_add_ln22_unr14_stage6_stallmux_q_8_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N1518_n_21851), .o(delay_add_ln22_unr14_stage6_stallmux_q_9_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_26150), .o(delay_add_ln22_unr17_stage7_stallmux_q_0_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_27090), .o(delay_add_ln22_unr17_stage7_stallmux_q_10_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_27160), .o(delay_add_ln22_unr17_stage7_stallmux_q_11_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_27278), .o(delay_add_ln22_unr17_stage7_stallmux_q_12_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_27360), .o(delay_add_ln22_unr17_stage7_stallmux_q_13_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_27472), .o(delay_add_ln22_unr17_stage7_stallmux_q_14_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_27534), .o(delay_add_ln22_unr17_stage7_stallmux_q_15_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_27580), .o(delay_add_ln22_unr17_stage7_stallmux_q_16_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_27617), .o(delay_add_ln22_unr17_stage7_stallmux_q_17_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_27665), .o(delay_add_ln22_unr17_stage7_stallmux_q_18_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_27686), .o(delay_add_ln22_unr17_stage7_stallmux_q_19_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_26439), .o(delay_add_ln22_unr17_stage7_stallmux_q_1_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_27714), .o(delay_add_ln22_unr17_stage7_stallmux_q_20_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_27728), .o(delay_add_ln22_unr17_stage7_stallmux_q_21_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_27727), .o(delay_add_ln22_unr17_stage7_stallmux_q_22_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_27726), .o(delay_add_ln22_unr17_stage7_stallmux_q_23_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(FE_OCP_RBN6258_n_27743), .o(delay_add_ln22_unr17_stage7_stallmux_q_24_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_27800), .o(delay_add_ln22_unr17_stage7_stallmux_q_25_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_27772), .o(delay_add_ln22_unr17_stage7_stallmux_q_26_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_27835), .o(delay_add_ln22_unr17_stage7_stallmux_q_27_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_27771), .o(delay_add_ln22_unr17_stage7_stallmux_q_28_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_27805), .o(delay_add_ln22_unr17_stage7_stallmux_q_29_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_26477), .o(delay_add_ln22_unr17_stage7_stallmux_q_2_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_27804), .o(delay_add_ln22_unr17_stage7_stallmux_q_30_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_27799), .o(delay_add_ln22_unr17_stage7_stallmux_q_31_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_26536), .o(delay_add_ln22_unr17_stage7_stallmux_q_3_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_26668), .o(delay_add_ln22_unr17_stage7_stallmux_q_4_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_26731), .o(delay_add_ln22_unr17_stage7_stallmux_q_5_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_26810), .o(delay_add_ln22_unr17_stage7_stallmux_q_6_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_26881), .o(delay_add_ln22_unr17_stage7_stallmux_q_7_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_26969), .o(delay_add_ln22_unr17_stage7_stallmux_q_8_) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_27046), .o(delay_add_ln22_unr17_stage7_stallmux_q_9_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_30734), .o(delay_add_ln22_unr20_stage8_stallmux_q_0_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_31670), .o(delay_add_ln22_unr20_stage8_stallmux_q_10_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_31750), .o(delay_add_ln22_unr20_stage8_stallmux_q_11_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_31996), .o(delay_add_ln22_unr20_stage8_stallmux_q_12_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_31998), .o(delay_add_ln22_unr20_stage8_stallmux_q_13_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_31958), .o(delay_add_ln22_unr20_stage8_stallmux_q_14_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_31999), .o(delay_add_ln22_unr20_stage8_stallmux_q_15_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_32029), .o(delay_add_ln22_unr20_stage8_stallmux_q_16_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_32085), .o(delay_add_ln22_unr20_stage8_stallmux_q_17_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_32113), .o(delay_add_ln22_unr20_stage8_stallmux_q_18_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_32147), .o(delay_add_ln22_unr20_stage8_stallmux_q_19_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_31008), .o(delay_add_ln22_unr20_stage8_stallmux_q_1_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_32192), .o(delay_add_ln22_unr20_stage8_stallmux_q_20_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_32255), .o(delay_add_ln22_unr20_stage8_stallmux_q_21_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(FE_OCP_RBN3421_n_32254), .o(delay_add_ln22_unr20_stage8_stallmux_q_22_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_32311), .o(delay_add_ln22_unr20_stage8_stallmux_q_23_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(FE_OCP_RBN3432_n_32239), .o(delay_add_ln22_unr20_stage8_stallmux_q_24_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_32290), .o(delay_add_ln22_unr20_stage8_stallmux_q_25_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(FE_OCP_RBN3442_n_32266), .o(delay_add_ln22_unr20_stage8_stallmux_q_26_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_32340), .o(delay_add_ln22_unr20_stage8_stallmux_q_27_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_32305), .o(delay_add_ln22_unr20_stage8_stallmux_q_28_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_32339), .o(delay_add_ln22_unr20_stage8_stallmux_q_29_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_31051), .o(delay_add_ln22_unr20_stage8_stallmux_q_2_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_32338), .o(delay_add_ln22_unr20_stage8_stallmux_q_30_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_32310), .o(delay_add_ln22_unr20_stage8_stallmux_q_31_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_31110), .o(delay_add_ln22_unr20_stage8_stallmux_q_3_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_31182), .o(delay_add_ln22_unr20_stage8_stallmux_q_4_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_31267), .o(delay_add_ln22_unr20_stage8_stallmux_q_5_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_31363), .o(delay_add_ln22_unr20_stage8_stallmux_q_6_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_31405), .o(delay_add_ln22_unr20_stage8_stallmux_q_7_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_31470), .o(delay_add_ln22_unr20_stage8_stallmux_q_8_) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_31561), .o(delay_add_ln22_unr20_stage8_stallmux_q_9_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_35309), .o(delay_add_ln22_unr23_stage9_stallmux_q_0_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N1510_n_36387), .o(delay_add_ln22_unr23_stage9_stallmux_q_10_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_36421), .o(delay_add_ln22_unr23_stage9_stallmux_q_11_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_36388), .o(delay_add_ln22_unr23_stage9_stallmux_q_12_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_36422), .o(delay_add_ln22_unr23_stage9_stallmux_q_13_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_36310), .o(delay_add_ln22_unr23_stage9_stallmux_q_14_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_36423), .o(delay_add_ln22_unr23_stage9_stallmux_q_15_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_36407), .o(delay_add_ln22_unr23_stage9_stallmux_q_16_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_36440), .o(delay_add_ln22_unr23_stage9_stallmux_q_17_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_36455), .o(delay_add_ln22_unr23_stage9_stallmux_q_18_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_36469), .o(delay_add_ln22_unr23_stage9_stallmux_q_19_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_35409), .o(delay_add_ln22_unr23_stage9_stallmux_q_1_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(FE_OFN5081_n_36439), .o(delay_add_ln22_unr23_stage9_stallmux_q_20_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_36430), .o(delay_add_ln22_unr23_stage9_stallmux_q_21_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_36468), .o(delay_add_ln22_unr23_stage9_stallmux_q_22_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_36487), .o(delay_add_ln22_unr23_stage9_stallmux_q_23_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_36544), .o(delay_add_ln22_unr23_stage9_stallmux_q_24_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_36549), .o(delay_add_ln22_unr23_stage9_stallmux_q_25_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_36581), .o(delay_add_ln22_unr23_stage9_stallmux_q_26_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_36632), .o(delay_add_ln22_unr23_stage9_stallmux_q_27_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_36608), .o(delay_add_ln22_unr23_stage9_stallmux_q_28_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_36651), .o(delay_add_ln22_unr23_stage9_stallmux_q_29_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_35464), .o(delay_add_ln22_unr23_stage9_stallmux_q_2_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_36669), .o(delay_add_ln22_unr23_stage9_stallmux_q_30_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_36629), .o(delay_add_ln22_unr23_stage9_stallmux_q_31_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_35481), .o(delay_add_ln22_unr23_stage9_stallmux_q_3_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_35518), .o(delay_add_ln22_unr23_stage9_stallmux_q_4_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_35592), .o(delay_add_ln22_unr23_stage9_stallmux_q_5_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_35705), .o(delay_add_ln22_unr23_stage9_stallmux_q_6_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_35791), .o(delay_add_ln22_unr23_stage9_stallmux_q_7_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_35874), .o(delay_add_ln22_unr23_stage9_stallmux_q_8_) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_35990), .o(delay_add_ln22_unr23_stage9_stallmux_q_9_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_39708), .o(delay_add_ln22_unr27_stage10_stallmux_q_0_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_40419), .o(delay_add_ln22_unr27_stage10_stallmux_q_10_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_40452), .o(delay_add_ln22_unr27_stage10_stallmux_q_11_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_40441), .o(delay_add_ln22_unr27_stage10_stallmux_q_12_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_40459), .o(delay_add_ln22_unr27_stage10_stallmux_q_13_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_40458), .o(delay_add_ln22_unr27_stage10_stallmux_q_14_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_40469), .o(delay_add_ln22_unr27_stage10_stallmux_q_15_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_40457), .o(delay_add_ln22_unr27_stage10_stallmux_q_16_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_40490), .o(delay_add_ln22_unr27_stage10_stallmux_q_17_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_40489), .o(delay_add_ln22_unr27_stage10_stallmux_q_18_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_40488), .o(delay_add_ln22_unr27_stage10_stallmux_q_19_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_39786), .o(delay_add_ln22_unr27_stage10_stallmux_q_1_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_40487), .o(delay_add_ln22_unr27_stage10_stallmux_q_20_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_40486), .o(delay_add_ln22_unr27_stage10_stallmux_q_21_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_40512), .o(delay_add_ln22_unr27_stage10_stallmux_q_22_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_40530), .o(delay_add_ln22_unr27_stage10_stallmux_q_23_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_40549), .o(delay_add_ln22_unr27_stage10_stallmux_q_24_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_40560), .o(delay_add_ln22_unr27_stage10_stallmux_q_25_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_40559), .o(delay_add_ln22_unr27_stage10_stallmux_q_26_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_40567), .o(delay_add_ln22_unr27_stage10_stallmux_q_27_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_40585), .o(delay_add_ln22_unr27_stage10_stallmux_q_28_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_40593), .o(delay_add_ln22_unr27_stage10_stallmux_q_29_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_39855), .o(delay_add_ln22_unr27_stage10_stallmux_q_2_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(FE_OCP_RBN6236_n_40586), .o(delay_add_ln22_unr27_stage10_stallmux_q_30_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_40592), .o(delay_add_ln22_unr27_stage10_stallmux_q_31_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_39896), .o(delay_add_ln22_unr27_stage10_stallmux_q_3_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_39986), .o(delay_add_ln22_unr27_stage10_stallmux_q_4_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_40161), .o(delay_add_ln22_unr27_stage10_stallmux_q_5_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_40427), .o(delay_add_ln22_unr27_stage10_stallmux_q_6_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_40439), .o(delay_add_ln22_unr27_stage10_stallmux_q_7_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_40428), .o(delay_add_ln22_unr27_stage10_stallmux_q_8_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_40440), .o(delay_add_ln22_unr27_stage10_stallmux_q_9_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_1134), .o(delay_add_ln22_unr2_stage2_stallmux_q_10_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_1163), .o(delay_add_ln22_unr2_stage2_stallmux_q_11_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_1137), .o(delay_add_ln22_unr2_stage2_stallmux_q_12_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_1169), .o(delay_add_ln22_unr2_stage2_stallmux_q_13_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_1164), .o(delay_add_ln22_unr2_stage2_stallmux_q_14_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2931), .o(delay_add_ln22_unr2_stage2_stallmux_q_15_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_973), .o(delay_add_ln22_unr2_stage2_stallmux_q_16_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_1025), .o(delay_add_ln22_unr2_stage2_stallmux_q_17_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_1001), .o(delay_add_ln22_unr2_stage2_stallmux_q_18_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2933), .o(delay_add_ln22_unr2_stage2_stallmux_q_19_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_1122), .o(delay_add_ln22_unr2_stage2_stallmux_q_1_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_1102), .o(delay_add_ln22_unr2_stage2_stallmux_q_20_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_1168), .o(delay_add_ln22_unr2_stage2_stallmux_q_21_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2935), .o(delay_add_ln22_unr2_stage2_stallmux_q_22_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_1205), .o(delay_add_ln22_unr2_stage2_stallmux_q_23_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_1190), .o(delay_add_ln22_unr2_stage2_stallmux_q_24_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2937), .o(delay_add_ln22_unr2_stage2_stallmux_q_25_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2939), .o(delay_add_ln22_unr2_stage2_stallmux_q_26_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_1217), .o(delay_add_ln22_unr2_stage2_stallmux_q_27_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_1066), .o(delay_add_ln22_unr2_stage2_stallmux_q_28_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_1124), .o(delay_add_ln22_unr2_stage2_stallmux_q_29_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_835), .o(delay_add_ln22_unr2_stage2_stallmux_q_2_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2941), .o(delay_add_ln22_unr2_stage2_stallmux_q_30_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_1118), .o(delay_add_ln22_unr2_stage2_stallmux_q_31_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_966), .o(delay_add_ln22_unr2_stage2_stallmux_q_3_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_958), .o(delay_add_ln22_unr2_stage2_stallmux_q_4_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_1010), .o(delay_add_ln22_unr2_stage2_stallmux_q_5_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_886), .o(delay_add_ln22_unr2_stage2_stallmux_q_6_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_1018), .o(delay_add_ln22_unr2_stage2_stallmux_q_7_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_1019), .o(delay_add_ln22_unr2_stage2_stallmux_q_8_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_1129), .o(delay_add_ln22_unr2_stage2_stallmux_q_9_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_4180), .o(delay_add_ln22_unr5_stage3_stallmux_q_0_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_5569), .o(delay_add_ln22_unr5_stage3_stallmux_q_10_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_5645), .o(delay_add_ln22_unr5_stage3_stallmux_q_11_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_5724), .o(delay_add_ln22_unr5_stage3_stallmux_q_12_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_5840), .o(delay_add_ln22_unr5_stage3_stallmux_q_13_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_5972), .o(delay_add_ln22_unr5_stage3_stallmux_q_14_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_6047), .o(delay_add_ln22_unr5_stage3_stallmux_q_15_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_6063), .o(delay_add_ln22_unr5_stage3_stallmux_q_16_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_6154), .o(delay_add_ln22_unr5_stage3_stallmux_q_17_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_6233), .o(delay_add_ln22_unr5_stage3_stallmux_q_18_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_6297), .o(delay_add_ln22_unr5_stage3_stallmux_q_19_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_4491), .o(delay_add_ln22_unr5_stage3_stallmux_q_1_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_6267), .o(delay_add_ln22_unr5_stage3_stallmux_q_20_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_6313), .o(delay_add_ln22_unr5_stage3_stallmux_q_21_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_46994), .o(delay_add_ln22_unr5_stage3_stallmux_q_22_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_6376), .o(delay_add_ln22_unr5_stage3_stallmux_q_23_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(FE_OCP_RBN3435_n_6379), .o(delay_add_ln22_unr5_stage3_stallmux_q_24_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_46993), .o(delay_add_ln22_unr5_stage3_stallmux_q_25_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(FE_OCP_RBN6247_n_6477), .o(delay_add_ln22_unr5_stage3_stallmux_q_26_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_6529), .o(delay_add_ln22_unr5_stage3_stallmux_q_27_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(FE_OCP_RBN6250_n_6567), .o(delay_add_ln22_unr5_stage3_stallmux_q_28_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_6627), .o(delay_add_ln22_unr5_stage3_stallmux_q_29_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_4623), .o(delay_add_ln22_unr5_stage3_stallmux_q_2_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_6648), .o(delay_add_ln22_unr5_stage3_stallmux_q_30_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_6720), .o(delay_add_ln22_unr5_stage3_stallmux_q_31_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_4679), .o(delay_add_ln22_unr5_stage3_stallmux_q_3_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_4828), .o(delay_add_ln22_unr5_stage3_stallmux_q_4_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_4997), .o(delay_add_ln22_unr5_stage3_stallmux_q_5_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_5273), .o(delay_add_ln22_unr5_stage3_stallmux_q_6_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_5323), .o(delay_add_ln22_unr5_stage3_stallmux_q_7_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_5379), .o(delay_add_ln22_unr5_stage3_stallmux_q_8_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_5483), .o(delay_add_ln22_unr5_stage3_stallmux_q_9_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_9474), .o(delay_add_ln22_unr8_stage4_stallmux_q_0_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_10739), .o(delay_add_ln22_unr8_stage4_stallmux_q_10_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_10885), .o(delay_add_ln22_unr8_stage4_stallmux_q_11_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_10959), .o(delay_add_ln22_unr8_stage4_stallmux_q_12_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_11098), .o(delay_add_ln22_unr8_stage4_stallmux_q_13_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_11177), .o(delay_add_ln22_unr8_stage4_stallmux_q_14_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_11252), .o(delay_add_ln22_unr8_stage4_stallmux_q_15_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_11297), .o(delay_add_ln22_unr8_stage4_stallmux_q_16_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_11356), .o(delay_add_ln22_unr8_stage4_stallmux_q_17_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_11411), .o(delay_add_ln22_unr8_stage4_stallmux_q_18_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_11453), .o(delay_add_ln22_unr8_stage4_stallmux_q_19_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_9760), .o(delay_add_ln22_unr8_stage4_stallmux_q_1_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_11605), .o(delay_add_ln22_unr8_stage4_stallmux_q_20_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_11759), .o(delay_add_ln22_unr8_stage4_stallmux_q_21_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_11856), .o(delay_add_ln22_unr8_stage4_stallmux_q_22_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_11873), .o(delay_add_ln22_unr8_stage4_stallmux_q_23_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_12131), .o(delay_add_ln22_unr8_stage4_stallmux_q_24_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_12068), .o(delay_add_ln22_unr8_stage4_stallmux_q_25_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_12158), .o(delay_add_ln22_unr8_stage4_stallmux_q_26_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_12145), .o(delay_add_ln22_unr8_stage4_stallmux_q_27_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(FE_OCP_RBN6252_n_12067), .o(delay_add_ln22_unr8_stage4_stallmux_q_28_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_12212), .o(delay_add_ln22_unr8_stage4_stallmux_q_29_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_9842), .o(delay_add_ln22_unr8_stage4_stallmux_q_2_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_12211), .o(delay_add_ln22_unr8_stage4_stallmux_q_30_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_12240), .o(delay_add_ln22_unr8_stage4_stallmux_q_31_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_10000), .o(delay_add_ln22_unr8_stage4_stallmux_q_3_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_10088), .o(delay_add_ln22_unr8_stage4_stallmux_q_4_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_10222), .o(delay_add_ln22_unr8_stage4_stallmux_q_5_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_10392), .o(delay_add_ln22_unr8_stage4_stallmux_q_6_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_10496), .o(delay_add_ln22_unr8_stage4_stallmux_q_7_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_10530), .o(delay_add_ln22_unr8_stage4_stallmux_q_8_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_10705), .o(delay_add_ln22_unr8_stage4_stallmux_q_9_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_14732), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_0_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_16212), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_10_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_16362), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_11_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_16575), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_12_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_16601), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_13_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_16699), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_14_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_16757), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_15_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_46976), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_16_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_46975), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_17_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_17128), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_18_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_46973), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_19_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_15065), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_1_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_17440), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_17459), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_17550), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_22_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_17591), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_23_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(FE_OCP_RBN6246_n_17587), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_24_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_17686), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_17685), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_26_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_17697), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_27_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_17688), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_28_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_17723), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_29_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_15168), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_2_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_17725), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_30_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_17687), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_31_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_15406), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_3_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_15488), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_4_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_15603), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_5_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_15722), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_6_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_15842), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_7_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_15978), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_8_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_16105), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_9_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_20378), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_0_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_21920), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_10_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_21969), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_11_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_22044), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_12_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_22112), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_13_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_22236), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_14_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_22359), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_15_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_22425), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_16_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_22540), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_46965), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_18_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_22640), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_19_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_20970), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_1_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_22635), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_20_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_22684), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_22718), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_22_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_22778), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_23_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(FE_OCP_RBN3451_n_22710), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_24_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_22806), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_25_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_22829), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_26_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_22914), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_27_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(FE_OCP_RBN4492_n_22755), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_28_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_22875), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_29_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_21066), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_2_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_22874), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_30_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_22835), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_31_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_21124), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_3_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_21276), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_4_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_21426), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_5_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_21541), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_6_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_21613), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_7_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N1516_n_21706), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_8_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_21810), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_9_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_26111), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_0_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_27059), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_10_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_27129), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_11_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_27279), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_12_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_27365), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_13_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_27364), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_14_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_27443), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_15_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_27576), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_27584), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_27622), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_18_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_27643), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_19_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_26365), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_1_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_27653), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_20_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_27655), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_21_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_27693), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_22_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_27720), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_23_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_27768), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_24_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_27782), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_25_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_27739), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_26_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_27785), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_27_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_27755), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_28_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_27784), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_29_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N1508_n_26491), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_2_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_27783), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_30_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_27781), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_31_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N1512_n_26582), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_3_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_26693), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_4_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N1520_n_26761), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_5_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N1522_n_26807), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_6_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_26853), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_7_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_26968), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_8_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_27029), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_9_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_30813), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_31878), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_10_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_31955), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_11_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_32251), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_12_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_32252), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_13_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_32234), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_14_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_32259), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_15_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_32235), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_32263), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_17_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_32262), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_18_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_32281), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_19_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_31176), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_32325), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_20_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_32384), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_21_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_32428), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_22_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_32471), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_23_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_32463), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_24_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_32517), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_25_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(FE_OCP_RBN5058_n_32427), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_26_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_32546), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_27_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_32468), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_28_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_32518), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_29_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_31193), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_2_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_32519), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_32516), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_31_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_31326), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_3_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_31397), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_4_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(FE_OCP_DRV_N1524_n_31435), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_5_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_31514), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_6_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_31673), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_7_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_31715), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_8_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_31806), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_9_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_35210), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_0_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_36337), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_10_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_36389), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_11_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_36340), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_12_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_36371), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_13_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_36345), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_14_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_36396), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_15_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_36377), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_36415), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_36442), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_18_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_36460), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_19_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_35378), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_1_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_36414), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_20_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_36433), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_21_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_36432), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_22_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_36449), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_23_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(FE_OCP_RBN1872_n_36489), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_24_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_36520), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_25_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_36569), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_26_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_36594), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_27_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_36553), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_28_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_36592), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_29_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_35419), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_2_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_36615), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_30_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_36567), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_31_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_35426), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_3_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_35474), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_4_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_35507), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_5_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_35557), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_6_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_35626), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_7_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_35757), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_35922), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_39716), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_0_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_40350), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_10_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_40404), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_11_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_40403), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_12_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_40421), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_13_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_40385), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_14_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_40405), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_15_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_40433), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_40465), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_17_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_40464), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_18_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_40477), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_19_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_39779), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_1_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_40498), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_20_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_40507), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_21_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_40506), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_22_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_40525), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_23_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_40544), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_24_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_40554), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_25_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_40553), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_26_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_40552), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_27_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_40576), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_28_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_40577), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_29_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_39847), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_2_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_40578), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_30_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_40579), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_31_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_39848), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_3_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_39958), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_40410), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_5_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_40198), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_6_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_40416), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_7_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_40411), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_40420), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_46055), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_0_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_990), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_10_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_1099), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_12_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(FE_OFN759_n_45813), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_13_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_938), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_15_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_1022), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_16_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_1040), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_17_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_1092), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_18_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_1132), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_19_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_1007), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_1_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_1127), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_20_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_1152), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_21_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_1144), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_22_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_1165), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_23_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_1005), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_24_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_1048), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_25_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_981), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_26_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2943), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_27_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(FE_OFN4811_n_902), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_28_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2945), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_29_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_1021), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_2_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_1167), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_3_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(FE_OFN4818_n_920), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_4_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_1017), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_5_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_934), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_6_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_1004), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_7_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_928), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_8_) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_934), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_9_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_4157), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_0_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_5618), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_10_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_5748), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_11_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_5841), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_12_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_5913), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_13_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_5971), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_14_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_46997), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_15_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_6105), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_16_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_6146), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_17_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_46995), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_18_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_6243), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_19_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_4600), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_1_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_6248), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_20_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_6301), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_21_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_6419), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_22_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_6476), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_23_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_6435), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_24_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_6500), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_25_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(FE_OCP_RBN3455_n_6557), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_26_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_6643), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_27_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_6670), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_6719), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_4590), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_2_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_6739), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_30_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_6774), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_31_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_4793), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_3_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_4857), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_4_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_4992), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_5_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_5244), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_6_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_5363), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_7_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_5408), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_8_) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_5527), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_9_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_9428), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_0_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_10783), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_10_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_10848), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_11_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_46988), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_12_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_11061), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_13_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_11212), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_14_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_11278), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_15_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_11307), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_16_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_11369), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_17_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_46986), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_18_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_11494), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_19_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_9878), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_1_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_11490), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_20_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_11655), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_21_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_11731), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_22_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_11778), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_23_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_12150), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_24_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_12144), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_25_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_12117), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_26_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_12217), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_27_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_12114), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_28_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_12196), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_29_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_9916), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_2_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_12197), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_30_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_12162), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_31_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_9958), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_3_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_10085), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_4_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_10213), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_5_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_10389), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_6_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_10490), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_7_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_10524), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_8_) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_10680), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_9_) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_36766), .o(delay_sub_ln21_unr24_stage9_stallmux_q_1_) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_36776), .o(delay_sub_ln21_unr24_stage9_stallmux_q_2_) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_36830), .o(delay_sub_ln21_unr24_stage9_stallmux_q_3_) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_36829), .o(delay_sub_ln21_unr24_stage9_stallmux_q_4_) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_36866), .o(delay_sub_ln21_unr24_stage9_stallmux_q_5_) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_36885), .o(delay_sub_ln21_unr24_stage9_stallmux_q_6_) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_36895), .o(delay_sub_ln21_unr24_stage9_stallmux_q_7_) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_36896), .o(delay_sub_ln21_unr24_stage9_stallmux_q_8_) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_36658), .o(delay_sub_ln22_unr24_stage9_stallmux_q_0_) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_36741), .o(delay_sub_ln22_unr24_stage9_stallmux_q_1_) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_36782), .o(delay_sub_ln22_unr24_stage9_stallmux_q_2_) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_36792), .o(delay_sub_ln22_unr24_stage9_stallmux_q_3_) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_36800), .o(delay_sub_ln22_unr24_stage9_stallmux_q_4_) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_36845), .o(delay_sub_ln22_unr24_stage9_stallmux_q_5_) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_36874), .o(delay_sub_ln22_unr24_stage9_stallmux_q_6_) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_36890), .o(delay_sub_ln22_unr24_stage9_stallmux_q_7_) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_36891), .o(n_46254) );
ms00f80 delay_sub_ln23_0_unr11_stage5_stallmux_q_reg ( .ck(ispd_clk), .d(FE_OCP_RBN3197_n_15599), .o(n_44365) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(FE_OCP_RBN5394_cordic_combinational_sub_ln23_0_unr12_z_0_), .o(cordic_combinational_sub_ln23_0_unr16_z_0_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_16550), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_10_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_16593), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_11_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_16592), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_12_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_16616), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_13_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_16721), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_14_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_16744), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_15_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_16767), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_16_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_16815), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_17_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_16847), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_18_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_16926), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_19_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_16409), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_1_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_16846), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_20_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_16925), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_21_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_16927), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_22_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_16924), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_23_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_16849), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_24_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_16967), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_25_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_17017), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_26_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_17058), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_27_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_17014), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_28_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_17103), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_29_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_16408), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_2_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_17102), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_30_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_16888), .o(n_17093) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_16410), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_3_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_16411), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_4_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_16412), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_5_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_16413), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_6_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_16414), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_7_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_16523), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_8_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_16549), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_) );
ms00f80 delay_sub_ln23_0_unr14_stage6_stallmux_q_reg ( .ck(ispd_clk), .d(n_20252), .o(n_44061) );
ms00f80 delay_sub_ln23_0_unr15_stage6_stallmux_q_reg ( .ck(ispd_clk), .d(n_21691), .o(delay_sub_ln23_0_unr15_stage6_stallmux_q) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(cordic_combinational_sub_ln23_0_unr20_z_0_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_22115), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_10_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_22116), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_11_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_22031), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_12_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_22118), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_13_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_22144), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_14_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_22245), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_15_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_22244), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_16_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_22362), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_17_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_22361), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_18_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_22398), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_19_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_21338), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_22521), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_20_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_22567), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_21_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_22522), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_22_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_22568), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_23_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_22545), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_24_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_22587), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_25_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_22548), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_26_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_22588), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_27_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_22606), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_28_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_22659), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_29_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_21929), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_2_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_22689), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_30_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_22550), .o(n_22641) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_21930), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_3_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_21931), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_4_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_21932), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_5_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_21802), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_6_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_21933), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_7_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_21994), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_8_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_22055), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_9_) );
ms00f80 delay_sub_ln23_0_unr17_stage7_stallmux_q_reg ( .ck(ispd_clk), .d(n_24188), .o(n_44722) );
ms00f80 delay_sub_ln23_0_unr18_stage7_stallmux_q_reg ( .ck(ispd_clk), .d(n_25160), .o(n_25834) );
ms00f80 delay_sub_ln23_0_unr19_stage7_stallmux_q_reg ( .ck(ispd_clk), .d(n_26896), .o(n_27014) );
ms00f80 delay_sub_ln23_0_unr1_stage2_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_50), .o(delay_sub_ln23_0_unr1_stage2_stallmux_q_0_) );
ms00f80 delay_sub_ln23_0_unr1_stage2_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_600), .o(delay_sub_ln23_0_unr1_stage2_stallmux_q_1_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_186) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_27016), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_10_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_27094), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_11_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_27015), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_27093), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_27092), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_14_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_27134), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_15_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_27107), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_27165), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_27200), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_18_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_27247), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_19_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_26997), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_1_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_27318), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_20_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_27323), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_21_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_27448), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_22_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_27479), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_23_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_27447), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_24_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_27539), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_25_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_27574), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_26_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_27588), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_27_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_27625), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_28_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_27656), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_29_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_26996), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_2_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_27676), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_30_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_27678), .o(n_27923) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_26998), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_3_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_26999), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_4_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_27000), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_5_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_26796), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_6_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_26973), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_7_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_27001), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_8_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_27002), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_9_) );
ms00f80 delay_sub_ln23_0_unr20_stage8_stallmux_q_reg ( .ck(ispd_clk), .d(FE_OFN622_n_28336), .o(n_44962) );
ms00f80 delay_sub_ln23_0_unr21_stage8_stallmux_q_reg ( .ck(ispd_clk), .d(n_28897), .o(delay_sub_ln23_0_unr21_stage8_stallmux_q) );
ms00f80 delay_sub_ln23_0_unr22_stage8_stallmux_q_reg ( .ck(ispd_clk), .d(n_30156), .o(delay_sub_ln23_0_unr22_stage8_stallmux_q) );
ms00f80 delay_sub_ln23_0_unr23_stage8_stallmux_q_reg ( .ck(ispd_clk), .d(n_31530), .o(delay_sub_ln23_0_unr23_stage8_stallmux_q) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_186), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_31976), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_10_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_32005), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_11_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_32004), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_12_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_32065), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_13_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_32064), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_14_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_32093), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_15_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_32173), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_32229), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_32247), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_18_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_32257), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_19_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_31226), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_1_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_32228), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_20_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_32258), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_21_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_32248), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_22_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_32274), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_23_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_32256), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_24_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_32294), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_25_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_32291), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_26_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_32342), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_27_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_32341), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_28_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_32379), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_29_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_31293), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_2_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_32378), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_30_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(n_32293), .o(delay_sub_ln23_unr25_stage8_stallmux_q_3_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_31689), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_31690), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_4_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_31691), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_5_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_31671), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_6_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_31779), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_7_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_31856), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_31960), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_) );
ms00f80 delay_sub_ln23_0_unr24_stage9_stallmux_q_reg ( .ck(ispd_clk), .d(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(delay_sub_ln23_0_unr24_stage9_stallmux_q) );
ms00f80 delay_sub_ln23_0_unr25_stage9_stallmux_q_reg ( .ck(ispd_clk), .d(n_33571), .o(delay_sub_ln23_0_unr25_stage9_stallmux_q) );
ms00f80 delay_sub_ln23_0_unr26_stage9_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(delay_sub_ln23_0_unr26_stage9_stallmux_q_0_) );
ms00f80 delay_sub_ln23_0_unr26_stage9_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_33337), .o(delay_sub_ln23_0_unr26_stage9_stallmux_q_1_) );
ms00f80 delay_sub_ln23_0_unr26_stage9_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_34666), .o(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_) );
ms00f80 delay_sub_ln23_0_unr27_stage10_stallmux_q_reg ( .ck(ispd_clk), .d(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n_44610) );
ms00f80 delay_sub_ln23_0_unr27_stage9_stallmux_q_reg ( .ck(ispd_clk), .d(FE_OCP_RBN3303_n_35539), .o(delay_sub_ln23_0_unr27_stage10_stallmux_z) );
ms00f80 delay_sub_ln23_0_unr28_stage10_stallmux_q_reg ( .ck(ispd_clk), .d(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(delay_sub_ln23_0_unr28_stage10_stallmux_q) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(FE_OFN231_n_35655), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_0_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_36453), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_10_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_36452), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_36496), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_36528), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_13_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_36527), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_36542), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_36573), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_36641), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_17_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_36640), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_18_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_36666), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_19_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_35726), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_1_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_36661), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_20_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_36699), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_21_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_36680), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_22_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_36714), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_36663), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_36700), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_25_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_36698), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_26_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_36729), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_27_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_36726), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_36728), .o(delay_sub_ln23_unr29_stage9_stallmux_q_2_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_36281), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_2_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_36282), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_36285), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_36330), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_5_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_36286), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_6_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_36384), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_7_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_36418), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_8_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_36454), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_9_) );
ms00f80 delay_sub_ln23_0_unr29_stage10_stallmux_q_reg ( .ck(ispd_clk), .d(n_45891), .o(delay_sub_ln23_0_unr29_stage10_stallmux_q) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_419), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_0_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_1082), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_10_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_1136), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_11_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_1166), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_12_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_1187), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_13_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_1207), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_14_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_1219), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_15_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_1224), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_16_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_1237), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_17_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_1234), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_18_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_1241), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_19_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_1140), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_1_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_1244), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_20_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_1249), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_21_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_1257), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_22_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_1261), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_23_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_1260), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_1273), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_25_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_1272), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_26_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_1274), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_27_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_1275), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_28_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_44624), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_729), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_738), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_3_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_740), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_4_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_1133), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_5_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_791), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_6_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_854), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_7_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_1112), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_8_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_1135), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_9_) );
ms00f80 delay_sub_ln23_0_unr30_stage10_stallmux_q_reg ( .ck(ispd_clk), .d(TIMEBOOST_net_2947), .o(delay_sub_ln23_0_unr30_stage10_stallmux_q) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_151), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_0_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_5211), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_10_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_5371), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_11_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_5399), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_12_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_5498), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_5578), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_5664), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_15_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_5753), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_16_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_5853), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_17_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_5929), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_18_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_5915), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_19_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_4031), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_5922), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_20_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_5992), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_21_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_6042), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_22_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_6159), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_23_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_6085), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_24_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_6183), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_25_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_6229), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_26_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_6286), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_27_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_6323), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_28_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_6384), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_29_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_4089), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_2_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(n_6405), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_30_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_31_ ( .ck(ispd_clk), .d(FE_OFN4789_n_46137), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_4192), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_4380), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_4_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_4526), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_5_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_4631), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_6_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_4775), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_7_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_4987), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_8_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_5151), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_9_) );
ms00f80 delay_sub_ln23_0_unr7_stage4_stallmux_q_reg ( .ck(ispd_clk), .d(n_167), .o(cordic_combinational_sub_ln23_0_unr12_z_0_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_9324), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_0_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_10301), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_10_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_10420), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_11_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_10549), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_12_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_10632), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_13_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_10652), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_14_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_10744), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_10717), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_10815), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_17_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_10840), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_18_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_10868), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_19_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_9437), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_1_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_10913), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_20_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_10981), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_21_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_11068), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_22_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_11153), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_23_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_11261), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_24_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_11286), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_25_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_11305), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_26_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_11344), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_27_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_11402), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_28_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_29_ ( .ck(ispd_clk), .d(n_11433), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_29_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_9518), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_2_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_30_ ( .ck(ispd_clk), .d(FE_OCP_RBN6166_n_46337), .o(n_45224) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_9653), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_9832), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_4_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_9957), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_5_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_9917), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_6_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_10044), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_10168), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_10295), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_9_) );
ms00f80 delay_sub_ln23_unr13_stage5_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_16887), .o(delay_sub_ln23_unr13_stage5_stallmux_q_1_) );
ms00f80 delay_sub_ln23_unr17_stage6_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_22549), .o(delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
ms00f80 delay_sub_ln23_unr21_stage7_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_27677), .o(delay_sub_ln23_unr21_stage7_stallmux_q_1_) );
ms00f80 delay_sub_ln23_unr25_stage8_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_32292), .o(delay_sub_ln23_unr25_stage8_stallmux_q_1_) );
ms00f80 delay_sub_ln23_unr9_stage4_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(FE_OCP_RBN6863_n_46285), .o(delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_16633), .o(n_44847) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_17654), .o(delay_xor_ln21_unr12_stage5_stallmux_q_10_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_17731), .o(delay_xor_ln21_unr12_stage5_stallmux_q_11_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_17777), .o(delay_xor_ln21_unr12_stage5_stallmux_q_12_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_17832), .o(delay_xor_ln21_unr12_stage5_stallmux_q_13_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_17829), .o(delay_xor_ln21_unr12_stage5_stallmux_q_14_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_17855), .o(delay_xor_ln21_unr12_stage5_stallmux_q_15_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_17808), .o(delay_xor_ln21_unr12_stage5_stallmux_q_16_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_17880), .o(delay_xor_ln21_unr12_stage5_stallmux_q_17_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_17879), .o(delay_xor_ln21_unr12_stage5_stallmux_q_18_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_17878), .o(delay_xor_ln21_unr12_stage5_stallmux_q_19_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_16700), .o(n_44721) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_16730), .o(delay_xor_ln21_unr12_stage5_stallmux_q_2_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_16789), .o(delay_xor_ln21_unr12_stage5_stallmux_q_3_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(FE_OFN4669_n_16873), .o(delay_xor_ln21_unr12_stage5_stallmux_q_4_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_17004), .o(delay_xor_ln21_unr12_stage5_stallmux_q_5_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_17144), .o(delay_xor_ln21_unr12_stage5_stallmux_q_6_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_17291), .o(delay_xor_ln21_unr12_stage5_stallmux_q_7_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_17418), .o(delay_xor_ln21_unr12_stage5_stallmux_q_8_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_17567), .o(delay_xor_ln21_unr12_stage5_stallmux_q_9_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_22449), .o(delay_xor_ln21_unr15_stage6_stallmux_q_0_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_22894), .o(delay_xor_ln21_unr15_stage6_stallmux_q_10_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_22893), .o(delay_xor_ln21_unr15_stage6_stallmux_q_11_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_22963), .o(delay_xor_ln21_unr15_stage6_stallmux_q_12_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_22892), .o(delay_xor_ln21_unr15_stage6_stallmux_q_13_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_22962), .o(delay_xor_ln21_unr15_stage6_stallmux_q_14_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_22960), .o(delay_xor_ln21_unr15_stage6_stallmux_q_15_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_22957), .o(delay_xor_ln21_unr15_stage6_stallmux_q_16_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_22535), .o(delay_xor_ln21_unr15_stage6_stallmux_q_1_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_22629), .o(delay_xor_ln21_unr15_stage6_stallmux_q_2_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_22704), .o(delay_xor_ln21_unr15_stage6_stallmux_q_3_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_22770), .o(delay_xor_ln21_unr15_stage6_stallmux_q_4_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_22742), .o(delay_xor_ln21_unr15_stage6_stallmux_q_5_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_22794), .o(delay_xor_ln21_unr15_stage6_stallmux_q_6_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_22766), .o(delay_xor_ln21_unr15_stage6_stallmux_q_7_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_22826), .o(delay_xor_ln21_unr15_stage6_stallmux_q_8_) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_22815), .o(delay_xor_ln21_unr15_stage6_stallmux_q_9_) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_27708), .o(n_44695) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_27819), .o(delay_xor_ln21_unr18_stage7_stallmux_q_10_) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_27863), .o(delay_xor_ln21_unr18_stage7_stallmux_q_11_) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_27862), .o(delay_xor_ln21_unr18_stage7_stallmux_q_12_) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_27855), .o(delay_xor_ln21_unr18_stage7_stallmux_q_13_) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_27725), .o(n_44422) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_27737), .o(delay_xor_ln21_unr18_stage7_stallmux_q_2_) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_27750), .o(delay_xor_ln21_unr18_stage7_stallmux_q_3_) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_27749), .o(n_45202) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_27748), .o(delay_xor_ln21_unr18_stage7_stallmux_q_5_) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_27815), .o(delay_xor_ln21_unr18_stage7_stallmux_q_6_) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_27858), .o(delay_xor_ln21_unr18_stage7_stallmux_q_7_) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_27818), .o(delay_xor_ln21_unr18_stage7_stallmux_q_8_) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_27894), .o(delay_xor_ln21_unr18_stage7_stallmux_q_9_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_32289), .o(delay_xor_ln21_unr21_stage8_stallmux_q_0_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_32353), .o(delay_xor_ln21_unr21_stage8_stallmux_q_10_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_32304), .o(delay_xor_ln21_unr21_stage8_stallmux_q_1_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_32352), .o(delay_xor_ln21_unr21_stage8_stallmux_q_2_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_32288), .o(delay_xor_ln21_unr21_stage8_stallmux_q_3_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_32337), .o(delay_xor_ln21_unr21_stage8_stallmux_q_4_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_32334), .o(delay_xor_ln21_unr21_stage8_stallmux_q_5_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_32374), .o(delay_xor_ln21_unr21_stage8_stallmux_q_6_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_32350), .o(delay_xor_ln21_unr21_stage8_stallmux_q_7_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_32370), .o(delay_xor_ln21_unr21_stage8_stallmux_q_8_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_32373), .o(delay_xor_ln21_unr21_stage8_stallmux_q_9_) );
ms00f80 delay_xor_ln21_unr28_stage10_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_40591), .o(delay_xor_ln21_unr28_stage10_stallmux_q_0_) );
ms00f80 delay_xor_ln21_unr28_stage10_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_40599), .o(delay_xor_ln21_unr28_stage10_stallmux_q_1_) );
ms00f80 delay_xor_ln21_unr28_stage10_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_40600), .o(delay_xor_ln21_unr28_stage10_stallmux_q_2_) );
ms00f80 delay_xor_ln21_unr28_stage10_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_40597), .o(delay_xor_ln21_unr28_stage10_stallmux_q_3_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_1327), .o(delay_xor_ln21_unr3_stage2_stallmux_q_0_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_1322), .o(delay_xor_ln21_unr3_stage2_stallmux_q_10_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_1298), .o(delay_xor_ln21_unr3_stage2_stallmux_q_11_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_1329), .o(delay_xor_ln21_unr3_stage2_stallmux_q_12_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_1288), .o(delay_xor_ln21_unr3_stage2_stallmux_q_13_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_1300), .o(delay_xor_ln21_unr3_stage2_stallmux_q_14_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_1332), .o(delay_xor_ln21_unr3_stage2_stallmux_q_15_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2949), .o(delay_xor_ln21_unr3_stage2_stallmux_q_16_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_1343), .o(delay_xor_ln21_unr3_stage2_stallmux_q_17_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_1333), .o(delay_xor_ln21_unr3_stage2_stallmux_q_18_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2951), .o(delay_xor_ln21_unr3_stage2_stallmux_q_19_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_1307), .o(delay_xor_ln21_unr3_stage2_stallmux_q_1_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2953), .o(delay_xor_ln21_unr3_stage2_stallmux_q_20_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_1302), .o(delay_xor_ln21_unr3_stage2_stallmux_q_21_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_1312), .o(delay_xor_ln21_unr3_stage2_stallmux_q_22_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2955), .o(delay_xor_ln21_unr3_stage2_stallmux_q_23_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_1336), .o(delay_xor_ln21_unr3_stage2_stallmux_q_24_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_1346), .o(delay_xor_ln21_unr3_stage2_stallmux_q_25_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_1303), .o(delay_xor_ln21_unr3_stage2_stallmux_q_26_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(TIMEBOOST_net_2957), .o(delay_xor_ln21_unr3_stage2_stallmux_q_27_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_1289), .o(delay_xor_ln21_unr3_stage2_stallmux_q_28_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_1301), .o(delay_xor_ln21_unr3_stage2_stallmux_q_2_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_1291), .o(delay_xor_ln21_unr3_stage2_stallmux_q_3_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_1345), .o(delay_xor_ln21_unr3_stage2_stallmux_q_4_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_1320), .o(delay_xor_ln21_unr3_stage2_stallmux_q_5_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_1287), .o(delay_xor_ln21_unr3_stage2_stallmux_q_6_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_1324), .o(delay_xor_ln21_unr3_stage2_stallmux_q_7_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_1315), .o(delay_xor_ln21_unr3_stage2_stallmux_q_8_) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_1306), .o(delay_xor_ln21_unr3_stage2_stallmux_q_9_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_46165), .o(delay_xor_ln21_unr6_stage3_stallmux_q_0_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_46160), .o(delay_xor_ln21_unr6_stage3_stallmux_q_10_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_46159), .o(delay_xor_ln21_unr6_stage3_stallmux_q_11_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_46167), .o(delay_xor_ln21_unr6_stage3_stallmux_q_12_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_46166), .o(delay_xor_ln21_unr6_stage3_stallmux_q_13_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_46155), .o(delay_xor_ln21_unr6_stage3_stallmux_q_14_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_46157), .o(delay_xor_ln21_unr6_stage3_stallmux_q_15_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_46149), .o(delay_xor_ln21_unr6_stage3_stallmux_q_16_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_46147), .o(delay_xor_ln21_unr6_stage3_stallmux_q_17_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_46178), .o(delay_xor_ln21_unr6_stage3_stallmux_q_18_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_46181), .o(delay_xor_ln21_unr6_stage3_stallmux_q_19_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_46174), .o(delay_xor_ln21_unr6_stage3_stallmux_q_1_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_46182), .o(delay_xor_ln21_unr6_stage3_stallmux_q_20_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_46184), .o(delay_xor_ln21_unr6_stage3_stallmux_q_21_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_46186), .o(delay_xor_ln21_unr6_stage3_stallmux_q_22_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_46187), .o(delay_xor_ln21_unr6_stage3_stallmux_q_23_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_46188), .o(delay_xor_ln21_unr6_stage3_stallmux_q_24_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_46192), .o(delay_xor_ln21_unr6_stage3_stallmux_q_25_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_46141), .o(delay_xor_ln21_unr6_stage3_stallmux_q_2_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_46156), .o(delay_xor_ln21_unr6_stage3_stallmux_q_3_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_46146), .o(delay_xor_ln21_unr6_stage3_stallmux_q_4_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_46176), .o(delay_xor_ln21_unr6_stage3_stallmux_q_5_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_46170), .o(delay_xor_ln21_unr6_stage3_stallmux_q_6_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_46163), .o(delay_xor_ln21_unr6_stage3_stallmux_q_7_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_46171), .o(delay_xor_ln21_unr6_stage3_stallmux_q_8_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_46152), .o(delay_xor_ln21_unr6_stage3_stallmux_q_9_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_46381), .o(delay_xor_ln21_unr9_stage4_stallmux_q_0_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_46367), .o(delay_xor_ln21_unr9_stage4_stallmux_q_10_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_46365), .o(delay_xor_ln21_unr9_stage4_stallmux_q_11_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_46362), .o(delay_xor_ln21_unr9_stage4_stallmux_q_12_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_46360), .o(delay_xor_ln21_unr9_stage4_stallmux_q_13_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_46359), .o(delay_xor_ln21_unr9_stage4_stallmux_q_14_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_46355), .o(delay_xor_ln21_unr9_stage4_stallmux_q_15_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_46354), .o(delay_xor_ln21_unr9_stage4_stallmux_q_16_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_46348), .o(delay_xor_ln21_unr9_stage4_stallmux_q_17_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_46353), .o(delay_xor_ln21_unr9_stage4_stallmux_q_18_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_46358), .o(delay_xor_ln21_unr9_stage4_stallmux_q_19_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_46384), .o(delay_xor_ln21_unr9_stage4_stallmux_q_1_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_46345), .o(delay_xor_ln21_unr9_stage4_stallmux_q_20_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_46342), .o(delay_xor_ln21_unr9_stage4_stallmux_q_21_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_46340), .o(delay_xor_ln21_unr9_stage4_stallmux_q_22_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_46373), .o(delay_xor_ln21_unr9_stage4_stallmux_q_2_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_46379), .o(delay_xor_ln21_unr9_stage4_stallmux_q_3_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_46385), .o(delay_xor_ln21_unr9_stage4_stallmux_q_4_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_46377), .o(delay_xor_ln21_unr9_stage4_stallmux_q_5_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_46372), .o(delay_xor_ln21_unr9_stage4_stallmux_q_6_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_46378), .o(delay_xor_ln21_unr9_stage4_stallmux_q_7_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_46374), .o(delay_xor_ln21_unr9_stage4_stallmux_q_8_) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_46386), .o(delay_xor_ln21_unr9_stage4_stallmux_q_9_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_16619), .o(delay_xor_ln22_unr12_stage5_stallmux_q_0_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_17585), .o(delay_xor_ln22_unr12_stage5_stallmux_q_10_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_17647), .o(delay_xor_ln22_unr12_stage5_stallmux_q_11_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_17677), .o(delay_xor_ln22_unr12_stage5_stallmux_q_12_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_17755), .o(delay_xor_ln22_unr12_stage5_stallmux_q_13_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_17754), .o(delay_xor_ln22_unr12_stage5_stallmux_q_14_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_17776), .o(delay_xor_ln22_unr12_stage5_stallmux_q_15_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_17750), .o(delay_xor_ln22_unr12_stage5_stallmux_q_16_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_17770), .o(delay_xor_ln22_unr12_stage5_stallmux_q_17_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_17769), .o(delay_xor_ln22_unr12_stage5_stallmux_q_18_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_17752), .o(delay_xor_ln22_unr12_stage5_stallmux_q_19_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_16636), .o(delay_xor_ln22_unr12_stage5_stallmux_q_1_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_16747), .o(delay_xor_ln22_unr12_stage5_stallmux_q_2_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_16804), .o(delay_xor_ln22_unr12_stage5_stallmux_q_3_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_16863), .o(delay_xor_ln22_unr12_stage5_stallmux_q_4_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_17029), .o(delay_xor_ln22_unr12_stage5_stallmux_q_5_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_17224), .o(delay_xor_ln22_unr12_stage5_stallmux_q_6_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_17337), .o(delay_xor_ln22_unr12_stage5_stallmux_q_7_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_17476), .o(delay_xor_ln22_unr12_stage5_stallmux_q_8_) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_17552), .o(delay_xor_ln22_unr12_stage5_stallmux_q_9_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_22424), .o(delay_xor_ln22_unr15_stage6_stallmux_q_0_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_22872), .o(delay_xor_ln22_unr15_stage6_stallmux_q_10_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_22908), .o(delay_xor_ln22_unr15_stage6_stallmux_q_11_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_22973), .o(delay_xor_ln22_unr15_stage6_stallmux_q_12_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_22834), .o(delay_xor_ln22_unr15_stage6_stallmux_q_13_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_22949), .o(delay_xor_ln22_unr15_stage6_stallmux_q_14_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_22947), .o(delay_xor_ln22_unr15_stage6_stallmux_q_15_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_22913), .o(delay_xor_ln22_unr15_stage6_stallmux_q_16_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_22480), .o(n_45204) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_22581), .o(delay_xor_ln22_unr15_stage6_stallmux_q_2_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_22671), .o(delay_xor_ln22_unr15_stage6_stallmux_q_3_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_22716), .o(delay_xor_ln22_unr15_stage6_stallmux_q_4_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_22712), .o(delay_xor_ln22_unr15_stage6_stallmux_q_5_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_22758), .o(delay_xor_ln22_unr15_stage6_stallmux_q_6_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_22777), .o(delay_xor_ln22_unr15_stage6_stallmux_q_7_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_22832), .o(delay_xor_ln22_unr15_stage6_stallmux_q_8_) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_22802), .o(delay_xor_ln22_unr15_stage6_stallmux_q_9_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_27652), .o(delay_xor_ln22_unr18_stage7_stallmux_q_0_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_27780), .o(delay_xor_ln22_unr18_stage7_stallmux_q_10_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_27846), .o(delay_xor_ln22_unr18_stage7_stallmux_q_11_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_27844), .o(delay_xor_ln22_unr18_stage7_stallmux_q_12_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_27838), .o(delay_xor_ln22_unr18_stage7_stallmux_q_13_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_27671), .o(delay_xor_ln22_unr18_stage7_stallmux_q_1_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_27687), .o(delay_xor_ln22_unr18_stage7_stallmux_q_2_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_27700), .o(delay_xor_ln22_unr18_stage7_stallmux_q_3_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_27731), .o(delay_xor_ln22_unr18_stage7_stallmux_q_4_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_27741), .o(delay_xor_ln22_unr18_stage7_stallmux_q_5_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_27797), .o(delay_xor_ln22_unr18_stage7_stallmux_q_6_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_27836), .o(delay_xor_ln22_unr18_stage7_stallmux_q_7_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_27779), .o(delay_xor_ln22_unr18_stage7_stallmux_q_8_) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_27843), .o(delay_xor_ln22_unr18_stage7_stallmux_q_9_) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_32431), .o(delay_xor_ln22_unr21_stage8_stallmux_q_0_) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_32567), .o(delay_xor_ln22_unr21_stage8_stallmux_q_10_) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_32467), .o(delay_xor_ln22_unr21_stage8_stallmux_q_1_) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_32545), .o(delay_xor_ln22_unr21_stage8_stallmux_q_2_) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_32511), .o(delay_xor_ln22_unr21_stage8_stallmux_q_3_) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_32565), .o(delay_xor_ln22_unr21_stage8_stallmux_q_4_) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_32541), .o(delay_xor_ln22_unr21_stage8_stallmux_q_5_) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_32594), .o(delay_xor_ln22_unr21_stage8_stallmux_q_6_) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_32515), .o(delay_xor_ln22_unr21_stage8_stallmux_q_7_) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_32571), .o(delay_xor_ln22_unr21_stage8_stallmux_q_8_) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_32569), .o(delay_xor_ln22_unr21_stage8_stallmux_q_9_) );
ms00f80 delay_xor_ln22_unr28_stage10_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_40580), .o(delay_xor_ln22_unr28_stage10_stallmux_q_0_) );
ms00f80 delay_xor_ln22_unr28_stage10_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_40589), .o(delay_xor_ln22_unr28_stage10_stallmux_q_1_) );
ms00f80 delay_xor_ln22_unr28_stage10_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_40588), .o(delay_xor_ln22_unr28_stage10_stallmux_q_2_) );
ms00f80 delay_xor_ln22_unr28_stage10_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_40587), .o(delay_xor_ln22_unr28_stage10_stallmux_q_3_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_1314), .o(delay_xor_ln22_unr3_stage2_stallmux_q_0_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_1325), .o(delay_xor_ln22_unr3_stage2_stallmux_q_10_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_44624), .o(delay_xor_ln22_unr3_stage2_stallmux_q_11_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_1337), .o(delay_xor_ln22_unr3_stage2_stallmux_q_12_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_1355), .o(delay_xor_ln22_unr3_stage2_stallmux_q_13_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_1348), .o(delay_xor_ln22_unr3_stage2_stallmux_q_14_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_1292), .o(delay_xor_ln22_unr3_stage2_stallmux_q_15_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_1350), .o(delay_xor_ln22_unr3_stage2_stallmux_q_16_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_1338), .o(delay_xor_ln22_unr3_stage2_stallmux_q_17_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_1311), .o(delay_xor_ln22_unr3_stage2_stallmux_q_18_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_1351), .o(delay_xor_ln22_unr3_stage2_stallmux_q_19_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_1340), .o(delay_xor_ln22_unr3_stage2_stallmux_q_1_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_1295), .o(delay_xor_ln22_unr3_stage2_stallmux_q_20_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_1297), .o(delay_xor_ln22_unr3_stage2_stallmux_q_21_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_1309), .o(delay_xor_ln22_unr3_stage2_stallmux_q_22_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_1357), .o(delay_xor_ln22_unr3_stage2_stallmux_q_23_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_1308), .o(delay_xor_ln22_unr3_stage2_stallmux_q_24_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_1356), .o(delay_xor_ln22_unr3_stage2_stallmux_q_25_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_26_ ( .ck(ispd_clk), .d(n_1286), .o(delay_xor_ln22_unr3_stage2_stallmux_q_26_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_27_ ( .ck(ispd_clk), .d(n_44624), .o(delay_xor_ln22_unr3_stage2_stallmux_q_27_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_28_ ( .ck(ispd_clk), .d(n_44624), .o(delay_xor_ln22_unr3_stage2_stallmux_q_28_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_1335), .o(delay_xor_ln22_unr3_stage2_stallmux_q_2_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_1360), .o(delay_xor_ln22_unr3_stage2_stallmux_q_3_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_1328), .o(delay_xor_ln22_unr3_stage2_stallmux_q_4_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_1316), .o(delay_xor_ln22_unr3_stage2_stallmux_q_5_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_1360), .o(delay_xor_ln22_unr3_stage2_stallmux_q_6_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_1285), .o(delay_xor_ln22_unr3_stage2_stallmux_q_7_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_44624), .o(delay_xor_ln22_unr3_stage2_stallmux_q_8_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_1294), .o(delay_xor_ln22_unr3_stage2_stallmux_q_9_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_46172), .o(delay_xor_ln22_unr6_stage3_stallmux_q_0_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_46158), .o(delay_xor_ln22_unr6_stage3_stallmux_q_10_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_46150), .o(delay_xor_ln22_unr6_stage3_stallmux_q_11_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_46161), .o(delay_xor_ln22_unr6_stage3_stallmux_q_12_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_46175), .o(delay_xor_ln22_unr6_stage3_stallmux_q_13_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_46151), .o(delay_xor_ln22_unr6_stage3_stallmux_q_14_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_46154), .o(delay_xor_ln22_unr6_stage3_stallmux_q_15_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_46177), .o(delay_xor_ln22_unr6_stage3_stallmux_q_16_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_46180), .o(delay_xor_ln22_unr6_stage3_stallmux_q_17_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_46179), .o(delay_xor_ln22_unr6_stage3_stallmux_q_18_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_46183), .o(delay_xor_ln22_unr6_stage3_stallmux_q_19_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_46169), .o(delay_xor_ln22_unr6_stage3_stallmux_q_1_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_46185), .o(delay_xor_ln22_unr6_stage3_stallmux_q_20_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_46189), .o(delay_xor_ln22_unr6_stage3_stallmux_q_21_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_46190), .o(delay_xor_ln22_unr6_stage3_stallmux_q_22_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_23_ ( .ck(ispd_clk), .d(n_46194), .o(delay_xor_ln22_unr6_stage3_stallmux_q_23_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_24_ ( .ck(ispd_clk), .d(n_46191), .o(delay_xor_ln22_unr6_stage3_stallmux_q_24_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_25_ ( .ck(ispd_clk), .d(n_46193), .o(delay_xor_ln22_unr6_stage3_stallmux_q_25_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_46148), .o(delay_xor_ln22_unr6_stage3_stallmux_q_2_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_46145), .o(delay_xor_ln22_unr6_stage3_stallmux_q_3_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_46162), .o(delay_xor_ln22_unr6_stage3_stallmux_q_4_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_46153), .o(delay_xor_ln22_unr6_stage3_stallmux_q_5_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_46164), .o(delay_xor_ln22_unr6_stage3_stallmux_q_6_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_46143), .o(delay_xor_ln22_unr6_stage3_stallmux_q_7_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_46168), .o(delay_xor_ln22_unr6_stage3_stallmux_q_8_) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_46173), .o(delay_xor_ln22_unr6_stage3_stallmux_q_9_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_0_ ( .ck(ispd_clk), .d(n_46380), .o(n_45209) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_10_ ( .ck(ispd_clk), .d(n_46366), .o(delay_xor_ln22_unr9_stage4_stallmux_q_10_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_11_ ( .ck(ispd_clk), .d(n_46369), .o(delay_xor_ln22_unr9_stage4_stallmux_q_11_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_12_ ( .ck(ispd_clk), .d(n_46364), .o(delay_xor_ln22_unr9_stage4_stallmux_q_12_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_13_ ( .ck(ispd_clk), .d(n_46363), .o(delay_xor_ln22_unr9_stage4_stallmux_q_13_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_14_ ( .ck(ispd_clk), .d(n_46361), .o(delay_xor_ln22_unr9_stage4_stallmux_q_14_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_15_ ( .ck(ispd_clk), .d(n_46356), .o(delay_xor_ln22_unr9_stage4_stallmux_q_15_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_16_ ( .ck(ispd_clk), .d(n_46351), .o(delay_xor_ln22_unr9_stage4_stallmux_q_16_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_17_ ( .ck(ispd_clk), .d(n_46352), .o(delay_xor_ln22_unr9_stage4_stallmux_q_17_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_18_ ( .ck(ispd_clk), .d(n_46344), .o(delay_xor_ln22_unr9_stage4_stallmux_q_18_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_19_ ( .ck(ispd_clk), .d(n_46357), .o(delay_xor_ln22_unr9_stage4_stallmux_q_19_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_1_ ( .ck(ispd_clk), .d(n_46387), .o(n_45622) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_20_ ( .ck(ispd_clk), .d(n_46347), .o(delay_xor_ln22_unr9_stage4_stallmux_q_20_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_21_ ( .ck(ispd_clk), .d(n_46350), .o(delay_xor_ln22_unr9_stage4_stallmux_q_21_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_22_ ( .ck(ispd_clk), .d(n_46349), .o(delay_xor_ln22_unr9_stage4_stallmux_q_22_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_2_ ( .ck(ispd_clk), .d(n_46382), .o(delay_xor_ln22_unr9_stage4_stallmux_q_2_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_3_ ( .ck(ispd_clk), .d(n_46383), .o(delay_xor_ln22_unr9_stage4_stallmux_q_3_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_4_ ( .ck(ispd_clk), .d(n_46375), .o(delay_xor_ln22_unr9_stage4_stallmux_q_4_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_5_ ( .ck(ispd_clk), .d(n_46370), .o(delay_xor_ln22_unr9_stage4_stallmux_q_5_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_6_ ( .ck(ispd_clk), .d(n_46376), .o(delay_xor_ln22_unr9_stage4_stallmux_q_6_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_7_ ( .ck(ispd_clk), .d(n_46371), .o(delay_xor_ln22_unr9_stage4_stallmux_q_7_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_8_ ( .ck(ispd_clk), .d(n_46388), .o(delay_xor_ln22_unr9_stage4_stallmux_q_8_) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_9_ ( .ck(ispd_clk), .d(n_46368), .o(delay_xor_ln22_unr9_stage4_stallmux_q_9_) );
ms00f80 delay_xor_ln23_unr3_stage2_stallmux_q_reg ( .ck(ispd_clk), .d(n_44626), .o(delay_xor_ln23_unr3_stage2_stallmux_q) );
ms00f80 delay_xor_ln23_unr6_stage3_stallmux_q_reg ( .ck(ispd_clk), .d(FE_OCP_RBN6198_FE_OFN789_n_46195), .o(delay_xor_ln23_unr6_stage3_stallmux_q) );
in01s02 drc ( .a(n_45809), .o(n_45812) );
in01s01 drc2 ( .a(n_45808), .o(n_45809) );
in01s03 drc28 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_46204) );
in01s02 drc784076 ( .a(n_45820), .o(n_45821) );
in01s02 drc784079 ( .a(n_45821), .o(n_45824) );
in01s04 drc784094 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_45840) );
in01s01 drc784098 ( .a(n_45844), .o(n_45845) );
in01s01 drc784099 ( .a(n_45843), .o(n_45844) );
in01s01 drc784123 ( .a(n_45873), .o(n_45874) );
in01s01 drc784124 ( .a(n_45872), .o(n_45873) );
in01s02 drc784129 ( .a(n_45879), .o(n_45880) );
in01s01 drc784130 ( .a(n_45878), .o(n_45879) );
in01s01 drc784142 ( .a(n_45890), .o(n_45891) );
in01s01 drc784145 ( .a(n_45891), .o(n_45894) );
in01s01 drc784748 ( .a(n_30633), .o(n_47233) );
in01s04 drc784749 ( .a(FE_OCPN1681_n_30614), .o(n_30633) );
in01s02 fopt ( .a(n_47187), .o(n_47186) );
in01s80 fopt782682 ( .a(FE_OCP_RBN3968_n_44061), .o(n_44083) );
in01m20 fopt782724 ( .a(FE_OCP_RBN2689_n_44100), .o(n_44102) );
in01m08 fopt782729 ( .a(n_34066), .o(n_44100) );
in01m02 fopt782732 ( .a(n_29316), .o(n_44139) );
in01s02 fopt782738 ( .a(n_17685), .o(n_44147) );
in01s02 fopt782742 ( .a(n_17686), .o(n_44153) );
in01s03 fopt782743 ( .a(n_22677), .o(n_44155) );
in01s02 fopt782745 ( .a(n_21119), .o(n_44158) );
in01s02 fopt782746 ( .a(n_44162), .o(n_44160) );
in01s01 fopt782748 ( .a(n_44163), .o(n_44162) );
in01f02 fopt782749 ( .a(n_20545), .o(n_44163) );
in01s02 fopt782750 ( .a(n_44166), .o(n_44165) );
in01s02 fopt782751 ( .a(n_38788), .o(n_44166) );
in01f04 fopt782752 ( .a(n_36535), .o(n_44168) );
in01s02 fopt782793 ( .a(n_32360), .o(n_44213) );
in01m02 fopt782795 ( .a(n_32290), .o(n_44216) );
in01s01 fopt782796 ( .a(n_44219), .o(n_44218) );
in01m10 fopt782821 ( .a(FE_OCP_RBN4905_n_44256), .o(n_44222) );
in01m08 fopt782831 ( .a(n_35550), .o(n_44256) );
in01f04 fopt782834 ( .a(n_33693), .o(n_44259) );
in01s01 fopt782836 ( .a(n_34890), .o(n_44262) );
in01s06 fopt782839 ( .a(n_27620), .o(n_44265) );
in01f06 fopt782845 ( .a(n_44275), .o(n_44267) );
in01s06 fopt782851 ( .a(n_44275), .o(n_44277) );
in01f04 fopt782852 ( .a(n_21973), .o(n_44275) );
in01m02 fopt782857 ( .a(n_44288), .o(n_44287) );
in01m01 fopt782858 ( .a(n_22028), .o(n_44288) );
in01m02 fopt782864 ( .a(n_21985), .o(n_44296) );
in01s01 fopt782874 ( .a(n_44311), .o(n_44309) );
in01s01 fopt782876 ( .a(n_44312), .o(n_44311) );
in01f08 fopt782877 ( .a(n_39290), .o(n_44312) );
in01s01 fopt782888 ( .a(n_22874), .o(n_44327) );
in01s01 fopt782889 ( .a(n_22875), .o(n_44329) );
in01s01 fopt782892 ( .a(n_17759), .o(n_44334) );
in01s01 fopt782900 ( .a(n_2308), .o(n_44344) );
in01s01 fopt782902 ( .a(n_44347), .o(n_44346) );
in01s01 fopt782903 ( .a(n_32966), .o(n_44347) );
in01s04 fopt782906 ( .a(n_8231), .o(n_44352) );
in01s01 fopt782907 ( .a(n_44355), .o(n_44354) );
in01s02 fopt782908 ( .a(n_44356), .o(n_44355) );
in01m06 fopt782909 ( .a(n_11726), .o(n_44356) );
in01s01 fopt782911 ( .a(n_27688), .o(n_44360) );
in01m40 fopt782960 ( .a(n_44422), .o(n_44420) );
in01m02 fopt782962 ( .a(n_24990), .o(n_44423) );
in01s01 fopt782963 ( .a(n_44426), .o(n_44425) );
in01f06 fopt782966 ( .a(n_44429), .o(n_44428) );
in01f06 fopt782967 ( .a(n_44430), .o(n_44429) );
in01f06 fopt782968 ( .a(n_41311), .o(n_44430) );
in01m02 fopt782969 ( .a(n_32338), .o(n_44432) );
in01s02 fopt782970 ( .a(n_32339), .o(n_44434) );
in01s01 fopt782972 ( .a(n_44438), .o(n_44437) );
in01s01 fopt782973 ( .a(n_44439), .o(n_44438) );
in01f02 fopt782974 ( .a(n_30451), .o(n_44439) );
in01s01 fopt782975 ( .a(n_25507), .o(n_44441) );
in01s01 fopt782976 ( .a(n_26208), .o(n_44443) );
in01s02 fopt782977 ( .a(n_24992), .o(n_44445) );
in01s01 fopt782978 ( .a(n_17729), .o(n_44447) );
in01s01 fopt782980 ( .a(n_44451), .o(n_44450) );
in01s01 fopt782981 ( .a(n_12065), .o(n_44451) );
in01m02 fopt782983 ( .a(n_44453), .o(n_44454) );
in01s02 fopt783041 ( .a(n_44511), .o(n_44516) );
in01s03 fopt783049 ( .a(FE_OFN4801_n_44498), .o(n_44511) );
in01s06 fopt783050 ( .a(FE_OFN4779_n_44490), .o(n_44498) );
in01s06 fopt783060 ( .a(FE_OFN4779_n_44490), .o(n_44492) );
in01s20 fopt783061 ( .a(FE_OFN756_n_44464), .o(n_44490) );
in01m08 fopt783094 ( .a(n_8875), .o(n_44570) );
in01s06 fopt783107 ( .a(n_44576), .o(n_44579) );
in01s10 fopt783110 ( .a(n_44575), .o(n_44576) );
in01m10 fopt783111 ( .a(n_44592), .o(n_44575) );
in01s10 fopt783125 ( .a(n_44575), .o(n_44594) );
in01m08 fopt783127 ( .a(n_8875), .o(n_44592) );
in01f04 fopt783135 ( .a(n_24862), .o(n_44621) );
in01s04 fopt783136 ( .a(n_44626), .o(n_44624) );
in01s06 fopt783137 ( .a(n_44623), .o(n_44626) );
in01m10 fopt783138 ( .a(n_44636), .o(n_44623) );
in01f06 fopt783139 ( .a(n_1282), .o(n_44636) );
in01s10 fopt783141 ( .a(n_44672), .o(n_44637) );
in01s01 fopt783144 ( .a(FE_OCPN5099_n_1282), .o(n_44650) );
in01s02 fopt783146 ( .a(n_44659), .o(n_44661) );
in01s06 fopt783149 ( .a(n_1282), .o(n_44659) );
in01s08 fopt783150 ( .a(n_1282), .o(n_44672) );
in01s06 fopt783151 ( .a(n_1282), .o(n_44652) );
in01m02 fopt783156 ( .a(n_40578), .o(n_44687) );
in01f02 fopt783158 ( .a(n_40577), .o(n_44690) );
in01s02 fopt783159 ( .a(n_40532), .o(n_44692) );
in01m80 fopt783161 ( .a(n_44695), .o(n_44696) );
in01s02 fopt783173 ( .a(n_44711), .o(n_44710) );
in01s06 fopt783174 ( .a(n_6487), .o(n_44711) );
in01f02 fopt783175 ( .a(n_35221), .o(n_44713) );
in01m02 fopt783177 ( .a(n_44718), .o(n_44717) );
in01m02 fopt783178 ( .a(n_21164), .o(n_44718) );
in01s40 fopt783179 ( .a(n_44721), .o(n_44720) );
in01s40 fopt783183 ( .a(FE_OCP_RBN7127_n_44722), .o(n_44723) );
in01m06 fopt783207 ( .a(FE_OCP_RBN7127_n_44722), .o(n_44759) );
in01s40 fopt783209 ( .a(FE_OCP_RBN7127_n_44722), .o(n_44761) );
in01s02 fopt783231 ( .a(n_44775), .o(n_44776) );
in01s10 fopt783235 ( .a(FE_OCP_RBN2443_n_44798), .o(n_44775) );
in01f20 fopt783240 ( .a(FE_OCP_RBN2433_FE_RN_107_0), .o(n_44798) );
in01m20 fopt783244 ( .a(FE_OCP_RBN2433_FE_RN_107_0), .o(n_44804) );
in01s02 fopt783247 ( .a(n_36669), .o(n_44809) );
in01s01 fopt783248 ( .a(n_44812), .o(n_44811) );
in01s01 fopt783249 ( .a(n_1863), .o(n_44812) );
in01f02 fopt783250 ( .a(n_44815), .o(n_44814) );
in01f04 fopt783251 ( .a(n_33547), .o(n_44815) );
in01m02 fopt783255 ( .a(n_9411), .o(n_44821) );
in01f02 fopt783256 ( .a(n_6720), .o(n_44823) );
in01s01 fopt783257 ( .a(n_44826), .o(n_44825) );
in01s01 fopt783258 ( .a(n_44827), .o(n_44826) );
in01m04 fopt783259 ( .a(n_28556), .o(n_44827) );
in01s01 fopt783260 ( .a(n_44829), .o(n_44828) );
in01s01 fopt783261 ( .a(n_7659), .o(n_44829) );
in01s01 fopt783262 ( .a(n_36410), .o(n_44831) );
in01f08 fopt783266 ( .a(n_36410), .o(n_44835) );
in01f02 fopt783276 ( .a(n_44849), .o(n_44850) );
in01f01 fopt783277 ( .a(n_14508), .o(n_44849) );
in01m06 fopt783278 ( .a(n_44853), .o(n_44852) );
in01m04 fopt783279 ( .a(n_10599), .o(n_44853) );
in01m06 fopt783280 ( .a(n_11146), .o(n_44855) );
in01s02 fopt783288 ( .a(n_44867), .o(n_44866) );
in01m06 fopt783289 ( .a(n_44869), .o(n_44867) );
in01s06 fopt783291 ( .a(n_44871), .o(n_44872) );
in01f06 fopt783292 ( .a(n_44869), .o(n_44871) );
in01s03 fopt783317 ( .a(FE_OCP_RBN2549_n_44881), .o(n_44887) );
in01m10 fopt783329 ( .a(n_44877), .o(n_44875) );
in01m10 fopt783333 ( .a(n_44920), .o(n_44877) );
in01m08 fopt783334 ( .a(n_44869), .o(n_44920) );
in01f08 fopt783335 ( .a(n_37850), .o(n_44869) );
in01m04 fopt783338 ( .a(n_38830), .o(n_44921) );
in01s08 fopt783356 ( .a(n_44925), .o(n_44926) );
in01s10 fopt783357 ( .a(n_44944), .o(n_44925) );
in01s10 fopt783359 ( .a(n_44944), .o(n_44946) );
in01f10 fopt783364 ( .a(n_38830), .o(n_44944) );
in01m06 fopt783366 ( .a(n_44955), .o(n_44954) );
in01m06 fopt783367 ( .a(n_38830), .o(n_44955) );
in01m02 fopt783369 ( .a(n_40579), .o(n_44958) );
in01s01 fopt783397 ( .a(n_44996), .o(n_44995) );
in01s01 fopt783405 ( .a(n_45010), .o(n_45008) );
in01s06 fopt783424 ( .a(n_45024), .o(n_45026) );
in01s01 fopt783427 ( .a(n_45024), .o(n_45023) );
in01m03 fopt783437 ( .a(n_45032), .o(n_45024) );
in01s06 fopt783438 ( .a(n_45013), .o(n_45032) );
in01s06 fopt783444 ( .a(n_45010), .o(n_45013) );
in01s03 fopt783446 ( .a(n_45012), .o(n_45050) );
in01s03 fopt783450 ( .a(n_45012), .o(n_45010) );
in01s06 fopt783451 ( .a(FE_OCPN869_n_45003), .o(n_45012) );
in01s01 fopt783454 ( .a(FE_OCPN869_n_45003), .o(n_45060) );
in01s03 fopt783465 ( .a(n_45073), .o(n_45072) );
in01s02 fopt783475 ( .a(n_45080), .o(n_45081) );
in01s06 fopt783477 ( .a(n_45073), .o(n_45080) );
in01s06 fopt783478 ( .a(n_45070), .o(n_45073) );
in01s06 fopt783481 ( .a(n_45091), .o(n_45070) );
in01s06 fopt783484 ( .a(n_45069), .o(n_45091) );
in01s03 fopt783489 ( .a(n_45066), .o(n_45069) );
in01s01 fopt783491 ( .a(n_45066), .o(n_45067) );
in01m01 fopt783493 ( .a(n_45066), .o(n_45101) );
in01m03 fopt783496 ( .a(n_45065), .o(n_45066) );
in01s03 fopt783499 ( .a(FE_OCPN869_n_45003), .o(n_45065) );
in01s06 fopt783507 ( .a(n_45002), .o(n_45003) );
in01s06 fopt783509 ( .a(FE_OCP_RBN2517_n_45120), .o(n_45002) );
in01s01 fopt783514 ( .a(FE_OCP_RBN2517_n_45120), .o(n_45118) );
in01m10 fopt783517 ( .a(n_18421), .o(n_45120) );
in01s01 fopt783522 ( .a(n_27805), .o(n_45132) );
in01f01 fopt783523 ( .a(n_15510), .o(n_45134) );
in01s01 fopt783524 ( .a(FE_OCP_RBN3041_n_45139), .o(n_45135) );
in01f06 fopt783528 ( .a(n_15510), .o(n_45139) );
in01s10 fopt783533 ( .a(FE_OCP_RBN5546_n_45145), .o(n_45146) );
in01s06 fopt783556 ( .a(n_45153), .o(n_45155) );
in01s20 fopt783560 ( .a(n_45149), .o(n_45153) );
in01s20 fopt783561 ( .a(n_45180), .o(n_45149) );
in01s20 fopt783562 ( .a(n_45180), .o(n_45181) );
in01s40 fopt783563 ( .a(n_45145), .o(n_45180) );
in01m40 fopt783564 ( .a(n_40662), .o(n_45145) );
in01m04 fopt783566 ( .a(n_34768), .o(n_45185) );
in01f02 fopt783567 ( .a(n_29451), .o(n_45186) );
in01f02 fopt783568 ( .a(n_39648), .o(n_45188) );
in01s02 fopt783569 ( .a(n_3161), .o(n_45190) );
in01m02 fopt783570 ( .a(n_38660), .o(n_45192) );
in01s01 fopt783571 ( .a(n_2408), .o(n_45194) );
in01s04 fopt783573 ( .a(n_40561), .o(n_45198) );
in01m40 fopt783574 ( .a(n_45202), .o(n_45200) );
in01s02 fopt783582 ( .a(n_45213), .o(n_45212) );
in01s01 fopt783583 ( .a(n_8405), .o(n_45213) );
in01s04 fopt783584 ( .a(n_6328), .o(n_45214) );
in01m02 fopt783586 ( .a(n_45216), .o(n_45217) );
in01m02 fopt783587 ( .a(n_6328), .o(n_45216) );
in01s01 fopt783655 ( .a(n_45301), .o(n_45300) );
in01s01 fopt783658 ( .a(n_45304), .o(n_45301) );
in01s02 fopt783659 ( .a(n_10742), .o(n_45304) );
in01s01 fopt783660 ( .a(n_40306), .o(n_45306) );
in01s02 fopt783662 ( .a(n_27782), .o(n_45309) );
in01m08 fopt783663 ( .a(FE_OCP_RBN5541_n_23044), .o(n_45311) );
in01s01 fopt783667 ( .a(n_2314), .o(n_45317) );
in01f01 fopt783669 ( .a(n_5031), .o(n_45319) );
in01m02 fopt783670 ( .a(n_45322), .o(n_45321) );
in01f02 fopt783671 ( .a(n_45323), .o(n_45322) );
in01f02 fopt783672 ( .a(n_5272), .o(n_45323) );
in01m06 fopt783675 ( .a(n_35275), .o(n_45327) );
in01f02 fopt783676 ( .a(n_25964), .o(n_45329) );
in01s02 fopt783796 ( .a(n_45474), .o(n_45475) );
in01s08 fopt783797 ( .a(n_45479), .o(n_45474) );
in01f06 fopt783798 ( .a(n_6214), .o(n_45479) );
in01m02 fopt783802 ( .a(n_5192), .o(n_45484) );
in01m01 fopt783804 ( .a(n_45488), .o(n_45487) );
in01s04 fopt783810 ( .a(FE_OCP_RBN2650_n_29470), .o(n_45489) );
in01m06 fopt783812 ( .a(n_45496), .o(n_45497) );
in01s06 fopt783813 ( .a(n_45498), .o(n_45496) );
in01m04 fopt783814 ( .a(n_22542), .o(n_45498) );
in01s02 fopt783815 ( .a(n_22542), .o(n_45499) );
in01s01 fopt783916 ( .a(n_7594), .o(n_45616) );
in01f02 fopt783917 ( .a(n_36447), .o(n_45617) );
in01s01 fopt783918 ( .a(n_27715), .o(n_45619) );
in01f04 fopt783920 ( .a(n_38671), .o(n_45623) );
in01s02 fopt783921 ( .a(n_36508), .o(n_45625) );
in01f02 fopt783922 ( .a(n_33492), .o(n_45627) );
in01m04 fopt783924 ( .a(n_45631), .o(n_45630) );
in01f06 fopt783925 ( .a(n_30302), .o(n_45631) );
in01s01 fopt783927 ( .a(FE_OCP_RBN5722_n_24506), .o(n_45633) );
in01s10 fopt783971 ( .a(FE_OCP_RBN2393_n_45697), .o(n_45685) );
in01s40 fopt783981 ( .a(FE_OCP_RBN6314_n_45224), .o(n_45697) );
in01s01 fopt783993 ( .a(n_45717), .o(n_45716) );
in01s01 fopt783994 ( .a(n_45718), .o(n_45717) );
in01f04 fopt784007 ( .a(n_45739), .o(n_45738) );
in01f06 fopt784008 ( .a(n_45740), .o(n_45739) );
in01m10 fopt784010 ( .a(n_32680), .o(n_45741) );
in01s01 fopt784012 ( .a(n_30263), .o(n_45744) );
in01s02 fopt784013 ( .a(n_27582), .o(n_45745) );
in01s04 fopt784014 ( .a(n_45748), .o(n_45747) );
in01m06 fopt784015 ( .a(n_11914), .o(n_45748) );
in01m02 fopt784019 ( .a(n_45755), .o(n_45754) );
in01m06 fopt784020 ( .a(n_32280), .o(n_45755) );
in01s02 fopt784023 ( .a(FE_OCP_RBN2635_n_29371), .o(n_45758) );
in01s03 fopt784288 ( .a(n_7), .o(n_46055) );
in01s06 fopt784300 ( .a(beta_31), .o(n_7) );
in01s06 fopt784327 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_46107) );
in01s01 fopt784701 ( .a(n_47180), .o(n_47181) );
in01m02 fopt784710 ( .a(n_21558), .o(n_47187) );
in01s01 fopt784716 ( .a(n_17835), .o(n_47195) );
in01m02 fopt784717 ( .a(n_5524), .o(n_47197) );
in01m02 fopt784718 ( .a(n_47200), .o(n_47199) );
in01f02 fopt784719 ( .a(n_11035), .o(n_47200) );
in01m40 fopt784721 ( .a(n_45508), .o(n_47203) );
in01s01 fopt784724 ( .a(n_22682), .o(n_47207) );
oa12s04 g2 ( .a(FE_OCP_RBN2430_FE_RN_107_0), .b(n_40737), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_6_), .o(n_44026) );
oa12f02 g736251 ( .a(n_333), .b(n_43912), .c(TIMEBOOST_net_1795), .o(n_43920) );
oa12f02 g736252 ( .a(n_294), .b(n_43911), .c(TIMEBOOST_net_1803), .o(n_43919) );
oa12f02 g736256 ( .a(n_295), .b(n_43907), .c(FE_OFN4653_n_43918), .o(n_43916) );
oa12f02 g736257 ( .a(n_293), .b(n_43908), .c(TIMEBOOST_net_1805), .o(n_43917) );
oa12f02 g736263 ( .a(n_302), .b(n_43901), .c(TIMEBOOST_net_1807), .o(n_43915) );
oa12f02 g736264 ( .a(n_322), .b(n_43900), .c(TIMEBOOST_net_1809), .o(n_43914) );
oa12f02 g736265 ( .a(n_331), .b(n_43902), .c(TIMEBOOST_net_1811), .o(n_43913) );
oa12s02 g736271 ( .a(n_289), .b(n_43861), .c(FE_OFN5_n_43918), .o(n_43903) );
oa12s02 g736272 ( .a(n_290), .b(n_43863), .c(FE_OFN5_n_43918), .o(n_43899) );
oa12s02 g736273 ( .a(n_310), .b(n_43862), .c(FE_OFN5_n_43918), .o(n_43898) );
oa12f02 g736274 ( .a(n_296), .b(n_43887), .c(TIMEBOOST_net_1813), .o(n_43910) );
oa12s01 g736275 ( .a(n_328), .b(n_43864), .c(FE_OFN5_n_43918), .o(n_43896) );
ao22f02 g736276 ( .a(n_43882), .b(n_43612), .c(FE_OCP_RBN6230_n_43882), .d(n_43611), .o(n_43908) );
in01f02 g736282 ( .a(n_43894), .o(n_43895) );
ao12f04 g736283 ( .a(n_43422), .b(n_43885), .c(n_43520), .o(n_43894) );
in01f02 g736284 ( .a(n_43892), .o(n_43893) );
ao12f04 g736285 ( .a(n_43471), .b(n_43885), .c(n_43384), .o(n_43892) );
oa12s01 g736286 ( .a(n_324), .b(n_43858), .c(FE_OFN4651_n_43918), .o(n_43890) );
oa12s02 g736287 ( .a(n_288), .b(n_43857), .c(FE_OFN5_n_43918), .o(n_43889) );
ao22f02 g736289 ( .a(n_43875), .b(n_43542), .c(n_43874), .d(n_43541), .o(n_43902) );
ao12f04 g736297 ( .a(FE_OCPN1226_n_43357), .b(n_43859), .c(n_43645), .o(n_43882) );
oa12f04 g736299 ( .a(n_43644), .b(n_43846), .c(n_43562), .o(n_43880) );
oa12f02 g736300 ( .a(n_297), .b(n_43879), .c(FE_OFN2_n_43918), .o(n_43909) );
oa12f02 g736301 ( .a(n_292), .b(n_43868), .c(TIMEBOOST_net_1801), .o(n_43897) );
ao22s02 g736303 ( .a(FE_RN_1622_0), .b(n_43544), .c(FE_OCP_RBN3424_FE_RN_1622_0), .d(n_43543), .o(n_43863) );
ao22s02 g736304 ( .a(n_43828), .b(n_43397), .c(n_43827), .d(n_43396), .o(n_43862) );
ao22s02 g736305 ( .a(n_43832), .b(n_43613), .c(n_43831), .d(n_43614), .o(n_43861) );
ao22f02 g736306 ( .a(n_43855), .b(n_43394), .c(n_43854), .d(n_43395), .o(n_43887) );
oa12f02 g736307 ( .a(n_308), .b(n_43867), .c(FE_OFN2_n_43918), .o(n_43906) );
oa12s02 g736308 ( .a(n_305), .b(n_43866), .c(FE_OFN4_n_43918), .o(n_43905) );
in01f02 g736314 ( .a(n_43876), .o(n_43877) );
na02f04 g736315 ( .a(n_43859), .b(n_43641), .o(n_43876) );
in01f02 g736316 ( .a(n_43874), .o(n_43875) );
oa12m02 g736318 ( .a(n_339), .b(n_43845), .c(TIMEBOOST_net_1797), .o(n_43886) );
oa12m02 g736319 ( .a(n_337), .b(n_43853), .c(FE_OFN2_n_43918), .o(n_43891) );
oa12s01 g736320 ( .a(n_332), .b(n_43823), .c(FE_OFN5_n_43918), .o(n_43873) );
ao22s01 g736321 ( .a(n_43808), .b(n_43619), .c(n_43807), .d(n_43620), .o(n_43858) );
oa12f02 g736322 ( .a(n_316), .b(n_43878), .c(TIMEBOOST_net_1799), .o(n_43904) );
ao22s02 g736323 ( .a(FE_OCP_RBN3411_n_43811), .b(n_43318), .c(n_43811), .d(n_43319), .o(n_43857) );
in01f02 g736325 ( .a(n_43871), .o(n_43872) );
in01f02 g736326 ( .a(n_43885), .o(n_43871) );
na02s02 TIMEBOOST_cell_1240 ( .a(n_28770), .b(TIMEBOOST_net_234), .o(n_28788) );
na02f08 g736336 ( .a(n_43833), .b(n_43432), .o(n_43859) );
in01f02 g736337 ( .a(n_43854), .o(n_43855) );
in01f02 g736338 ( .a(n_43846), .o(n_43854) );
no02f06 g736339 ( .a(n_43833), .b(n_43646), .o(n_43846) );
na02s01 TIMEBOOST_cell_6031 ( .a(FE_OCP_RBN6570_n_44875), .b(n_37598), .o(TIMEBOOST_net_1867) );
in01s01 g736341 ( .a(n_43831), .o(n_43832) );
oa12s02 g736342 ( .a(n_43566), .b(FE_OCP_RBN3402_n_43775), .c(n_43437), .o(n_43831) );
oa12s02 g736344 ( .a(n_43326), .b(n_43789), .c(n_43361), .o(n_43829) );
in01s01 g736345 ( .a(n_43827), .o(n_43828) );
oa12s02 g736346 ( .a(n_43525), .b(FE_OCP_RBN3402_n_43775), .c(n_43360), .o(n_43827) );
oa12f02 g736349 ( .a(n_291), .b(n_43847), .c(FE_OFN2_n_43918), .o(n_43884) );
oa12m02 g736350 ( .a(n_347), .b(n_43839), .c(FE_OFN2_n_43918), .o(n_43870) );
oa12m02 g736351 ( .a(n_298), .b(n_43838), .c(FE_OFN2_n_43918), .o(n_43869) );
ao22f02 g736352 ( .a(n_43849), .b(n_43602), .c(n_43848), .d(FE_OCPN1230_n_43601), .o(n_43879) );
oa12s01 g736353 ( .a(n_340), .b(n_43774), .c(FE_OFN4651_n_43918), .o(n_43813) );
ao22f02 g736354 ( .a(n_43840), .b(n_43600), .c(n_43841), .d(n_43599), .o(n_43868) );
ao22f02 g736355 ( .a(n_43836), .b(n_43598), .c(FE_OCP_RBN3464_n_43836), .d(n_43597), .o(n_43867) );
oa12s02 g736357 ( .a(n_342), .b(n_43835), .c(FE_OFN2_n_43918), .o(n_43865) );
na02s02 g736362 ( .a(n_43789), .b(n_43291), .o(n_43811) );
na02s02 g736364 ( .a(FE_OCP_RBN3402_n_43775), .b(n_43440), .o(n_43809) );
in01s01 g736365 ( .a(n_43807), .o(n_43808) );
oa12s02 g736366 ( .a(FE_OCPN1224_n_43521), .b(n_43772), .c(n_43255), .o(n_43807) );
in01f06 g736368 ( .a(n_43788), .o(n_43833) );
na02f08 g736369 ( .a(n_43775), .b(n_43408), .o(n_43788) );
ao22m02 g736370 ( .a(n_43799), .b(n_43604), .c(n_43798), .d(n_43603), .o(n_43845) );
ao22s02 g736371 ( .a(n_43820), .b(n_43516), .c(n_43821), .d(n_43517), .o(n_43853) );
oa12s02 g736372 ( .a(n_349), .b(n_43771), .c(FE_OFN4651_n_43918), .o(n_43805) );
oa12s01 g736373 ( .a(n_300), .b(n_43770), .c(FE_OFN5_n_43918), .o(n_43804) );
oa12s01 g736374 ( .a(n_312), .b(n_43785), .c(FE_OFN4651_n_43918), .o(n_43824) );
ao22s01 g736375 ( .a(n_43772), .b(n_43561), .c(n_43759), .d(n_43560), .o(n_43823) );
oa12f02 g736377 ( .a(n_329), .b(n_43794), .c(FE_OFN1_n_43918), .o(n_43852) );
oa12f02 g736378 ( .a(n_315), .b(n_43793), .c(FE_OFN1_n_43918), .o(n_43851) );
oa12s02 g736379 ( .a(n_350), .b(n_43795), .c(FE_OFN4_n_43918), .o(n_43850) );
oa12s01 g736380 ( .a(n_309), .b(n_43784), .c(FE_OFN4_n_43918), .o(n_43844) );
oa12s02 g736381 ( .a(n_338), .b(n_43815), .c(FE_OFN2_n_43918), .o(n_43860) );
na02s06 g736386 ( .a(n_43759), .b(n_43433), .o(n_43789) );
in01f02 g736389 ( .a(n_43840), .o(n_43841) );
ao12f04 g736390 ( .a(n_43684), .b(n_43822), .c(n_43429), .o(n_43840) );
in01m02 g736391 ( .a(n_43848), .o(n_43849) );
na02m04 g736392 ( .a(n_43801), .b(n_43658), .o(n_43848) );
no02f08 g736394 ( .a(n_43747), .b(n_43434), .o(n_43775) );
ao22s02 g736396 ( .a(FE_OCP_RBN3449_n_43777), .b(n_43606), .c(n_43777), .d(FE_OCPN1228_n_43605), .o(n_43838) );
ao22m02 g736397 ( .a(n_43783), .b(n_43425), .c(n_43792), .d(n_43426), .o(n_43847) );
oa12s02 g736398 ( .a(n_327), .b(n_43758), .c(FE_OFN5_n_43918), .o(n_43803) );
oa12s01 g736399 ( .a(n_325), .b(n_43757), .c(FE_OFN4651_n_43918), .o(n_43802) );
ao22s01 g736400 ( .a(n_43731), .b(n_43546), .c(n_43732), .d(n_43545), .o(n_43774) );
oa12s01 g736401 ( .a(n_320), .b(n_43730), .c(FE_OFN4651_n_43918), .o(n_43773) );
ao12f04 g736403 ( .a(n_43683), .b(n_43822), .c(n_43466), .o(n_43836) );
na02m04 g736409 ( .a(n_43800), .b(n_43420), .o(n_43801) );
in01s02 g736410 ( .a(n_43820), .o(n_43821) );
no02s04 g736411 ( .a(n_43800), .b(n_43657), .o(n_43820) );
na02s02 g736412 ( .a(n_43790), .b(n_43682), .o(n_43819) );
no02m04 g736413 ( .a(n_43791), .b(n_43678), .o(n_43834) );
in01s01 g736416 ( .a(n_43759), .o(n_43772) );
in01s02 g736417 ( .a(n_43747), .o(n_43759) );
ao12f08 g736418 ( .a(n_43443), .b(n_43721), .c(FE_OCP_DRV_N1406_n_43514), .o(n_43747) );
in01s02 g736419 ( .a(n_43798), .o(n_43799) );
oa12m04 g736420 ( .a(n_43649), .b(n_43768), .c(n_43390), .o(n_43798) );
ao22s02 g736421 ( .a(n_43729), .b(n_43550), .c(n_43728), .d(n_43549), .o(n_43771) );
ao22s01 g736422 ( .a(n_43727), .b(n_43548), .c(n_43726), .d(n_43547), .o(n_43770) );
ao22s01 g736423 ( .a(n_43744), .b(n_43354), .c(n_43745), .d(n_43353), .o(n_43785) );
oa12s01 g736424 ( .a(n_303), .b(n_43749), .c(FE_OFN4_n_43918), .o(n_43797) );
oa12s01 g736425 ( .a(n_346), .b(n_43748), .c(FE_OFN4_n_43918), .o(n_43796) );
oa12s01 g736426 ( .a(n_344), .b(n_43761), .c(FE_OFN4_n_43918), .o(n_43818) );
ao22s02 g736427 ( .a(n_43754), .b(n_43584), .c(n_43755), .d(n_43583), .o(n_43795) );
oa12s02 g736428 ( .a(n_336), .b(n_43760), .c(FE_OFN1_n_43918), .o(n_43817) );
ao22f02 g736429 ( .a(n_43752), .b(n_43631), .c(n_43753), .d(n_43630), .o(n_43794) );
ao22f02 g736430 ( .a(n_43750), .b(n_43310), .c(n_43751), .d(n_43309), .o(n_43793) );
ao22s01 g736431 ( .a(n_43740), .b(n_43582), .c(n_43739), .d(n_43581), .o(n_43784) );
no02m08 g736434 ( .a(n_43435), .b(n_43768), .o(n_43800) );
no02s02 g736435 ( .a(n_43762), .b(n_43636), .o(n_43783) );
na02m04 g736436 ( .a(n_43763), .b(n_43642), .o(n_43792) );
in01s01 g736437 ( .a(n_43731), .o(n_43732) );
no02s01 g736438 ( .a(n_43444), .b(n_43721), .o(n_43731) );
in01s02 g736439 ( .a(n_43781), .o(n_43782) );
oa12s02 g736440 ( .a(n_43480), .b(n_43716), .c(n_43225), .o(n_43781) );
in01s02 g736441 ( .a(n_43779), .o(n_43780) );
oa12s02 g736442 ( .a(n_43414), .b(n_43716), .c(n_43214), .o(n_43779) );
oa12s02 g736444 ( .a(n_43527), .b(n_43716), .c(n_43331), .o(n_43777) );
in01m02 g736445 ( .a(n_43790), .o(n_43791) );
in01m03 g736446 ( .a(n_43822), .o(n_43790) );
ao22s01 g736448 ( .a(n_43720), .b(n_43221), .c(n_43719), .d(n_43220), .o(n_43758) );
ao22s01 g736449 ( .a(n_43718), .b(n_43321), .c(n_43717), .d(n_43322), .o(n_43757) );
oa12s01 g736450 ( .a(n_335), .b(n_43704), .c(FE_OFN5_n_43918), .o(n_43746) );
ao22s01 g736451 ( .a(n_43690), .b(n_43537), .c(n_43689), .d(n_43536), .o(n_43730) );
oa12s02 g736452 ( .a(n_314), .b(n_43724), .c(FE_OFN1_n_43918), .o(n_43767) );
oa12s01 g736453 ( .a(n_348), .b(n_43737), .c(FE_OFN4_n_43918), .o(n_43776) );
oa12s01 g736454 ( .a(n_330), .b(n_43723), .c(FE_OFN4_n_43918), .o(n_43766) );
in01s01 g736457 ( .a(n_43744), .o(n_43745) );
na03s08 TIMEBOOST_cell_7128 ( .a(n_17894), .b(n_17827), .c(n_17848), .o(n_17895) );
in01s01 g736460 ( .a(n_43764), .o(n_43765) );
na02s02 g736461 ( .a(n_43716), .b(n_43368), .o(n_43764) );
in01m02 g736463 ( .a(n_43762), .o(n_43763) );
in01m04 g736464 ( .a(n_43768), .o(n_43762) );
in01m10 g736465 ( .a(n_43742), .o(n_43768) );
no02m10 g736466 ( .a(n_43716), .b(n_43330), .o(n_43742) );
in01s01 g736467 ( .a(n_43728), .o(n_43729) );
na02s02 g736468 ( .a(n_43691), .b(n_43227), .o(n_43728) );
in01s01 g736469 ( .a(n_43754), .o(n_43755) );
oa12s02 g736470 ( .a(n_43245), .b(n_43722), .c(n_43311), .o(n_43754) );
in01f02 g736471 ( .a(n_43752), .o(n_43753) );
ao12m04 g736472 ( .a(n_43168), .b(n_43741), .c(n_43515), .o(n_43752) );
in01s01 g736473 ( .a(n_43726), .o(n_43727) );
oa12s01 g736474 ( .a(n_43375), .b(n_43664), .c(n_43272), .o(n_43726) );
in01f02 g736475 ( .a(n_43750), .o(n_43751) );
ao12m04 g736476 ( .a(n_43372), .b(n_43741), .c(n_43273), .o(n_43750) );
oa12s01 g736477 ( .a(n_323), .b(n_43672), .c(FE_OFN5_n_43918), .o(n_43707) );
ao22s01 g736478 ( .a(n_43715), .b(n_43588), .c(n_43714), .d(n_43587), .o(n_43749) );
ao22s01 g736479 ( .a(n_43713), .b(n_43586), .c(n_43712), .d(n_43585), .o(n_43748) );
ao22s01 g736480 ( .a(n_43735), .b(n_43344), .c(n_43722), .d(n_43345), .o(n_43761) );
ao22m01 g736481 ( .a(n_43711), .b(n_43552), .c(n_43741), .d(n_43551), .o(n_43760) );
in01s01 g736482 ( .a(n_43739), .o(n_43740) );
oa12s01 g736483 ( .a(n_43373), .b(n_43711), .c(n_43366), .o(n_43739) );
in01s01 g736487 ( .a(n_43719), .o(n_43720) );
na02s02 g736488 ( .a(n_43676), .b(n_43164), .o(n_43719) );
na02s02 g736489 ( .a(n_43675), .b(n_43183), .o(n_43691) );
in01s01 g736490 ( .a(n_43717), .o(n_43718) );
na02s01 g736491 ( .a(n_43664), .b(n_43333), .o(n_43717) );
na02s02 TIMEBOOST_cell_7612 ( .a(n_2320), .b(n_2870), .o(TIMEBOOST_net_2437) );
in01s01 g736493 ( .a(n_43689), .o(n_43690) );
oa12s01 g736494 ( .a(n_43519), .b(n_43665), .c(n_43108), .o(n_43689) );
na02m10 g736498 ( .a(n_43701), .b(n_43367), .o(n_43716) );
oa12s01 g736499 ( .a(n_326), .b(n_43653), .c(FE_OFN5_n_43918), .o(n_43677) );
ao22s01 g736500 ( .a(n_43665), .b(n_43557), .c(n_43670), .d(n_43556), .o(n_43704) );
oa12s01 g736501 ( .a(n_313), .b(n_43708), .c(FE_OFN4_n_43918), .o(n_43738) );
ao22m02 g736502 ( .a(n_43696), .b(n_43590), .c(n_43697), .d(n_43589), .o(n_43724) );
ao22s02 g736503 ( .a(n_43699), .b(n_43264), .c(n_43700), .d(n_43263), .o(n_43723) );
ao22s01 g736504 ( .a(n_43710), .b(n_43261), .c(n_43709), .d(n_43262), .o(n_43737) );
in01s01 g736506 ( .a(n_43675), .o(n_43676) );
no02s01 g736507 ( .a(n_43665), .b(n_43234), .o(n_43675) );
in01s01 g736508 ( .a(n_43714), .o(n_43715) );
na02s02 g736509 ( .a(n_43687), .b(n_43277), .o(n_43714) );
in01s01 g736510 ( .a(n_43712), .o(n_43713) );
oa12s01 g736511 ( .a(n_43478), .b(n_43661), .c(n_43223), .o(n_43712) );
na02f08 g736515 ( .a(n_43654), .b(n_43235), .o(n_43664) );
oa12s01 g736516 ( .a(n_311), .b(n_43663), .c(FE_OFN5_n_43918), .o(n_43703) );
ao22s01 g736517 ( .a(n_43640), .b(n_43607), .c(n_43639), .d(n_43608), .o(n_43672) );
oa12s01 g736518 ( .a(n_319), .b(n_43652), .c(FE_OFN4_n_43918), .o(n_43688) );
oa12s01 g736519 ( .a(n_287), .b(n_43662), .c(FE_OFN4_n_43918), .o(n_43702) );
in01s01 g736521 ( .a(n_43722), .o(n_43735) );
oa12s02 g736522 ( .a(n_43477), .b(n_43661), .c(n_43275), .o(n_43722) );
in01f04 g736525 ( .a(n_43711), .o(n_43741) );
in01f02 g736526 ( .a(n_43701), .o(n_43711) );
oa12f10 g736527 ( .a(n_43411), .b(n_43661), .c(n_43328), .o(n_43701) );
in01s01 g736529 ( .a(n_43699), .o(n_43700) );
no02s02 g736530 ( .a(n_43686), .b(n_43276), .o(n_43699) );
na02s02 g736531 ( .a(n_43686), .b(n_43217), .o(n_43687) );
in01s01 g736532 ( .a(n_43709), .o(n_43710) );
na02s01 g736533 ( .a(n_43661), .b(n_43409), .o(n_43709) );
in01s02 g736534 ( .a(n_43696), .o(n_43697) );
ao12s04 g736535 ( .a(n_43489), .b(n_43659), .c(n_43553), .o(n_43696) );
in01s01 g736537 ( .a(n_43665), .o(n_43670) );
in01s01 g736538 ( .a(n_43654), .o(n_43665) );
oa12f08 g736539 ( .a(FE_OCP_DRV_N3520_n_43153), .b(n_43629), .c(FE_OCP_DRV_N3522_n_43538), .o(n_43654) );
ao22s01 g736540 ( .a(n_43573), .b(n_43146), .c(n_43574), .d(n_43145), .o(n_43653) );
oa12s01 g736541 ( .a(n_341), .b(n_43660), .c(FE_OFN4_n_43918), .o(n_43695) );
ao22s01 g736542 ( .a(n_43651), .b(n_43622), .c(n_43659), .d(n_43621), .o(n_43708) );
no02s02 g736544 ( .a(n_43651), .b(n_43285), .o(n_43686) );
in01s01 g736545 ( .a(n_43639), .o(n_43640) );
na02s01 g736546 ( .a(n_43629), .b(n_43091), .o(n_43639) );
ao22s01 g736547 ( .a(n_43572), .b(n_43615), .c(n_43571), .d(n_43616), .o(n_43663) );
oa12s02 g736548 ( .a(n_318), .b(n_43650), .c(FE_OFN1_n_43918), .o(n_43685) );
ao22s01 g736549 ( .a(n_43569), .b(n_43178), .c(n_43570), .d(n_43177), .o(n_43652) );
ao22s01 g736550 ( .a(n_43567), .b(n_43592), .c(n_43568), .d(n_43591), .o(n_43662) );
na02f10 g736554 ( .a(n_43638), .b(n_43286), .o(n_43661) );
na02f08 g736557 ( .a(n_43532), .b(n_43111), .o(n_43629) );
in01s01 g736558 ( .a(n_43573), .o(n_43574) );
no02s01 g736559 ( .a(n_43152), .b(n_43532), .o(n_43573) );
oa12s01 g736560 ( .a(n_345), .b(n_43656), .c(FE_OFN4_n_43918), .o(n_43694) );
ao22s01 g736561 ( .a(n_43628), .b(n_43594), .c(n_43627), .d(n_43593), .o(n_43660) );
in01s02 g736564 ( .a(n_43651), .o(n_43659) );
in01s01 g736565 ( .a(n_43638), .o(n_43651) );
na02s01 TIMEBOOST_cell_3909 ( .a(n_38270), .b(FE_OCP_RBN4026_n_37577), .o(TIMEBOOST_net_1045) );
no02s02 TIMEBOOST_cell_6879 ( .a(n_40909), .b(n_40908), .o(TIMEBOOST_net_2198) );
no02f08 g736568 ( .a(n_43450), .b(FE_OCPN1715_n_43449), .o(n_43532) );
in01s01 g736569 ( .a(n_43571), .o(n_43572) );
na02s01 g736570 ( .a(n_43450), .b(n_43518), .o(n_43571) );
na02m04 g736571 ( .a(n_43682), .b(n_43424), .o(n_43684) );
na02m04 g736572 ( .a(n_43682), .b(n_43473), .o(n_43683) );
na02s02 g736573 ( .a(n_43682), .b(n_43563), .o(n_43681) );
in01s01 g736574 ( .a(n_43569), .o(n_43570) );
ao12s01 g736575 ( .a(n_43162), .b(n_43446), .c(n_43529), .o(n_43569) );
in01s01 g736576 ( .a(n_43567), .o(n_43568) );
no02s01 g736577 ( .a(n_43528), .b(n_43224), .o(n_43567) );
oa12s01 g736578 ( .a(n_304), .b(n_43648), .c(FE_OFN4653_n_43918), .o(n_43680) );
ao22s02 g736579 ( .a(n_43378), .b(n_43555), .c(n_43379), .d(n_43554), .o(n_43650) );
oa12s01 g736580 ( .a(n_301), .b(n_43655), .c(FE_OFN4_n_43918), .o(n_43693) );
na02f08 g736583 ( .a(n_43335), .b(n_43385), .o(n_43450) );
no02s02 g736584 ( .a(n_43657), .b(n_43464), .o(n_43658) );
in01m01 g736586 ( .a(n_43682), .o(n_43678) );
no02m08 g736587 ( .a(n_43657), .b(n_43431), .o(n_43682) );
no02f10 g736588 ( .a(n_43417), .b(n_43114), .o(n_43528) );
in01s01 g736589 ( .a(n_43627), .o(n_43628) );
na02s01 g736590 ( .a(n_43447), .b(n_43495), .o(n_43627) );
ao22s01 g736591 ( .a(n_43376), .b(n_43633), .c(n_43377), .d(n_43632), .o(n_43656) );
no02s03 g736592 ( .a(n_43636), .b(n_43391), .o(n_43649) );
na02m08 g736593 ( .a(n_43626), .b(n_43404), .o(n_43657) );
in01s01 g736594 ( .a(n_43446), .o(n_43447) );
in01s01 g736595 ( .a(n_43417), .o(n_43446) );
na02f08 g736596 ( .a(n_43334), .b(n_43084), .o(n_43417) );
oa12s01 g736597 ( .a(n_306), .b(n_43191), .c(FE_OFN4653_n_43918), .o(n_43337) );
ao22s01 g736598 ( .a(n_43241), .b(n_43578), .c(n_43240), .d(n_43577), .o(n_43648) );
oa12s01 g736599 ( .a(n_343), .b(n_43236), .c(FE_OFN4_n_43918), .o(n_43381) );
ao22s01 g736600 ( .a(n_43238), .b(n_43596), .c(n_43239), .d(n_43595), .o(n_43655) );
in01s01 g736601 ( .a(n_43378), .o(n_43379) );
in01s01 g736602 ( .a(n_43335), .o(n_43378) );
oa12f06 g736603 ( .a(n_43159), .b(n_43157), .c(FE_OCP_RBN3310_n_43022), .o(n_43335) );
na02m04 g736606 ( .a(n_43623), .b(n_43625), .o(n_43637) );
no02s02 g736608 ( .a(n_43646), .b(n_43564), .o(n_43645) );
no02s02 g736609 ( .a(n_43624), .b(n_43467), .o(n_43644) );
in01s02 g736611 ( .a(n_43636), .o(n_43642) );
in01s02 g736612 ( .a(n_43626), .o(n_43636) );
na02s02 TIMEBOOST_cell_6338 ( .a(TIMEBOOST_net_2020), .b(n_32051), .o(n_32120) );
no02s02 g736614 ( .a(n_43646), .b(n_43406), .o(n_43641) );
in01s01 g736615 ( .a(n_43376), .o(n_43377) );
in01s01 g736616 ( .a(n_43334), .o(n_43376) );
no02s01 TIMEBOOST_cell_3068 ( .a(n_7582), .b(n_8840), .o(TIMEBOOST_net_825) );
na02s01 g736620 ( .a(n_43442), .b(n_43320), .o(n_43444) );
no02s01 g736621 ( .a(n_43565), .b(n_43316), .o(n_43566) );
in01s01 g736622 ( .a(n_43240), .o(n_43241) );
na02s01 g736623 ( .a(n_43118), .b(n_43054), .o(n_43240) );
in01s01 g736624 ( .a(n_43238), .o(n_43239) );
no02s01 g736625 ( .a(n_43193), .b(n_43067), .o(n_43238) );
no02f06 TIMEBOOST_cell_6214 ( .a(TIMEBOOST_net_1958), .b(n_35122), .o(n_35178) );
na02f06 g736627 ( .a(n_43156), .b(n_43158), .o(n_43159) );
no02s02 g736628 ( .a(n_43479), .b(n_43266), .o(n_43527) );
na02s08 g736629 ( .a(n_43442), .b(n_43284), .o(n_43443) );
in01s03 g736630 ( .a(n_43625), .o(n_43646) );
no02s06 g736631 ( .a(n_43565), .b(n_43407), .o(n_43625) );
no02f06 g736632 ( .a(n_43156), .b(n_43045), .o(n_43157) );
in01s01 g736633 ( .a(n_43623), .o(n_43624) );
oa12s02 g736634 ( .a(FE_OCP_RBN3312_n_43022), .b(n_43564), .c(n_43298), .o(n_43623) );
no02m10 TIMEBOOST_cell_1186 ( .a(n_41294), .b(TIMEBOOST_net_207), .o(n_41314) );
oa12s01 g736636 ( .a(n_299), .b(n_43115), .c(FE_OFN4653_n_43918), .o(n_43237) );
ao22s01 g736637 ( .a(n_43096), .b(n_43069), .c(n_43095), .d(n_43068), .o(n_43191) );
ao22s01 g736638 ( .a(n_43117), .b(n_43089), .c(n_43116), .d(n_43090), .o(n_43236) );
oa12s01 g736639 ( .a(n_321), .b(n_43151), .c(FE_OFN1_n_43918), .o(n_43288) );
in01s01 g736640 ( .a(n_43156), .o(n_43118) );
no02f08 g736641 ( .a(n_43075), .b(n_43035), .o(n_43156) );
no02s01 g736642 ( .a(n_43413), .b(n_43215), .o(n_43414) );
no02f04 g736643 ( .a(n_43094), .b(n_43066), .o(n_43193) );
no02s01 g736644 ( .a(n_43374), .b(n_43271), .o(n_43375) );
no02s01 g736645 ( .a(n_43475), .b(n_43352), .o(n_43526) );
in01s01 g736646 ( .a(n_43479), .o(n_43480) );
in01s01 g736647 ( .a(n_43441), .o(n_43479) );
no02s06 g736648 ( .a(n_43413), .b(n_43370), .o(n_43441) );
no02s01 g736649 ( .a(n_43369), .b(n_43216), .o(n_43478) );
in01s01 g736650 ( .a(n_43442), .o(n_43412) );
no02s06 g736651 ( .a(n_43374), .b(n_43233), .o(n_43442) );
in01s01 g736652 ( .a(n_43565), .o(n_43525) );
na02m04 g736653 ( .a(n_43440), .b(n_43365), .o(n_43565) );
no02s01 g736654 ( .a(n_43369), .b(n_43283), .o(n_43477) );
na02s02 g736655 ( .a(n_43474), .b(FE_OCP_RBN6191_n_43103), .o(n_43563) );
no02s10 g736656 ( .a(n_43332), .b(n_43369), .o(n_43411) );
oa12s01 g736657 ( .a(n_334), .b(n_43074), .c(FE_OFN4653_n_43918), .o(n_43155) );
oa12s01 g736658 ( .a(n_317), .b(n_43073), .c(FE_OFN4653_n_43918), .o(n_43154) );
na02s02 g736659 ( .a(n_43405), .b(n_43393), .o(n_43564) );
no02s01 g736660 ( .a(n_43372), .b(n_43166), .o(n_43373) );
no02s06 TIMEBOOST_cell_1185 ( .a(n_41293), .b(FE_OCPN3556_n_40986), .o(TIMEBOOST_net_207) );
ao12m02 g736662 ( .a(n_43152), .b(FE_OCP_RBN3306_n_43022), .c(n_43071), .o(n_43153) );
in01s01 g736663 ( .a(n_43374), .o(n_43333) );
na02s04 g736664 ( .a(n_43190), .b(n_43164), .o(n_43374) );
in01s01 g736666 ( .a(n_43440), .o(n_43475) );
no02s06 g736667 ( .a(n_43327), .b(n_43325), .o(n_43440) );
na02s02 g736668 ( .a(n_43473), .b(n_43006), .o(n_43474) );
ao12m08 g736669 ( .a(n_43162), .b(n_43171), .c(n_43143), .o(n_43287) );
in01s01 g736673 ( .a(n_43369), .o(n_43409) );
no03s02 TIMEBOOST_cell_8276 ( .a(FE_RN_303_0), .b(FE_RN_304_0), .c(n_2605), .o(n_47025) );
in01s01 g736676 ( .a(n_43413), .o(n_43368) );
na02s06 g736677 ( .a(n_43281), .b(n_43229), .o(n_43413) );
in01s01 g736678 ( .a(n_43095), .o(n_43096) );
in01s01 g736679 ( .a(n_43075), .o(n_43095) );
ao12f04 g736680 ( .a(n_43023), .b(n_43028), .c(n_43043), .o(n_43075) );
in01s01 g736681 ( .a(n_43116), .o(n_43117) );
in01s01 g736682 ( .a(n_43094), .o(n_43116) );
ao12f02 g736683 ( .a(n_43033), .b(n_43039), .c(n_43051), .o(n_43094) );
na02s02 g736684 ( .a(n_43469), .b(n_43472), .o(n_43562) );
ao22s01 g736686 ( .a(n_43055), .b(n_43041), .c(n_43056), .d(n_43040), .o(n_43115) );
ao22s01 g736687 ( .a(n_43065), .b(n_43072), .c(n_43064), .d(n_43050), .o(n_43151) );
na02s01 g736688 ( .a(n_43401), .b(n_43350), .o(n_43437) );
no02s01 g736689 ( .a(n_43471), .b(n_43470), .o(n_43472) );
na02s01 g736690 ( .a(n_43278), .b(n_43315), .o(n_43331) );
no02s01 g736692 ( .a(n_43465), .b(n_43451), .o(n_43522) );
no02s03 g736693 ( .a(n_43366), .b(n_43292), .o(n_43367) );
no02s06 g736694 ( .a(n_43234), .b(n_43150), .o(n_43235) );
na02s06 g736695 ( .a(n_43363), .b(n_43433), .o(n_43434) );
no02s03 g736696 ( .a(n_43323), .b(n_43360), .o(n_43408) );
in01s01 g736697 ( .a(n_43468), .o(n_43469) );
na02s02 g736698 ( .a(n_43432), .b(n_43358), .o(n_43468) );
in01s02 g736699 ( .a(n_43329), .o(n_43330) );
no02m06 g736700 ( .a(n_43225), .b(n_43188), .o(n_43329) );
no02s06 g736701 ( .a(n_43285), .b(n_43185), .o(n_43286) );
na02s08 g736702 ( .a(n_43222), .b(n_43274), .o(n_43328) );
no02s06 TIMEBOOST_cell_3204 ( .a(n_39551), .b(n_45840), .o(TIMEBOOST_net_893) );
no02s01 TIMEBOOST_cell_8472 ( .a(n_6816), .b(n_6828), .o(TIMEBOOST_net_2723) );
na02s02 g736705 ( .a(n_43182), .b(FE_OCPN878_n_43022), .o(n_43284) );
no03m08 TIMEBOOST_cell_8217 ( .a(TIMEBOOST_net_600), .b(n_37609), .c(TIMEBOOST_net_2379), .o(n_37707) );
na02s02 g736707 ( .a(n_43269), .b(FE_OCPN878_n_43022), .o(n_43365) );
na02s01 TIMEBOOST_cell_1024 ( .a(TIMEBOOST_net_126), .b(n_1869), .o(n_1928) );
in01s01 g736709 ( .a(n_43405), .o(n_43406) );
na02f06 TIMEBOOST_cell_7957 ( .a(TIMEBOOST_net_2609), .b(n_10665), .o(n_10666) );
no02s20 TIMEBOOST_cell_1026 ( .a(TIMEBOOST_net_127), .b(n_12401), .o(n_12445) );
na02s03 TIMEBOOST_cell_980 ( .a(TIMEBOOST_net_104), .b(n_23313), .o(n_23336) );
no03f06 TIMEBOOST_cell_2374 ( .a(FE_RN_752_0), .b(n_38063), .c(FE_RN_757_0), .o(FE_RN_759_0) );
na02m01 g736714 ( .a(n_43314), .b(FE_OCP_RBN6191_n_43103), .o(n_43404) );
no02s02 g736715 ( .a(n_43346), .b(FE_OCP_RBN4478_FE_OCPN913_n_43230), .o(n_43431) );
na02s02 g736716 ( .a(n_43313), .b(FE_OCP_RBN6191_n_43103), .o(n_43473) );
na02m01 TIMEBOOST_cell_6311 ( .a(n_36032), .b(n_36033), .o(TIMEBOOST_net_2007) );
na02s10 TIMEBOOST_cell_8461 ( .a(n_6619), .b(TIMEBOOST_net_2717), .o(TIMEBOOST_net_2) );
in01s01 g736719 ( .a(n_43282), .o(n_43283) );
no02s02 TIMEBOOST_cell_4500 ( .a(TIMEBOOST_net_1340), .b(n_11620), .o(n_11749) );
na02f08 TIMEBOOST_cell_7439 ( .a(TIMEBOOST_net_2350), .b(FE_OCP_RBN2443_n_44798), .o(n_40852) );
in01s01 g736722 ( .a(n_43281), .o(n_43372) );
na02s03 g736723 ( .a(n_43139), .b(n_43228), .o(n_43281) );
na02s03 g736724 ( .a(n_43138), .b(n_43228), .o(n_43229) );
no02s01 g736725 ( .a(n_43042), .b(n_43029), .o(n_43074) );
no02s01 g736726 ( .a(n_43072), .b(n_43027), .o(n_43073) );
na02s06 g736727 ( .a(n_43092), .b(n_43087), .o(n_43234) );
no02s01 g736728 ( .a(n_43200), .b(n_43136), .o(n_43227) );
na02s02 g736729 ( .a(n_43183), .b(n_43149), .o(n_43150) );
na02s02 g736730 ( .a(n_43213), .b(n_43226), .o(n_43692) );
no02s02 g736731 ( .a(n_43280), .b(n_43255), .o(n_43433) );
no02s01 g736732 ( .a(n_43325), .b(n_43270), .o(n_43326) );
no02s01 g736733 ( .a(n_43361), .b(n_43362), .o(n_43363) );
in01s01 g736735 ( .a(n_43360), .o(n_43401) );
na02s02 g736736 ( .a(n_43306), .b(n_43324), .o(n_43360) );
na02s01 g736737 ( .a(n_43350), .b(n_43303), .o(n_43323) );
no02s02 g736738 ( .a(n_43342), .b(n_43359), .o(n_43432) );
no02s02 g736739 ( .a(n_43357), .b(n_43356), .o(n_43358) );
na02s02 g736740 ( .a(n_43389), .b(n_43400), .o(n_43471) );
no02s01 g736741 ( .a(n_43152), .b(n_43085), .o(n_43091) );
in01s01 g736743 ( .a(n_43225), .o(n_43278) );
na02s02 g736744 ( .a(n_43165), .b(n_43189), .o(n_43225) );
na02m04 g736745 ( .a(n_43187), .b(n_43315), .o(n_43188) );
na02s06 g736746 ( .a(n_43355), .b(n_43339), .o(n_43435) );
in01s01 g736747 ( .a(n_43465), .o(n_43466) );
na02s02 g736748 ( .a(n_43430), .b(n_43429), .o(n_43465) );
na02s01 g736749 ( .a(n_43197), .b(n_43144), .o(n_43224) );
na02s02 g736750 ( .a(n_43553), .b(n_43186), .o(n_43285) );
na02s06 g736751 ( .a(n_43529), .b(n_43113), .o(n_43114) );
no02s01 g736752 ( .a(n_43276), .b(n_43174), .o(n_43277) );
na02s06 g736753 ( .a(n_43184), .b(n_43217), .o(n_43185) );
in01s01 g736754 ( .a(n_43274), .o(n_43275) );
no02s03 g736755 ( .a(n_43205), .b(n_43223), .o(n_43274) );
no02s04 g736756 ( .a(n_43202), .b(n_43204), .o(n_43222) );
na02s06 g736757 ( .a(n_43273), .b(n_43260), .o(n_43366) );
in01s01 g736758 ( .a(n_43220), .o(n_43221) );
na02s01 g736759 ( .a(n_43110), .b(n_43183), .o(n_43220) );
na02m04 g736760 ( .a(n_43054), .b(n_46943), .o(n_43045) );
na02s04 g736761 ( .a(n_43062), .b(n_43070), .o(n_43071) );
no02f08 TIMEBOOST_cell_3203 ( .a(TIMEBOOST_net_892), .b(FE_OCP_RBN4363_n_39584), .o(n_39633) );
in01s01 g736763 ( .a(n_43321), .o(n_43322) );
no02s01 g736764 ( .a(n_43272), .b(n_43271), .o(n_43321) );
in01s01 g736765 ( .a(n_43353), .o(n_43354) );
na02s01 g736766 ( .a(FE_RN_1819_0), .b(n_43320), .o(n_43353) );
na02s04 TIMEBOOST_cell_6033 ( .a(FE_RN_852_0), .b(FE_RN_851_0), .o(TIMEBOOST_net_1868) );
na02s01 g736768 ( .a(n_43320), .b(n_43181), .o(n_43182) );
in01s01 g736769 ( .a(n_43560), .o(n_43561) );
na02s01 g736770 ( .a(n_43521), .b(n_43307), .o(n_43560) );
in01s01 g736771 ( .a(n_43318), .o(n_43319) );
no02s01 g736772 ( .a(n_43361), .b(n_43270), .o(n_43318) );
in01s01 g736773 ( .a(n_43055), .o(n_43056) );
na02s01 g736774 ( .a(n_43043), .b(n_43024), .o(n_43055) );
no02s01 g736776 ( .a(n_43352), .b(n_43351), .o(n_43398) );
na02m06 TIMEBOOST_cell_7788 ( .a(n_34282), .b(n_34728), .o(TIMEBOOST_net_2525) );
na02s02 g736778 ( .a(n_43254), .b(n_43251), .o(n_43269) );
in01s01 g736779 ( .a(n_43396), .o(n_43397) );
na02s01 g736780 ( .a(n_43305), .b(n_43350), .o(n_43396) );
in01s01 g736781 ( .a(n_43394), .o(n_43395) );
no02s01 g736782 ( .a(n_43359), .b(n_43349), .o(n_43394) );
na02s01 TIMEBOOST_cell_1023 ( .a(n_1601), .b(n_1580), .o(TIMEBOOST_net_126) );
in01s01 g736784 ( .a(n_43427), .o(n_43428) );
na02s01 g736785 ( .a(n_43341), .b(n_43393), .o(n_43427) );
na02m04 TIMEBOOST_cell_5527 ( .a(TIMEBOOST_net_1711), .b(n_6053), .o(n_6146) );
in01s01 g736787 ( .a(n_43558), .o(n_43559) );
na02s01 g736788 ( .a(n_43389), .b(n_43520), .o(n_43558) );
in01s01 g736789 ( .a(n_43556), .o(n_43557) );
na02s01 g736790 ( .a(n_43519), .b(n_43087), .o(n_43556) );
in01s01 g736791 ( .a(n_43068), .o(n_43069) );
na02s01 g736792 ( .a(n_43054), .b(n_43036), .o(n_43068) );
no02s10 TIMEBOOST_cell_1025 ( .a(n_12136), .b(n_12402), .o(TIMEBOOST_net_127) );
in01s01 g736794 ( .a(n_43554), .o(n_43555) );
na02s01 g736795 ( .a(n_43518), .b(n_43385), .o(n_43554) );
in01s01 g736796 ( .a(n_43145), .o(n_43146) );
na02s01 g736797 ( .a(n_43111), .b(n_43062), .o(n_43145) );
na02s01 TIMEBOOST_cell_979 ( .a(n_23031), .b(n_23335), .o(TIMEBOOST_net_104) );
in01s01 g736799 ( .a(n_43347), .o(n_43348) );
na02s01 g736800 ( .a(n_43247), .b(n_43315), .o(n_43347) );
no02f02 TIMEBOOST_cell_2133 ( .a(n_5773), .b(n_5836), .o(TIMEBOOST_net_681) );
in01s01 g736802 ( .a(n_43425), .o(n_43426) );
no02s01 g736803 ( .a(n_43391), .b(n_43390), .o(n_43425) );
in01s01 g736804 ( .a(n_43516), .o(n_43517) );
no02s01 g736805 ( .a(n_43464), .b(n_43387), .o(n_43516) );
na02s01 g736806 ( .a(n_43297), .b(n_46936), .o(n_43314) );
no02s01 g736807 ( .a(n_43464), .b(n_43001), .o(n_43346) );
in01s01 g736808 ( .a(n_43462), .o(n_43463) );
na02s01 g736809 ( .a(n_43424), .b(n_43429), .o(n_43462) );
in01s01 g736810 ( .a(n_43089), .o(n_43090) );
no02s01 g736811 ( .a(n_43067), .b(n_43066), .o(n_43089) );
na02s01 g736812 ( .a(n_43424), .b(n_46935), .o(n_43313) );
in01s01 g736813 ( .a(n_43177), .o(n_43178) );
na02s01 g736814 ( .a(n_43144), .b(n_43113), .o(n_43177) );
in01s01 g736815 ( .a(n_43621), .o(n_43622) );
na02s01 g736816 ( .a(n_43490), .b(n_43553), .o(n_43621) );
in01s01 g736817 ( .a(n_43263), .o(n_43264) );
na02s01 g736818 ( .a(n_43133), .b(n_43217), .o(n_43263) );
na02s06 g736819 ( .a(n_43048), .b(n_43052), .o(n_43053) );
na02m08 g736820 ( .a(n_43144), .b(n_43130), .o(n_43143) );
na02s06 g736821 ( .a(n_43133), .b(n_43129), .o(n_43142) );
in01s01 g736822 ( .a(n_43261), .o(n_43262) );
no02s01 g736823 ( .a(n_43223), .b(n_43216), .o(n_43261) );
no02s04 TIMEBOOST_cell_5299 ( .a(TIMEBOOST_net_1597), .b(n_4125), .o(n_4294) );
in01s01 g736825 ( .a(n_43344), .o(n_43345) );
no02s01 g736826 ( .a(n_43204), .b(n_43311), .o(n_43344) );
na02s04 g736827 ( .a(n_43127), .b(n_42906), .o(n_43140) );
in01s01 g736828 ( .a(n_43551), .o(n_43552) );
na02s01 g736829 ( .a(n_43515), .b(n_43126), .o(n_43551) );
na02s02 g736830 ( .a(n_43126), .b(n_46940), .o(n_43139) );
in01s01 g736831 ( .a(n_43309), .o(n_43310) );
na02s01 g736832 ( .a(n_43260), .b(n_43125), .o(n_43309) );
in01s01 g736833 ( .a(n_43064), .o(n_43065) );
na02s01 g736834 ( .a(n_43034), .b(n_43051), .o(n_43064) );
na02s02 g736835 ( .a(n_43125), .b(n_46939), .o(n_43138) );
in01s01 g736836 ( .a(n_43258), .o(n_43259) );
no02s01 g736837 ( .a(n_43215), .b(n_43214), .o(n_43258) );
no02s01 g736838 ( .a(FE_OCP_RBN4402_n_43013), .b(n_43016), .o(n_43029) );
no02s01 g736839 ( .a(n_43018), .b(n_42249), .o(n_43042) );
in01s01 g736840 ( .a(n_43040), .o(n_43041) );
in01s01 g736841 ( .a(n_43028), .o(n_43040) );
no02f02 g736842 ( .a(n_43013), .b(n_43016), .o(n_43028) );
no02s01 g736843 ( .a(n_43026), .b(n_43025), .o(n_43027) );
in01s01 g736844 ( .a(n_43072), .o(n_43050) );
in01s01 g736845 ( .a(n_43039), .o(n_43072) );
na02f02 g736846 ( .a(n_43026), .b(n_43025), .o(n_43039) );
in01s01 g736847 ( .a(n_43549), .o(n_43550) );
na02s01 g736848 ( .a(n_43461), .b(n_43149), .o(n_43549) );
in01s01 g736849 ( .a(n_43547), .o(n_43548) );
na02s01 g736850 ( .a(n_43460), .b(n_43226), .o(n_43547) );
in01s01 g736851 ( .a(n_43545), .o(n_43546) );
na02s01 g736852 ( .a(n_43514), .b(n_43458), .o(n_43545) );
in01s01 g736853 ( .a(n_43619), .o(n_43620) );
no02s01 g736854 ( .a(n_43280), .b(n_43511), .o(n_43619) );
in01s01 g736855 ( .a(n_43617), .o(n_43618) );
na03f08 TIMEBOOST_cell_8432 ( .a(n_6386), .b(n_6354), .c(FE_OCP_RBN3404_n_6205), .o(n_6416) );
in01s01 g736857 ( .a(n_43543), .o(n_43544) );
na02s01 g736858 ( .a(n_43324), .b(n_43456), .o(n_43543) );
in01s01 g736859 ( .a(n_43615), .o(n_43616) );
no02s01 g736860 ( .a(n_43504), .b(n_43449), .o(n_43615) );
in01s01 g736861 ( .a(n_43613), .o(n_43614) );
no02s01 g736862 ( .a(n_43304), .b(n_43508), .o(n_43613) );
in01s01 g736863 ( .a(n_43541), .o(n_43542) );
na02s01 g736864 ( .a(n_43343), .b(n_43455), .o(n_43541) );
in01s01 g736865 ( .a(n_43611), .o(n_43612) );
no02s01 g736866 ( .a(n_43356), .b(n_43505), .o(n_43611) );
in01s01 g736867 ( .a(n_43539), .o(n_43540) );
na02s01 g736868 ( .a(n_43400), .b(n_43454), .o(n_43539) );
in01s01 g736869 ( .a(n_43609), .o(n_43610) );
no02m04 TIMEBOOST_cell_4459 ( .a(n_21573), .b(FE_OCP_RBN3245_n_21351), .o(TIMEBOOST_net_1320) );
in01s01 g736871 ( .a(n_43607), .o(n_43608) );
no02s01 g736872 ( .a(n_43507), .b(n_43538), .o(n_43607) );
in01s01 g736873 ( .a(n_43536), .o(n_43537) );
na02s01 g736874 ( .a(n_43453), .b(n_43092), .o(n_43536) );
in01s01 g736875 ( .a(FE_OCPN1228_n_43605), .o(n_43606) );
no02s04 TIMEBOOST_cell_5376 ( .a(n_21742), .b(n_21552), .o(TIMEBOOST_net_1636) );
in01s01 g736877 ( .a(n_43603), .o(n_43604) );
na02s01 g736878 ( .a(n_43355), .b(n_43501), .o(n_43603) );
in01s01 g736879 ( .a(n_43601), .o(n_43602) );
na02s01 g736880 ( .a(n_43523), .b(n_43500), .o(n_43601) );
in01s01 g736881 ( .a(n_43599), .o(n_43600) );
na02s01 g736882 ( .a(n_43430), .b(n_43499), .o(n_43599) );
in01s01 g736883 ( .a(n_43597), .o(n_43598) );
na02s01 g736884 ( .a(n_43452), .b(n_43497), .o(n_43597) );
in01s01 g736885 ( .a(n_43595), .o(n_43596) );
oa12s01 g736886 ( .a(n_43192), .b(FE_OCP_RBN4478_FE_OCPN913_n_43230), .c(n_43052), .o(n_43595) );
in01s01 g736887 ( .a(n_43593), .o(n_43594) );
na02s01 g736888 ( .a(n_43493), .b(n_43529), .o(n_43593) );
in01s01 g736889 ( .a(n_43591), .o(n_43592) );
na02s01 g736890 ( .a(n_43492), .b(n_43530), .o(n_43591) );
in01s01 g736891 ( .a(n_43589), .o(n_43590) );
na02s01 g736892 ( .a(n_43488), .b(n_43186), .o(n_43589) );
in01s01 g736893 ( .a(n_43587), .o(n_43588) );
na02s01 g736894 ( .a(n_43486), .b(n_43184), .o(n_43587) );
in01s01 g736895 ( .a(n_43585), .o(n_43586) );
na02s01 g736896 ( .a(n_43485), .b(n_43206), .o(n_43585) );
in01s01 g736897 ( .a(n_43583), .o(n_43584) );
na02s01 g736898 ( .a(n_43203), .b(n_43484), .o(n_43583) );
in01s01 g736899 ( .a(n_43581), .o(n_43582) );
na02s01 g736900 ( .a(n_43293), .b(n_43483), .o(n_43581) );
in01s01 g736901 ( .a(n_43579), .o(n_43580) );
na02s01 g736902 ( .a(n_43189), .b(n_43482), .o(n_43579) );
in01s01 g736903 ( .a(n_43533), .o(n_43534) );
oa22s01 g736904 ( .a(FE_OCP_RBN3312_n_43022), .b(n_42967), .c(FE_OCP_RBN3315_n_43022), .d(FE_OCP_RBN3321_n_42959), .o(n_43533) );
in01s01 g736905 ( .a(n_43577), .o(n_43578) );
oa22s01 g736906 ( .a(FE_OCP_RBN3312_n_43022), .b(n_43158), .c(FE_OCP_RBN3315_n_43022), .d(n_46943), .o(n_43577) );
in01s01 g736907 ( .a(n_43634), .o(n_43635) );
oa22s01 g736908 ( .a(FE_OCP_RBN6191_n_43103), .b(n_42946), .c(FE_OCP_RBN4478_FE_OCPN913_n_43230), .d(n_42961), .o(n_43634) );
in01s01 g736909 ( .a(n_43632), .o(n_43633) );
oa22s01 g736910 ( .a(FE_OCP_RBN6191_n_43103), .b(n_43494), .c(FE_OCP_RBN4479_FE_OCPN913_n_43230), .d(n_43121), .o(n_43632) );
in01s01 g736911 ( .a(n_43630), .o(n_43631) );
oa22s01 g736912 ( .a(FE_OCP_RBN6192_n_43103), .b(n_42936), .c(FE_OCP_RBN4476_FE_OCPN913_n_43230), .d(n_46940), .o(n_43630) );
in01s01 g736914 ( .a(n_43110), .o(n_43136) );
na02s02 g736915 ( .a(FE_OCP_RBN3306_n_43022), .b(n_42802), .o(n_43110) );
na02s02 g736916 ( .a(FE_OCP_RBN3311_n_43022), .b(n_42803), .o(n_43183) );
no02s01 g736917 ( .a(FE_OCP_RBN3306_n_43022), .b(n_42748), .o(n_43538) );
no02s06 g736918 ( .a(FE_OCP_RBN3306_n_43022), .b(n_42730), .o(n_43449) );
na02s06 g736919 ( .a(FE_OCP_RBN3310_n_43022), .b(n_43037), .o(n_43385) );
in01s01 g736920 ( .a(n_43023), .o(n_43024) );
no02m04 g736921 ( .a(n_43015), .b(n_43014), .o(n_43023) );
in01s01 g736922 ( .a(n_43035), .o(n_43036) );
no02s06 g736923 ( .a(n_43022), .b(n_43021), .o(n_43035) );
na02m04 g736924 ( .a(n_43015), .b(n_43014), .o(n_43043) );
na02s04 g736925 ( .a(n_43022), .b(n_43021), .o(n_43054) );
na02s06 g736926 ( .a(FE_OCP_RBN3309_n_43022), .b(n_42668), .o(n_43111) );
in01s01 g736928 ( .a(n_43087), .o(n_43108) );
na02s02 g736929 ( .a(FE_OCP_RBN3311_n_43022), .b(n_42792), .o(n_43087) );
in01s01 g736931 ( .a(n_43062), .o(n_43085) );
na02s06 g736932 ( .a(FE_OCP_RBN3306_n_43022), .b(n_46944), .o(n_43062) );
na02s02 g736933 ( .a(FE_OCP_RBN3311_n_43022), .b(n_46942), .o(n_43092) );
na02s02 g736934 ( .a(FE_OCP_RBN3311_n_43022), .b(n_43106), .o(n_43149) );
na02s01 g736935 ( .a(FE_OCP_RBN4446_n_43022), .b(n_42805), .o(n_43461) );
in01s01 g736936 ( .a(n_43213), .o(n_43272) );
na02s02 g736937 ( .a(FE_OCP_RBN3311_n_43022), .b(n_46941), .o(n_43213) );
no02s02 g736938 ( .a(FE_OCP_RBN3311_n_43022), .b(n_46941), .o(n_43271) );
na02s01 g736939 ( .a(FE_OCP_RBN4446_n_43022), .b(n_43147), .o(n_43460) );
na02s02 g736940 ( .a(FE_OCP_RBN3311_n_43022), .b(n_42829), .o(n_43226) );
no02s01 g736942 ( .a(FE_OCPN878_n_43022), .b(n_43135), .o(n_43256) );
na02s01 g736943 ( .a(FE_OCP_RBN3306_n_43022), .b(n_43135), .o(n_43320) );
na02s01 g736944 ( .a(FE_OCP_RBN4446_n_43022), .b(n_42883), .o(n_43458) );
na02s01 g736945 ( .a(FE_OCP_RBN3311_n_43022), .b(n_43181), .o(n_43514) );
in01s01 g736947 ( .a(n_43255), .o(n_43307) );
no02s02 g736948 ( .a(FE_OCPN878_n_43022), .b(n_43211), .o(n_43255) );
na02s01 g736949 ( .a(FE_OCP_RBN4446_n_43022), .b(n_43211), .o(n_43521) );
no02s01 g736950 ( .a(FE_OCPN878_n_43022), .b(n_42941), .o(n_43280) );
no02s01 g736951 ( .a(FE_OCP_RBN3307_n_43022), .b(n_42926), .o(n_43511) );
no02s02 g736952 ( .a(FE_OCP_RBN3311_n_43022), .b(n_42924), .o(n_43270) );
no02s01 g736953 ( .a(FE_OCPN878_n_43022), .b(n_42925), .o(n_43361) );
no02s02 TIMEBOOST_cell_7651 ( .a(TIMEBOOST_net_2456), .b(n_2957), .o(n_3076) );
no02s02 g736955 ( .a(FE_OCPN878_n_43022), .b(n_46938), .o(n_43362) );
na02s01 g736956 ( .a(FE_OCP_RBN3312_n_43022), .b(n_42714), .o(n_43518) );
in01s01 g736957 ( .a(n_43254), .o(n_43352) );
na02s01 g736958 ( .a(FE_OCPN878_n_43022), .b(n_42922), .o(n_43254) );
in01s01 g736959 ( .a(n_43306), .o(n_43351) );
na02s01 g736960 ( .a(FE_OCP_RBN3311_n_43022), .b(n_42923), .o(n_43306) );
na02s02 g736961 ( .a(FE_OCP_RBN3307_n_43022), .b(n_43251), .o(n_43324) );
na02s01 g736962 ( .a(FE_OCP_RBN4446_n_43022), .b(n_42969), .o(n_43456) );
in01s01 g736963 ( .a(n_43316), .o(n_43305) );
no02s01 g736964 ( .a(FE_OCP_RBN3307_n_43022), .b(n_43250), .o(n_43316) );
na02s01 g736965 ( .a(FE_OCP_RBN3307_n_43022), .b(n_43250), .o(n_43350) );
in01s01 g736966 ( .a(n_43303), .o(n_43304) );
na02s01 g736967 ( .a(FE_OCP_RBN3307_n_43022), .b(n_42968), .o(n_43303) );
no02s01 g736968 ( .a(FE_OCP_RBN3307_n_43022), .b(n_42968), .o(n_43508) );
in01s01 g736969 ( .a(n_43248), .o(n_43349) );
na02s01 g736970 ( .a(FE_OCPN878_n_43022), .b(n_43208), .o(n_43248) );
no02s01 g736971 ( .a(FE_OCPN878_n_43022), .b(n_43208), .o(n_43359) );
in01s01 g736972 ( .a(n_43342), .o(n_43343) );
no02s01 g736973 ( .a(FE_OCPN878_n_43022), .b(n_43300), .o(n_43342) );
na02s01 g736974 ( .a(FE_OCP_RBN3312_n_43022), .b(n_43300), .o(n_43455) );
in01s01 g736975 ( .a(n_43357), .o(n_43341) );
no02s01 g736976 ( .a(FE_OCPN878_n_43022), .b(n_43299), .o(n_43357) );
na02s01 g736977 ( .a(FE_OCPN878_n_43022), .b(n_43299), .o(n_43393) );
no02s01 g736978 ( .a(FE_OCP_RBN3307_n_43022), .b(n_43070), .o(n_43507) );
no02s01 g736979 ( .a(FE_OCP_RBN3307_n_43022), .b(n_42972), .o(n_43505) );
no02s01 g736980 ( .a(FE_OCP_RBN3312_n_43022), .b(n_43298), .o(n_43356) );
no02s01 g736981 ( .a(FE_OCP_RBN3307_n_43022), .b(n_43061), .o(n_43504) );
in01s01 g736983 ( .a(n_43389), .o(n_43422) );
na02s01 g736984 ( .a(FE_OCP_RBN3308_n_43022), .b(n_42982), .o(n_43389) );
na02s01 g736985 ( .a(FE_OCP_RBN3312_n_43022), .b(n_43002), .o(n_43520) );
na02s01 g736986 ( .a(FE_OCP_RBN3312_n_43022), .b(n_43003), .o(n_43454) );
na02s02 g736987 ( .a(FE_OCP_RBN3308_n_43022), .b(n_42997), .o(n_43400) );
na02s01 g736988 ( .a(FE_OCP_RBN4446_n_43022), .b(n_42774), .o(n_43453) );
na02m08 TIMEBOOST_cell_4458 ( .a(TIMEBOOST_net_1319), .b(n_21703), .o(n_21786) );
no02s01 g736990 ( .a(n_43388), .b(FE_OCP_RBN3312_n_43022), .o(n_43470) );
na02s01 g736991 ( .a(FE_OCP_RBN4446_n_43022), .b(n_42771), .o(n_43519) );
in01s01 g736992 ( .a(n_43266), .o(n_43247) );
no02s02 g736993 ( .a(FE_OCP_RBN3375_n_43046), .b(n_43134), .o(n_43266) );
na02s02 g736994 ( .a(FE_OCP_RBN3375_n_43046), .b(n_43134), .o(n_43315) );
no02m08 TIMEBOOST_cell_5382 ( .a(FE_OCP_RBN6077_n_16084), .b(n_14730), .o(TIMEBOOST_net_1639) );
na02m02 g736996 ( .a(FE_OCP_RBN4456_n_43103), .b(n_42989), .o(n_43187) );
in01s01 g736997 ( .a(n_43297), .o(n_43391) );
na02s06 g736998 ( .a(FE_OCP_RBN6191_n_43103), .b(n_42954), .o(n_43297) );
in01s01 g736999 ( .a(n_43339), .o(n_43390) );
na02s01 g737000 ( .a(FE_OCP_RBN4456_n_43103), .b(n_42955), .o(n_43339) );
na02s01 g737001 ( .a(FE_OCP_RBN6191_n_43103), .b(n_42994), .o(n_43501) );
na02s06 g737002 ( .a(FE_OCP_RBN4479_FE_OCPN913_n_43230), .b(n_46936), .o(n_43355) );
no02s01 g737003 ( .a(FE_OCP_RBN4456_n_43103), .b(n_42992), .o(n_43464) );
in01s01 g737005 ( .a(n_43387), .o(n_43420) );
no02m01 g737006 ( .a(n_42993), .b(FE_OCP_RBN6191_n_43103), .o(n_43387) );
na02s01 g737007 ( .a(FE_OCP_RBN6191_n_43103), .b(n_43001), .o(n_43500) );
na02m01 g737008 ( .a(n_43007), .b(FE_OCP_RBN4478_FE_OCPN913_n_43230), .o(n_43523) );
na02m01 g737009 ( .a(n_42991), .b(FE_OCP_RBN4478_FE_OCPN913_n_43230), .o(n_43429) );
na02s01 g737010 ( .a(FE_OCP_RBN6191_n_43103), .b(n_43010), .o(n_43499) );
na02s01 g737011 ( .a(FE_OCP_RBN4478_FE_OCPN913_n_43230), .b(n_46935), .o(n_43430) );
na02s01 g737012 ( .a(FE_OCP_RBN6191_n_43103), .b(n_43418), .o(n_43497) );
in01s01 g737013 ( .a(n_43451), .o(n_43452) );
no02s01 g737014 ( .a(FE_OCP_RBN6191_n_43103), .b(n_43418), .o(n_43451) );
na02s01 g737015 ( .a(FE_OCP_RBN6191_n_43103), .b(n_43494), .o(n_43495) );
na02s01 g737016 ( .a(FE_OCP_RBN6191_n_43103), .b(n_42596), .o(n_43493) );
na02s01 g737017 ( .a(FE_OCP_RBN6192_n_43103), .b(n_42666), .o(n_43492) );
in01s01 g737018 ( .a(n_43489), .o(n_43490) );
no02s01 g737019 ( .a(FE_OCP_RBN4477_FE_OCPN913_n_43230), .b(n_43132), .o(n_43489) );
na02s01 g737020 ( .a(FE_OCP_RBN6192_n_43103), .b(n_42750), .o(n_43488) );
in01s01 g737022 ( .a(n_43133), .o(n_43174) );
na02s03 g737023 ( .a(n_43103), .b(n_42772), .o(n_43133) );
na02s06 g737024 ( .a(FE_OCP_RBN4456_n_43103), .b(n_42773), .o(n_43217) );
na02s02 g737025 ( .a(n_43030), .b(n_42780), .o(n_43186) );
na02s02 g737026 ( .a(n_43030), .b(n_43132), .o(n_43553) );
no02s02 g737027 ( .a(n_43032), .b(n_43031), .o(n_43066) );
in01s01 g737028 ( .a(n_43033), .o(n_43034) );
no02s02 g737029 ( .a(n_43020), .b(n_43019), .o(n_43033) );
na02s02 g737030 ( .a(n_43020), .b(n_43019), .o(n_43051) );
na02s06 g737031 ( .a(n_43030), .b(n_43052), .o(n_43192) );
na02s02 g737032 ( .a(FE_OCP_RBN3373_n_43046), .b(n_43121), .o(n_43084) );
na02s02 g737033 ( .a(n_43030), .b(n_43083), .o(n_43529) );
na02s06 g737034 ( .a(FE_OCP_RBN3373_n_43046), .b(n_42597), .o(n_43113) );
in01s01 g737035 ( .a(n_43048), .o(n_43067) );
na02s04 g737036 ( .a(n_43032), .b(n_43031), .o(n_43048) );
na02s03 g737037 ( .a(FE_OCP_RBN3372_n_43046), .b(n_43130), .o(n_43530) );
na02s08 g737038 ( .a(n_43046), .b(n_42598), .o(n_43144) );
na02s01 g737039 ( .a(FE_OCP_RBN6192_n_43103), .b(n_42804), .o(n_43486) );
na02s02 g737040 ( .a(FE_OCP_RBN3372_n_43046), .b(n_43129), .o(n_43184) );
in01s01 g737041 ( .a(n_43128), .o(n_43216) );
na02s02 g737042 ( .a(n_43046), .b(n_43104), .o(n_43128) );
no02s02 g737043 ( .a(n_43171), .b(n_43104), .o(n_43223) );
na02s01 g737044 ( .a(FE_OCP_RBN6192_n_43103), .b(n_43172), .o(n_43485) );
in01s01 g737045 ( .a(n_43205), .o(n_43206) );
no02s02 g737046 ( .a(n_43171), .b(n_43172), .o(n_43205) );
in01s01 g737047 ( .a(n_43127), .o(n_43311) );
na02s03 g737048 ( .a(n_43103), .b(n_43102), .o(n_43127) );
in01s01 g737050 ( .a(n_43204), .o(n_43245) );
no02s02 g737051 ( .a(n_43171), .b(n_43102), .o(n_43204) );
na02s01 g737052 ( .a(FE_OCP_RBN6192_n_43103), .b(n_43170), .o(n_43484) );
in01s01 g737053 ( .a(n_43202), .o(n_43203) );
no02s02 g737054 ( .a(n_43171), .b(n_43170), .o(n_43202) );
in01s01 g737056 ( .a(n_43126), .o(n_43168) );
na02s02 g737057 ( .a(n_43046), .b(n_42956), .o(n_43126) );
na02s03 g737058 ( .a(FE_OCP_RBN4476_FE_OCPN913_n_43230), .b(n_42878), .o(n_43515) );
in01s01 g737060 ( .a(n_43125), .o(n_43166) );
na02s02 g737061 ( .a(n_43046), .b(n_42910), .o(n_43125) );
na02s02 g737062 ( .a(FE_OCP_RBN3374_n_43046), .b(n_42911), .o(n_43260) );
na02m01 g737063 ( .a(FE_OCP_RBN6191_n_43103), .b(n_42990), .o(n_43424) );
na02s01 g737064 ( .a(FE_OCP_RBN6192_n_43103), .b(n_43243), .o(n_43483) );
in01s01 g737065 ( .a(n_43292), .o(n_43293) );
no02s02 g737066 ( .a(n_43243), .b(FE_OCP_RBN6192_n_43103), .o(n_43292) );
no02s02 g737067 ( .a(FE_OCP_RBN3374_n_43046), .b(n_43123), .o(n_43215) );
in01s01 g737068 ( .a(n_43165), .o(n_43214) );
na02s02 g737069 ( .a(FE_OCP_RBN4456_n_43103), .b(n_43123), .o(n_43165) );
na02s01 g737070 ( .a(FE_OCP_RBN6192_n_43103), .b(n_43179), .o(n_43482) );
na02s02 g737071 ( .a(FE_OCP_RBN3374_n_43046), .b(n_46937), .o(n_43189) );
in01s01 g737073 ( .a(n_43164), .o(n_43200) );
na02s02 g737074 ( .a(FE_OCP_RBN3306_n_43022), .b(n_42794), .o(n_43164) );
ao12s02 g737075 ( .a(FE_OCP_RBN3310_n_43022), .b(n_43061), .c(n_43037), .o(n_43152) );
in01s01 g737076 ( .a(n_43325), .o(n_43291) );
no02s02 g737077 ( .a(FE_OCP_RBN3307_n_43022), .b(n_42942), .o(n_43325) );
in01s01 g737078 ( .a(n_43383), .o(n_43384) );
no02s01 TIMEBOOST_cell_5516 ( .a(n_36009), .b(n_36010), .o(TIMEBOOST_net_1706) );
in01s01 g737080 ( .a(n_43199), .o(n_43276) );
na02s02 g737081 ( .a(n_43103), .b(n_42781), .o(n_43199) );
in01s01 g737083 ( .a(n_43162), .o(n_43197) );
na02s02 g737085 ( .a(FE_OCP_RBN4456_n_43103), .b(n_42957), .o(n_43273) );
in01s01 g737086 ( .a(FE_OCP_RBN4402_n_43013), .o(n_43018) );
oa22f01 g737088 ( .a(FE_OCP_RBN3258_n_42998), .b(delay_sub_ln23_0_unr30_stage10_stallmux_q), .c(n_42998), .d(n_43012), .o(n_43013) );
ao22f01 g737089 ( .a(n_43011), .b(n_43012), .c(n_43000), .d(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n_43026) );
in01s04 g737128 ( .a(n_43015), .o(n_43022) );
na02m06 g737129 ( .a(FE_OCP_RBN3257_n_42998), .b(n_43012), .o(n_43015) );
in01s03 g737131 ( .a(n_43030), .o(n_43171) );
in01s01 g737138 ( .a(FE_OCP_RBN3374_n_43046), .o(n_43228) );
in01s10 g737168 ( .a(n_43030), .o(n_43103) );
in01s10 g737170 ( .a(n_43030), .o(n_43046) );
in01s10 g737171 ( .a(n_43032), .o(n_43030) );
in01s08 g737172 ( .a(n_43020), .o(n_43032) );
no02s08 g737173 ( .a(n_43011), .b(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n_43020) );
no02s06 TIMEBOOST_cell_6366 ( .a(TIMEBOOST_net_2034), .b(n_17195), .o(n_17343) );
in01s01 g737176 ( .a(n_43001), .o(n_43007) );
oa22s01 g737177 ( .a(n_42974), .b(n_42693), .c(n_42973), .d(n_42694), .o(n_43001) );
in01s01 g737178 ( .a(n_46935), .o(n_43010) );
in01s01 g737180 ( .a(n_43006), .o(n_43418) );
ao22s01 g737181 ( .a(n_42984), .b(n_42692), .c(n_42983), .d(n_42691), .o(n_43006) );
no02s01 g737183 ( .a(n_42985), .b(n_42708), .o(n_42996) );
in01s01 g737184 ( .a(n_42989), .o(n_43265) );
ao22s01 g737185 ( .a(n_42934), .b(n_42622), .c(n_42933), .d(n_42623), .o(n_42989) );
no02f06 g737187 ( .a(n_42978), .b(n_42965), .o(n_42998) );
in01s01 g737188 ( .a(n_43003), .o(n_42997) );
na02s01 g737189 ( .a(n_42976), .b(n_42964), .o(n_43003) );
in01s01 g737190 ( .a(n_43388), .o(n_43005) );
no03m06 TIMEBOOST_cell_8404 ( .a(n_11312), .b(n_11482), .c(n_11484), .o(TIMEBOOST_net_571) );
in01f04 g737192 ( .a(n_43000), .o(n_43011) );
na02f06 g737193 ( .a(n_42977), .b(n_42988), .o(n_43000) );
no02f04 g737194 ( .a(n_42947), .b(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n_42965) );
no02f04 g737195 ( .a(n_42946), .b(n_43012), .o(n_42978) );
na02f06 g737196 ( .a(FE_OCP_RBN3320_n_42959), .b(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n_42988) );
na02s04 g737197 ( .a(n_42959), .b(n_43012), .o(n_42977) );
na02s01 g737198 ( .a(n_42948), .b(n_42815), .o(n_42964) );
no02s06 TIMEBOOST_cell_8684 ( .a(FE_OCP_RBN3221_n_21242), .b(n_45070), .o(TIMEBOOST_net_2829) );
no02m08 TIMEBOOST_cell_7621 ( .a(TIMEBOOST_net_2441), .b(n_29319), .o(n_29440) );
na02s01 g737201 ( .a(n_42949), .b(n_42816), .o(n_42976) );
oa12s01 g737203 ( .a(n_42656), .b(n_42975), .c(n_42606), .o(n_42985) );
in01s01 g737204 ( .a(n_42983), .o(n_42984) );
oa12s01 g737205 ( .a(n_42351), .b(n_42975), .c(n_42342), .o(n_42983) );
in01s01 g737206 ( .a(n_42973), .o(n_42974) );
oa12s01 g737207 ( .a(n_42417), .b(n_42927), .c(n_42279), .o(n_42973) );
in01s01 g737208 ( .a(n_46936), .o(n_42994) );
in01s01 g737210 ( .a(n_42992), .o(n_42993) );
ao22s01 g737211 ( .a(n_42938), .b(n_42354), .c(n_42927), .d(n_42353), .o(n_42992) );
in01s01 g737212 ( .a(n_43298), .o(n_42972) );
na02s02 g737213 ( .a(n_42935), .b(n_42920), .o(n_43298) );
in01s01 g737214 ( .a(n_42990), .o(n_42991) );
oa22s01 g737215 ( .a(n_42940), .b(n_42677), .c(n_42975), .d(n_42678), .o(n_42990) );
na02s01 g737216 ( .a(n_42907), .b(n_42797), .o(n_42920) );
na02s01 g737217 ( .a(n_42908), .b(n_42798), .o(n_42935) );
no02s01 g737219 ( .a(n_42928), .b(n_42673), .o(n_42950) );
in01s01 g737220 ( .a(n_42948), .o(n_42949) );
oa12s01 g737221 ( .a(n_42801), .b(n_42902), .c(n_42755), .o(n_42948) );
in01s01 g737222 ( .a(n_42970), .o(n_42971) );
oa12s01 g737223 ( .a(n_42522), .b(n_42902), .c(n_42526), .o(n_42970) );
in01s01 g737224 ( .a(n_42933), .o(n_42934) );
oa12s01 g737225 ( .a(n_42363), .b(n_42888), .c(n_42280), .o(n_42933) );
ao22s01 g737226 ( .a(n_42900), .b(n_42356), .c(n_42888), .d(n_42355), .o(n_43134) );
in01s01 g737227 ( .a(n_43002), .o(n_42982) );
na02s01 g737228 ( .a(n_42932), .b(n_42945), .o(n_43002) );
in01s01 g737229 ( .a(n_43251), .o(n_42969) );
no02s01 g737230 ( .a(n_42931), .b(n_42919), .o(n_43251) );
in01s01 g737232 ( .a(n_42968), .o(n_42980) );
ao22s01 g737233 ( .a(n_42912), .b(n_42800), .c(n_42913), .d(n_42799), .o(n_42968) );
in01s01 g737234 ( .a(n_42962), .o(n_43300) );
ao22s01 g737235 ( .a(n_42894), .b(n_42759), .c(n_42895), .d(n_42758), .o(n_42962) );
in01s01 g737236 ( .a(n_42946), .o(n_42961) );
in01f04 g737238 ( .a(n_42947), .o(n_42946) );
in01s01 g737240 ( .a(FE_OCP_RBN3321_n_42959), .o(n_42967) );
in01s01 g737244 ( .a(n_46937), .o(n_43179) );
na02s01 g737246 ( .a(n_42916), .b(n_42817), .o(n_42932) );
na02s01 g737247 ( .a(n_42902), .b(n_42818), .o(n_42945) );
no02s01 g737248 ( .a(n_42898), .b(n_42765), .o(n_42919) );
no02s01 g737249 ( .a(n_42899), .b(n_42764), .o(n_42931) );
no02s01 g737251 ( .a(n_42914), .b(n_42610), .o(n_42930) );
no02s01 g737252 ( .a(n_42941), .b(n_43211), .o(n_42942) );
na02s01 g737253 ( .a(n_42936), .b(n_42956), .o(n_42957) );
in01s01 g737254 ( .a(n_42975), .o(n_42940) );
no02s01 g737255 ( .a(n_42905), .b(n_42401), .o(n_42975) );
in01s01 g737256 ( .a(n_42907), .o(n_42908) );
oa12s01 g737257 ( .a(n_42486), .b(n_42857), .c(n_42549), .o(n_42907) );
oa12s01 g737259 ( .a(n_42657), .b(n_42918), .c(n_42608), .o(n_42928) );
in01s01 g737261 ( .a(n_42927), .o(n_42938) );
oa12s01 g737262 ( .a(n_42295), .b(n_42918), .c(n_42344), .o(n_42927) );
in01s01 g737263 ( .a(n_42954), .o(n_42955) );
oa22s01 g737264 ( .a(n_42876), .b(n_42679), .c(n_42918), .d(n_42680), .o(n_42954) );
in01s01 g737265 ( .a(n_46938), .o(n_42953) );
oa22s01 g737267 ( .a(n_42871), .b(n_42525), .c(n_42857), .d(n_42524), .o(n_43299) );
in01s01 g737268 ( .a(n_42906), .o(n_43170) );
ao22s01 g737269 ( .a(n_42844), .b(n_42618), .c(n_42845), .d(n_42619), .o(n_42906) );
in01s01 g737270 ( .a(n_46939), .o(n_43243) );
no02s01 g737272 ( .a(n_42918), .b(n_42440), .o(n_42905) );
na02s01 g737274 ( .a(n_42881), .b(n_42760), .o(n_42904) );
no02s01 g737276 ( .a(n_42869), .b(n_42616), .o(n_42890) );
in01s01 g737278 ( .a(n_42902), .o(n_42916) );
ao12s01 g737279 ( .a(n_42591), .b(n_42889), .c(n_42592), .o(n_42902) );
in01s01 g737281 ( .a(n_42888), .o(n_42900) );
oa12s01 g737282 ( .a(n_42299), .b(n_42842), .c(n_42297), .o(n_42888) );
oa12s01 g737284 ( .a(n_42624), .b(n_42842), .c(n_42556), .o(n_42914) );
in01s01 g737285 ( .a(n_42898), .o(n_42899) );
ao12s01 g737286 ( .a(n_42418), .b(n_42847), .c(n_42746), .o(n_42898) );
in01f04 g737287 ( .a(n_42896), .o(n_42897) );
no02s06 TIMEBOOST_cell_816 ( .a(TIMEBOOST_net_22), .b(n_6745), .o(n_6802) );
in01s01 g737289 ( .a(n_42912), .o(n_42913) );
ao12s01 g737290 ( .a(n_42420), .b(n_42864), .c(n_42463), .o(n_42912) );
in01s01 g737291 ( .a(n_42894), .o(n_42895) );
ao12s01 g737292 ( .a(n_42724), .b(n_42889), .c(n_42766), .o(n_42894) );
in01f06 g737293 ( .a(n_42886), .o(n_42887) );
oa12f08 g737294 ( .a(n_42512), .b(n_42860), .c(n_42462), .o(n_42886) );
in01s01 g737295 ( .a(n_42941), .o(n_42926) );
na02s01 g737296 ( .a(n_42885), .b(n_42875), .o(n_42941) );
in01s01 g737297 ( .a(n_42924), .o(n_42925) );
ao22s01 g737298 ( .a(n_42867), .b(n_42490), .c(n_42868), .d(n_42489), .o(n_42924) );
in01s01 g737299 ( .a(n_42922), .o(n_42923) );
oa22s01 g737300 ( .a(n_42847), .b(n_42767), .c(n_42862), .d(n_42768), .o(n_42922) );
no02s01 g737301 ( .a(n_42891), .b(n_42909), .o(n_43250) );
oa22s01 g737302 ( .a(n_42889), .b(n_42788), .c(n_42855), .d(n_42789), .o(n_43208) );
in01s01 g737305 ( .a(n_46940), .o(n_42936) );
in01s01 g737307 ( .a(n_42910), .o(n_42911) );
na02s01 g737308 ( .a(n_42873), .b(n_42859), .o(n_42910) );
ao22s01 g737309 ( .a(n_42842), .b(n_42642), .c(n_42852), .d(n_42641), .o(n_43123) );
in01s01 g737312 ( .a(n_42876), .o(n_42918) );
na02s01 g737314 ( .a(n_42860), .b(n_42473), .o(n_42876) );
na02s01 g737315 ( .a(n_42850), .b(n_42756), .o(n_42875) );
na02s01 g737316 ( .a(n_42851), .b(n_42757), .o(n_42885) );
no02s01 g737318 ( .a(n_42848), .b(n_42612), .o(n_42874) );
na02s01 g737319 ( .a(n_42840), .b(n_42408), .o(n_42873) );
na02s01 g737320 ( .a(n_42839), .b(n_42409), .o(n_42859) );
no02s01 g737321 ( .a(n_42864), .b(n_42488), .o(n_42909) );
no02s01 g737322 ( .a(n_42879), .b(n_42487), .o(n_42891) );
in01s01 g737323 ( .a(n_42844), .o(n_42845) );
ao12s01 g737324 ( .a(n_42300), .b(n_42812), .c(n_42327), .o(n_42844) );
no03s08 TIMEBOOST_cell_815 ( .a(n_6716), .b(n_6523), .c(n_6715), .o(TIMEBOOST_net_22) );
in01s01 g737327 ( .a(n_42857), .o(n_42871) );
ao12s01 g737328 ( .a(n_42648), .b(n_42834), .c(n_42503), .o(n_42857) );
na02s01 g737330 ( .a(n_42831), .b(n_42329), .o(n_42869) );
in01s01 g737331 ( .a(n_43181), .o(n_42883) );
no02s01 g737332 ( .a(n_42841), .b(n_42832), .o(n_43181) );
ao12s01 g737334 ( .a(n_42450), .b(n_42854), .c(n_42464), .o(n_42881) );
in01s01 g737335 ( .a(n_42856), .o(n_43172) );
ao22s01 g737336 ( .a(n_42813), .b(n_42615), .c(n_42814), .d(n_42614), .o(n_42856) );
oa22s01 g737337 ( .a(n_42823), .b(n_42348), .c(n_42812), .d(n_42349), .o(n_43102) );
na02f08 g737338 ( .a(n_42833), .b(n_42388), .o(n_42860) );
in01s01 g737339 ( .a(n_42889), .o(n_42855) );
in01s01 g737340 ( .a(n_42843), .o(n_42889) );
no02f08 g737341 ( .a(n_42834), .b(n_42594), .o(n_42843) );
in01s01 g737342 ( .a(n_42867), .o(n_42868) );
no02s01 g737343 ( .a(n_42854), .b(n_42433), .o(n_42867) );
in01s01 g737347 ( .a(n_42842), .o(n_42852) );
no02s02 g737348 ( .a(n_42833), .b(n_42399), .o(n_42842) );
no02s01 g737349 ( .a(n_42821), .b(n_42763), .o(n_42832) );
no02s01 g737350 ( .a(n_42822), .b(n_42762), .o(n_42841) );
in01s01 g737351 ( .a(n_42839), .o(n_42840) );
no02s01 g737352 ( .a(n_42830), .b(n_42368), .o(n_42839) );
na02s01 g737353 ( .a(n_42830), .b(n_42414), .o(n_42831) );
in01s01 g737355 ( .a(n_42864), .o(n_42879) );
ao12s01 g737356 ( .a(n_42551), .b(n_42808), .c(n_42530), .o(n_42864) );
in01s01 g737357 ( .a(n_42850), .o(n_42851) );
oa12s01 g737358 ( .a(n_42747), .b(n_42838), .c(n_42727), .o(n_42850) );
oa12s01 g737360 ( .a(n_42580), .b(n_42807), .c(n_42514), .o(n_42848) );
in01s01 g737362 ( .a(n_42847), .o(n_42862) );
oa12s01 g737363 ( .a(n_42511), .b(n_42838), .c(n_42529), .o(n_42847) );
in01s01 g737364 ( .a(n_42829), .o(n_43147) );
ao22s01 g737365 ( .a(n_42779), .b(n_42729), .c(n_42778), .d(n_42728), .o(n_42829) );
na02s01 g737366 ( .a(n_42846), .b(n_42861), .o(n_43211) );
in01s01 g737367 ( .a(n_42956), .o(n_42878) );
na02s01 g737368 ( .a(n_42828), .b(n_42837), .o(n_42956) );
no02s01 g737369 ( .a(n_42838), .b(n_42468), .o(n_42854) );
na02s01 g737370 ( .a(n_42808), .b(n_42769), .o(n_42861) );
na02s01 g737371 ( .a(n_42838), .b(n_42770), .o(n_42846) );
no02s01 g737372 ( .a(n_42340), .b(n_42811), .o(n_42830) );
na02s01 g737373 ( .a(n_42806), .b(n_42625), .o(n_42837) );
na02s01 g737374 ( .a(n_42807), .b(n_42626), .o(n_42828) );
in01s01 g737376 ( .a(n_42813), .o(n_42814) );
ao12s01 g737377 ( .a(n_42559), .b(n_42796), .c(n_42581), .o(n_42813) );
in01s01 g737379 ( .a(n_42812), .o(n_42823) );
ao12s02 g737380 ( .a(n_42370), .b(n_42796), .c(n_42359), .o(n_42812) );
in01s01 g737382 ( .a(n_42821), .o(n_42822) );
no02s02 TIMEBOOST_cell_6921 ( .a(n_7863), .b(n_7900), .o(TIMEBOOST_net_2219) );
na02s01 g737384 ( .a(n_42783), .b(n_42791), .o(n_43135) );
na02s01 g737385 ( .a(n_42810), .b(n_42795), .o(n_43104) );
na02s01 g737386 ( .a(n_42796), .b(n_42627), .o(n_42810) );
na02s01 g737387 ( .a(n_42775), .b(n_42628), .o(n_42795) );
no02s04 TIMEBOOST_cell_2089 ( .a(n_30530), .b(n_30201), .o(TIMEBOOST_net_659) );
na02s01 g737389 ( .a(n_46942), .b(n_42792), .o(n_42794) );
na02s01 g737390 ( .a(n_42782), .b(n_42466), .o(n_42783) );
na02s01 g737391 ( .a(n_42751), .b(n_42465), .o(n_42791) );
na02s01 g737392 ( .a(n_42780), .b(n_43132), .o(n_42781) );
in01s02 g737397 ( .a(n_42808), .o(n_42838) );
in01m01 g737398 ( .a(n_42790), .o(n_42808) );
in01s01 g737400 ( .a(n_42778), .o(n_42779) );
oa12s01 g737401 ( .a(n_42700), .b(n_42738), .c(n_42660), .o(n_42778) );
in01s01 g737404 ( .a(n_42806), .o(n_42807) );
in01s01 g737405 ( .a(n_42811), .o(n_42806) );
in01s01 g737407 ( .a(n_43106), .o(n_42805) );
ao22s01 g737408 ( .a(n_42732), .b(n_42698), .c(n_42731), .d(n_42699), .o(n_43106) );
in01s01 g737410 ( .a(n_43129), .o(n_42804) );
no02s02 g737411 ( .a(n_42753), .b(n_42740), .o(n_43129) );
no02s01 g737412 ( .a(n_42718), .b(n_42621), .o(n_42740) );
no02s01 g737413 ( .a(n_42719), .b(n_42620), .o(n_42753) );
no02s01 g737415 ( .a(n_42734), .b(n_42712), .o(n_42752) );
in01s01 g737417 ( .a(n_42796), .o(n_42775) );
na02m01 g737418 ( .a(n_42428), .b(n_42736), .o(n_42796) );
in01s01 g737421 ( .a(n_42802), .o(n_42803) );
na02s01 g737422 ( .a(n_42749), .b(n_42733), .o(n_42802) );
in01s01 g737423 ( .a(n_46942), .o(n_42774) );
in01s01 g737425 ( .a(n_42782), .o(n_42751) );
na02s01 g737426 ( .a(n_42706), .b(n_42495), .o(n_42782) );
in01s01 g737427 ( .a(n_42772), .o(n_42773) );
oa12s01 g737428 ( .a(n_42723), .b(n_42722), .c(n_42721), .o(n_42772) );
in01s01 g737429 ( .a(n_42780), .o(n_42750) );
no02s01 g737430 ( .a(n_42707), .b(n_42690), .o(n_42780) );
no02s01 g737431 ( .a(n_42671), .b(n_42575), .o(n_42690) );
no02s01 g737432 ( .a(n_42672), .b(n_42574), .o(n_42707) );
na02s01 g737433 ( .a(n_42705), .b(n_42451), .o(n_42706) );
in01s01 g737435 ( .a(n_42738), .o(n_42734) );
no02f08 g737436 ( .a(n_42705), .b(n_42494), .o(n_42738) );
na02f08 g737437 ( .a(n_42703), .b(n_42577), .o(n_42736) );
na02s01 g737438 ( .a(n_42716), .b(n_42425), .o(n_42733) );
na02s01 g737439 ( .a(n_42717), .b(n_42426), .o(n_42749) );
na02s01 g737440 ( .a(n_42722), .b(n_42721), .o(n_42723) );
no02s01 g737442 ( .a(n_42687), .b(n_42681), .o(n_42704) );
in01s01 g737443 ( .a(n_42718), .o(n_42719) );
no02s01 g737444 ( .a(n_42703), .b(n_42357), .o(n_42718) );
in01s01 g737445 ( .a(n_42731), .o(n_42732) );
na02s01 g737446 ( .a(n_42689), .b(n_42427), .o(n_42731) );
no02s01 g737447 ( .a(n_42655), .b(n_42372), .o(n_42722) );
no02f08 g737448 ( .a(n_42654), .b(FE_OCPN1713_n_42306), .o(n_42703) );
in01s01 g737449 ( .a(n_42716), .o(n_42717) );
na02s01 g737450 ( .a(n_42670), .b(n_42386), .o(n_42716) );
na02s01 g737451 ( .a(n_42669), .b(n_42402), .o(n_42689) );
in01s01 g737452 ( .a(n_42671), .o(n_42672) );
ao12s01 g737453 ( .a(n_42545), .b(n_42639), .c(n_42582), .o(n_42671) );
oa12s01 g737456 ( .a(n_42663), .b(n_42637), .c(n_42583), .o(n_42687) );
in01s01 g737457 ( .a(n_42792), .o(n_42771) );
no02s01 g737458 ( .a(n_42702), .b(n_42715), .o(n_42792) );
no02s01 g737459 ( .a(n_42638), .b(n_42653), .o(n_43132) );
in01s01 g737460 ( .a(n_42654), .o(n_42655) );
no02s01 g737462 ( .a(n_42639), .b(n_42629), .o(n_42638) );
no02s01 g737463 ( .a(n_42599), .b(n_42630), .o(n_42653) );
no02s01 g737464 ( .a(n_42637), .b(n_42684), .o(n_42715) );
no02s01 g737465 ( .a(n_42650), .b(n_42683), .o(n_42702) );
in01s01 g737466 ( .a(n_42669), .o(n_42670) );
in01s01 g737467 ( .a(n_42652), .o(n_42669) );
in01s01 g737469 ( .a(n_43070), .o(n_42748) );
no02s01 g737470 ( .a(n_42686), .b(n_42701), .o(n_43070) );
in01s01 g737471 ( .a(n_46944), .o(n_42668) );
in01s01 g737473 ( .a(n_43130), .o(n_42666) );
ao12s02 g737474 ( .a(n_42604), .b(n_42603), .c(n_42602), .o(n_43130) );
no02s01 g737475 ( .a(n_42603), .b(n_42602), .o(n_42604) );
no02s01 g737476 ( .a(n_42565), .b(n_42661), .o(n_42686) );
no02s01 g737477 ( .a(n_42564), .b(n_42662), .o(n_42701) );
na02s01 g737479 ( .a(n_42552), .b(n_42314), .o(n_42567) );
in01s01 g737481 ( .a(n_42637), .o(n_42650) );
in01s01 g737482 ( .a(n_42600), .o(n_42637) );
ao12f08 g737483 ( .a(n_42566), .b(n_42554), .c(n_42378), .o(n_42600) );
in01s01 g737484 ( .a(n_42639), .o(n_42599) );
ao12f08 g737485 ( .a(n_42247), .b(n_42555), .c(n_42259), .o(n_42639) );
in01s01 g737486 ( .a(n_43061), .o(n_42730) );
no02s01 g737487 ( .a(n_42665), .b(n_42685), .o(n_43061) );
no02s01 g737488 ( .a(n_42635), .b(n_42645), .o(n_42685) );
no02s01 g737489 ( .a(n_42636), .b(n_42644), .o(n_42665) );
na02s01 g737490 ( .a(n_42215), .b(n_42555), .o(n_42603) );
in01s01 g737491 ( .a(n_42564), .o(n_42565) );
na02s01 g737492 ( .a(n_42554), .b(n_42316), .o(n_42564) );
ao12s01 g737494 ( .a(n_42377), .b(n_42541), .c(n_42540), .o(n_42552) );
in01s01 g737495 ( .a(n_42597), .o(n_42598) );
ao12s01 g737496 ( .a(n_42539), .b(n_42538), .c(n_42537), .o(n_42597) );
in01s01 g737497 ( .a(n_42635), .o(n_42636) );
no02s01 g737498 ( .a(n_42541), .b(n_42589), .o(n_42635) );
no02s01 g737499 ( .a(n_42538), .b(n_42537), .o(n_42539) );
ao12f08 g737500 ( .a(n_42497), .b(n_42498), .c(n_42225), .o(n_42555) );
in01s01 g737502 ( .a(n_43037), .o(n_42714) );
no02s02 g737503 ( .a(n_42664), .b(n_42649), .o(n_43037) );
in01s01 g737504 ( .a(n_43083), .o(n_42596) );
ao12s01 g737505 ( .a(n_42536), .b(n_42535), .c(n_42534), .o(n_43083) );
no02s01 g737506 ( .a(n_42535), .b(n_42534), .o(n_42536) );
no02f08 g737507 ( .a(n_42475), .b(n_42474), .o(n_42541) );
no02s01 g737508 ( .a(n_42498), .b(n_42497), .o(n_42538) );
no02s01 g737509 ( .a(n_42475), .b(n_42631), .o(n_42649) );
no02s01 g737510 ( .a(n_42454), .b(n_42632), .o(n_42664) );
na02s01 g737511 ( .a(n_42595), .b(n_42520), .o(n_42648) );
no02f08 g737512 ( .a(n_42455), .b(n_42213), .o(n_42498) );
na02s01 g737513 ( .a(n_42455), .b(n_42496), .o(n_42535) );
in01s01 g737514 ( .a(n_46943), .o(n_43158) );
in01s01 g737516 ( .a(n_43121), .o(n_43494) );
ao12s01 g737517 ( .a(n_42533), .b(n_42532), .c(n_42531), .o(n_43121) );
in01s01 g737518 ( .a(n_42475), .o(n_42454) );
no02f08 g737519 ( .a(n_42381), .b(n_42336), .o(n_42475) );
na02f08 g737520 ( .a(n_42532), .b(n_42403), .o(n_42455) );
in01s01 g737521 ( .a(n_42594), .o(n_42595) );
na02m04 g737522 ( .a(n_42550), .b(n_42491), .o(n_42594) );
no02s01 g737523 ( .a(n_42532), .b(n_42531), .o(n_42533) );
ao12f06 g737524 ( .a(n_42203), .b(n_42337), .c(n_42242), .o(n_42381) );
no02s01 g737526 ( .a(n_42379), .b(n_42587), .o(n_42634) );
ao12m04 g737527 ( .a(n_42453), .b(n_42472), .c(n_42461), .o(n_42512) );
na02s01 g737529 ( .a(n_42337), .b(n_42253), .o(n_42379) );
no02s01 g737530 ( .a(n_42494), .b(n_42435), .o(n_42495) );
no02s06 g737531 ( .a(n_42337), .b(n_42335), .o(n_42336) );
in01s01 g737532 ( .a(n_42550), .o(n_42551) );
no02m04 g737533 ( .a(n_42510), .b(n_42447), .o(n_42550) );
na02s02 g737534 ( .a(n_42291), .b(n_42318), .o(n_43021) );
ao12s02 g737535 ( .a(n_42509), .b(n_42508), .c(n_42507), .o(n_43052) );
oa12f06 g737536 ( .a(n_42268), .b(n_42265), .c(n_42192), .o(n_42532) );
no02s01 g737537 ( .a(n_42529), .b(n_42470), .o(n_42530) );
na02s02 g737538 ( .a(n_42590), .b(n_42563), .o(n_42633) );
na02f08 g737539 ( .a(n_42290), .b(n_42254), .o(n_42337) );
na02s01 g737540 ( .a(n_42290), .b(n_42262), .o(n_42291) );
na02s01 g737541 ( .a(n_42264), .b(n_42263), .o(n_42318) );
oa12s02 g737543 ( .a(n_42386), .b(n_42375), .c(n_42367), .o(n_42494) );
no02s06 g737544 ( .a(n_42317), .b(n_42377), .o(n_42378) );
in01s01 g737545 ( .a(n_42510), .o(n_42511) );
oa12s02 g737546 ( .a(n_42449), .b(n_42422), .c(n_42367), .o(n_42510) );
no02s01 g737547 ( .a(n_42508), .b(n_42507), .o(n_42509) );
na02s02 g737549 ( .a(n_42592), .b(n_42528), .o(n_42593) );
in01s01 g737550 ( .a(n_42472), .o(n_42473) );
oa12m02 g737551 ( .a(n_42373), .b(n_42398), .c(n_42387), .o(n_42472) );
ao22s01 g737552 ( .a(n_42252), .b(n_42218), .c(n_42251), .d(n_42208), .o(n_43014) );
no02s01 g737553 ( .a(n_42504), .b(n_42549), .o(n_42592) );
in01s01 g737554 ( .a(n_42590), .o(n_42591) );
no02s02 g737555 ( .a(n_42521), .b(n_42505), .o(n_42590) );
na02f06 g737556 ( .a(n_42266), .b(n_42267), .o(n_42268) );
no02s01 g737557 ( .a(n_42266), .b(n_42221), .o(n_42508) );
na02s04 g737558 ( .a(n_42400), .b(n_42412), .o(n_42453) );
in01s01 g737561 ( .a(n_42492), .o(n_42529) );
in01s01 TIMEBOOST_cell_8907 ( .a(TIMEBOOST_net_2950), .o(TIMEBOOST_net_2951) );
no02s03 TIMEBOOST_cell_2085 ( .a(n_34982), .b(n_30588), .o(TIMEBOOST_net_657) );
no02s06 g737564 ( .a(n_42261), .b(n_42285), .o(n_42317) );
na02m01 g737565 ( .a(n_42442), .b(n_42216), .o(n_42491) );
no02f06 g737566 ( .a(n_42266), .b(n_42210), .o(n_42265) );
in01s01 g737568 ( .a(n_42290), .o(n_42264) );
na02s01 TIMEBOOST_cell_7562 ( .a(n_25253), .b(n_25254), .o(TIMEBOOST_net_2412) );
oa12s01 g737570 ( .a(n_42238), .b(n_42240), .c(n_42237), .o(n_43031) );
no02s01 g737571 ( .a(n_42377), .b(n_42287), .o(n_42316) );
na02s01 g737572 ( .a(n_42449), .b(n_42448), .o(n_42450) );
no02s01 g737573 ( .a(n_42410), .b(n_42334), .o(n_42427) );
no02s01 g737574 ( .a(n_42527), .b(n_42526), .o(n_42528) );
na02s02 g737577 ( .a(n_42446), .b(n_42445), .o(n_42447) );
no02s01 g737579 ( .a(n_42288), .b(n_42287), .o(n_42314) );
in01s01 g737580 ( .a(n_42425), .o(n_42426) );
na02s01 g737581 ( .a(n_42402), .b(n_42364), .o(n_42425) );
na02s01 g737583 ( .a(n_42700), .b(n_42659), .o(n_42712) );
in01s01 g737584 ( .a(n_42769), .o(n_42770) );
na02s01 g737585 ( .a(n_42747), .b(n_42726), .o(n_42769) );
in01s01 g737586 ( .a(n_42767), .o(n_42768) );
na02s01 g737587 ( .a(n_42746), .b(n_42445), .o(n_42767) );
in01s01 g737588 ( .a(n_42683), .o(n_42684) );
na02s01 g737589 ( .a(n_42663), .b(n_42584), .o(n_42683) );
in01s01 g737590 ( .a(n_42788), .o(n_42789) );
na02s01 g737591 ( .a(n_42766), .b(n_42725), .o(n_42788) );
in01s01 g737592 ( .a(n_42524), .o(n_42525) );
no02s01 g737593 ( .a(n_42505), .b(n_42549), .o(n_42524) );
in01s01 g737594 ( .a(n_42817), .o(n_42818) );
na02s01 g737595 ( .a(n_42754), .b(n_42801), .o(n_42817) );
in01s01 g737596 ( .a(n_42631), .o(n_42632) );
no02s01 g737597 ( .a(n_42589), .b(n_42474), .o(n_42631) );
no02s04 TIMEBOOST_cell_2084 ( .a(TIMEBOOST_net_656), .b(n_19566), .o(n_19642) );
in01s01 g737599 ( .a(n_42465), .o(n_42466) );
no02s01 g737600 ( .a(n_42444), .b(n_42443), .o(n_42465) );
in01s01 g737601 ( .a(n_42489), .o(n_42490) );
na02s01 g737602 ( .a(n_42464), .b(n_42448), .o(n_42489) );
in01s01 g737603 ( .a(n_42262), .o(n_42263) );
na02s01 g737604 ( .a(n_42254), .b(n_42253), .o(n_42262) );
no02s02 g737606 ( .a(n_42334), .b(n_42374), .o(n_42375) );
no02s04 g737607 ( .a(n_42222), .b(n_42241), .o(n_42242) );
no02s02 g737608 ( .a(n_42287), .b(n_42286), .o(n_42261) );
no02s01 g737609 ( .a(n_42389), .b(n_42421), .o(n_42422) );
na02s02 g737610 ( .a(n_42463), .b(n_42441), .o(n_42442) );
no02f08 g737611 ( .a(n_42240), .b(n_42220), .o(n_42266) );
in01s01 g737612 ( .a(n_42487), .o(n_42488) );
na02s01 g737613 ( .a(n_42437), .b(n_42463), .o(n_42487) );
ao12s02 g737614 ( .a(n_42298), .b(n_42311), .c(FE_OCPN873_n_42202), .o(n_42373) );
in01s01 g737615 ( .a(n_42251), .o(n_42252) );
na02s01 g737616 ( .a(n_42239), .b(n_42223), .o(n_42251) );
in01s01 g737617 ( .a(n_42400), .o(n_42401) );
ao12s02 g737618 ( .a(n_42294), .b(n_42308), .c(n_42270), .o(n_42400) );
na02s02 TIMEBOOST_cell_7561 ( .a(TIMEBOOST_net_2411), .b(n_25288), .o(FE_RN_701_0) );
na02s01 g737620 ( .a(n_42240), .b(n_42237), .o(n_42238) );
no02m04 g737621 ( .a(n_42330), .b(n_42372), .o(n_42428) );
in01s01 g737623 ( .a(n_42398), .o(n_42399) );
ao12s02 g737624 ( .a(n_42368), .b(n_42303), .c(FE_OCPN873_n_42202), .o(n_42398) );
in01s02 g737625 ( .a(n_42461), .o(n_42462) );
no02s02 g737626 ( .a(n_42385), .b(n_42440), .o(n_42461) );
in01s01 g737627 ( .a(n_42661), .o(n_42662) );
ao12s01 g737628 ( .a(n_42566), .b(n_42392), .c(n_42286), .o(n_42661) );
in01s01 g737629 ( .a(n_42644), .o(n_42645) );
oa12s01 g737630 ( .a(n_42540), .b(FE_OCPN1044_n_42367), .c(n_41909), .o(n_42644) );
in01s01 g737631 ( .a(n_42698), .o(n_42699) );
ao12s01 g737632 ( .a(n_42333), .b(n_42392), .c(n_42374), .o(n_42698) );
in01s01 g737633 ( .a(n_42764), .o(n_42765) );
oa12s01 g737634 ( .a(n_42446), .b(n_42392), .c(n_42391), .o(n_42764) );
in01s01 g737635 ( .a(n_42762), .o(n_42763) );
ao12s01 g737636 ( .a(n_42396), .b(n_42392), .c(n_42423), .o(n_42762) );
ao12s01 g737638 ( .a(n_42467), .b(n_42392), .c(n_42421), .o(n_42760) );
in01s01 g737639 ( .a(n_42825), .o(n_42826) );
ao12s01 g737640 ( .a(n_42527), .b(n_42392), .c(n_42112), .o(n_42825) );
in01s01 g737641 ( .a(n_42799), .o(n_42800) );
no02s01 g737642 ( .a(n_42742), .b(n_42469), .o(n_42799) );
no02f06 TIMEBOOST_cell_5347 ( .a(TIMEBOOST_net_1621), .b(n_21013), .o(n_21230) );
na02s02 TIMEBOOST_cell_2942 ( .a(FE_OCP_RBN4038_n_2059), .b(n_2081), .o(TIMEBOOST_net_762) );
oa22s01 g737646 ( .a(FE_OCPN1044_n_42367), .b(n_42335), .c(n_42392), .d(n_42241), .o(n_42587) );
oa22s01 g737648 ( .a(FE_OCPN1044_n_42367), .b(n_41936), .c(n_42392), .d(n_42358), .o(n_42681) );
in01s01 g737649 ( .a(n_42728), .o(n_42729) );
oa22s01 g737650 ( .a(n_42392), .b(n_41983), .c(FE_OCPN1044_n_42367), .d(n_41993), .o(n_42728) );
in01s01 g737651 ( .a(n_42758), .o(n_42759) );
oa22s01 g737652 ( .a(FE_OCPN1044_n_42367), .b(n_42093), .c(n_42392), .d(n_42072), .o(n_42758) );
in01s01 g737653 ( .a(n_42797), .o(n_42798) );
oa22s01 g737654 ( .a(FE_OCPN1044_n_42367), .b(n_42459), .c(n_42392), .d(n_42483), .o(n_42797) );
in01s01 g737655 ( .a(n_42815), .o(n_42816) );
oa22s01 g737656 ( .a(FE_OCPN1044_n_42367), .b(n_42116), .c(n_42392), .d(n_42101), .o(n_42815) );
in01s01 g737657 ( .a(n_42756), .o(n_42757) );
oa22s01 g737658 ( .a(FE_OCPN1044_n_42367), .b(n_42066), .c(n_42392), .d(n_42048), .o(n_42756) );
ao12s01 g737659 ( .a(n_42236), .b(n_42235), .c(n_42234), .o(n_43019) );
in01s01 g737660 ( .a(n_42585), .o(n_42586) );
na02s02 g737661 ( .a(n_42519), .b(n_42502), .o(n_42585) );
in01s01 g737662 ( .a(n_42583), .o(n_42584) );
no02s01 g737663 ( .a(n_42392), .b(n_42562), .o(n_42583) );
no02s01 g737664 ( .a(FE_OCPN1044_n_42367), .b(n_41884), .o(n_42589) );
in01s01 g737665 ( .a(n_42659), .o(n_42660) );
na02s01 g737666 ( .a(FE_OCPN1044_n_42367), .b(n_41992), .o(n_42659) );
in01s01 g737667 ( .a(n_42726), .o(n_42727) );
na02s01 g737668 ( .a(FE_OCPN1044_n_42367), .b(n_42065), .o(n_42726) );
na02s01 g737669 ( .a(n_42392), .b(n_42562), .o(n_42663) );
no02s01 g737670 ( .a(FE_OCPN1044_n_42367), .b(n_42441), .o(n_42742) );
na02s01 g737671 ( .a(FE_OCPN1044_n_42367), .b(n_42710), .o(n_42766) );
in01s01 g737672 ( .a(n_42724), .o(n_42725) );
no02s01 g737673 ( .a(FE_OCPN1044_n_42367), .b(n_42710), .o(n_42724) );
na02s01 g737674 ( .a(n_42392), .b(n_41982), .o(n_42700) );
in01s01 g737675 ( .a(n_42754), .o(n_42755) );
na02s01 g737676 ( .a(FE_OCPN1044_n_42367), .b(n_42115), .o(n_42754) );
na02s01 g737677 ( .a(n_42392), .b(n_42049), .o(n_42801) );
na02s01 g737678 ( .a(n_42392), .b(n_42069), .o(n_42519) );
in01s01 g737679 ( .a(n_42505), .o(n_42486) );
no02s01 g737680 ( .a(n_42285), .b(n_42053), .o(n_42505) );
no02s01 TIMEBOOST_cell_4023 ( .a(FE_OCP_RBN4351_n_20456), .b(FE_OCP_RBN2721_n_19601), .o(TIMEBOOST_net_1102) );
no02s01 g737682 ( .a(n_42216), .b(n_42052), .o(n_42549) );
no02s01 g737683 ( .a(n_42392), .b(n_42112), .o(n_42527) );
na02m04 TIMEBOOST_cell_2941 ( .a(TIMEBOOST_net_761), .b(n_19599), .o(TIMEBOOST_net_281) );
no02s06 g737685 ( .a(n_42367), .b(n_42366), .o(n_42443) );
in01s01 g737686 ( .a(n_42397), .o(n_42444) );
na02s01 g737687 ( .a(n_42367), .b(n_42366), .o(n_42397) );
in01s01 g737688 ( .a(n_42395), .o(n_42396) );
na02s01 g737689 ( .a(n_42367), .b(n_41991), .o(n_42395) );
in01s01 g737691 ( .a(n_42334), .o(n_42364) );
no02s02 g737692 ( .a(n_42285), .b(n_42312), .o(n_42334) );
no02s02 g737693 ( .a(n_42216), .b(n_42286), .o(n_42566) );
no02s02 g737694 ( .a(n_42216), .b(n_41797), .o(n_42288) );
in01s01 g737695 ( .a(n_42260), .o(n_42540) );
no02s02 g737696 ( .a(n_42216), .b(n_41916), .o(n_42260) );
no02s02 g737697 ( .a(n_42216), .b(n_41915), .o(n_42474) );
na02s06 g737698 ( .a(n_42203), .b(n_42211), .o(n_42254) );
in01s01 g737699 ( .a(n_42222), .o(n_42253) );
no02s02 g737700 ( .a(n_42198), .b(n_42211), .o(n_42222) );
no02s02 g737701 ( .a(n_42203), .b(n_41796), .o(n_42287) );
na02s01 g737702 ( .a(n_42285), .b(n_42312), .o(n_42402) );
in01s01 g737703 ( .a(n_42332), .o(n_42333) );
na02s01 g737704 ( .a(n_42285), .b(n_41956), .o(n_42332) );
in01s01 g737706 ( .a(n_42420), .o(n_42437) );
no02s01 g737707 ( .a(n_42394), .b(n_42390), .o(n_42420) );
in01s01 g737708 ( .a(n_42419), .o(n_42464) );
no02s01 g737709 ( .a(n_42216), .b(n_42077), .o(n_42419) );
no02s02 g737710 ( .a(n_42394), .b(n_42172), .o(n_42469) );
no02s01 g737711 ( .a(n_42392), .b(n_42421), .o(n_42467) );
na02s01 g737712 ( .a(n_42394), .b(n_42391), .o(n_42446) );
in01s01 g737713 ( .a(n_42445), .o(n_42418) );
na02s01 g737714 ( .a(n_42392), .b(n_42124), .o(n_42445) );
na02s02 g737715 ( .a(n_42394), .b(n_42390), .o(n_42463) );
in01s01 g737716 ( .a(n_42389), .o(n_42448) );
no02s01 g737717 ( .a(n_42285), .b(n_42076), .o(n_42389) );
na02s01 g737718 ( .a(n_42392), .b(n_41988), .o(n_42747) );
na02s01 g737719 ( .a(n_42367), .b(n_42050), .o(n_42502) );
na02s01 g737720 ( .a(FE_OCPN1044_n_42367), .b(n_42158), .o(n_42746) );
na02m06 g737721 ( .a(n_42195), .b(n_41505), .o(n_42239) );
na02f04 g737722 ( .a(n_42194), .b(n_41504), .o(n_42223) );
no02s01 g737723 ( .a(n_42235), .b(n_42234), .o(n_42236) );
in01s01 g737724 ( .a(n_42387), .o(n_42388) );
no03m08 TIMEBOOST_cell_6456 ( .a(TIMEBOOST_net_1237), .b(FE_OCP_RBN2636_n_29371), .c(FE_OFN775_n_25834), .o(n_29527) );
na03s02 g737726 ( .a(n_42417), .b(n_42343), .c(n_42416), .o(n_42440) );
na02s01 g737729 ( .a(n_42392), .b(n_42094), .o(n_42520) );
na02s02 g737730 ( .a(n_42352), .b(n_42270), .o(n_42412) );
na02s01 g737731 ( .a(n_42392), .b(n_42117), .o(n_42522) );
na02s01 g737732 ( .a(n_42285), .b(n_42073), .o(n_42503) );
no02s01 g737733 ( .a(n_42392), .b(n_42114), .o(n_42526) );
in01s01 g737734 ( .a(n_42434), .o(n_42435) );
na02s01 g737735 ( .a(n_42392), .b(n_41994), .o(n_42434) );
na02s01 g737736 ( .a(n_42285), .b(n_41984), .o(n_42451) );
in01s01 g737738 ( .a(n_42386), .o(n_42410) );
oa12s01 g737739 ( .a(n_42216), .b(n_42358), .c(n_42562), .o(n_42386) );
no02s06 g737740 ( .a(n_42285), .b(n_41917), .o(n_42377) );
no02s02 g737742 ( .a(n_42394), .b(n_42159), .o(n_42470) );
no02s01 g737743 ( .a(n_42216), .b(n_42067), .o(n_42468) );
in01s01 g737744 ( .a(n_42449), .o(n_42433) );
na02s01 g737745 ( .a(n_42216), .b(n_42064), .o(n_42449) );
na02s04 g737746 ( .a(n_42202), .b(n_42233), .o(n_42259) );
na02s06 TIMEBOOST_cell_8464 ( .a(n_36887), .b(n_36886), .o(TIMEBOOST_net_2719) );
in01s01 g737748 ( .a(n_43016), .o(n_42249) );
ao12s01 g737749 ( .a(n_42206), .b(n_42205), .c(n_42204), .o(n_43016) );
na02s01 g737751 ( .a(n_42341), .b(n_42384), .o(n_42385) );
na02s01 g737752 ( .a(n_42293), .b(n_42258), .o(n_42357) );
no02s01 g737753 ( .a(n_42368), .b(n_42274), .o(n_42329) );
in01s01 g737754 ( .a(n_42355), .o(n_42356) );
na02s01 g737755 ( .a(n_42363), .b(n_42310), .o(n_42355) );
in01s01 g737756 ( .a(n_42679), .o(n_42680) );
na02s01 g737757 ( .a(n_42657), .b(n_42609), .o(n_42679) );
na02s02 g737758 ( .a(n_42310), .b(n_42309), .o(n_42311) );
in01s01 g737759 ( .a(n_42353), .o(n_42354) );
na02s01 g737760 ( .a(n_42307), .b(n_42417), .o(n_42353) );
na02s01 g737761 ( .a(n_42307), .b(n_42323), .o(n_42308) );
in01s01 g737762 ( .a(n_42677), .o(n_42678) );
na02s01 g737763 ( .a(n_42656), .b(n_42607), .o(n_42677) );
na02s02 g737764 ( .a(n_42351), .b(n_42350), .o(n_42352) );
na02s02 g737765 ( .a(n_42215), .b(n_42232), .o(n_42233) );
na02m04 g737766 ( .a(n_42193), .b(n_42209), .o(n_42210) );
no02s01 g737767 ( .a(n_42283), .b(n_42306), .o(n_42721) );
in01s01 g737768 ( .a(n_42629), .o(n_42630) );
na02s01 g737769 ( .a(n_42546), .b(n_42582), .o(n_42629) );
no02s01 g737770 ( .a(n_42221), .b(n_42220), .o(n_42237) );
na02s01 g737771 ( .a(n_42496), .b(n_42403), .o(n_42531) );
no02s01 g737772 ( .a(n_42227), .b(n_42226), .o(n_42537) );
in01s01 g737773 ( .a(n_42627), .o(n_42628) );
na02s01 g737774 ( .a(n_42558), .b(n_42581), .o(n_42627) );
no02m04 TIMEBOOST_cell_5510 ( .a(n_21847), .b(FE_OCP_RBN6131_n_21736), .o(TIMEBOOST_net_1703) );
in01s01 g737776 ( .a(n_42348), .o(n_42349) );
na02s01 g737777 ( .a(n_42328), .b(n_42327), .o(n_42348) );
in01s01 g737778 ( .a(n_42625), .o(n_42626) );
na02s01 g737779 ( .a(n_42580), .b(n_42515), .o(n_42625) );
in01s01 g737781 ( .a(n_42408), .o(n_42409) );
na02s01 g737782 ( .a(n_42414), .b(n_42302), .o(n_42408) );
na02s01 g737783 ( .a(n_42302), .b(n_42321), .o(n_42303) );
in01s01 g737784 ( .a(n_42641), .o(n_42642) );
na02s01 g737785 ( .a(n_42624), .b(n_42557), .o(n_42641) );
in01s01 g737787 ( .a(n_42208), .o(n_42218) );
no02m04 g737788 ( .a(n_42187), .b(n_42204), .o(n_42208) );
no02s01 g737790 ( .a(n_42199), .b(n_42207), .o(n_42235) );
no02s01 g737791 ( .a(n_42205), .b(n_42204), .o(n_42206) );
in01s10 g737827 ( .a(n_42367), .o(n_42392) );
in01s06 g737828 ( .a(n_42216), .o(n_42367) );
in01s02 g737837 ( .a(n_42285), .o(n_42394) );
in01s06 g737842 ( .a(n_42216), .o(n_42285) );
in01s06 g737845 ( .a(n_42203), .o(n_42216) );
oa12s08 g737846 ( .a(n_42197), .b(n_42178), .c(n_42196), .o(n_42203) );
oa12s02 g737847 ( .a(n_42197), .b(n_42178), .c(n_42196), .o(n_42198) );
in01s01 g737848 ( .a(n_42622), .o(n_42623) );
oa12s01 g737849 ( .a(n_42362), .b(n_42547), .c(n_42309), .o(n_42622) );
in01s01 g737850 ( .a(n_42693), .o(n_42694) );
oa12s01 g737851 ( .a(n_42416), .b(n_42547), .c(n_42323), .o(n_42693) );
in01s01 g737852 ( .a(n_42691), .o(n_42692) );
oa12s01 g737853 ( .a(n_42384), .b(n_42547), .c(n_42350), .o(n_42691) );
oa12s01 g737854 ( .a(n_42214), .b(n_42201), .c(n_42212), .o(n_42534) );
oa12s01 g737855 ( .a(n_42248), .b(n_42547), .c(n_42232), .o(n_42602) );
in01s01 g737856 ( .a(n_42620), .o(n_42621) );
oa12s01 g737857 ( .a(n_42577), .b(n_42201), .c(n_42276), .o(n_42620) );
in01s01 g737858 ( .a(n_42618), .o(n_42619) );
oa12s01 g737859 ( .a(n_42360), .b(n_42547), .c(n_42304), .o(n_42618) );
oa12s01 g737861 ( .a(n_42413), .b(n_42547), .c(n_42321), .o(n_42616) );
oa22s01 g737863 ( .a(n_42270), .b(n_42137), .c(n_42547), .d(n_42113), .o(n_42673) );
oa22s01 g737865 ( .a(n_42270), .b(n_42160), .c(n_42547), .d(n_42151), .o(n_42708) );
in01s01 g737866 ( .a(n_42480), .o(n_42481) );
na02s02 g737867 ( .a(n_42406), .b(n_42383), .o(n_42480) );
in01m02 g737868 ( .a(n_42194), .o(n_42195) );
in01s01 g737870 ( .a(n_42574), .o(n_42575) );
oa22s01 g737871 ( .a(n_42270), .b(n_41949), .c(n_42547), .d(n_41923), .o(n_42574) );
ao22s01 g737872 ( .a(n_42201), .b(n_42209), .c(n_42270), .d(n_42267), .o(n_42507) );
in01s01 g737873 ( .a(n_42614), .o(n_42615) );
oa22s01 g737874 ( .a(n_42270), .b(n_41953), .c(n_42201), .d(n_42272), .o(n_42614) );
oa22s01 g737876 ( .a(n_42270), .b(n_42046), .c(n_42201), .d(n_42026), .o(n_42612) );
oa22s01 g737878 ( .a(n_42270), .b(n_42107), .c(n_42201), .d(n_42081), .o(n_42610) );
in01s01 g737879 ( .a(n_42310), .o(n_42280) );
na02s01 g737880 ( .a(n_42202), .b(n_42103), .o(n_42310) );
na02s02 g737881 ( .a(n_42201), .b(n_42104), .o(n_42363) );
na02s02 g737882 ( .a(n_42201), .b(n_42309), .o(n_42362) );
na02s01 g737883 ( .a(n_42270), .b(n_42570), .o(n_42657) );
in01s01 g737884 ( .a(n_42608), .o(n_42609) );
no02s01 g737885 ( .a(n_42270), .b(n_42570), .o(n_42608) );
in01s01 g737886 ( .a(n_42307), .o(n_42279) );
na02s02 g737887 ( .a(FE_OCPN873_n_42202), .b(n_42130), .o(n_42307) );
na02s01 g737888 ( .a(n_42201), .b(n_42131), .o(n_42417) );
na02s01 g737889 ( .a(n_42201), .b(n_42323), .o(n_42416) );
na02s01 g737890 ( .a(n_42270), .b(n_42569), .o(n_42656) );
in01s01 g737891 ( .a(n_42606), .o(n_42607) );
no02s01 g737892 ( .a(n_42270), .b(n_42569), .o(n_42606) );
na02s01 g737893 ( .a(n_42201), .b(n_42350), .o(n_42384) );
na02s01 g737894 ( .a(n_42270), .b(n_42122), .o(n_42406) );
na02s01 g737895 ( .a(n_42201), .b(n_42139), .o(n_42383) );
in01s01 g737896 ( .a(n_42247), .o(n_42248) );
no02s02 g737897 ( .a(n_42202), .b(n_41911), .o(n_42247) );
in01s01 g737899 ( .a(n_42215), .o(n_42227) );
na02s02 g737900 ( .a(n_42202), .b(n_41867), .o(n_42215) );
in01s01 g737901 ( .a(n_42225), .o(n_42226) );
na02s03 g737902 ( .a(n_42201), .b(n_41868), .o(n_42225) );
no02s06 g737903 ( .a(n_42189), .b(n_42188), .o(n_42220) );
in01s01 g737904 ( .a(n_42193), .o(n_42221) );
na02m02 g737905 ( .a(n_42189), .b(n_42188), .o(n_42193) );
na02s02 g737906 ( .a(n_42192), .b(n_42191), .o(n_42403) );
in01s01 g737907 ( .a(n_42213), .o(n_42214) );
no02s06 g737908 ( .a(n_42202), .b(n_41910), .o(n_42213) );
no02s01 g737909 ( .a(n_42202), .b(n_41922), .o(n_42306) );
in01s01 g737910 ( .a(n_42283), .o(n_42258) );
no02m01 g737911 ( .a(n_42201), .b(n_41921), .o(n_42283) );
in01s01 g737912 ( .a(n_42545), .o(n_42546) );
no02s01 g737913 ( .a(n_42201), .b(n_42478), .o(n_42545) );
na02s01 g737914 ( .a(n_42201), .b(n_42478), .o(n_42582) );
na02s01 g737915 ( .a(n_42270), .b(n_41886), .o(n_42496) );
na02s02 g737916 ( .a(n_42277), .b(n_42276), .o(n_42577) );
in01s01 g737917 ( .a(n_42558), .o(n_42559) );
na02s01 g737918 ( .a(n_42270), .b(n_41952), .o(n_42558) );
na02s01 g737919 ( .a(n_42547), .b(n_42271), .o(n_42581) );
na02s01 g737920 ( .a(n_42202), .b(n_41960), .o(n_42327) );
in01s01 g737921 ( .a(n_42328), .o(n_42300) );
na02s01 g737922 ( .a(n_42201), .b(n_41961), .o(n_42328) );
na02s01 g737923 ( .a(n_42201), .b(n_42304), .o(n_42360) );
na02s01 g737924 ( .a(n_42270), .b(n_42500), .o(n_42580) );
in01s01 g737925 ( .a(n_42514), .o(n_42515) );
no02s01 g737926 ( .a(n_42270), .b(n_42500), .o(n_42514) );
in01s01 g737927 ( .a(n_42302), .o(n_42274) );
na02s01 g737928 ( .a(n_42202), .b(n_42035), .o(n_42302) );
na02s01 g737929 ( .a(n_42201), .b(n_42036), .o(n_42414) );
na02s01 g737930 ( .a(n_42201), .b(n_42321), .o(n_42413) );
na02s01 g737931 ( .a(n_42270), .b(n_42542), .o(n_42624) );
in01s01 g737932 ( .a(n_42556), .o(n_42557) );
no02s01 g737933 ( .a(n_42270), .b(n_42542), .o(n_42556) );
no02f06 g737934 ( .a(n_42180), .b(n_41516), .o(n_42207) );
no02f06 g737935 ( .a(n_42179), .b(n_41515), .o(n_42199) );
in01s01 g737936 ( .a(n_42298), .o(n_42299) );
no02s01 g737937 ( .a(n_42201), .b(n_42108), .o(n_42298) );
in01s01 g737938 ( .a(n_42296), .o(n_42297) );
na02s01 g737939 ( .a(n_42277), .b(n_42106), .o(n_42296) );
in01s01 g737940 ( .a(n_42294), .o(n_42295) );
no02s01 g737941 ( .a(n_42277), .b(n_42136), .o(n_42294) );
in01s01 g737942 ( .a(n_42343), .o(n_42344) );
na02s01 g737943 ( .a(n_42201), .b(n_42138), .o(n_42343) );
na02s01 g737944 ( .a(n_42270), .b(n_42152), .o(n_42351) );
in01s01 g737945 ( .a(n_42341), .o(n_42342) );
na02s01 TIMEBOOST_cell_4135 ( .a(n_10821), .b(n_10713), .o(TIMEBOOST_net_1158) );
ao12s02 g737948 ( .a(n_42192), .b(n_42212), .c(n_42191), .o(n_42497) );
in01s01 g737949 ( .a(n_42372), .o(n_42293) );
no02s01 g737950 ( .a(n_42201), .b(n_41948), .o(n_42372) );
na02s01 g737951 ( .a(n_42201), .b(n_41954), .o(n_42359) );
ao12s02 g737952 ( .a(n_42201), .b(n_42272), .c(n_42271), .o(n_42370) );
no02s01 g737953 ( .a(n_42201), .b(n_42045), .o(n_42368) );
in01s01 g737954 ( .a(n_42339), .o(n_42340) );
na02s01 g737955 ( .a(n_42201), .b(n_42047), .o(n_42339) );
in01s01 g737956 ( .a(n_42187), .o(n_42205) );
oa12s01 g737958 ( .a(n_42183), .b(n_42182), .c(n_42181), .o(n_43025) );
no02m08 g737962 ( .a(n_42169), .b(n_42196), .o(n_42178) );
na02f04 g737963 ( .a(FE_OCP_RBN5845_n_42169), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42177) );
na02s01 g737964 ( .a(n_42182), .b(n_42181), .o(n_42183) );
no02f06 g737965 ( .a(n_42182), .b(n_41369), .o(n_42234) );
in01s01 g737971 ( .a(n_42202), .o(n_42277) );
in01s01 g737981 ( .a(n_42270), .o(n_42547) );
in01s03 g737999 ( .a(n_42201), .o(n_42270) );
in01s10 g738006 ( .a(n_42202), .o(n_42201) );
in01s08 g738007 ( .a(n_42192), .o(n_42202) );
in01s04 g738008 ( .a(n_42189), .o(n_42192) );
na02s06 TIMEBOOST_cell_7492 ( .a(n_23605), .b(n_23599), .o(TIMEBOOST_net_2377) );
in01f02 g738010 ( .a(n_42175), .o(n_42176) );
na02f06 g738011 ( .a(n_42167), .b(n_42165), .o(n_42175) );
in01f02 g738012 ( .a(n_42179), .o(n_42180) );
no03s04 TIMEBOOST_cell_8319 ( .a(FE_OCP_RBN5810_n_3645), .b(n_3576), .c(n_3646), .o(n_3784) );
na02f04 g738015 ( .a(n_42149), .b(n_42196), .o(n_42167) );
na02s04 g738016 ( .a(n_42150), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42165) );
in01s01 g738017 ( .a(n_42172), .o(n_42441) );
oa12s01 g738018 ( .a(n_42164), .b(n_42163), .c(n_42162), .o(n_42172) );
na02f08 g738023 ( .a(n_42153), .b(n_42146), .o(n_42169) );
na02s04 g738024 ( .a(n_42144), .b(n_42196), .o(n_42146) );
in01f06 g738025 ( .a(n_42166), .o(n_42173) );
no02f08 g738026 ( .a(n_42147), .b(n_42196), .o(n_42166) );
na02f06 g738027 ( .a(n_42143), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42153) );
na02s01 g738028 ( .a(n_42163), .b(n_42162), .o(n_42164) );
na02s01 g738029 ( .a(n_42151), .b(n_42102), .o(n_42152) );
na02s01 TIMEBOOST_cell_4134 ( .a(n_36335), .b(TIMEBOOST_net_1157), .o(n_36369) );
no02s01 g738031 ( .a(n_42148), .b(n_42158), .o(n_42159) );
in01s02 g738032 ( .a(n_42150), .o(n_42197) );
in01f02 g738033 ( .a(n_42150), .o(n_42149) );
no02s02 TIMEBOOST_cell_8146 ( .a(n_18791), .b(n_18746), .o(TIMEBOOST_net_2704) );
in01f03 g738035 ( .a(n_42156), .o(n_42157) );
no03m04 TIMEBOOST_cell_8382 ( .a(n_20582), .b(n_20583), .c(n_20735), .o(TIMEBOOST_net_1615) );
no02f08 TIMEBOOST_cell_8593 ( .a(TIMEBOOST_net_2783), .b(n_15241), .o(n_15387) );
na02s01 g738039 ( .a(n_42137), .b(n_42570), .o(n_42138) );
no02s01 g738040 ( .a(n_42137), .b(n_42570), .o(n_42136) );
ao12s01 g738041 ( .a(n_41687), .b(n_42145), .c(n_41602), .o(n_42163) );
no02s02 g738042 ( .a(n_42120), .b(n_42111), .o(n_42309) );
no02s02 g738043 ( .a(n_42119), .b(n_42110), .o(n_42323) );
in01s01 g738044 ( .a(n_42151), .o(n_42160) );
no02s01 g738045 ( .a(n_42118), .b(n_42109), .o(n_42151) );
in01s01 g738046 ( .a(n_42148), .o(n_42391) );
ao12s01 g738047 ( .a(n_42134), .b(n_42133), .c(n_42132), .o(n_42148) );
oa12s01 g738048 ( .a(n_42142), .b(n_42145), .c(n_42141), .o(n_42390) );
in01s04 g738049 ( .a(n_42154), .o(n_42155) );
in01m04 g738050 ( .a(n_42147), .o(n_42154) );
no02m03 TIMEBOOST_cell_5928 ( .a(n_46254), .b(TIMEBOOST_net_1815), .o(n_37014) );
in01s01 g738052 ( .a(n_42144), .o(n_42350) );
in01f02 g738053 ( .a(n_42144), .o(n_42143) );
na02f08 g738055 ( .a(n_42099), .b(n_42196), .o(n_42135) );
na02s02 TIMEBOOST_cell_3947 ( .a(n_9090), .b(n_8362), .o(TIMEBOOST_net_1064) );
no02s01 g738057 ( .a(n_42133), .b(n_42132), .o(n_42134) );
no02s02 g738058 ( .a(n_42092), .b(n_41906), .o(n_42120) );
no02s01 g738059 ( .a(n_42091), .b(n_41907), .o(n_42111) );
no02s01 g738060 ( .a(n_42089), .b(n_41903), .o(n_42110) );
no02s01 g738061 ( .a(n_42090), .b(n_41902), .o(n_42119) );
no02s01 g738062 ( .a(n_42087), .b(n_41881), .o(n_42109) );
no02s01 g738063 ( .a(n_42088), .b(n_41882), .o(n_42118) );
na02s01 g738064 ( .a(n_42145), .b(n_42141), .o(n_42142) );
na02s01 g738065 ( .a(n_42116), .b(n_42115), .o(n_42117) );
no02s01 g738066 ( .a(n_42116), .b(n_42115), .o(n_42114) );
in01s01 g738067 ( .a(n_42137), .o(n_42113) );
na02s01 g738068 ( .a(n_42074), .b(n_42060), .o(n_42137) );
in01s01 g738069 ( .a(n_42130), .o(n_42131) );
oa12s01 g738070 ( .a(n_42097), .b(n_42096), .c(n_42095), .o(n_42130) );
in01f02 g738071 ( .a(n_42122), .o(n_42139) );
in01s01 g738073 ( .a(n_42459), .o(n_42483) );
ao12s01 g738074 ( .a(n_42063), .b(n_42062), .c(n_42061), .o(n_42459) );
in01f06 g738075 ( .a(n_42128), .o(n_42129) );
no03s03 TIMEBOOST_cell_2814 ( .a(TIMEBOOST_net_91), .b(n_76), .c(n_160), .o(TIMEBOOST_net_698) );
no02f08 g738078 ( .a(n_42050), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42098) );
no02s06 TIMEBOOST_cell_2047 ( .a(n_29594), .b(n_29630), .o(TIMEBOOST_net_638) );
no02s01 g738080 ( .a(n_42062), .b(n_42061), .o(n_42063) );
na02s01 g738081 ( .a(n_42096), .b(n_42095), .o(n_42097) );
na02s01 g738082 ( .a(n_42042), .b(n_41904), .o(n_42074) );
na02s01 g738083 ( .a(n_42041), .b(n_41905), .o(n_42060) );
no02f06 TIMEBOOST_cell_4952 ( .a(FE_RN_1960_0), .b(FE_RN_1961_0), .o(TIMEBOOST_net_1424) );
no02s01 g738085 ( .a(n_42107), .b(n_42542), .o(n_42108) );
na02s01 g738086 ( .a(n_42107), .b(n_42542), .o(n_42106) );
na02s01 g738087 ( .a(n_42093), .b(n_42710), .o(n_42094) );
na02s01 g738088 ( .a(n_42072), .b(n_42013), .o(n_42073) );
oa12s01 g738089 ( .a(n_41875), .b(n_42105), .c(n_41532), .o(n_42133) );
in01s01 g738090 ( .a(n_42091), .o(n_42092) );
oa12s01 g738091 ( .a(n_41677), .b(n_42071), .c(n_41586), .o(n_42091) );
in01s01 g738092 ( .a(n_42089), .o(n_42090) );
ao12s01 g738093 ( .a(n_41710), .b(n_42059), .c(n_41592), .o(n_42089) );
in01s01 g738094 ( .a(n_42087), .o(n_42088) );
oa12s01 g738095 ( .a(n_41731), .b(n_42070), .c(n_41670), .o(n_42087) );
in01f03 g738096 ( .a(n_42085), .o(n_42086) );
ao12f06 g738097 ( .a(n_41772), .b(n_42070), .c(n_41751), .o(n_42085) );
in01s01 g738098 ( .a(n_42103), .o(n_42104) );
oa22s01 g738099 ( .a(n_42071), .b(n_41703), .c(n_42037), .d(n_41704), .o(n_42103) );
in01s01 g738100 ( .a(n_42102), .o(n_42569) );
ao12s01 g738101 ( .a(n_42055), .b(n_42070), .c(n_42054), .o(n_42102) );
in01s01 g738102 ( .a(n_42116), .o(n_42101) );
ao12s01 g738103 ( .a(n_42058), .b(n_42057), .c(n_42056), .o(n_42116) );
in01s01 g738105 ( .a(n_42112), .o(n_42125) );
in01s01 g738106 ( .a(n_42100), .o(n_42112) );
in01f04 g738107 ( .a(n_42100), .o(n_42099) );
in01s01 g738109 ( .a(n_42158), .o(n_42124) );
ao12s01 g738110 ( .a(n_42084), .b(n_42105), .c(n_42083), .o(n_42158) );
no02s01 g738111 ( .a(n_42059), .b(n_41735), .o(n_42096) );
no02s01 g738112 ( .a(n_42056), .b(n_42057), .o(n_42058) );
no02s01 g738113 ( .a(n_42105), .b(n_42083), .o(n_42084) );
no02s01 g738114 ( .a(n_42070), .b(n_42054), .o(n_42055) );
na02s01 g738115 ( .a(n_42046), .b(n_42500), .o(n_42047) );
no02s01 g738116 ( .a(n_42046), .b(n_42500), .o(n_42045) );
ao12s01 g738117 ( .a(n_41722), .b(n_42031), .c(n_41657), .o(n_42062) );
ao12f06 g738119 ( .a(n_41885), .b(n_42030), .c(n_41791), .o(n_42043) );
na02f06 TIMEBOOST_cell_2044 ( .a(n_41924), .b(TIMEBOOST_net_636), .o(n_41976) );
in01s01 g738121 ( .a(n_42041), .o(n_42042) );
ao12s01 g738122 ( .a(n_41809), .b(n_42030), .c(n_41830), .o(n_42041) );
oa22s01 g738123 ( .a(n_42016), .b(n_41856), .c(n_42029), .d(n_41857), .o(n_42570) );
in01s01 g738124 ( .a(n_42052), .o(n_42053) );
oa12s01 g738125 ( .a(n_42024), .b(n_42031), .c(n_42023), .o(n_42052) );
in01s01 g738126 ( .a(n_42072), .o(n_42093) );
oa12s01 g738127 ( .a(n_42022), .b(n_42021), .c(n_42020), .o(n_42072) );
oa12s01 g738128 ( .a(n_42080), .b(n_42079), .c(n_42078), .o(n_42421) );
in01s01 g738129 ( .a(n_42050), .o(n_42069) );
in01f04 g738131 ( .a(n_42051), .o(n_42050) );
ao12s01 g738133 ( .a(n_42019), .b(n_42018), .c(n_42017), .o(n_42321) );
in01s01 g738134 ( .a(n_42107), .o(n_42081) );
na02s01 g738135 ( .a(n_42040), .b(n_42028), .o(n_42107) );
na02s01 g738136 ( .a(n_42031), .b(n_42023), .o(n_42024) );
na02s01 g738137 ( .a(n_42021), .b(n_42020), .o(n_42022) );
no02s01 g738138 ( .a(n_42029), .b(n_41708), .o(n_42059) );
no02s01 g738139 ( .a(n_42018), .b(n_42017), .o(n_42019) );
na02s01 g738140 ( .a(n_42012), .b(n_41853), .o(n_42040) );
na02s01 g738141 ( .a(n_42011), .b(n_41854), .o(n_42028) );
na02s01 g738142 ( .a(n_42079), .b(n_42078), .o(n_42080) );
no02s01 g738143 ( .a(n_42066), .b(n_42065), .o(n_42067) );
na02s01 g738144 ( .a(n_42066), .b(n_42065), .o(n_42064) );
oa12s01 g738145 ( .a(n_41721), .b(n_42027), .c(n_41658), .o(n_42057) );
ao12f08 g738147 ( .a(n_41741), .b(n_42027), .c(n_41762), .o(n_42038) );
no02s01 g738148 ( .a(n_42025), .b(n_41770), .o(n_42105) );
in01s01 g738149 ( .a(n_42071), .o(n_42037) );
na02s01 g738150 ( .a(n_42004), .b(n_41793), .o(n_42071) );
in01s01 g738151 ( .a(n_42115), .o(n_42049) );
ao12s01 g738152 ( .a(n_42015), .b(n_42027), .c(n_42014), .o(n_42115) );
in01s01 g738153 ( .a(n_42076), .o(n_42077) );
ao12s01 g738154 ( .a(n_42034), .b(n_42033), .c(n_42032), .o(n_42076) );
na02f08 g738155 ( .a(n_42005), .b(n_41908), .o(n_42070) );
in01s01 g738156 ( .a(n_42046), .o(n_42026) );
oa22s01 g738157 ( .a(n_41981), .b(n_41851), .c(n_41980), .d(n_41852), .o(n_42046) );
in01s01 g738158 ( .a(n_42035), .o(n_42036) );
oa12s01 g738159 ( .a(n_42000), .b(n_41999), .c(n_41998), .o(n_42035) );
oa12s01 g738160 ( .a(n_42002), .b(n_42003), .c(n_42001), .o(n_42542) );
in01s01 g738161 ( .a(n_42029), .o(n_42016) );
in01s01 g738162 ( .a(n_42030), .o(n_42029) );
no02m02 TIMEBOOST_cell_8835 ( .a(TIMEBOOST_net_2904), .b(n_5221), .o(n_5458) );
na02s01 g738165 ( .a(n_42003), .b(n_41706), .o(n_42004) );
na02s01 g738166 ( .a(n_42003), .b(n_42001), .o(n_42002) );
no02s01 g738167 ( .a(n_42006), .b(n_41912), .o(n_42025) );
no02s01 g738168 ( .a(n_42033), .b(n_42032), .o(n_42034) );
na02s01 g738169 ( .a(n_41999), .b(n_41998), .o(n_42000) );
no02s01 g738170 ( .a(n_42027), .b(n_42014), .o(n_42015) );
ao12s01 g738171 ( .a(n_41788), .b(n_41995), .c(n_41761), .o(n_42031) );
in01f02 g738172 ( .a(n_41996), .o(n_41997) );
ao12f06 g738173 ( .a(n_41858), .b(n_41995), .c(n_41810), .o(n_41996) );
ao12s01 g738174 ( .a(n_41878), .b(n_41995), .c(n_41901), .o(n_42021) );
no02s06 TIMEBOOST_cell_1896 ( .a(TIMEBOOST_net_562), .b(n_40251), .o(n_40332) );
oa12s01 g738176 ( .a(n_41775), .b(n_41985), .c(n_41667), .o(n_42018) );
in01s01 g738177 ( .a(n_42013), .o(n_42710) );
oa12s01 g738178 ( .a(n_41987), .b(n_41995), .c(n_41986), .o(n_42013) );
in01s01 g738179 ( .a(n_42066), .o(n_42048) );
ao12s01 g738180 ( .a(n_42010), .b(n_42009), .c(n_42008), .o(n_42066) );
ao12s01 g738181 ( .a(n_41970), .b(n_41969), .c(n_41968), .o(n_42304) );
in01s01 g738182 ( .a(n_42011), .o(n_42012) );
ao12s01 g738183 ( .a(n_41863), .b(n_41973), .c(n_41694), .o(n_42011) );
no02s01 g738184 ( .a(n_41969), .b(n_41968), .o(n_41970) );
na02s01 g738185 ( .a(n_41995), .b(n_41986), .o(n_41987) );
na02s01 g738186 ( .a(n_41974), .b(n_41862), .o(n_42003) );
no02s01 g738187 ( .a(n_42009), .b(n_42008), .o(n_42010) );
in01s01 g738188 ( .a(n_42006), .o(n_42007) );
na02s01 g738189 ( .a(n_41989), .b(n_41662), .o(n_42006) );
na02s01 g738190 ( .a(n_41990), .b(n_41729), .o(n_42033) );
na02s01 g738191 ( .a(n_41985), .b(n_41792), .o(n_41999) );
na02s01 g738192 ( .a(n_41993), .b(n_41992), .o(n_41994) );
na02s01 g738193 ( .a(n_41983), .b(n_41982), .o(n_41984) );
no02s01 TIMEBOOST_cell_3044 ( .a(n_2946), .b(n_2849), .o(TIMEBOOST_net_813) );
in01s01 g738195 ( .a(n_41980), .o(n_41981) );
ao12s01 g738196 ( .a(n_41585), .b(n_41977), .c(n_41814), .o(n_41980) );
na02f08 g738197 ( .a(n_41976), .b(n_41859), .o(n_42027) );
in01s01 g738198 ( .a(n_41991), .o(n_42423) );
ao12s01 g738199 ( .a(n_41967), .b(n_41966), .c(n_41965), .o(n_41991) );
oa12s01 g738200 ( .a(n_41964), .b(n_41977), .c(n_41963), .o(n_42500) );
na02s08 TIMEBOOST_cell_7986 ( .a(n_30936), .b(FE_OCP_RBN5335_FE_RN_1144_0), .o(TIMEBOOST_net_2624) );
no02s01 g738203 ( .a(n_41966), .b(n_41965), .o(n_41967) );
in01s01 g738204 ( .a(n_41989), .o(n_41990) );
no02s01 g738205 ( .a(n_41971), .b(n_41828), .o(n_41989) );
no02s01 g738206 ( .a(n_41972), .b(n_41803), .o(n_42009) );
na02s01 g738207 ( .a(n_41977), .b(n_41749), .o(n_41985) );
na02s01 g738208 ( .a(n_41977), .b(n_41963), .o(n_41964) );
na02s01 g738209 ( .a(n_41953), .b(n_41952), .o(n_41954) );
oa12s01 g738210 ( .a(n_41674), .b(n_41946), .c(n_41510), .o(n_41969) );
in01f06 g738212 ( .a(n_41974), .o(n_41973) );
in01f04 g738213 ( .a(n_41962), .o(n_41974) );
in01s01 g738215 ( .a(n_41983), .o(n_41993) );
oa12s01 g738216 ( .a(n_41945), .b(n_41944), .c(n_41943), .o(n_41983) );
in01s01 g738217 ( .a(n_42065), .o(n_41988) );
ao12s01 g738218 ( .a(n_41958), .b(n_41924), .c(n_41957), .o(n_42065) );
in01s01 g738219 ( .a(n_41960), .o(n_41961) );
oa12s01 g738220 ( .a(n_41934), .b(n_41946), .c(n_41933), .o(n_41960) );
na02s01 g738221 ( .a(n_41944), .b(n_41943), .o(n_41945) );
na02s01 g738222 ( .a(n_41946), .b(n_41933), .o(n_41934) );
in01s01 g738223 ( .a(n_41971), .o(n_41972) );
na02s01 g738224 ( .a(n_41924), .b(n_41850), .o(n_41971) );
no02s01 g738225 ( .a(n_41924), .b(n_41957), .o(n_41958) );
no02s01 g738228 ( .a(n_41949), .b(n_41947), .o(n_41948) );
oa12s01 g738230 ( .a(n_41663), .b(n_41940), .c(n_41558), .o(n_41966) );
in01s01 g738231 ( .a(n_41939), .o(n_41977) );
no03s01 TIMEBOOST_cell_7460 ( .a(TIMEBOOST_net_1387), .b(n_32608), .c(n_32561), .o(TIMEBOOST_net_2361) );
ao12s01 g738233 ( .a(n_41926), .b(n_41940), .c(n_41925), .o(n_42366) );
in01s01 g738234 ( .a(n_41956), .o(n_42374) );
ao12s01 g738235 ( .a(n_41929), .b(n_41928), .c(n_41927), .o(n_41956) );
in01s01 g738236 ( .a(n_41955), .o(n_42276) );
oa12s01 g738237 ( .a(n_41932), .b(n_41931), .c(n_41930), .o(n_41955) );
in01s01 g738238 ( .a(n_41953), .o(n_42272) );
oa12s01 g738239 ( .a(n_41900), .b(n_41899), .c(n_41898), .o(n_41953) );
na02s01 g738240 ( .a(n_41896), .b(n_41753), .o(n_41946) );
na02s01 g738241 ( .a(n_41931), .b(n_41930), .o(n_41932) );
na02s01 g738242 ( .a(n_41899), .b(n_41898), .o(n_41900) );
no02s01 g738243 ( .a(n_41928), .b(n_41927), .o(n_41929) );
no02s01 g738244 ( .a(n_41940), .b(n_41925), .o(n_41926) );
oa12s01 g738245 ( .a(n_41826), .b(n_41919), .c(n_41879), .o(n_41944) );
no02m04 TIMEBOOST_cell_7459 ( .a(TIMEBOOST_net_2360), .b(n_23038), .o(TIMEBOOST_net_132) );
oa12f10 g738250 ( .a(n_41693), .b(n_41919), .c(n_41666), .o(n_41924) );
in01s01 g738251 ( .a(n_41982), .o(n_41992) );
oa12s01 g738252 ( .a(n_41920), .b(n_41919), .c(n_41918), .o(n_41982) );
in01s01 g738253 ( .a(n_42358), .o(n_41936) );
oa12s01 g738254 ( .a(n_41895), .b(n_41894), .c(n_41893), .o(n_42358) );
ao12s01 g738255 ( .a(n_41892), .b(n_41891), .c(n_41890), .o(n_42312) );
in01s01 g738256 ( .a(n_41949), .o(n_41923) );
oa12s01 g738257 ( .a(n_41871), .b(n_41870), .c(n_41869), .o(n_41949) );
in01s01 g738258 ( .a(n_41921), .o(n_41922) );
ao12s01 g738259 ( .a(n_41874), .b(n_41873), .c(n_41872), .o(n_41921) );
in01s01 g738260 ( .a(n_41952), .o(n_42271) );
oa12s01 g738261 ( .a(n_41847), .b(n_41846), .c(n_41845), .o(n_41952) );
no02s01 g738262 ( .a(n_41873), .b(n_41872), .o(n_41874) );
na02s01 g738263 ( .a(n_41870), .b(n_41869), .o(n_41871) );
na02s01 g738264 ( .a(n_41919), .b(n_41918), .o(n_41920) );
na02s01 g738265 ( .a(n_41894), .b(n_41893), .o(n_41895) );
no02s01 g738266 ( .a(n_41891), .b(n_41890), .o(n_41892) );
na02s01 g738267 ( .a(n_41846), .b(n_41845), .o(n_41847) );
na02f08 g738268 ( .a(n_41846), .b(n_41641), .o(n_41896) );
oa12s01 g738269 ( .a(n_41512), .b(n_41776), .c(n_41548), .o(n_41931) );
oa12s01 g738270 ( .a(n_41712), .b(n_41801), .c(n_41640), .o(n_41899) );
ao12s01 g738271 ( .a(n_41673), .b(n_41844), .c(n_41577), .o(n_41928) );
oa12s01 g738272 ( .a(n_41734), .b(n_41824), .c(n_41619), .o(n_41940) );
no02s01 g738273 ( .a(n_41777), .b(n_41595), .o(n_41873) );
no02f10 g738274 ( .a(n_41823), .b(n_41733), .o(n_41919) );
no02s01 g738275 ( .a(n_41844), .b(n_41620), .o(n_41891) );
na02f08 g738276 ( .a(n_41801), .b(n_41646), .o(n_41846) );
ao12s01 g738277 ( .a(n_41786), .b(n_41888), .c(n_41825), .o(n_41870) );
oa12s01 g738278 ( .a(n_41502), .b(n_41865), .c(n_41807), .o(n_41894) );
oa12s01 g738279 ( .a(n_41866), .b(n_41865), .c(n_41864), .o(n_42562) );
in01s01 g738280 ( .a(n_41947), .o(n_42478) );
oa12s01 g738281 ( .a(n_41889), .b(n_41888), .c(n_41887), .o(n_41947) );
in01s01 g738282 ( .a(n_42232), .o(n_41911) );
ao12s01 g738283 ( .a(n_41843), .b(n_41842), .c(n_41841), .o(n_42232) );
in01s01 g738284 ( .a(n_41867), .o(n_41868) );
oa12s01 g738285 ( .a(n_41800), .b(n_41799), .c(n_41798), .o(n_41867) );
in01s01 g738286 ( .a(n_42212), .o(n_41910) );
ao12s01 g738287 ( .a(n_41840), .b(n_41839), .c(n_41838), .o(n_42212) );
no02s01 g738288 ( .a(n_41842), .b(n_41841), .o(n_41843) );
no02s01 g738289 ( .a(n_41839), .b(n_41838), .o(n_41840) );
in01s01 g738290 ( .a(n_41776), .o(n_41777) );
na02s01 g738291 ( .a(n_41888), .b(n_41550), .o(n_41776) );
na02s01 g738292 ( .a(n_41799), .b(n_41798), .o(n_41800) );
no02s01 g738293 ( .a(n_41865), .b(n_41480), .o(n_41844) );
na02s01 g738294 ( .a(n_41865), .b(n_41864), .o(n_41866) );
na02s01 g738295 ( .a(n_41888), .b(n_41887), .o(n_41889) );
no02s01 g738296 ( .a(n_41916), .b(n_41915), .o(n_41917) );
in01s01 g738297 ( .a(n_41823), .o(n_41824) );
no02f10 g738298 ( .a(n_41865), .b(n_41578), .o(n_41823) );
na02f08 g738299 ( .a(n_41888), .b(n_41594), .o(n_41801) );
oa12s01 g738300 ( .a(n_41837), .b(n_41836), .c(n_41835), .o(n_42286) );
na02s01 g738301 ( .a(n_41836), .b(n_41835), .o(n_41837) );
oa12f08 g738302 ( .a(n_41485), .b(n_41757), .c(n_41593), .o(n_41865) );
oa12s01 g738303 ( .a(n_41424), .b(n_41648), .c(n_41455), .o(n_41799) );
oa12f08 g738304 ( .a(n_41522), .b(n_41648), .c(n_41524), .o(n_41888) );
oa12s01 g738305 ( .a(n_41744), .b(n_41648), .c(n_41769), .o(n_41839) );
oa12s01 g738306 ( .a(n_41454), .b(n_41648), .c(n_41477), .o(n_41842) );
in01s01 g738307 ( .a(n_41796), .o(n_41797) );
ao12s01 g738308 ( .a(n_41738), .b(n_41737), .c(n_41736), .o(n_41796) );
in01s01 g738309 ( .a(n_41916), .o(n_41909) );
oa12s01 g738310 ( .a(n_41834), .b(n_41833), .c(n_41832), .o(n_41916) );
in01s01 g738311 ( .a(n_42191), .o(n_41886) );
ao12s01 g738312 ( .a(n_41822), .b(n_41648), .c(n_41820), .o(n_42191) );
no02s01 g738313 ( .a(n_41737), .b(n_41736), .o(n_41738) );
no02s01 g738314 ( .a(n_41648), .b(n_41820), .o(n_41822) );
na02s01 g738315 ( .a(n_41833), .b(n_41832), .o(n_41834) );
no02f04 TIMEBOOST_cell_1828 ( .a(TIMEBOOST_net_528), .b(n_15951), .o(n_16047) );
oa12s01 g738318 ( .a(n_41541), .b(n_41818), .c(n_41683), .o(n_41737) );
no02s06 g738319 ( .a(n_41861), .b(n_41756), .o(n_41908) );
na02s04 g738320 ( .a(n_41831), .b(n_41755), .o(n_41885) );
oa12f08 g738324 ( .a(n_41475), .b(n_41596), .c(n_41426), .o(n_41648) );
oa12s01 g738325 ( .a(n_41445), .b(n_41818), .c(n_41760), .o(n_41833) );
in01s01 g738326 ( .a(n_41915), .o(n_41884) );
oa12s01 g738327 ( .a(n_41819), .b(n_41818), .c(n_41817), .o(n_41915) );
in01s01 g738328 ( .a(n_42209), .o(n_42267) );
ao12s01 g738329 ( .a(n_41553), .b(n_41596), .c(n_41552), .o(n_42209) );
na02s01 g738330 ( .a(n_41862), .b(n_41699), .o(n_41863) );
na02s01 g738331 ( .a(n_41818), .b(n_41817), .o(n_41819) );
no02s01 g738332 ( .a(n_41647), .b(n_41624), .o(n_41712) );
no02s01 g738333 ( .a(n_41596), .b(n_41552), .o(n_41553) );
in01s02 g738334 ( .a(n_41860), .o(n_41861) );
no02m06 g738335 ( .a(n_41816), .b(n_41794), .o(n_41860) );
na03m08 TIMEBOOST_cell_7368 ( .a(n_34113), .b(n_34026), .c(n_34126), .o(n_34223) );
na02f06 g738337 ( .a(n_41476), .b(n_41523), .o(n_41524) );
no02s01 g738338 ( .a(n_41732), .b(n_41668), .o(n_41775) );
no02m08 g738339 ( .a(n_41790), .b(n_41813), .o(n_41859) );
ao12m06 g738340 ( .a(n_41453), .b(n_41434), .c(FE_OCP_RBN5639_n_41381), .o(n_41522) );
no03f06 TIMEBOOST_cell_8333 ( .a(n_15464), .b(n_15421), .c(n_15535), .o(n_15679) );
in01s02 g738342 ( .a(n_41755), .o(n_41756) );
ao12s02 g738343 ( .a(n_41735), .b(n_41639), .c(FE_OCP_RBN5676_n_41420), .o(n_41755) );
na02s04 g738344 ( .a(n_41793), .b(n_41711), .o(n_41794) );
in01s01 g738345 ( .a(n_41816), .o(n_41862) );
na03s02 TIMEBOOST_cell_2754 ( .a(FE_OCP_RBN6223_n_27110), .b(n_27210), .c(n_27211), .o(n_27351) );
na02s06 g738348 ( .a(n_41753), .b(n_41645), .o(n_41754) );
in01s01 g738349 ( .a(n_41646), .o(n_41647) );
ao12m04 g738350 ( .a(n_41595), .b(n_41474), .c(FE_OCP_RBN5674_n_41420), .o(n_41646) );
oa12f08 g738351 ( .a(n_41449), .b(n_41551), .c(n_41399), .o(n_41818) );
no02m04 g738352 ( .a(n_41773), .b(n_41752), .o(n_41791) );
oa12f08 g738353 ( .a(n_41408), .b(n_41517), .c(n_41452), .o(n_41596) );
in01s01 g738354 ( .a(n_42241), .o(n_42335) );
oa12s01 g738355 ( .a(n_41521), .b(n_41551), .c(n_41520), .o(n_42241) );
oa12s01 g738356 ( .a(n_41519), .b(n_41518), .c(n_41517), .o(n_42188) );
in01s01 g738357 ( .a(n_41476), .o(n_41477) );
no02f06 g738358 ( .a(n_41455), .b(n_41410), .o(n_41476) );
na02s04 g738359 ( .a(n_41751), .b(n_41745), .o(n_41752) );
no02s01 g738360 ( .a(n_41733), .b(n_41692), .o(n_41734) );
na02s01 g738361 ( .a(n_41520), .b(n_41551), .o(n_41521) );
na02s01 g738362 ( .a(n_41518), .b(n_41517), .o(n_41519) );
no02s06 g738364 ( .a(n_41549), .b(n_41514), .o(n_41594) );
in01s02 g738365 ( .a(n_41773), .o(n_41774) );
na02s06 g738366 ( .a(n_41709), .b(n_41643), .o(n_41773) );
no02s06 g738367 ( .a(n_41705), .b(n_41678), .o(n_41978) );
in01s01 g738368 ( .a(n_41771), .o(n_41772) );
no02s02 TIMEBOOST_cell_4117 ( .a(FE_RN_2139_0), .b(FE_OCP_RBN2907_n_25238), .o(TIMEBOOST_net_1149) );
na02s02 g738370 ( .a(n_41700), .b(FE_OCP_RBN5673_n_41420), .o(n_41793) );
na02s02 g738371 ( .a(n_41636), .b(FE_OCP_RBN5673_n_41420), .o(n_41711) );
in01s01 g738372 ( .a(n_41792), .o(n_41732) );
na02s04 g738373 ( .a(n_41633), .b(FE_OCP_RBN5674_n_41420), .o(n_41792) );
na04s10 TIMEBOOST_cell_8199 ( .a(FE_RN_2530_0), .b(n_17579), .c(FE_RN_2529_0), .d(FE_RN_969_0), .o(n_17762) );
na02s06 g738375 ( .a(n_41630), .b(FE_OCP_RBN5674_n_41420), .o(n_41753) );
na02s06 g738376 ( .a(n_41547), .b(FE_OCP_RBN5674_n_41420), .o(n_41645) );
in01m04 g738377 ( .a(n_41789), .o(n_41790) );
no02m08 g738378 ( .a(n_41727), .b(n_41770), .o(n_41789) );
na03f02 TIMEBOOST_cell_7768 ( .a(n_9707), .b(n_9840), .c(n_9706), .o(TIMEBOOST_net_2515) );
in01s01 g738380 ( .a(n_41515), .o(n_41516) );
oa12s01 g738381 ( .a(n_41432), .b(n_41431), .c(n_41430), .o(n_41515) );
na02s02 g738383 ( .a(n_41513), .b(n_41472), .o(n_41514) );
in01s01 g738384 ( .a(n_41549), .o(n_41550) );
na02s04 g738385 ( .a(n_41470), .b(n_41825), .o(n_41549) );
no02s02 g738386 ( .a(n_41642), .b(n_41588), .o(n_41643) );
na02s01 g738387 ( .a(n_41621), .b(n_41638), .o(n_41710) );
na02f04 g738388 ( .a(n_41416), .b(n_41391), .o(n_41455) );
in01s02 g738389 ( .a(n_41708), .o(n_41709) );
na02s02 g738390 ( .a(n_41680), .b(n_41830), .o(n_41708) );
no02s03 g738391 ( .a(n_41707), .b(n_41671), .o(n_41751) );
no02s01 g738392 ( .a(n_41453), .b(n_41428), .o(n_41454) );
no02s01 g738393 ( .a(n_41595), .b(n_41511), .o(n_41512) );
in01s01 g738394 ( .a(n_41705), .o(n_41706) );
na02s06 g738395 ( .a(n_41679), .b(n_41694), .o(n_41705) );
na02s03 g738396 ( .a(n_41677), .b(n_41676), .o(n_41678) );
na02s06 g738397 ( .a(n_41622), .b(n_41674), .o(n_41675) );
no02s02 g738398 ( .a(n_41580), .b(n_41640), .o(n_41641) );
in01s01 g738399 ( .a(n_41703), .o(n_41704) );
na02s01 g738400 ( .a(n_41677), .b(n_41635), .o(n_41703) );
in01s01 g738401 ( .a(n_41856), .o(n_41857) );
na02s01 g738402 ( .a(n_41830), .b(n_41808), .o(n_41856) );
na02m04 g738403 ( .a(n_41414), .b(n_41433), .o(n_41434) );
no02s01 g738404 ( .a(n_41642), .b(n_41587), .o(n_42095) );
no02m01 TIMEBOOST_cell_4116 ( .a(TIMEBOOST_net_1148), .b(n_36036), .o(n_36194) );
na02s01 g738406 ( .a(n_41731), .b(n_41701), .o(n_42054) );
na02s01 g738407 ( .a(n_41787), .b(n_41825), .o(n_41887) );
na02s01 g738408 ( .a(n_41411), .b(n_41414), .o(n_41798) );
na02s01 g738409 ( .a(n_41475), .b(n_41427), .o(n_41552) );
no02s01 g738410 ( .a(n_41743), .b(n_41769), .o(n_41820) );
no02s01 g738411 ( .a(n_41511), .b(n_41548), .o(n_41872) );
na02s01 g738412 ( .a(n_41638), .b(n_41637), .o(n_41639) );
na02s01 g738413 ( .a(n_41579), .b(n_41583), .o(n_41845) );
na02s02 g738414 ( .a(n_41699), .b(n_41698), .o(n_41700) );
na02s02 g738415 ( .a(n_41635), .b(n_41634), .o(n_41636) );
na02s01 g738416 ( .a(n_41674), .b(n_41546), .o(n_41933) );
na02s02 g738417 ( .a(n_41632), .b(n_41631), .o(n_41633) );
na02f08 TIMEBOOST_cell_7787 ( .a(TIMEBOOST_net_2524), .b(n_42239), .o(n_42290) );
na02s01 g738419 ( .a(n_41814), .b(n_41632), .o(n_41963) );
na02s01 g738420 ( .a(n_41730), .b(n_41696), .o(n_41998) );
na02s06 g738421 ( .a(n_41583), .b(n_41629), .o(n_41630) );
na02s06 g738422 ( .a(n_41546), .b(n_41545), .o(n_41547) );
na02s01 g738423 ( .a(n_41694), .b(n_41699), .o(n_42001) );
na02m04 g738424 ( .a(n_41450), .b(n_41473), .o(n_41474) );
na02s01 g738425 ( .a(n_41672), .b(n_41499), .o(n_41673) );
na02m02 TIMEBOOST_cell_8602 ( .a(n_15898), .b(n_14730), .o(TIMEBOOST_net_2788) );
oa12m06 g738427 ( .a(n_41729), .b(FE_OCP_RBN6585_n_41491), .c(n_41615), .o(n_41770) );
in01s03 g738428 ( .a(n_41812), .o(n_41813) );
no02s06 g738429 ( .a(n_41742), .b(n_41788), .o(n_41812) );
oa12m04 g738430 ( .a(n_41598), .b(n_41478), .c(n_41612), .o(n_41727) );
ao12m08 g738431 ( .a(n_41692), .b(FE_OCP_RBN6590_n_41491), .c(n_41566), .o(n_41693) );
na02f08 g738432 ( .a(n_41541), .b(n_41506), .o(n_41593) );
na02m08 g738433 ( .a(n_41672), .b(n_41573), .o(n_41733) );
na02s01 g738434 ( .a(n_41431), .b(n_41430), .o(n_41432) );
no02s01 g738435 ( .a(n_41452), .b(n_41409), .o(n_41518) );
in01s01 g738436 ( .a(n_41906), .o(n_41907) );
oa12s01 g738437 ( .a(n_41676), .b(FE_OCPN884_n_41540), .c(n_41634), .o(n_41906) );
in01s01 g738438 ( .a(n_41904), .o(n_41905) );
oa12s01 g738439 ( .a(n_41680), .b(FE_OCPN884_n_41540), .c(n_41590), .o(n_41904) );
in01s01 g738440 ( .a(n_41902), .o(n_41903) );
oa12s01 g738441 ( .a(n_41589), .b(FE_OCPN884_n_41540), .c(n_41637), .o(n_41902) );
in01s01 g738442 ( .a(n_41766), .o(n_41767) );
na02s01 g738443 ( .a(n_41691), .b(n_41745), .o(n_41766) );
in01s01 g738444 ( .a(n_41881), .o(n_41882) );
ao12s01 g738445 ( .a(n_41707), .b(n_41660), .c(n_41310), .o(n_41881) );
ao12s01 g738446 ( .a(n_41471), .b(n_41660), .c(n_41156), .o(n_41869) );
oa12s01 g738447 ( .a(n_41523), .b(FE_OCPN884_n_41540), .c(n_41433), .o(n_41841) );
oa12s01 g738448 ( .a(n_41416), .b(FE_OCPN884_n_41540), .c(n_41407), .o(n_41838) );
oa12s01 g738449 ( .a(n_41513), .b(FE_OCPN884_n_41540), .c(n_41473), .o(n_41930) );
oa12s01 g738450 ( .a(n_41581), .b(FE_OCPN884_n_41540), .c(n_41629), .o(n_41898) );
ao12s01 g738451 ( .a(n_41623), .b(n_41660), .c(n_41180), .o(n_41968) );
oa12s01 g738452 ( .a(n_41748), .b(FE_OCPN884_n_41540), .c(n_41695), .o(n_42017) );
in01s01 g738453 ( .a(n_41853), .o(n_41854) );
oa12s01 g738454 ( .a(n_41679), .b(FE_OCPN884_n_41540), .c(n_41698), .o(n_41853) );
no02s04 g738455 ( .a(n_41784), .b(n_41763), .o(n_41810) );
no02f08 g738456 ( .a(n_41380), .b(n_41388), .o(n_41517) );
ao12s01 g738457 ( .a(n_41509), .b(n_41508), .c(n_41507), .o(n_42211) );
oa12f06 g738458 ( .a(n_41443), .b(n_41405), .c(n_41397), .o(n_41551) );
in01s01 g738459 ( .a(n_41851), .o(n_41852) );
oa22s01 g738460 ( .a(n_41660), .b(n_41275), .c(FE_OCPN884_n_41540), .d(n_41631), .o(n_41851) );
in01s01 g738461 ( .a(n_41764), .o(n_41765) );
na02s01 g738462 ( .a(n_41669), .b(n_41690), .o(n_41764) );
na02m04 g738463 ( .a(n_41762), .b(n_41759), .o(n_41763) );
na02s02 g738464 ( .a(FE_OCP_RBN5637_n_41381), .b(n_41473), .o(n_41513) );
in01s01 g738465 ( .a(n_41472), .o(n_41548) );
na02s02 g738466 ( .a(FE_OCP_RBN5637_n_41381), .b(n_41173), .o(n_41472) );
in01s01 g738467 ( .a(n_41470), .o(n_41471) );
na02s02 g738468 ( .a(FE_OCP_RBN5637_n_41381), .b(n_41153), .o(n_41470) );
na02s02 g738469 ( .a(FE_OCP_RBN5637_n_41381), .b(n_41415), .o(n_41825) );
in01s01 g738471 ( .a(n_41414), .o(n_41428) );
na02m02 g738472 ( .a(FE_OCP_RBN4115_n_41381), .b(n_41392), .o(n_41414) );
in01s01 g738473 ( .a(n_41808), .o(n_41809) );
na02s01 g738474 ( .a(n_41660), .b(n_41320), .o(n_41808) );
in01s01 g738475 ( .a(n_41426), .o(n_41427) );
no02s06 g738476 ( .a(FE_OCP_RBN6619_n_41381), .b(n_41412), .o(n_41426) );
na02s03 g738477 ( .a(FE_OCP_RBN6618_n_41381), .b(n_41412), .o(n_41475) );
in01s01 g738478 ( .a(n_41642), .o(n_41592) );
no02s01 g738479 ( .a(FE_OCP_RBN5673_n_41420), .b(n_41543), .o(n_41642) );
in01s01 g738480 ( .a(n_41410), .o(n_41411) );
no02s02 g738481 ( .a(FE_OCP_RBN4115_n_41381), .b(n_41392), .o(n_41410) );
na02s02 g738482 ( .a(n_41381), .b(n_41407), .o(n_41416) );
na02s02 g738483 ( .a(n_41582), .b(n_41292), .o(n_41830) );
in01s01 g738484 ( .a(n_41391), .o(n_41769) );
na02f01 g738485 ( .a(n_41381), .b(n_41406), .o(n_41391) );
na02s02 g738486 ( .a(n_41582), .b(n_41590), .o(n_41680) );
in01s01 g738487 ( .a(n_41588), .o(n_41589) );
no02s01 g738488 ( .a(FE_OCP_RBN5673_n_41420), .b(n_41347), .o(n_41588) );
na02s02 g738489 ( .a(FE_OCP_RBN5637_n_41381), .b(n_41433), .o(n_41523) );
no02m01 g738490 ( .a(FE_OCP_RBN5676_n_41420), .b(n_41310), .o(n_41707) );
in01s01 g738491 ( .a(n_41671), .o(n_41731) );
no02s02 g738492 ( .a(FE_OCP_RBN5676_n_41420), .b(n_41628), .o(n_41671) );
in01s01 g738493 ( .a(n_41701), .o(n_41670) );
na02s02 g738494 ( .a(FE_OCP_RBN5676_n_41420), .b(n_41628), .o(n_41701) );
na02s01 g738495 ( .a(n_41660), .b(n_41330), .o(n_41691) );
na02s01 g738496 ( .a(n_41540), .b(n_41345), .o(n_41745) );
na02s01 g738497 ( .a(n_41540), .b(n_41298), .o(n_41669) );
na02s01 g738498 ( .a(FE_OCP_RBN5676_n_41420), .b(FE_OCP_RBN4046_n_41298), .o(n_41690) );
in01s01 g738499 ( .a(n_41786), .o(n_41787) );
no02s01 g738500 ( .a(FE_OCPN884_n_41540), .b(n_41415), .o(n_41786) );
in01s01 g738501 ( .a(n_41743), .o(n_41744) );
no02s01 g738502 ( .a(FE_OCPN884_n_41540), .b(n_41406), .o(n_41743) );
in01s01 g738503 ( .a(n_41638), .o(n_41587) );
na02s02 g738504 ( .a(FE_OCP_RBN5673_n_41420), .b(n_41543), .o(n_41638) );
na02s02 g738505 ( .a(FE_OCP_RBN5673_n_41420), .b(n_41290), .o(n_41699) );
in01s01 g738506 ( .a(n_41635), .o(n_41586) );
na02s02 g738507 ( .a(FE_OCP_RBN5673_n_41420), .b(n_41317), .o(n_41635) );
in01s01 g738508 ( .a(n_41632), .o(n_41585) );
na02s04 g738509 ( .a(FE_OCP_RBN5674_n_41420), .b(n_41219), .o(n_41632) );
na02s01 g738510 ( .a(FE_OCPN884_n_41540), .b(n_41576), .o(n_41814) );
in01s01 g738511 ( .a(n_41696), .o(n_41668) );
na02s02 g738512 ( .a(FE_OCP_RBN5674_n_41420), .b(n_41626), .o(n_41696) );
na02s02 g738513 ( .a(n_41582), .b(n_41291), .o(n_41694) );
na02s03 g738514 ( .a(n_41540), .b(n_41698), .o(n_41679) );
na02s01 g738515 ( .a(n_41420), .b(n_41316), .o(n_41677) );
na02s02 g738516 ( .a(n_41420), .b(n_41634), .o(n_41676) );
in01s01 g738517 ( .a(n_41667), .o(n_41730) );
no02s01 g738518 ( .a(FE_OCP_RBN5674_n_41420), .b(n_41626), .o(n_41667) );
na02s01 g738519 ( .a(n_41695), .b(n_41582), .o(n_41748) );
in01s01 g738521 ( .a(n_41583), .o(n_41624) );
na02s06 g738522 ( .a(FE_OCP_RBN5674_n_41420), .b(n_41542), .o(n_41583) );
na02s03 g738523 ( .a(n_41582), .b(n_41176), .o(n_41674) );
in01s01 g738524 ( .a(n_41546), .o(n_41510) );
na02s06 g738525 ( .a(FE_OCP_RBN5674_n_41420), .b(n_41175), .o(n_41546) );
in01s01 g738526 ( .a(n_41622), .o(n_41623) );
na02s06 g738527 ( .a(n_41582), .b(n_41545), .o(n_41622) );
in01s01 g738528 ( .a(n_41580), .o(n_41581) );
no02s02 g738529 ( .a(FE_OCP_RBN5674_n_41420), .b(n_41218), .o(n_41580) );
in01s01 g738530 ( .a(n_41640), .o(n_41579) );
no02s02 g738531 ( .a(FE_OCP_RBN5674_n_41420), .b(n_41542), .o(n_41640) );
in01s01 g738532 ( .a(n_41450), .o(n_41511) );
na02s02 g738533 ( .a(FE_OCP_RBN5638_n_41381), .b(n_41174), .o(n_41450) );
in01s01 g738534 ( .a(n_41408), .o(n_41409) );
na02s04 g738535 ( .a(n_41390), .b(n_41389), .o(n_41408) );
no02f04 g738536 ( .a(n_41390), .b(n_41389), .o(n_41452) );
no02f04 g738537 ( .a(n_41379), .b(n_41430), .o(n_41380) );
no02s01 g738538 ( .a(n_41508), .b(n_41507), .o(n_41509) );
no02s01 g738539 ( .a(n_41379), .b(n_41388), .o(n_41431) );
in01s04 g738541 ( .a(n_41784), .o(n_41785) );
na02s06 g738542 ( .a(n_41761), .b(n_41723), .o(n_41784) );
na02f08 g738543 ( .a(n_41618), .b(n_41572), .o(n_41666) );
no02s02 g738544 ( .a(n_41420), .b(n_41157), .o(n_41595) );
in01s01 g738545 ( .a(n_41453), .o(n_41424) );
in01s01 g738547 ( .a(n_41735), .o(n_41621) );
no02s01 g738548 ( .a(n_41582), .b(n_41321), .o(n_41735) );
oa12s01 g738549 ( .a(n_41420), .b(n_41631), .c(n_41576), .o(n_41749) );
na02s06 TIMEBOOST_cell_3888 ( .a(n_1921), .b(TIMEBOOST_net_1034), .o(n_1987) );
na02s02 TIMEBOOST_cell_7770 ( .a(n_42129), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(TIMEBOOST_net_2516) );
in01s01 g738553 ( .a(n_41541), .o(n_41574) );
na02f06 g738554 ( .a(n_41446), .b(n_41382), .o(n_41541) );
na02m04 g738555 ( .a(n_41500), .b(n_41483), .o(n_41573) );
in01s01 g738556 ( .a(n_41672), .o(n_41620) );
no03m08 TIMEBOOST_cell_8383 ( .a(n_10505), .b(FE_OCP_RBN3182_n_10477), .c(n_44492), .o(n_10612) );
in01s02 g738558 ( .a(n_41740), .o(n_41741) );
na02m01 TIMEBOOST_cell_8603 ( .a(TIMEBOOST_net_2788), .b(n_16048), .o(n_16113) );
in01s01 g738560 ( .a(n_41504), .o(n_41505) );
ao12s01 g738561 ( .a(n_41423), .b(n_41422), .c(n_41421), .o(n_41504) );
no02s06 g738564 ( .a(n_41604), .b(n_41725), .o(n_41761) );
no02s06 g738565 ( .a(n_41607), .b(n_41724), .o(n_41762) );
no02s06 g738566 ( .a(n_41685), .b(n_41722), .o(n_41723) );
in01s01 g738567 ( .a(n_41618), .o(n_41619) );
no02m04 g738568 ( .a(n_41534), .b(n_41879), .o(n_41618) );
no02s06 g738569 ( .a(n_41571), .b(n_41533), .o(n_41572) );
na02s01 g738570 ( .a(n_41616), .b(n_41557), .o(n_41617) );
no02f04 TIMEBOOST_cell_6740 ( .a(TIMEBOOST_net_2127), .b(n_14628), .o(n_14709) );
no02m06 g738576 ( .a(n_41614), .b(n_41613), .o(n_41615) );
no02s01 g738577 ( .a(n_41688), .b(n_41722), .o(n_42023) );
na02s01 g738578 ( .a(n_41877), .b(n_41901), .o(n_41986) );
no02s06 g738579 ( .a(n_41560), .b(n_41481), .o(n_41612) );
na02s01 g738580 ( .a(n_41721), .b(n_41608), .o(n_42014) );
no02s01 g738581 ( .a(n_41827), .b(n_41879), .o(n_41918) );
na02s01 g738582 ( .a(n_41536), .b(n_41663), .o(n_41925) );
no02s01 g738583 ( .a(n_41807), .b(n_41457), .o(n_41864) );
no02s01 g738584 ( .a(n_41487), .b(n_41458), .o(n_41890) );
na02m08 g738585 ( .a(n_41536), .b(n_41187), .o(n_41566) );
na02s01 g738586 ( .a(n_41461), .b(n_41419), .o(n_41736) );
no02s01 g738587 ( .a(n_41760), .b(n_41418), .o(n_41817) );
na02s01 g738588 ( .a(n_41400), .b(n_41449), .o(n_41520) );
no02s01 g738589 ( .a(n_41876), .b(n_41532), .o(n_42083) );
no02s01 g738590 ( .a(n_41560), .b(n_41687), .o(n_42141) );
na02s01 g738591 ( .a(n_41561), .b(n_41662), .o(n_42032) );
no02s01 TIMEBOOST_cell_4497 ( .a(FE_OCP_RBN1034_n_25844), .b(n_27170), .o(TIMEBOOST_net_1339) );
na02s01 g738593 ( .a(n_41804), .b(n_41850), .o(n_41957) );
na02f04 g738594 ( .a(n_41445), .b(n_41444), .o(n_41446) );
na02s02 TIMEBOOST_cell_7563 ( .a(TIMEBOOST_net_2412), .b(n_25199), .o(FE_RN_702_0) );
na02m02 g738596 ( .a(n_41499), .b(n_41462), .o(n_41500) );
na02m04 TIMEBOOST_cell_4068 ( .a(TIMEBOOST_net_1124), .b(n_11004), .o(TIMEBOOST_net_920) );
no02s06 g738598 ( .a(n_41365), .b(n_40930), .o(n_41388) );
no02f02 g738599 ( .a(n_41364), .b(n_40929), .o(n_41379) );
no02s01 g738600 ( .a(n_41422), .b(n_41421), .o(n_41423) );
na02s01 g738601 ( .a(n_41443), .b(n_41398), .o(n_41508) );
ao12s01 g738602 ( .a(n_41725), .b(n_41716), .c(n_41656), .o(n_42020) );
oa12s01 g738603 ( .a(n_41686), .b(n_41713), .c(n_41326), .o(n_42061) );
ao12s01 g738604 ( .a(n_41724), .b(n_41716), .c(n_41339), .o(n_42056) );
in01s02 g738605 ( .a(n_41782), .o(n_41783) );
na02s02 g738606 ( .a(n_41759), .b(n_41717), .o(n_41782) );
oa12s01 g738607 ( .a(n_41535), .b(n_41713), .c(n_41526), .o(n_41943) );
ao12s01 g738608 ( .a(n_41571), .b(n_41716), .c(n_41492), .o(n_41965) );
ao12s01 g738609 ( .a(n_41489), .b(n_41716), .c(n_41140), .o(n_41927) );
ao12s01 g738610 ( .a(n_41486), .b(n_41716), .c(n_41062), .o(n_41835) );
oa12s01 g738611 ( .a(n_41616), .b(n_41713), .c(n_41263), .o(n_42132) );
oa12s01 g738612 ( .a(n_41528), .b(n_41713), .c(n_41286), .o(n_42162) );
ao12s01 g738613 ( .a(n_41828), .b(n_41716), .c(n_41484), .o(n_42008) );
ao12s01 g738614 ( .a(n_41912), .b(n_41716), .c(n_41613), .o(n_42078) );
na03m08 TIMEBOOST_cell_8251 ( .a(n_2419), .b(FE_OCP_RBN4071_n_2289), .c(n_2394), .o(n_2453) );
oa22s01 g738616 ( .a(n_41716), .b(n_41124), .c(n_41713), .d(n_41501), .o(n_41893) );
oa22s01 g738617 ( .a(n_41716), .b(n_41050), .c(n_41713), .d(n_41444), .o(n_41832) );
in01s01 g738618 ( .a(n_41405), .o(n_41507) );
no02s02 TIMEBOOST_cell_6062 ( .a(TIMEBOOST_net_1882), .b(TIMEBOOST_net_1496), .o(n_30703) );
in01s01 g738638 ( .a(n_41540), .o(n_41660) );
in01m03 g738642 ( .a(FE_OCP_RBN5676_n_41420), .o(n_41540) );
in01s06 g738647 ( .a(FE_OCP_RBN5673_n_41420), .o(n_41582) );
in01m40 g738662 ( .a(FE_OCP_RBN5638_n_41381), .o(n_41420) );
ao12f08 g738666 ( .a(n_41360), .b(n_41367), .c(n_41372), .o(n_41381) );
in01s01 g738667 ( .a(n_41779), .o(n_41780) );
na02s02 g738668 ( .a(n_41684), .b(n_41715), .o(n_41779) );
in01s01 g738670 ( .a(n_41608), .o(n_41658) );
na02s02 g738671 ( .a(n_41525), .b(FE_OFN4755_n_41563), .o(n_41608) );
in01s01 g738672 ( .a(n_41688), .o(n_41657) );
no02s02 g738673 ( .a(n_41478), .b(n_41296), .o(n_41688) );
in01s01 g738674 ( .a(n_41607), .o(n_41721) );
no02s04 g738675 ( .a(FE_OCP_RBN6592_n_41491), .b(n_41563), .o(n_41607) );
no02s03 g738676 ( .a(n_41525), .b(n_41339), .o(n_41724) );
no02s06 g738677 ( .a(n_41525), .b(n_41656), .o(n_41725) );
na02s01 g738678 ( .a(n_41478), .b(n_41605), .o(n_41759) );
in01s01 g738679 ( .a(n_41604), .o(n_41901) );
no02s06 g738680 ( .a(FE_OCP_RBN6592_n_41491), .b(n_41562), .o(n_41604) );
in01s01 g738681 ( .a(n_41685), .o(n_41686) );
no02s04 g738682 ( .a(n_41525), .b(n_41654), .o(n_41685) );
no02s04 g738683 ( .a(n_41525), .b(n_41297), .o(n_41722) );
in01s01 g738684 ( .a(n_41614), .o(n_41561) );
no02s06 g738685 ( .a(FE_OCP_RBN6587_n_41491), .b(n_41212), .o(n_41614) );
in01s01 g738686 ( .a(n_41877), .o(n_41878) );
na02s01 g738687 ( .a(n_41716), .b(n_41562), .o(n_41877) );
na02s02 g738688 ( .a(n_41716), .b(FE_OCP_RBN4054_n_41325), .o(n_41717) );
in01s01 g738689 ( .a(n_41826), .o(n_41827) );
na02s01 g738690 ( .a(n_41716), .b(n_41494), .o(n_41826) );
in01s01 g738692 ( .a(n_41560), .o(n_41602) );
no02s06 g738693 ( .a(FE_OCP_RBN6586_n_41491), .b(n_41255), .o(n_41560) );
no02s01 g738694 ( .a(n_41716), .b(n_41438), .o(n_41807) );
in01s01 g738696 ( .a(n_41536), .o(n_41558) );
na02m06 g738697 ( .a(n_41491), .b(n_41490), .o(n_41536) );
no02s01 g738698 ( .a(n_41716), .b(n_41401), .o(n_41760) );
in01s01 g738699 ( .a(n_41534), .o(n_41535) );
no02m01 g738700 ( .a(n_41382), .b(n_41141), .o(n_41534) );
no02f01 g738701 ( .a(n_41382), .b(n_41494), .o(n_41879) );
no02s03 g738702 ( .a(n_41483), .b(n_41492), .o(n_41571) );
in01s01 g738703 ( .a(n_41533), .o(n_41663) );
no02s04 g738704 ( .a(n_41491), .b(n_41490), .o(n_41533) );
in01s01 g738705 ( .a(n_41488), .o(n_41489) );
na02s04 g738706 ( .a(n_41456), .b(n_41462), .o(n_41488) );
in01s01 g738707 ( .a(n_41577), .o(n_41487) );
in01s01 g738709 ( .a(n_41875), .o(n_41876) );
na02s01 g738710 ( .a(n_41716), .b(n_41482), .o(n_41875) );
in01s01 g738711 ( .a(n_41803), .o(n_41804) );
no02s01 g738712 ( .a(n_41713), .b(n_41198), .o(n_41803) );
in01s01 g738714 ( .a(n_41419), .o(n_41440) );
na02f04 g738715 ( .a(n_41378), .b(n_41402), .o(n_41419) );
in01s01 g738716 ( .a(n_41445), .o(n_41418) );
na02f04 g738717 ( .a(n_41378), .b(n_41401), .o(n_41445) );
in01s01 g738718 ( .a(n_41460), .o(n_41461) );
no02f04 g738719 ( .a(n_41382), .b(n_41402), .o(n_41460) );
na02f04 g738720 ( .a(n_41386), .b(n_41385), .o(n_41449) );
in01s01 g738721 ( .a(n_41485), .o(n_41486) );
na02s06 g738722 ( .a(n_41435), .b(n_41447), .o(n_41485) );
in01s01 g738723 ( .a(n_41399), .o(n_41400) );
no02f04 g738724 ( .a(n_41386), .b(n_41385), .o(n_41399) );
in01s01 g738725 ( .a(n_41499), .o(n_41458) );
na02m02 g738726 ( .a(n_41382), .b(n_41121), .o(n_41499) );
in01s01 g738727 ( .a(n_41502), .o(n_41457) );
na02s02 g738728 ( .a(n_41382), .b(n_41438), .o(n_41502) );
no02m02 g738729 ( .a(n_41483), .b(n_41484), .o(n_41828) );
in01s01 g738731 ( .a(n_41532), .o(n_41557) );
no02s03 g738732 ( .a(n_41483), .b(n_41482), .o(n_41532) );
no02m02 g738733 ( .a(n_41483), .b(n_41613), .o(n_41912) );
in01s01 g738734 ( .a(n_41531), .o(n_41662) );
no02s02 g738735 ( .a(n_41483), .b(FE_OCPN1222_n_41211), .o(n_41531) );
in01s01 g738736 ( .a(n_41530), .o(n_41616) );
no02s02 g738737 ( .a(n_41483), .b(n_41228), .o(n_41530) );
in01s01 g738738 ( .a(n_41529), .o(n_41850) );
no02s02 g738739 ( .a(n_41483), .b(n_41142), .o(n_41529) );
in01s01 g738740 ( .a(n_41527), .o(n_41528) );
no02s02 g738741 ( .a(n_41483), .b(n_41481), .o(n_41527) );
no02s02 g738742 ( .a(n_41483), .b(n_41254), .o(n_41687) );
na02s01 g738743 ( .a(FE_OCP_RBN6592_n_41491), .b(n_41366), .o(n_41715) );
na02s01 g738744 ( .a(FE_OCP_RBN6595_n_41491), .b(n_41372), .o(n_41684) );
no02m02 g738745 ( .a(n_41372), .b(n_41355), .o(n_41361) );
no02s06 TIMEBOOST_cell_7409 ( .a(n_37160), .b(TIMEBOOST_net_2335), .o(n_37219) );
na02s01 g738747 ( .a(n_41375), .b(n_41371), .o(n_41422) );
na02f04 g738748 ( .a(n_41384), .b(n_41383), .o(n_41443) );
na02s01 TIMEBOOST_cell_4493 ( .a(n_5895), .b(n_5621), .o(TIMEBOOST_net_1337) );
in01s01 g738750 ( .a(n_41397), .o(n_41398) );
no02f04 g738751 ( .a(n_41384), .b(n_41383), .o(n_41397) );
no02s02 g738752 ( .a(n_41478), .b(n_41328), .o(n_41788) );
in01s01 g738753 ( .a(n_41729), .o(n_41600) );
na02s06 g738754 ( .a(FE_OCP_RBN6591_n_41491), .b(n_41199), .o(n_41729) );
in01s01 g738755 ( .a(n_41598), .o(n_41599) );
na02s03 g738756 ( .a(n_41525), .b(n_41264), .o(n_41598) );
ao12s03 g738757 ( .a(n_41478), .b(n_41526), .c(n_41123), .o(n_41692) );
in01s01 g738758 ( .a(n_41479), .o(n_41480) );
na02s04 g738759 ( .a(n_41456), .b(n_41125), .o(n_41479) );
no02f04 g738760 ( .a(n_41382), .b(n_41063), .o(n_41683) );
in01s02 g738761 ( .a(n_41364), .o(n_41365) );
no02m08 g738763 ( .a(n_41372), .b(n_41337), .o(n_41360) );
in01s01 g738764 ( .a(n_41374), .o(n_41375) );
no02f06 g738765 ( .a(n_41358), .b(n_40864), .o(n_41374) );
in01s01 g738766 ( .a(n_41370), .o(n_41371) );
no02f04 g738767 ( .a(n_41357), .b(FE_OCPN1220_n_40863), .o(n_41370) );
in01f06 g738768 ( .a(n_41355), .o(n_41367) );
no02m06 TIMEBOOST_cell_1916 ( .a(TIMEBOOST_net_572), .b(n_11410), .o(n_11480) );
in01s01 g738770 ( .a(n_41369), .o(n_42181) );
ao22s01 g738771 ( .a(n_41339), .b(n_41343), .c(n_41324), .d(n_40658), .o(n_41369) );
na02f04 g738772 ( .a(n_41362), .b(n_41359), .o(n_41384) );
in01f02 g738773 ( .a(n_41386), .o(n_41378) );
in01m08 g738775 ( .a(n_41435), .o(n_41483) );
in01m06 g738778 ( .a(n_41382), .o(n_41435) );
in01s01 g738792 ( .a(n_41716), .o(n_41713) );
in01s06 g738793 ( .a(FE_OCP_RBN6594_n_41491), .o(n_41716) );
in01m08 g738800 ( .a(n_41456), .o(n_41491) );
in01s06 g738803 ( .a(n_41478), .o(n_41525) );
in01s03 g738809 ( .a(n_41382), .o(n_41478) );
in01m04 g738811 ( .a(n_41382), .o(n_41456) );
in01f08 g738817 ( .a(n_41386), .o(n_41382) );
oa12f08 g738818 ( .a(n_41333), .b(n_41356), .c(FE_OCP_RBN4044_n_41298), .o(n_41386) );
no03m08 TIMEBOOST_cell_8726 ( .a(FE_OCP_RBN2479_n_47245), .b(TIMEBOOST_net_1418), .c(n_23166), .o(TIMEBOOST_net_2850) );
in01f01 g738820 ( .a(n_41353), .o(n_41344) );
na02f06 g738821 ( .a(n_41312), .b(delay_sub_ln23_0_unr28_stage10_stallmux_q), .o(n_41353) );
no02s02 g738822 ( .a(n_41324), .b(n_41343), .o(n_41430) );
oa12f02 g738824 ( .a(n_41298), .b(n_41349), .c(n_44429), .o(n_41359) );
in01f02 g738825 ( .a(n_41357), .o(n_41358) );
na02f04 g738826 ( .a(n_41342), .b(n_41341), .o(n_41357) );
in01s02 g738827 ( .a(n_41372), .o(n_41366) );
no02m10 g738828 ( .a(n_41327), .b(n_41314), .o(n_41372) );
na02f03 g738829 ( .a(n_44430), .b(n_41302), .o(n_41342) );
na02f02 g738830 ( .a(n_41311), .b(n_41301), .o(n_41341) );
no02s01 g738831 ( .a(n_41656), .b(n_41562), .o(n_41328) );
na02s01 TIMEBOOST_cell_4903 ( .a(TIMEBOOST_net_1399), .b(n_1787), .o(TIMEBOOST_net_249) );
na02f08 g738834 ( .a(n_44428), .b(n_41348), .o(n_41356) );
in01s01 g738835 ( .a(n_41654), .o(n_41326) );
oa12s02 g738836 ( .a(n_41289), .b(n_41288), .c(n_41287), .o(n_41654) );
in01s01 g738838 ( .a(FE_OCP_RBN4054_n_41325), .o(n_41605) );
in01m02 g738840 ( .a(n_41313), .o(n_41325) );
oa22f06 g738841 ( .a(n_41258), .b(n_40953), .c(FE_OCP_RBN4043_n_41258), .d(n_40952), .o(n_41313) );
ao22s01 g738842 ( .a(n_41300), .b(n_41309), .c(n_41310), .d(n_40657), .o(n_42204) );
in01s01 g738846 ( .a(n_41324), .o(n_41339) );
in01s01 g738847 ( .a(n_41312), .o(n_41324) );
na02s02 g738849 ( .a(n_41288), .b(n_41287), .o(n_41289) );
in01f06 g738851 ( .a(n_41349), .o(n_41348) );
no02f08 g738852 ( .a(n_41319), .b(n_41337), .o(n_41349) );
no02f06 g738857 ( .a(n_41285), .b(n_41337), .o(n_41311) );
na02f08 g738858 ( .a(FE_OCP_RBN4044_n_41298), .b(delay_sub_ln23_0_unr28_stage10_stallmux_q), .o(n_41333) );
na02s01 g738859 ( .a(n_41263), .b(n_41217), .o(n_41264) );
in01s01 g738860 ( .a(n_41322), .o(n_41421) );
na02s04 g738861 ( .a(n_41310), .b(n_41309), .o(n_41322) );
no02s01 g738862 ( .a(n_41299), .b(n_41320), .o(n_41321) );
oa22s01 g738863 ( .a(n_41253), .b(n_40906), .c(n_41252), .d(n_40907), .o(n_41563) );
oa12s02 g738864 ( .a(n_41274), .b(n_41273), .c(n_41272), .o(n_41656) );
in01s01 g738865 ( .a(n_41296), .o(n_41297) );
ao12s01 g738866 ( .a(n_41262), .b(n_41261), .c(n_41260), .o(n_41296) );
in01s01 g738867 ( .a(n_41481), .o(n_41286) );
oa12s02 g738868 ( .a(n_41232), .b(n_41231), .c(n_41230), .o(n_41481) );
na02s02 TIMEBOOST_cell_1840 ( .a(TIMEBOOST_net_534), .b(n_16912), .o(n_17007) );
in01s01 g738870 ( .a(n_41347), .o(n_41637) );
oa12s01 g738871 ( .a(n_41308), .b(n_41307), .c(n_41306), .o(n_41347) );
ao12s01 g738872 ( .a(n_41305), .b(n_41304), .c(n_41303), .o(n_41634) );
na02s01 g738873 ( .a(n_41273), .b(n_41272), .o(n_41274) );
no02s01 g738874 ( .a(n_41261), .b(n_41260), .o(n_41262) );
na02s01 g738875 ( .a(n_41231), .b(n_41230), .o(n_41232) );
na02s01 g738876 ( .a(n_41307), .b(n_41306), .o(n_41308) );
no02s01 g738877 ( .a(n_41304), .b(n_41303), .o(n_41305) );
ao12s01 g738879 ( .a(n_41015), .b(n_41196), .c(n_40886), .o(n_41288) );
oa12f08 g738881 ( .a(n_41047), .b(n_41194), .c(n_41229), .o(n_41258) );
in01m02 g738882 ( .a(n_41256), .o(n_41257) );
na03s08 TIMEBOOST_cell_7249 ( .a(FE_RN_1276_0), .b(FE_OCP_RBN6802_n_15156), .c(TIMEBOOST_net_2267), .o(TIMEBOOST_net_864) );
oa12s02 g738884 ( .a(n_41250), .b(n_41249), .c(n_41248), .o(n_41562) );
in01s01 g738885 ( .a(n_41263), .o(n_41228) );
ao22s01 g738886 ( .a(n_41163), .b(n_41079), .c(n_41164), .d(n_41080), .o(n_41263) );
in01s01 g738888 ( .a(n_41330), .o(n_41345) );
in01s01 g738890 ( .a(n_41319), .o(n_41330) );
in01f04 g738891 ( .a(n_41302), .o(n_41319) );
in01f01 g738892 ( .a(n_41302), .o(n_41301) );
in01s01 g738894 ( .a(n_41254), .o(n_41255) );
oa12s01 g738895 ( .a(n_41203), .b(n_41202), .c(n_41201), .o(n_41254) );
in01s01 g738898 ( .a(n_41310), .o(n_41300) );
in01m01 g738899 ( .a(n_41285), .o(n_41310) );
in01s01 g738901 ( .a(n_41299), .o(n_41590) );
oa12s01 g738902 ( .a(n_41271), .b(n_41270), .c(n_41269), .o(n_41299) );
oa12s01 g738903 ( .a(n_41284), .b(n_41283), .c(n_41282), .o(n_41543) );
ao12s01 g738904 ( .a(n_41281), .b(n_41280), .c(n_41279), .o(n_41698) );
in01s01 g738905 ( .a(n_41316), .o(n_41317) );
ao12s01 g738906 ( .a(n_41278), .b(n_41277), .c(n_41276), .o(n_41316) );
ao12s01 g738907 ( .a(n_41268), .b(n_41267), .c(n_41266), .o(n_41695) );
no02f08 g738911 ( .a(n_41265), .b(n_41251), .o(n_41298) );
in01s01 g738912 ( .a(n_41252), .o(n_41253) );
no02s01 g738913 ( .a(n_41215), .b(n_41048), .o(n_41252) );
na02s01 g738914 ( .a(n_41195), .b(n_41014), .o(n_41261) );
no02m06 g738915 ( .a(n_41223), .b(n_40983), .o(n_41251) );
na02s01 g738916 ( .a(n_41202), .b(n_41201), .o(n_41203) );
na02s01 g738917 ( .a(n_41270), .b(n_41269), .o(n_41271) );
na02s01 g738918 ( .a(n_41283), .b(n_41282), .o(n_41284) );
no02s01 g738919 ( .a(n_41280), .b(n_41279), .o(n_41281) );
no02s01 g738920 ( .a(n_41267), .b(n_41266), .o(n_41268) );
no02f08 g738921 ( .a(n_41224), .b(n_40984), .o(n_41265) );
no02s01 g738922 ( .a(n_41277), .b(n_41276), .o(n_41278) );
no02s02 TIMEBOOST_cell_8481 ( .a(TIMEBOOST_net_2727), .b(TIMEBOOST_net_2346), .o(n_6914) );
na02s01 g738924 ( .a(n_41249), .b(n_41248), .o(n_41250) );
na02s01 g738925 ( .a(n_41190), .b(n_41198), .o(n_41199) );
no02s02 TIMEBOOST_cell_7100 ( .a(TIMEBOOST_net_2308), .b(n_27223), .o(n_27353) );
no02s01 g738927 ( .a(n_41247), .b(n_41027), .o(n_41307) );
ao12s01 g738928 ( .a(n_40961), .b(n_41221), .c(n_40841), .o(n_41304) );
oa12s01 g738930 ( .a(n_41245), .b(n_41244), .c(n_41243), .o(n_41628) );
oa12s02 g738931 ( .a(n_41170), .b(n_41169), .c(n_41168), .o(n_41613) );
in01s01 g738932 ( .a(n_41217), .o(n_41482) );
ao12s01 g738933 ( .a(n_41167), .b(n_41166), .c(n_41165), .o(n_41217) );
in01s01 g738934 ( .a(n_41320), .o(n_41292) );
oa12s01 g738935 ( .a(n_41242), .b(n_41241), .c(n_41240), .o(n_41320) );
in01s01 g738936 ( .a(n_41290), .o(n_41291) );
oa12s01 g738937 ( .a(n_41239), .b(n_41238), .c(n_41237), .o(n_41290) );
in01s01 g738938 ( .a(n_41631), .o(n_41275) );
ao12s01 g738939 ( .a(n_41227), .b(n_41226), .c(n_41225), .o(n_41631) );
oa12s01 g738940 ( .a(n_41236), .b(n_41235), .c(n_41234), .o(n_41626) );
no02f06 TIMEBOOST_cell_1810 ( .a(TIMEBOOST_net_519), .b(n_15702), .o(n_15799) );
na02s01 g738942 ( .a(n_41171), .b(n_40943), .o(n_41202) );
no02s02 TIMEBOOST_cell_1820 ( .a(TIMEBOOST_net_524), .b(n_10401), .o(n_10506) );
no02s01 g738944 ( .a(n_41246), .b(n_40850), .o(n_41247) );
na02s01 g738945 ( .a(n_41246), .b(n_41026), .o(n_41283) );
no02s01 g738946 ( .a(n_41159), .b(n_40962), .o(n_41249) );
in01s01 g738947 ( .a(n_41195), .o(n_41196) );
na02s02 g738948 ( .a(n_41159), .b(n_40911), .o(n_41195) );
na02s01 g738949 ( .a(n_41244), .b(n_41243), .o(n_41245) );
na02s01 g738950 ( .a(n_41169), .b(n_41168), .o(n_41170) );
no02s01 g738951 ( .a(n_41166), .b(n_41165), .o(n_41167) );
na02s01 g738952 ( .a(n_41241), .b(n_41240), .o(n_41242) );
no02s01 g738953 ( .a(n_41226), .b(n_41225), .o(n_41227) );
na02s01 g738954 ( .a(n_41220), .b(n_40960), .o(n_41277) );
na02s01 g738955 ( .a(n_41238), .b(n_41237), .o(n_41239) );
na02s01 g738956 ( .a(n_41235), .b(n_41234), .o(n_41236) );
in01f04 g738957 ( .a(n_41223), .o(n_41224) );
oa12f08 g738958 ( .a(n_41061), .b(n_41186), .c(n_40935), .o(n_41223) );
ao12f02 g738959 ( .a(n_41060), .b(n_41155), .c(n_41208), .o(n_41222) );
no02s01 TIMEBOOST_cell_6979 ( .a(FE_OFN742_delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n_21975), .o(TIMEBOOST_net_2248) );
in01s06 g738962 ( .a(n_41194), .o(n_41215) );
in01f06 g738963 ( .a(n_41191), .o(n_41194) );
no02f08 g738964 ( .a(n_41154), .b(n_40912), .o(n_41191) );
ao12f06 g738966 ( .a(n_40996), .b(n_41155), .c(n_40872), .o(n_41213) );
ao12s01 g738967 ( .a(n_40978), .b(n_41207), .c(n_40718), .o(n_41270) );
in01s01 g738968 ( .a(n_41211), .o(n_41212) );
oa12s01 g738969 ( .a(n_41162), .b(n_41161), .c(n_41160), .o(n_41211) );
in01s01 g738970 ( .a(n_41190), .o(n_41484) );
ao12s01 g738971 ( .a(n_41148), .b(n_41147), .c(n_41146), .o(n_41190) );
in01s01 g738972 ( .a(n_41163), .o(n_41164) );
ao12s01 g738973 ( .a(n_41012), .b(n_41149), .c(n_40758), .o(n_41163) );
no02s01 TIMEBOOST_cell_1757 ( .a(n_5299), .b(n_5331), .o(TIMEBOOST_net_493) );
ao12s01 g738975 ( .a(n_40768), .b(n_41204), .c(n_40858), .o(n_41267) );
no02s01 g738976 ( .a(n_41155), .b(n_40993), .o(n_41244) );
no02s01 g738977 ( .a(n_41149), .b(n_40914), .o(n_41166) );
na02s01 g738978 ( .a(n_41149), .b(n_40827), .o(n_41171) );
no02s01 TIMEBOOST_cell_8796 ( .a(FE_OCP_RBN2759_n_13796), .b(FE_OCP_RBN4200_n_13796), .o(TIMEBOOST_net_2885) );
no02s01 g738980 ( .a(n_41207), .b(n_40989), .o(n_41241) );
na02s01 g738981 ( .a(n_41207), .b(n_40934), .o(n_41246) );
no02s01 g738982 ( .a(n_41185), .b(n_40813), .o(n_41193) );
no02s01 g738983 ( .a(n_41205), .b(n_41206), .o(n_41238) );
in01s01 g738984 ( .a(n_41220), .o(n_41221) );
na02s01 g738985 ( .a(n_41205), .b(n_40856), .o(n_41220) );
no02s01 g738986 ( .a(n_41204), .b(n_40867), .o(n_41235) );
no02s01 g738987 ( .a(n_41147), .b(n_41146), .o(n_41148) );
na02s01 g738988 ( .a(n_41161), .b(n_41160), .o(n_41162) );
oa12s01 g738989 ( .a(n_41077), .b(n_41192), .c(n_41107), .o(n_41226) );
in01s01 g738992 ( .a(n_41154), .o(n_41159) );
na02f08 g738993 ( .a(n_41149), .b(n_40910), .o(n_41154) );
ao12s01 g738994 ( .a(n_40791), .b(n_41114), .c(n_40829), .o(n_41169) );
in01s01 g738995 ( .a(n_41492), .o(n_41187) );
oa12s02 g738996 ( .a(n_41145), .b(n_41144), .c(n_41143), .o(n_41492) );
in01s01 g738997 ( .a(n_41576), .o(n_41219) );
ao12s01 g738998 ( .a(n_41184), .b(n_41192), .c(n_41183), .o(n_41576) );
in01s01 g738999 ( .a(n_41186), .o(n_41207) );
na02f08 g739000 ( .a(n_41158), .b(n_40936), .o(n_41186) );
na02s01 g739001 ( .a(n_41144), .b(n_41143), .o(n_41145) );
in01s01 g739002 ( .a(n_41185), .o(n_41205) );
na02s01 g739003 ( .a(n_41158), .b(n_40884), .o(n_41185) );
no02s01 g739004 ( .a(n_41192), .b(n_40775), .o(n_41204) );
na02s01 g739005 ( .a(n_41098), .b(n_40869), .o(n_41161) );
no02s01 g739006 ( .a(n_41192), .b(n_41183), .o(n_41184) );
no02s01 g739007 ( .a(n_41156), .b(n_41126), .o(n_41157) );
no02f08 g739011 ( .a(n_41133), .b(n_46947), .o(n_41155) );
na02s01 g739012 ( .a(n_41124), .b(n_41438), .o(n_41125) );
no02f08 g739013 ( .a(n_41098), .b(n_40830), .o(n_41149) );
oa12s01 g739014 ( .a(n_41053), .b(n_41119), .c(n_41038), .o(n_41147) );
in01s01 g739015 ( .a(n_41198), .o(n_41142) );
ao22s01 g739016 ( .a(n_41119), .b(n_41071), .c(n_41085), .d(n_41070), .o(n_41198) );
in01s01 g739017 ( .a(n_41141), .o(n_41526) );
oa12s01 g739018 ( .a(n_41104), .b(n_41103), .c(n_41102), .o(n_41141) );
oa12s02 g739019 ( .a(n_41118), .b(n_41117), .c(n_41116), .o(n_41490) );
in01s01 g739020 ( .a(n_41462), .o(n_41140) );
ao12s01 g739021 ( .a(n_41101), .b(n_41100), .c(n_41099), .o(n_41462) );
in01s01 g739022 ( .a(n_41218), .o(n_41629) );
oa12s01 g739023 ( .a(n_41179), .b(n_41178), .c(n_41177), .o(n_41218) );
in01s01 g739024 ( .a(n_41545), .o(n_41180) );
ao12s02 g739025 ( .a(n_41139), .b(n_41138), .c(n_41137), .o(n_41545) );
ao12s01 g739026 ( .a(n_41136), .b(n_41135), .c(n_41134), .o(n_41473) );
na02s01 g739027 ( .a(n_41103), .b(n_41102), .o(n_41104) );
na02s01 g739028 ( .a(n_41117), .b(n_41116), .o(n_41118) );
no02s01 g739029 ( .a(n_41100), .b(n_41099), .o(n_41101) );
na02s01 g739030 ( .a(n_41178), .b(n_41177), .o(n_41179) );
no02s01 g739031 ( .a(n_41138), .b(n_41137), .o(n_41139) );
no02s01 g739032 ( .a(n_41135), .b(n_41134), .o(n_41136) );
in01s01 g739034 ( .a(n_41098), .o(n_41114) );
na02f08 g739035 ( .a(n_41073), .b(n_40757), .o(n_41098) );
no02s01 g739036 ( .a(n_41093), .b(n_41042), .o(n_41144) );
in01s01 g739037 ( .a(n_41158), .o(n_41192) );
in01f04 g739038 ( .a(n_41133), .o(n_41158) );
ao12f08 g739039 ( .a(n_40956), .b(n_41110), .c(FE_OCP_DRV_N3494_n_40837), .o(n_41133) );
in01s01 g739040 ( .a(n_41156), .o(n_41153) );
oa12s01 g739041 ( .a(n_41113), .b(n_41112), .c(n_41111), .o(n_41156) );
in01s01 g739042 ( .a(n_41494), .o(n_41123) );
oa12s01 g739043 ( .a(n_41091), .b(n_41090), .c(n_41089), .o(n_41494) );
in01s01 g739044 ( .a(n_41124), .o(n_41501) );
oa12s01 g739045 ( .a(n_41076), .b(n_41075), .c(n_41074), .o(n_41124) );
oa12s01 g739047 ( .a(n_41088), .b(n_41087), .c(n_41086), .o(n_41121) );
oa12s01 g739048 ( .a(n_41152), .b(n_41151), .c(n_41150), .o(n_41542) );
in01s01 g739049 ( .a(n_41175), .o(n_41176) );
oa12s01 g739050 ( .a(n_41132), .b(n_41131), .c(n_41130), .o(n_41175) );
in01s01 g739051 ( .a(n_41173), .o(n_41174) );
ao12s01 g739052 ( .a(n_41129), .b(n_41128), .c(n_41127), .o(n_41173) );
na02s01 g739053 ( .a(n_41092), .b(n_41041), .o(n_41117) );
no02s01 g739054 ( .a(n_41092), .b(n_40704), .o(n_41093) );
na02s01 g739055 ( .a(n_41112), .b(n_41111), .o(n_41113) );
na02s01 g739056 ( .a(n_41090), .b(n_41089), .o(n_41091) );
na02s01 g739057 ( .a(n_41075), .b(n_41074), .o(n_41076) );
na02s01 g739058 ( .a(n_41131), .b(n_41130), .o(n_41132) );
na02s01 g739059 ( .a(n_41087), .b(n_41086), .o(n_41088) );
na02s01 g739060 ( .a(n_41151), .b(n_41150), .o(n_41152) );
no02s01 g739061 ( .a(n_40959), .b(n_41110), .o(n_41138) );
no02s01 g739062 ( .a(n_41128), .b(n_41127), .o(n_41129) );
in01s01 g739063 ( .a(n_41119), .o(n_41085) );
in01s01 g739064 ( .a(n_41073), .o(n_41119) );
oa12f08 g739065 ( .a(n_40926), .b(n_41031), .c(n_40797), .o(n_41073) );
ao12s01 g739066 ( .a(n_41011), .b(n_41065), .c(n_40730), .o(n_41103) );
ao12s01 g739067 ( .a(n_40851), .b(n_41081), .c(n_40810), .o(n_41135) );
ao12s01 g739068 ( .a(n_40708), .b(n_41064), .c(n_40698), .o(n_41100) );
no02s06 TIMEBOOST_cell_1725 ( .a(n_25750), .b(n_25669), .o(TIMEBOOST_net_477) );
no02s01 g739070 ( .a(n_41065), .b(n_40868), .o(n_41090) );
na02s01 g739071 ( .a(n_41065), .b(n_40796), .o(n_41092) );
no02s01 g739072 ( .a(n_41096), .b(n_40811), .o(n_41109) );
no02s01 g739073 ( .a(n_41097), .b(n_41120), .o(n_41151) );
no02s01 g739074 ( .a(n_41064), .b(n_40834), .o(n_41087) );
na02s01 g739075 ( .a(n_41082), .b(n_40893), .o(n_41128) );
oa12s01 g739077 ( .a(n_40958), .b(n_41108), .c(n_41084), .o(n_41131) );
oa12s01 g739078 ( .a(n_41022), .b(n_41083), .c(n_41052), .o(n_41112) );
oa12s01 g739079 ( .a(n_40971), .b(n_41051), .c(n_40988), .o(n_41075) );
no02s02 g739080 ( .a(n_41444), .b(n_41028), .o(n_41063) );
in01s01 g739081 ( .a(n_41126), .o(n_41415) );
oa12s01 g739082 ( .a(n_41095), .b(n_41108), .c(n_41094), .o(n_41126) );
oa12s01 g739083 ( .a(n_41033), .b(n_41051), .c(n_41032), .o(n_41438) );
in01s01 g739084 ( .a(n_41096), .o(n_41097) );
na02s01 g739085 ( .a(n_41072), .b(n_40866), .o(n_41096) );
no02s01 g739086 ( .a(n_41051), .b(n_40749), .o(n_41064) );
in01s01 g739087 ( .a(n_41081), .o(n_41082) );
no02s01 g739088 ( .a(n_41083), .b(n_40826), .o(n_41081) );
na02s01 g739089 ( .a(n_41108), .b(n_41094), .o(n_41095) );
na02s01 g739090 ( .a(n_41051), .b(n_41032), .o(n_41033) );
in01s01 g739091 ( .a(n_41031), .o(n_41065) );
na02f08 g739092 ( .a(n_40997), .b(n_40751), .o(n_41031) );
ao12s02 g739093 ( .a(n_41059), .b(n_41058), .c(n_41057), .o(n_41433) );
in01s01 g739094 ( .a(n_41447), .o(n_41062) );
ao12s02 g739095 ( .a(n_41018), .b(n_41017), .c(n_41016), .o(n_41447) );
oa12s01 g739096 ( .a(n_41003), .b(n_41002), .c(n_41001), .o(n_41402) );
in01s01 g739097 ( .a(n_41444), .o(n_41050) );
ao12s02 g739098 ( .a(n_41000), .b(n_40999), .c(n_40998), .o(n_41444) );
no02s04 g739099 ( .a(n_41060), .b(n_40918), .o(n_41061) );
no02m04 g739100 ( .a(n_41048), .b(n_40845), .o(n_41049) );
no02s01 g739101 ( .a(n_41058), .b(n_41057), .o(n_41059) );
no02s03 g739102 ( .a(n_41048), .b(n_40939), .o(n_41047) );
no02s01 g739103 ( .a(n_41017), .b(n_41016), .o(n_41018) );
na02s01 g739104 ( .a(n_41002), .b(n_41001), .o(n_41003) );
no02s01 g739105 ( .a(n_40999), .b(n_40998), .o(n_41000) );
na02s06 g739106 ( .a(n_41029), .b(n_40940), .o(n_41293) );
oa12s01 g739107 ( .a(n_41056), .b(n_41055), .c(n_41054), .o(n_41392) );
ao12s01 g739108 ( .a(n_41045), .b(n_41044), .c(n_41043), .o(n_41407) );
in01s01 g739109 ( .a(n_40997), .o(n_41051) );
no03s02 TIMEBOOST_cell_4898 ( .a(n_6594), .b(n_6775), .c(n_6595), .o(TIMEBOOST_net_1397) );
in01s01 g739111 ( .a(n_41072), .o(n_41108) );
in01s01 g739112 ( .a(n_41083), .o(n_41072) );
ao12f08 g739113 ( .a(n_40782), .b(n_41030), .c(n_40803), .o(n_41083) );
no02s01 g739114 ( .a(n_41030), .b(n_40780), .o(n_41058) );
na02s01 g739115 ( .a(n_41014), .b(n_40887), .o(n_41015) );
no02s01 g739116 ( .a(n_40945), .b(n_40789), .o(n_41017) );
na02m04 g739117 ( .a(n_40979), .b(n_40805), .o(n_40996) );
in01s01 g739118 ( .a(n_41048), .o(n_41029) );
na02m08 g739119 ( .a(n_41014), .b(n_40865), .o(n_41048) );
na02s01 g739121 ( .a(n_41055), .b(n_41054), .o(n_41056) );
in01m04 g739122 ( .a(n_41060), .o(n_41046) );
na02m08 g739123 ( .a(n_40979), .b(n_40905), .o(n_41060) );
no02s01 g739124 ( .a(n_41044), .b(n_41043), .o(n_41045) );
oa12s01 g739125 ( .a(n_40787), .b(n_40964), .c(n_40919), .o(n_41002) );
oa12s01 g739126 ( .a(n_40933), .b(n_40964), .c(n_40902), .o(n_40999) );
in01s01 g739127 ( .a(n_41028), .o(n_41401) );
ao22s01 g739128 ( .a(n_40964), .b(n_40955), .c(n_40925), .d(n_40954), .o(n_41028) );
na02s01 g739129 ( .a(n_41026), .b(n_40823), .o(n_41027) );
na02s01 g739130 ( .a(n_40976), .b(n_40831), .o(n_40995) );
no02m08 g739131 ( .a(n_40962), .b(n_40832), .o(n_41014) );
na02s01 g739132 ( .a(n_40991), .b(n_41006), .o(n_41055) );
in01s01 g739134 ( .a(n_40979), .o(n_40993) );
no02s01 g739137 ( .a(n_40964), .b(n_40744), .o(n_40945) );
oa12s01 g739138 ( .a(n_41013), .b(n_40992), .c(n_40981), .o(n_41044) );
ao22s01 g739139 ( .a(n_40990), .b(n_41036), .c(n_40975), .d(n_41037), .o(n_41406) );
na02s01 g739140 ( .a(n_40943), .b(n_40885), .o(n_40944) );
na02s01 g739141 ( .a(n_41041), .b(n_41040), .o(n_41042) );
na02s01 g739142 ( .a(n_40957), .b(n_40822), .o(n_40978) );
in01s01 g739144 ( .a(n_40962), .o(n_40976) );
na02m08 g739145 ( .a(n_40943), .b(n_40794), .o(n_40962) );
na02s02 TIMEBOOST_cell_7394 ( .a(n_17158), .b(n_17015), .o(TIMEBOOST_net_2328) );
na02s01 g739147 ( .a(n_40990), .b(n_40712), .o(n_40991) );
no02s01 g739148 ( .a(n_40989), .b(n_40963), .o(n_41026) );
in01s01 g739149 ( .a(n_40964), .o(n_40925) );
in01s01 g739150 ( .a(n_40915), .o(n_40964) );
ao12f06 g739151 ( .a(n_40693), .b(n_40897), .c(n_40742), .o(n_40915) );
ao22s01 g739152 ( .a(n_40897), .b(n_40784), .c(n_40833), .d(n_40783), .o(n_41385) );
na02s01 g739153 ( .a(n_40960), .b(n_40882), .o(n_40961) );
na02s01 g739154 ( .a(n_40958), .b(n_40873), .o(n_40959) );
na02s01 g739155 ( .a(n_40895), .b(n_41009), .o(n_41012) );
na02s01 g739156 ( .a(n_40896), .b(n_41007), .o(n_41011) );
no02s06 TIMEBOOST_cell_1794 ( .a(TIMEBOOST_net_511), .b(n_10800), .o(n_10915) );
in01s01 g739158 ( .a(n_40913), .o(n_41041) );
na02m08 g739159 ( .a(n_40896), .b(n_40792), .o(n_40913) );
in01s01 g739160 ( .a(n_40957), .o(n_40989) );
no02s01 g739161 ( .a(n_40942), .b(n_40941), .o(n_40957) );
na02f08 g739162 ( .a(n_40958), .b(n_40853), .o(n_40956) );
oa12s02 g739163 ( .a(n_45155), .b(n_40939), .c(delay_add_ln22_unr27_stage10_stallmux_q_30_), .o(n_40940) );
in01s01 g739164 ( .a(n_40990), .o(n_40975) );
in01s01 g739165 ( .a(n_40992), .o(n_40990) );
oa12f08 g739166 ( .a(n_40848), .b(n_40938), .c(n_40753), .o(n_40992) );
ao12m01 g739167 ( .a(n_40924), .b(n_40938), .c(n_40923), .o(n_41412) );
no02s01 g739168 ( .a(n_40923), .b(n_40938), .o(n_40924) );
in01s01 g739170 ( .a(n_40914), .o(n_40895) );
na02m08 g739171 ( .a(n_40869), .b(n_40795), .o(n_40914) );
in01s01 g739172 ( .a(n_40896), .o(n_40868) );
na02s01 TIMEBOOST_cell_6925 ( .a(n_18140), .b(n_18230), .o(TIMEBOOST_net_2221) );
in01s01 g739174 ( .a(n_40942), .o(n_40960) );
no02f08 g739176 ( .a(n_41120), .b(n_40881), .o(n_40958) );
in01s01 g739177 ( .a(n_40897), .o(n_40833) );
ao12f08 g739178 ( .a(n_40672), .b(n_40801), .c(n_40735), .o(n_40897) );
oa12s01 g739179 ( .a(n_40800), .b(n_40801), .c(n_40799), .o(n_41383) );
na02s01 g739180 ( .a(n_40801), .b(n_40799), .o(n_40800) );
no02s02 TIMEBOOST_cell_1672 ( .a(TIMEBOOST_net_450), .b(n_3304), .o(n_5109) );
in01s01 g739182 ( .a(n_40894), .o(n_41206) );
ao12m04 g739183 ( .a(n_40867), .b(n_44804), .c(n_40767), .o(n_40894) );
na02f08 g739184 ( .a(n_40852), .b(n_40893), .o(n_41120) );
na02s06 g739186 ( .a(n_40911), .b(n_40860), .o(n_40912) );
na02s06 g739188 ( .a(n_40796), .b(n_40706), .o(n_40797) );
no02f06 TIMEBOOST_cell_7969 ( .a(TIMEBOOST_net_2615), .b(n_30597), .o(n_30723) );
no02m08 g739190 ( .a(n_40857), .b(n_40883), .o(n_40936) );
oa12f08 g739191 ( .a(n_40820), .b(n_40892), .c(n_40728), .o(n_40938) );
no02s01 TIMEBOOST_cell_7540 ( .a(FE_OCP_RBN2540_n_12880), .b(FE_OCP_RBN4092_n_12880), .o(TIMEBOOST_net_2401) );
ao12s06 g739193 ( .a(n_45153), .b(n_40831), .c(n_40575), .o(n_40832) );
no03f04 TIMEBOOST_cell_8431 ( .a(n_5754), .b(n_6228), .c(n_6371), .o(n_6425) );
no02m04 TIMEBOOST_cell_1759 ( .a(n_39481), .b(FE_OCPN1667_n_39207), .o(TIMEBOOST_net_494) );
oa12s06 g739196 ( .a(n_45149), .b(n_40700), .c(delay_add_ln22_unr27_stage10_stallmux_q_23_), .o(n_40794) );
oa12s02 g739197 ( .a(n_45149), .b(n_40763), .c(delay_add_ln22_unr27_stage10_stallmux_q_27_), .o(n_40865) );
ao12s02 g739198 ( .a(n_45153), .b(n_40888), .c(n_40891), .o(n_40939) );
na02s06 g739199 ( .a(n_40701), .b(n_45181), .o(n_40792) );
no02f04 TIMEBOOST_cell_1736 ( .a(TIMEBOOST_net_482), .b(n_26277), .o(n_26316) );
no02f08 TIMEBOOST_cell_8881 ( .a(TIMEBOOST_net_2927), .b(TIMEBOOST_net_904), .o(n_20907) );
oa22s01 g739202 ( .a(n_40840), .b(n_40846), .c(n_40892), .d(n_40847), .o(n_41389) );
in01s01 g739203 ( .a(FE_OCPN1220_n_40863), .o(n_40864) );
oa12s01 g739204 ( .a(n_40741), .b(n_40740), .c(n_40739), .o(n_40863) );
na02s01 g739205 ( .a(n_40869), .b(n_40790), .o(n_40791) );
na02s01 g739206 ( .a(n_40687), .b(n_40689), .o(n_40708) );
na02s02 g739207 ( .a(n_40889), .b(n_40890), .o(n_41229) );
no02s02 g739208 ( .a(n_40862), .b(n_40861), .o(n_40911) );
no02s01 g739209 ( .a(n_40859), .b(n_40843), .o(n_40860) );
na02s01 g739210 ( .a(n_40788), .b(n_40787), .o(n_40789) );
in01s01 g739211 ( .a(n_40743), .o(n_40744) );
no02s06 g739213 ( .a(n_40692), .b(n_40707), .o(n_40796) );
no02s06 g739214 ( .a(n_40704), .b(n_40705), .o(n_40706) );
na02s06 g739215 ( .a(n_40829), .b(n_40814), .o(n_40830) );
in01s01 g739216 ( .a(n_40827), .o(n_40828) );
no02s02 g739217 ( .a(n_40786), .b(n_40785), .o(n_40827) );
no02s01 TIMEBOOST_cell_4884 ( .a(n_32459), .b(n_32406), .o(TIMEBOOST_net_1390) );
ao12s06 g739219 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_21_), .b(n_45181), .c(delay_add_ln22_unr27_stage10_stallmux_q_20_), .o(n_40681) );
in01s01 g739220 ( .a(n_40783), .o(n_40784) );
na02s01 g739221 ( .a(n_40742), .b(n_40694), .o(n_40783) );
na02s01 g739222 ( .a(n_40740), .b(n_40739), .o(n_40741) );
na02s06 g739223 ( .a(n_44026), .b(n_40726), .o(n_40782) );
na02m04 TIMEBOOST_cell_5066 ( .a(n_13724), .b(n_13728), .o(TIMEBOOST_net_1481) );
na02m08 TIMEBOOST_cell_3952 ( .a(TIMEBOOST_net_1066), .b(n_24521), .o(n_24719) );
ao12s10 g739226 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_15_), .b(n_45146), .c(delay_add_ln22_unr27_stage10_stallmux_q_14_), .o(n_40679) );
in01s01 g739227 ( .a(n_40906), .o(n_40907) );
na02s01 g739228 ( .a(n_40890), .b(n_40888), .o(n_40906) );
no02s01 g739229 ( .a(n_40765), .b(n_40862), .o(n_41248) );
na02s01 g739230 ( .a(n_40887), .b(n_40886), .o(n_41260) );
na02s01 g739231 ( .a(n_40829), .b(n_40790), .o(n_41160) );
in01s01 g739232 ( .a(n_41070), .o(n_41071) );
na02s01 g739233 ( .a(n_41053), .b(n_41039), .o(n_41070) );
no02s01 g739234 ( .a(n_41010), .b(n_40785), .o(n_41165) );
na02s01 g739235 ( .a(n_40842), .b(n_40885), .o(n_41201) );
no02s01 g739236 ( .a(n_40692), .b(n_41008), .o(n_41089) );
na02s01 g739237 ( .a(n_41040), .b(n_40691), .o(n_41116) );
no02s01 g739238 ( .a(n_40972), .b(n_40988), .o(n_41032) );
no02s01 g739239 ( .a(n_40738), .b(n_40674), .o(n_41086) );
no02s01 g739240 ( .a(n_40781), .b(FE_RN_1244_0), .o(n_41016) );
oa12s01 g739241 ( .a(n_40788), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_6_), .o(n_41001) );
in01s01 g739242 ( .a(n_40954), .o(n_40955) );
na02s01 g739243 ( .a(n_40933), .b(n_40903), .o(n_40954) );
in01s01 g739244 ( .a(n_40921), .o(n_40922) );
oa12s01 g739245 ( .a(n_40889), .b(n_45153), .c(n_40891), .o(n_40921) );
ao12s01 g739246 ( .a(n_40861), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_25_), .o(n_41272) );
ao12s01 g739247 ( .a(n_40859), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_27_), .o(n_41287) );
ao12s01 g739249 ( .a(n_40815), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_19_), .o(n_41168) );
in01s01 g739250 ( .a(n_40883), .o(n_40884) );
na02s06 g739251 ( .a(n_40776), .b(n_40858), .o(n_40883) );
na02m04 g739252 ( .a(n_40856), .b(n_40772), .o(n_40857) );
in01s01 g739253 ( .a(n_41079), .o(n_41080) );
ao12s01 g739254 ( .a(n_40786), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_21_), .o(n_41079) );
ao12s01 g739255 ( .a(n_40909), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_23_), .o(n_41230) );
ao12s01 g739256 ( .a(n_40707), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_13_), .o(n_41102) );
ao12s01 g739257 ( .a(n_40705), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_15_), .o(n_41143) );
ao12s01 g739258 ( .a(n_40750), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_11_), .o(n_41099) );
oa12f08 g739260 ( .a(n_40669), .b(n_40699), .c(n_40739), .o(n_40801) );
in01s01 g739261 ( .a(n_40952), .o(n_40953) );
ao12s02 g739262 ( .a(n_40932), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_30_), .o(n_40952) );
ao12m04 g739263 ( .a(FE_OCP_RBN2441_n_44798), .b(n_40823), .c(n_40573), .o(n_40824) );
ao12m06 g739266 ( .a(FE_OCP_RBN2441_n_44798), .b(n_40882), .c(n_40558), .o(n_40941) );
oa12s06 g739267 ( .a(FE_OCP_RBN2442_n_44798), .b(n_40900), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_29_), .o(n_40905) );
na02m04 TIMEBOOST_cell_5669 ( .a(TIMEBOOST_net_1782), .b(n_17252), .o(n_17460) );
in01s01 TIMEBOOST_cell_6856 ( .a(TIMEBOOST_net_2186), .o(TIMEBOOST_net_2185) );
na02s02 TIMEBOOST_cell_7981 ( .a(TIMEBOOST_net_2621), .b(TIMEBOOST_net_1698), .o(n_5253) );
in01s01 g739271 ( .a(n_40929), .o(n_40930) );
oa12s01 g739272 ( .a(n_40877), .b(n_40876), .c(n_40875), .o(n_40929) );
oa22s01 g739273 ( .a(n_45153), .b(n_40756), .c(n_45155), .d(delay_add_ln22_unr27_stage10_stallmux_q_17_), .o(n_41146) );
oa22s01 g739274 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_9_), .c(n_45153), .d(n_40499), .o(n_41074) );
oa22s01 g739275 ( .a(n_45153), .b(n_40341), .c(n_45155), .d(delay_add_ln22_unr27_stage10_stallmux_q_5_), .o(n_40998) );
oa22s01 g739277 ( .a(n_45153), .b(n_40594), .c(n_45155), .d(delay_add_ln22_unr27_stage10_stallmux_q_31_), .o(n_40986) );
na02s01 g739278 ( .a(n_40893), .b(n_40809), .o(n_40851) );
in01s01 g739279 ( .a(n_44026), .o(n_40780) );
no02s04 g739282 ( .a(n_40775), .b(n_40774), .o(n_40776) );
no02s04 g739283 ( .a(n_40773), .b(n_40813), .o(n_40856) );
no02s02 g739284 ( .a(n_40771), .b(n_40723), .o(n_40772) );
no02s06 g739286 ( .a(n_40850), .b(n_40849), .o(n_40878) );
no02s02 g739288 ( .a(n_40770), .b(n_40769), .o(n_40934) );
no02s06 g739289 ( .a(n_40901), .b(n_40904), .o(n_41208) );
na02s01 g739290 ( .a(n_40713), .b(n_40766), .o(n_40768) );
na02s01 g739291 ( .a(n_40754), .b(n_40848), .o(n_40923) );
in01s01 g739292 ( .a(n_40846), .o(n_40847) );
na02s01 g739293 ( .a(n_40729), .b(n_40820), .o(n_40846) );
na02s01 g739294 ( .a(n_40876), .b(n_40875), .o(n_40877) );
in01s01 g739295 ( .a(n_41038), .o(n_41039) );
no02s01 g739296 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_16_), .o(n_41038) );
na02s01 g739297 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_16_), .o(n_41053) );
na02s04 g739298 ( .a(n_40766), .b(n_40508), .o(n_40767) );
in01s01 g739299 ( .a(n_40831), .o(n_40765) );
na02s06 g739300 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_24_), .o(n_40831) );
in01s01 g739302 ( .a(n_40971), .o(n_40972) );
na02s01 g739303 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_8_), .o(n_40971) );
no02s01 g739304 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_8_), .o(n_40988) );
na02s04 g739305 ( .a(n_45145), .b(delay_add_ln22_unr27_stage10_stallmux_q_18_), .o(n_40790) );
in01s01 g739306 ( .a(n_41009), .o(n_41010) );
na02s01 g739307 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_20_), .o(n_41009) );
na02s01 g739308 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_4_), .o(n_40933) );
in01s01 g739309 ( .a(n_40902), .o(n_40903) );
no02s01 g739310 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_4_), .o(n_40902) );
in01s06 g739311 ( .a(n_40885), .o(n_40700) );
na02s10 g739312 ( .a(n_45181), .b(delay_add_ln22_unr27_stage10_stallmux_q_22_), .o(n_40885) );
in01s02 g739313 ( .a(n_40887), .o(n_40763) );
na02s06 g739314 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_26_), .o(n_40887) );
in01s01 g739315 ( .a(n_40888), .o(n_40845) );
na02s01 g739316 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_28_), .o(n_40888) );
na02s01 g739317 ( .a(n_40673), .b(n_40735), .o(n_40799) );
na02s02 g739318 ( .a(n_45153), .b(n_40590), .o(n_40890) );
na02s01 g739319 ( .a(n_45153), .b(n_40891), .o(n_40889) );
no02s01 g739320 ( .a(n_40670), .b(n_40699), .o(n_40740) );
no02s01 g739321 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_24_), .o(n_40862) );
no02s01 g739322 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_25_), .o(n_40861) );
no02s01 g739323 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_27_), .o(n_40859) );
in01s01 g739324 ( .a(n_40843), .o(n_40886) );
no02s01 g739325 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_26_), .o(n_40843) );
no02s10 g739326 ( .a(FE_OCP_RBN6544_n_45145), .b(delay_add_ln22_unr27_stage10_stallmux_q_11_), .o(n_40750) );
in01s01 g739327 ( .a(n_40738), .o(n_40698) );
no02s10 g739328 ( .a(FE_OCP_RBN6544_n_45145), .b(delay_add_ln22_unr27_stage10_stallmux_q_10_), .o(n_40738) );
no02s06 g739329 ( .a(FE_OCP_RBN5544_n_45145), .b(n_40695), .o(n_40781) );
no03f04 TIMEBOOST_cell_8036 ( .a(n_31058), .b(n_30965), .c(FE_OCP_RBN6079_n_30965), .o(TIMEBOOST_net_2649) );
in01s01 g739331 ( .a(n_40734), .o(n_40788) );
no02s08 g739332 ( .a(FE_OCP_RBN5545_n_45145), .b(n_40696), .o(n_40734) );
na02s10 g739334 ( .a(n_45180), .b(n_40695), .o(n_40732) );
in01s01 g739335 ( .a(n_40693), .o(n_40694) );
no02m04 g739336 ( .a(n_40676), .b(delay_add_ln22_unr27_stage10_stallmux_q_3_), .o(n_40693) );
no02m08 TIMEBOOST_cell_3932 ( .a(TIMEBOOST_net_1056), .b(n_29405), .o(n_29470) );
na02m04 g739338 ( .a(n_40676), .b(delay_add_ln22_unr27_stage10_stallmux_q_3_), .o(n_40742) );
na02s01 TIMEBOOST_cell_7959 ( .a(TIMEBOOST_net_2610), .b(n_42971), .o(n_43388) );
in01s01 g739341 ( .a(n_40692), .o(n_40730) );
no02s06 g739342 ( .a(FE_OCP_RBN6543_n_45145), .b(delay_add_ln22_unr27_stage10_stallmux_q_12_), .o(n_40692) );
no02s06 g739343 ( .a(n_45146), .b(delay_add_ln22_unr27_stage10_stallmux_q_13_), .o(n_40707) );
no02s06 g739344 ( .a(FE_OCP_RBN6543_n_45145), .b(delay_add_ln22_unr27_stage10_stallmux_q_15_), .o(n_40705) );
in01s01 g739345 ( .a(n_40704), .o(n_40691) );
no02s06 g739346 ( .a(FE_OCP_RBN6543_n_45145), .b(delay_add_ln22_unr27_stage10_stallmux_q_14_), .o(n_40704) );
in01s01 g739347 ( .a(n_41007), .o(n_41008) );
no02f06 TIMEBOOST_cell_5065 ( .a(TIMEBOOST_net_1480), .b(FE_RN_1624_0), .o(n_13724) );
na02s01 g739349 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_12_), .o(n_41007) );
in01s01 g739351 ( .a(n_40674), .o(n_40689) );
no02s04 g739352 ( .a(n_40662), .b(n_40461), .o(n_40674) );
na02s01 g739353 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_14_), .o(n_41040) );
in01s01 g739354 ( .a(n_40814), .o(n_40815) );
na02s06 g739355 ( .a(n_45153), .b(n_40702), .o(n_40814) );
na02s06 g739356 ( .a(n_45153), .b(n_40514), .o(n_40829) );
no02s01 g739357 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_23_), .o(n_40909) );
in01s01 g739358 ( .a(n_40908), .o(n_40842) );
no02s02 g739359 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_22_), .o(n_40908) );
no02s02 g739360 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_21_), .o(n_40786) );
in01s01 g739361 ( .a(n_40785), .o(n_40758) );
no02s02 g739362 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_20_), .o(n_40785) );
no02s02 g739363 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_30_), .o(n_40932) );
no02s01 g739364 ( .a(n_41052), .b(n_41023), .o(n_41094) );
no02s01 g739365 ( .a(n_40727), .b(n_40802), .o(n_41057) );
oa12s01 g739366 ( .a(n_40717), .b(n_44775), .c(n_40299), .o(n_41054) );
in01s01 g739367 ( .a(n_41036), .o(n_41037) );
na02s01 g739368 ( .a(n_41013), .b(n_40982), .o(n_41036) );
no02s01 g739369 ( .a(n_40901), .b(n_40900), .o(n_41243) );
in01s01 g739370 ( .a(n_40949), .o(n_40950) );
na02s02 g739371 ( .a(n_40917), .b(n_40928), .o(n_40949) );
no02s01 g739372 ( .a(n_40769), .b(FE_RN_1248_0), .o(n_41240) );
na02s01 g739373 ( .a(n_40823), .b(n_40719), .o(n_41282) );
no02s01 g739374 ( .a(n_40813), .b(n_40812), .o(n_41237) );
na02s01 g739375 ( .a(n_40841), .b(n_40882), .o(n_41276) );
no02s01 g739376 ( .a(n_41107), .b(n_41078), .o(n_41183) );
no02s01 g739377 ( .a(n_40724), .b(n_40721), .o(n_41234) );
no02s01 g739378 ( .a(n_40816), .b(n_40811), .o(n_41150) );
na02s01 g739379 ( .a(n_40807), .b(n_40873), .o(n_41130) );
na02s01 g739380 ( .a(n_40810), .b(n_40809), .o(n_41127) );
in01s01 g739381 ( .a(n_40892), .o(n_40840) );
ao12f08 g739382 ( .a(n_40808), .b(n_40709), .c(n_40645), .o(n_40892) );
in01s01 g739383 ( .a(n_40969), .o(n_40970) );
ao12s02 g739384 ( .a(n_40904), .b(n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_29_), .o(n_40969) );
oa12s08 g739385 ( .a(n_45181), .b(delay_add_ln22_unr27_stage10_stallmux_q_17_), .c(delay_add_ln22_unr27_stage10_stallmux_q_16_), .o(n_40869) );
no02s10 g739386 ( .a(n_45181), .b(n_40500), .o(n_40749) );
in01s04 g739387 ( .a(n_40787), .o(n_40688) );
na02s08 g739388 ( .a(n_45145), .b(n_40342), .o(n_40787) );
ao12s01 g739389 ( .a(n_40770), .b(FE_OCPN882_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_25_), .o(n_41269) );
ao12s01 g739390 ( .a(n_40849), .b(FE_OCPN882_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_27_), .o(n_41306) );
ao12s01 g739391 ( .a(n_40773), .b(FE_OCPN882_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_21_), .o(n_41279) );
ao12s01 g739392 ( .a(n_40771), .b(FE_OCPN882_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_23_), .o(n_41303) );
no02s01 g739393 ( .a(n_45155), .b(n_40340), .o(n_40919) );
ao12s01 g739394 ( .a(n_40774), .b(FE_OCPN882_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_19_), .o(n_41266) );
in01s04 g739395 ( .a(n_40687), .o(n_40834) );
oa12s04 g739396 ( .a(n_45145), .b(delay_add_ln22_unr27_stage10_stallmux_q_8_), .c(delay_add_ln22_unr27_stage10_stallmux_q_9_), .o(n_40687) );
ao12s01 g739397 ( .a(n_40777), .b(FE_OCPN882_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_13_), .o(n_41177) );
oa12s06 g739398 ( .a(n_45153), .b(n_40756), .c(n_40494), .o(n_40757) );
ao12s01 g739399 ( .a(n_40838), .b(FE_OCPN882_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_15_), .o(n_41137) );
ao12s01 g739400 ( .a(n_40825), .b(FE_OCPN882_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_11_), .o(n_41134) );
oa22s01 g739401 ( .a(FE_OCPN882_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_), .c(n_44775), .d(n_40460), .o(n_41111) );
oa22s01 g739402 ( .a(FE_OCPN882_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_5_), .c(n_44775), .d(n_40480), .o(n_41043) );
oa22s01 g739403 ( .a(FE_OCPN882_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_17_), .c(n_44775), .d(n_40522), .o(n_41225) );
in01s01 g739404 ( .a(n_40983), .o(n_40984) );
oa22m01 g739405 ( .a(n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_31_), .c(n_44775), .d(n_40582), .o(n_40983) );
in01s01 g739406 ( .a(n_40728), .o(n_40729) );
no02f08 g739407 ( .a(n_40686), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_2_), .o(n_40728) );
no02s01 g739408 ( .a(FE_OCPN882_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_), .o(n_41052) );
in01s01 g739409 ( .a(n_41022), .o(n_41023) );
na02s01 g739410 ( .a(FE_OCPN882_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_), .o(n_41022) );
in01s01 g739411 ( .a(n_40981), .o(n_40982) );
no02s01 g739412 ( .a(FE_OCPN882_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_), .o(n_40981) );
na02s01 g739413 ( .a(FE_OCPN882_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_), .o(n_41013) );
in01s01 g739414 ( .a(n_40726), .o(n_40727) );
na02s03 g739415 ( .a(FE_OCP_RBN2430_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_7_), .o(n_40726) );
no02s01 g739416 ( .a(n_40710), .b(n_40808), .o(n_40876) );
in01s01 g739417 ( .a(n_40725), .o(n_40810) );
no02f10 g739418 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_10_), .o(n_40725) );
in01s01 g739419 ( .a(n_40917), .o(n_40918) );
na02s02 g739420 ( .a(n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_30_), .o(n_40917) );
no02f10 g739421 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_11_), .o(n_40825) );
no02m10 g739422 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_12_), .o(n_40811) );
in01s01 g739423 ( .a(n_40806), .o(n_40807) );
no02s10 g739424 ( .a(FE_OCP_RBN2443_n_44798), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_14_), .o(n_40806) );
no02m10 g739425 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_13_), .o(n_40777) );
in01s02 g739426 ( .a(n_40724), .o(n_40858) );
no02s02 g739427 ( .a(FE_OCP_RBN2431_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_18_), .o(n_40724) );
no02s02 g739428 ( .a(FE_OCP_RBN2431_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_19_), .o(n_40774) );
no02s02 g739429 ( .a(FE_OCP_RBN2431_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_21_), .o(n_40773) );
na02s04 g739430 ( .a(n_44798), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_26_), .o(n_40823) );
no02s02 g739431 ( .a(FE_OCP_RBN2431_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_20_), .o(n_40813) );
no02s02 g739432 ( .a(FE_OCP_RBN2429_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_23_), .o(n_40771) );
in01s01 g739433 ( .a(n_40723), .o(n_40841) );
no02s02 g739434 ( .a(FE_OCP_RBN2429_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_22_), .o(n_40723) );
na02m04 g739436 ( .a(FE_OCP_RBN2429_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_24_), .o(n_40822) );
in01s01 g739437 ( .a(n_40766), .o(n_40721) );
na02s04 g739438 ( .a(FE_OCP_RBN2431_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_18_), .o(n_40766) );
in01s01 g739439 ( .a(n_40720), .o(n_40812) );
na02s02 g739440 ( .a(FE_OCP_RBN2431_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_20_), .o(n_40720) );
na02s06 g739441 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_22_), .o(n_40882) );
in01s06 g739442 ( .a(n_40805), .o(n_40900) );
na02s08 g739443 ( .a(FE_OCP_RBN2442_n_44798), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_28_), .o(n_40805) );
in01s01 g739444 ( .a(n_40850), .o(n_40719) );
no02s03 g739445 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_26_), .o(n_40850) );
no02s02 g739446 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_27_), .o(n_40849) );
no02s02 g739447 ( .a(FE_OCP_RBN2429_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_25_), .o(n_40770) );
in01s01 g739448 ( .a(n_40769), .o(n_40718) );
no02s02 g739449 ( .a(FE_OCP_RBN2429_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_24_), .o(n_40769) );
na02s02 g739450 ( .a(n_44775), .b(n_40581), .o(n_40928) );
in01s01 g739451 ( .a(n_40901), .o(n_40872) );
no02s06 g739452 ( .a(FE_OCP_RBN2442_n_44798), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_28_), .o(n_40901) );
no02s06 g739453 ( .a(FE_OCP_RBN2442_n_44798), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_29_), .o(n_40904) );
na02s06 g739454 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_14_), .o(n_40873) );
na02m08 g739455 ( .a(FE_OCP_RBN2431_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_10_), .o(n_40809) );
in01s01 g739456 ( .a(n_40669), .o(n_40670) );
na02f06 g739457 ( .a(n_40663), .b(delay_add_ln22_unr27_stage10_stallmux_q_1_), .o(n_40669) );
no02m08 g739458 ( .a(n_40663), .b(delay_add_ln22_unr27_stage10_stallmux_q_1_), .o(n_40699) );
no02s06 g739459 ( .a(FE_OCP_RBN2433_FE_RN_107_0), .b(n_40454), .o(n_40816) );
na02m08 g739460 ( .a(n_40668), .b(n_40667), .o(n_40735) );
in01s01 g739461 ( .a(n_40837), .o(n_40838) );
na02s10 g739462 ( .a(n_44775), .b(n_40761), .o(n_40837) );
in01s01 g739463 ( .a(n_40672), .o(n_40673) );
no02f06 g739464 ( .a(n_40668), .b(n_40667), .o(n_40672) );
in01s01 g739465 ( .a(n_41077), .o(n_41078) );
na02s01 g739466 ( .a(FE_OCPN882_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_), .o(n_41077) );
no02s01 g739467 ( .a(FE_OCPN882_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_), .o(n_41107) );
in01s06 g739468 ( .a(n_40802), .o(n_40803) );
no02s06 g739469 ( .a(n_44798), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_7_), .o(n_40802) );
in01s01 g739470 ( .a(n_40716), .o(n_40717) );
no02s08 g739471 ( .a(FE_OCP_RBN2430_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_6_), .o(n_40716) );
na02f08 g739472 ( .a(n_40715), .b(n_40714), .o(n_40848) );
in01s01 g739473 ( .a(n_40753), .o(n_40754) );
no02f08 g739474 ( .a(n_40715), .b(n_40714), .o(n_40753) );
na02f08 g739475 ( .a(n_40686), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_2_), .o(n_40820) );
na02s01 g739476 ( .a(FE_OCPN882_n_44776), .b(n_40737), .o(n_41006) );
no02s02 g739478 ( .a(FE_OCP_RBN2431_FE_RN_107_0), .b(n_40523), .o(n_40775) );
in01s02 g739479 ( .a(n_40713), .o(n_40867) );
oa12s02 g739480 ( .a(FE_OCP_RBN2431_FE_RN_107_0), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_17_), .o(n_40713) );
in01s01 g739482 ( .a(n_40711), .o(n_40712) );
no02s08 g739483 ( .a(FE_OCP_RBN2430_FE_RN_107_0), .b(n_40479), .o(n_40711) );
oa12m40 g739512 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_3_), .b(FE_OCP_RBN6503_n_44610), .c(n_47203), .o(n_40662) );
no02f08 g739514 ( .a(n_40685), .b(n_40684), .o(n_40808) );
in01s01 g739515 ( .a(n_40709), .o(n_40710) );
na02f08 g739516 ( .a(n_40685), .b(n_40684), .o(n_40709) );
ao22f10 g739549 ( .a(n_40646), .b(n_40652), .c(n_40650), .d(n_40651), .o(n_40686) );
na02f10 g739552 ( .a(n_40660), .b(n_44027), .o(n_40685) );
in01s01 g739553 ( .a(n_41309), .o(n_40657) );
oa12s01 g739554 ( .a(n_40634), .b(n_40633), .c(delay_add_ln22_unr27_stage10_stallmux_q_0_), .o(n_41309) );
na02s06 TIMEBOOST_cell_3853 ( .a(n_23160), .b(n_23161), .o(TIMEBOOST_net_1017) );
na02s06 g739558 ( .a(n_45511), .b(n_40617), .o(n_40639) );
na02s01 g739561 ( .a(n_40633), .b(delay_add_ln22_unr27_stage10_stallmux_q_0_), .o(n_40634) );
na02s06 g739562 ( .a(n_40616), .b(delay_add_ln22_unr27_stage10_stallmux_q_0_), .o(n_40739) );
in01f10 g739563 ( .a(n_40651), .o(n_40652) );
na02f40 g739564 ( .a(n_40647), .b(n_40622), .o(n_40651) );
na02m10 g739566 ( .a(n_40609), .b(n_40617), .o(n_40631) );
in01m06 g739567 ( .a(n_40629), .o(n_40630) );
na02m10 g739568 ( .a(n_45513), .b(n_40608), .o(n_40629) );
in01s01 g739569 ( .a(n_41343), .o(n_40658) );
ao12s01 g739570 ( .a(n_40636), .b(n_40638), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_0_), .o(n_41343) );
in01m04 g739571 ( .a(n_40627), .o(n_40628) );
na02m08 g739572 ( .a(n_40610), .b(n_40612), .o(n_40627) );
no02f10 g739573 ( .a(n_40649), .b(n_40655), .o(n_40650) );
na02m10 g739574 ( .a(n_40653), .b(n_40654), .o(n_40646) );
na02f20 g739575 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_2_), .b(FE_OCP_RBN6501_n_44610), .o(n_40622) );
in01s01 g739576 ( .a(n_40645), .o(n_40875) );
na02m08 g739577 ( .a(n_40638), .b(n_39737), .o(n_40645) );
in01f08 g739578 ( .a(n_40647), .o(n_40637) );
na02f80 g739579 ( .a(n_40615), .b(n_44610), .o(n_40647) );
in01m20 g739583 ( .a(n_40617), .o(n_40619) );
na02m40 g739584 ( .a(n_40604), .b(n_44610), .o(n_40617) );
na02s03 g739585 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_3_), .b(FE_OCP_RBN6500_n_44610), .o(n_40610) );
na02m03 g739586 ( .a(n_40602), .b(n_44610), .o(n_40612) );
na02s10 g739587 ( .a(FE_OCP_RBN6499_n_44610), .b(delay_xor_ln22_unr28_stage10_stallmux_q_1_), .o(n_40609) );
na02s10 g739588 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_2_), .b(FE_OCP_RBN6499_n_44610), .o(n_40608) );
no02s01 g739589 ( .a(n_40638), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_0_), .o(n_40636) );
in01f06 g739590 ( .a(n_40643), .o(n_40644) );
oa22f10 g739591 ( .a(FE_OCP_RBN6500_n_44610), .b(delay_xor_ln21_unr28_stage10_stallmux_q_3_), .c(n_40624), .d(n_44610), .o(n_40643) );
na02s06 TIMEBOOST_cell_3852 ( .a(n_7335), .b(TIMEBOOST_net_1016), .o(n_7389) );
in01s01 g739593 ( .a(n_40616), .o(n_40633) );
ao22s06 g739594 ( .a(FE_OCP_RBN6499_n_44610), .b(n_40611), .c(n_44610), .d(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .o(n_40616) );
in01f80 g739595 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_2_), .o(n_40615) );
in01m40 g739599 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_1_), .o(n_40604) );
in01m03 g739602 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_3_), .o(n_40602) );
in01f10 g739604 ( .a(n_40654), .o(n_40649) );
na02f80 g739605 ( .a(n_40614), .b(n_44610), .o(n_40654) );
na02f20 g739606 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_1_), .b(FE_OCP_RBN6501_n_44610), .o(n_40641) );
na02f06 TIMEBOOST_cell_2937 ( .a(TIMEBOOST_net_759), .b(n_41419), .o(n_41506) );
no02s10 g739609 ( .a(FE_OCP_RBN6499_n_44610), .b(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .o(n_40601) );
ao22m08 g739611 ( .a(FE_OCP_RBN5498_n_44610), .b(n_40607), .c(n_44610), .d(delay_xor_ln21_unr28_stage10_stallmux_q_0_), .o(n_40638) );
in01f80 g739612 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_1_), .o(n_40614) );
in01m40 g739617 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_3_), .o(n_40624) );
no02f40 g739620 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_0_), .b(FE_OCP_RBN5498_n_44610), .o(n_40655) );
na02f80 g739621 ( .a(n_40607), .b(n_44610), .o(n_40653) );
oa22f02 g739622 ( .a(n_40586), .b(delay_sub_ln23_0_unr27_stage10_stallmux_z), .c(FE_OCP_RBN6236_n_40586), .d(n_40598), .o(n_40600) );
in01f40 g739626 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_0_), .o(n_40607) );
in01s01 g739629 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_31_), .o(n_40582) );
in01s01 g739631 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_30_), .o(n_40581) );
oa22m02 g739636 ( .a(n_40592), .b(n_40598), .c(n_40583), .d(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n_40597) );
in01s01 g739638 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_27_), .o(n_40573) );
in01s01 g739641 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_25_), .o(n_40572) );
in01s01 g739644 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_29_), .o(n_40891) );
in01s01 g739646 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_31_), .o(n_40594) );
oa22f02 g739648 ( .a(n_40585), .b(n_40598), .c(n_40574), .d(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n_40591) );
na02m06 TIMEBOOST_cell_4187 ( .a(FE_RN_1284_0), .b(n_27439), .o(TIMEBOOST_net_1184) );
no02f02 TIMEBOOST_cell_8061 ( .a(TIMEBOOST_net_2661), .b(n_40131), .o(TIMEBOOST_net_954) );
no02s01 TIMEBOOST_cell_1536 ( .a(TIMEBOOST_net_382), .b(n_14948), .o(n_15030) );
ao22f04 g739656 ( .a(n_40565), .b(n_40271), .c(FE_OCP_RBN6228_n_40565), .d(n_40272), .o(n_40586) );
in01s01 g739658 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_23_), .o(n_40558) );
in01s01 g739661 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_28_), .o(n_40590) );
na02s02 TIMEBOOST_cell_4026 ( .a(TIMEBOOST_net_1103), .b(n_4524), .o(n_4692) );
na02f04 g739664 ( .a(n_40537), .b(n_40249), .o(n_40557) );
na02m10 TIMEBOOST_cell_7427 ( .a(TIMEBOOST_net_2344), .b(FE_RN_1561_0), .o(FE_RN_1562_0) );
na02m04 g739666 ( .a(n_40535), .b(n_40224), .o(n_40556) );
no02s01 TIMEBOOST_cell_1535 ( .a(n_14947), .b(n_14338), .o(TIMEBOOST_net_382) );
na02m04 g739668 ( .a(n_44692), .b(n_40222), .o(n_40555) );
oa22f02 g739669 ( .a(n_40519), .b(n_40279), .c(n_40520), .d(n_40280), .o(n_40554) );
oa22s02 g739670 ( .a(n_40114), .b(n_40517), .c(n_40518), .d(n_40115), .o(n_40553) );
oa22m02 g739671 ( .a(n_40515), .b(n_40277), .c(n_40516), .d(n_40278), .o(n_40552) );
in01s02 g739672 ( .a(n_40568), .o(n_40576) );
in01f02 g739674 ( .a(n_40593), .o(n_40584) );
in01m02 g739676 ( .a(n_40592), .o(n_40583) );
oa22m06 g739677 ( .a(n_40561), .b(n_40304), .c(n_45198), .d(n_40305), .o(n_40592) );
in01s01 g739678 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_25_), .o(n_40575) );
oa22f02 g739684 ( .a(n_40491), .b(n_40281), .c(n_40492), .d(n_40282), .o(n_40525) );
in01f02 g739686 ( .a(n_40536), .o(n_40537) );
oa12f04 g739687 ( .a(n_40376), .b(n_40524), .c(n_40112), .o(n_40536) );
in01s02 g739688 ( .a(n_40534), .o(n_40535) );
oa12m04 g739689 ( .a(n_40375), .b(n_40524), .c(n_40138), .o(n_40534) );
oa12m06 g739691 ( .a(n_40373), .b(n_40524), .c(n_40191), .o(n_40532) );
oa22s02 g739692 ( .a(n_40540), .b(n_40354), .c(n_40541), .d(n_40353), .o(n_40567) );
in01f02 g739693 ( .a(n_40574), .o(n_40585) );
ao22m04 g739694 ( .a(n_40550), .b(n_40213), .c(n_40543), .d(n_40212), .o(n_40574) );
oa12m06 g739696 ( .a(n_40211), .b(n_40543), .c(n_40251), .o(n_40565) );
in01s01 g739697 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_19_), .o(n_40508) );
no02s01 g739702 ( .a(n_40471), .b(n_40522), .o(n_40523) );
no02s02 g739703 ( .a(n_40501), .b(n_40374), .o(n_40521) );
na02m04 g739704 ( .a(n_40502), .b(n_40371), .o(n_40531) );
oa22m02 g739705 ( .a(n_40473), .b(n_40283), .c(n_40474), .d(n_40284), .o(n_40507) );
oa22f02 g739706 ( .a(n_40475), .b(n_40146), .c(n_40476), .d(n_40145), .o(n_40506) );
in01m02 g739707 ( .a(n_40519), .o(n_40520) );
oa12m02 g739708 ( .a(n_40338), .b(n_40505), .c(n_40117), .o(n_40519) );
in01f02 g739709 ( .a(n_40517), .o(n_40518) );
oa12f02 g739710 ( .a(n_40337), .b(n_40505), .c(n_40113), .o(n_40517) );
in01m01 g739711 ( .a(n_40515), .o(n_40516) );
oa12s02 g739712 ( .a(n_40335), .b(n_40505), .c(n_40192), .o(n_40515) );
oa22m02 g739713 ( .a(n_40526), .b(n_40390), .c(n_40527), .d(n_40391), .o(n_40560) );
oa22m02 g739714 ( .a(n_40528), .b(n_40172), .c(n_40529), .d(n_40171), .o(n_40559) );
na02s02 TIMEBOOST_cell_6830 ( .a(TIMEBOOST_net_2172), .b(n_31683), .o(n_31684) );
no02s01 TIMEBOOST_cell_1372 ( .a(TIMEBOOST_net_300), .b(n_13136), .o(n_13306) );
in01s01 g739720 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_17_), .o(n_40522) );
in01m02 g739723 ( .a(n_40503), .o(n_40504) );
na02s02 g739724 ( .a(n_40505), .b(n_40257), .o(n_40503) );
in01m02 g739726 ( .a(n_40543), .o(n_40550) );
na02m08 g739727 ( .a(n_40511), .b(n_40409), .o(n_40543) );
na02f08 TIMEBOOST_cell_8039 ( .a(TIMEBOOST_net_2650), .b(n_31518), .o(n_31563) );
oa22m02 g739729 ( .a(n_40434), .b(n_40285), .c(n_40435), .d(n_40286), .o(n_40477) );
oa22s01 g739730 ( .a(n_40462), .b(n_40077), .c(n_40463), .d(n_40076), .o(n_40498) );
in01f01 g739731 ( .a(n_40491), .o(n_40492) );
oa12m01 g739732 ( .a(n_40229), .b(n_40466), .c(n_40119), .o(n_40491) );
in01s02 g739733 ( .a(n_40501), .o(n_40502) );
in01s04 g739734 ( .a(n_40524), .o(n_40501) );
oa22s02 g739736 ( .a(n_40496), .b(n_40408), .c(n_40497), .d(n_40407), .o(n_40530) );
oa22s01 g739737 ( .a(n_40509), .b(n_40174), .c(n_40510), .d(n_40173), .o(n_40549) );
in01s02 g739738 ( .a(n_40540), .o(n_40541) );
oa12s02 g739739 ( .a(n_40399), .b(n_40513), .c(n_40130), .o(n_40540) );
no02s01 TIMEBOOST_cell_1371 ( .a(n_12857), .b(n_12854), .o(TIMEBOOST_net_300) );
in01s01 g739741 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_19_), .o(n_40702) );
in01s01 g739743 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_18_), .o(n_40514) );
in01s01 g739745 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_17_), .o(n_40756) );
in01m01 g739749 ( .a(n_40475), .o(n_40476) );
na02s02 g739750 ( .a(n_40466), .b(n_40196), .o(n_40475) );
in01m02 g739751 ( .a(n_40528), .o(n_40529) );
na02m02 g739752 ( .a(n_40513), .b(n_40367), .o(n_40528) );
oa22s01 g739753 ( .a(n_40423), .b(n_40324), .c(n_40424), .d(n_40325), .o(n_40465) );
oa22s02 g739754 ( .a(n_40425), .b(n_40079), .c(n_40426), .d(n_40078), .o(n_40464) );
in01s02 g739755 ( .a(n_40473), .o(n_40474) );
oa12m02 g739756 ( .a(n_40197), .b(n_40456), .c(n_40042), .o(n_40473) );
in01s06 g739757 ( .a(n_40472), .o(n_40505) );
oa22s01 g739759 ( .a(n_40484), .b(n_40103), .c(n_40485), .d(n_40102), .o(n_40512) );
in01m01 g739760 ( .a(n_40526), .o(n_40527) );
oa12m01 g739761 ( .a(n_40368), .b(n_40468), .c(n_40132), .o(n_40526) );
in01f04 g739762 ( .a(n_40511), .o(n_40538) );
in01s01 g739764 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_), .o(n_40471) );
in01s06 g739766 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_15_), .o(n_40761) );
in01s01 g739769 ( .a(n_40462), .o(n_40463) );
na02s02 g739770 ( .a(n_40456), .b(n_40121), .o(n_40462) );
in01s01 g739771 ( .a(n_40509), .o(n_40510) );
na02s01 g739772 ( .a(n_40468), .b(n_40295), .o(n_40509) );
in01m01 g739773 ( .a(n_40434), .o(n_40435) );
oa12s01 g739774 ( .a(n_40017), .b(n_40406), .c(n_40043), .o(n_40434) );
oa22s01 g739776 ( .a(n_40450), .b(n_40394), .c(n_40451), .d(n_40395), .o(n_40490) );
oa22s02 g739777 ( .a(n_40448), .b(n_40311), .c(n_40449), .d(n_40312), .o(n_40489) );
oa22s01 g739778 ( .a(n_40446), .b(n_40392), .c(n_40447), .d(n_40393), .o(n_40488) );
oa22m01 g739779 ( .a(n_40444), .b(n_40062), .c(n_40445), .d(n_40061), .o(n_40487) );
oa22s01 g739780 ( .a(n_40442), .b(n_40356), .c(n_40443), .d(n_40355), .o(n_40486) );
in01s01 g739781 ( .a(n_40496), .o(n_40497) );
oa12s02 g739782 ( .a(n_40256), .b(n_40470), .c(n_40060), .o(n_40496) );
in01s01 g739783 ( .a(n_40495), .o(n_40513) );
no02f08 g739784 ( .a(n_40468), .b(n_40101), .o(n_40495) );
in01s01 g739785 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_16_), .o(n_40494) );
in01s02 g739789 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_11_), .o(n_40455) );
in01s01 g739792 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_13_), .o(n_40493) );
no02s06 g739795 ( .a(n_40467), .b(n_40499), .o(n_40500) );
in01s01 g739796 ( .a(n_40425), .o(n_40426) );
na02s01 g739797 ( .a(n_40406), .b(n_39976), .o(n_40425) );
in01s01 g739798 ( .a(n_40484), .o(n_40485) );
na02s02 g739799 ( .a(n_40470), .b(n_40225), .o(n_40484) );
oa22m02 g739800 ( .a(n_40301), .b(n_40287), .c(n_40302), .d(n_40288), .o(n_40405) );
oa22s01 g739801 ( .a(n_40383), .b(n_40330), .c(FE_OCP_RBN3420_n_40300), .d(n_40331), .o(n_40433) );
in01s02 g739802 ( .a(n_40423), .o(n_40424) );
oa12s01 g739803 ( .a(n_40292), .b(FE_OCP_RBN3420_n_40300), .c(n_40218), .o(n_40423) );
in01s01 g739804 ( .a(n_40422), .o(n_40456) );
oa22m02 g739806 ( .a(n_40429), .b(n_40358), .c(n_40430), .d(n_40357), .o(n_40469) );
na02f08 g739810 ( .a(n_40058), .b(n_40453), .o(n_40468) );
in01s01 g739811 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_9_), .o(n_40499) );
in01s01 g739813 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_10_), .o(n_40461) );
in01s01 g739815 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_), .o(n_40460) );
in01s01 g739818 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_12_), .o(n_40454) );
na02f08 g739821 ( .a(n_40300), .b(n_39944), .o(n_40406) );
in01s01 g739822 ( .a(n_40453), .o(n_40470) );
no02f08 g739823 ( .a(n_40431), .b(n_40308), .o(n_40453) );
oa22m02 g739824 ( .a(n_40261), .b(n_40289), .c(n_40262), .d(n_40290), .o(n_40404) );
oa22s02 g739825 ( .a(n_40347), .b(n_40327), .c(n_40348), .d(n_40326), .o(n_40421) );
oa22s01 g739826 ( .a(n_40263), .b(n_40019), .c(n_40264), .d(n_40018), .o(n_40385) );
oa22f02 g739827 ( .a(n_40381), .b(n_40396), .c(n_40382), .d(n_40397), .o(n_40452) );
oa22s02 g739828 ( .a(n_40414), .b(n_40360), .c(n_40415), .d(n_40359), .o(n_40459) );
oa22s01 g739829 ( .a(n_40417), .b(n_40315), .c(n_40418), .d(n_40314), .o(n_40458) );
oa22s01 g739830 ( .a(n_40412), .b(n_40365), .c(n_40432), .d(n_40366), .o(n_40457) );
in01s01 g739831 ( .a(n_40450), .o(n_40451) );
oa12s02 g739832 ( .a(n_40313), .b(n_40432), .c(n_40242), .o(n_40450) );
in01s02 g739833 ( .a(n_40448), .o(n_40449) );
oa12s02 g739834 ( .a(n_40064), .b(n_40432), .c(n_39931), .o(n_40448) );
in01s01 g739835 ( .a(n_40446), .o(n_40447) );
oa12s02 g739836 ( .a(n_40253), .b(n_40432), .c(n_39968), .o(n_40446) );
in01s01 g739837 ( .a(n_40444), .o(n_40445) );
oa12s01 g739838 ( .a(n_40136), .b(n_40432), .c(n_40066), .o(n_40444) );
in01s01 g739839 ( .a(n_40442), .o(n_40443) );
na02s01 g739840 ( .a(n_40431), .b(n_40226), .o(n_40442) );
oa22s01 g739842 ( .a(n_40234), .b(n_39984), .c(n_40235), .d(n_39985), .o(n_40350) );
oa22s01 g739843 ( .a(n_40232), .b(n_40294), .c(n_40233), .d(n_40293), .o(n_40403) );
in01m01 g739844 ( .a(n_40301), .o(n_40302) );
oa12m01 g739845 ( .a(n_40091), .b(n_40265), .c(n_39983), .o(n_40301) );
in01s01 g739847 ( .a(FE_OCP_RBN3420_n_40300), .o(n_40383) );
oa12f08 g739849 ( .a(n_40090), .b(n_40265), .c(n_39954), .o(n_40300) );
oa22s01 g739850 ( .a(n_40343), .b(n_40318), .c(n_40344), .d(n_40319), .o(n_40420) );
oa22s01 g739851 ( .a(n_40345), .b(n_39972), .c(n_40346), .d(n_39971), .o(n_40419) );
oa22s01 g739852 ( .a(n_40400), .b(n_40317), .c(n_40401), .d(n_40316), .o(n_40441) );
in01s02 g739853 ( .a(n_40429), .o(n_40430) );
oa12s02 g739854 ( .a(n_40194), .b(n_40402), .c(n_40273), .o(n_40429) );
na02f08 g739855 ( .a(n_40380), .b(n_40067), .o(n_40431) );
oa22s01 g739856 ( .a(n_40377), .b(n_40386), .c(n_40378), .d(n_40387), .o(n_40440) );
in01s01 g739857 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_8_), .o(n_40467) );
in01s06 g739859 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_7_), .o(n_40695) );
in01s01 g739862 ( .a(n_40263), .o(n_40264) );
na02s01 g739863 ( .a(n_40265), .b(n_40046), .o(n_40263) );
in01s01 g739864 ( .a(n_40417), .o(n_40418) );
na02s02 g739865 ( .a(n_40402), .b(n_40151), .o(n_40417) );
in01s02 g739866 ( .a(n_40261), .o(n_40262) );
oa12m02 g739867 ( .a(n_39908), .b(n_40200), .c(n_39902), .o(n_40261) );
in01s01 g739868 ( .a(n_40347), .o(n_40348) );
oa12s02 g739869 ( .a(n_40048), .b(n_40199), .c(n_40254), .o(n_40347) );
oa22s02 g739870 ( .a(n_40164), .b(n_40320), .c(n_40165), .d(n_40321), .o(n_40416) );
in01s02 g739871 ( .a(n_40381), .o(n_40382) );
oa12m02 g739872 ( .a(n_40039), .b(n_40298), .c(n_39973), .o(n_40381) );
in01m02 g739873 ( .a(n_40414), .o(n_40415) );
oa12s02 g739874 ( .a(n_40153), .b(n_40379), .c(n_40274), .o(n_40414) );
in01s01 g739876 ( .a(n_40432), .o(n_40412) );
in01m01 g739877 ( .a(n_40380), .o(n_40432) );
oa12f08 g739878 ( .a(n_40080), .b(n_40260), .c(n_39997), .o(n_40380) );
in01s01 g739879 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_6_), .o(n_40299) );
na02s01 g739881 ( .a(n_40478), .b(n_40480), .o(n_40737) );
no02s01 g739882 ( .a(n_40480), .b(n_40478), .o(n_40479) );
in01s01 g739883 ( .a(n_40234), .o(n_40235) );
na02s01 g739884 ( .a(n_40200), .b(n_39862), .o(n_40234) );
in01s01 g739885 ( .a(n_40232), .o(n_40233) );
na02s01 g739886 ( .a(n_40199), .b(FE_OCP_RBN3394_FE_RN_1094_0), .o(n_40232) );
in01s01 g739887 ( .a(n_40345), .o(n_40346) );
na02s01 g739888 ( .a(n_40298), .b(n_39975), .o(n_40345) );
in01s01 g739889 ( .a(n_40400), .o(n_40401) );
na02s02 g739890 ( .a(n_40379), .b(n_40068), .o(n_40400) );
na02s02 g739891 ( .a(n_40297), .b(n_39996), .o(n_40402) );
na02f08 g739892 ( .a(n_40124), .b(n_39922), .o(n_40265) );
oa22s01 g739893 ( .a(n_40092), .b(n_40328), .c(n_40123), .d(n_40329), .o(n_40411) );
in01s01 g739894 ( .a(n_40343), .o(n_40344) );
oa12s01 g739895 ( .a(n_40291), .b(n_40123), .c(n_40214), .o(n_40343) );
oa22s01 g739896 ( .a(n_40369), .b(n_40389), .c(n_40370), .d(n_40388), .o(n_40439) );
oa22s01 g739897 ( .a(n_40230), .b(n_40362), .c(n_40258), .d(n_40361), .o(n_40428) );
in01s01 g739898 ( .a(n_40377), .o(n_40378) );
oa12s01 g739899 ( .a(n_40309), .b(n_40230), .c(n_40238), .o(n_40377) );
in01m01 g739900 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_6_), .o(n_40696) );
in01s01 g739902 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_5_), .o(n_40480) );
na02s01 g739904 ( .a(n_40084), .b(n_40341), .o(n_40342) );
in01s01 g739905 ( .a(n_40339), .o(n_40340) );
na02s02 g739906 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_5_), .b(delay_add_ln22_unr27_stage10_stallmux_q_4_), .o(n_40339) );
na02f01 g739907 ( .a(n_40092), .b(n_39925), .o(n_40200) );
no02s04 g739908 ( .a(n_40374), .b(n_40111), .o(n_40376) );
no02s02 g739909 ( .a(n_40374), .b(n_40154), .o(n_40375) );
na02f08 TIMEBOOST_cell_6716 ( .a(TIMEBOOST_net_2115), .b(n_14583), .o(n_14716) );
na02m01 g739911 ( .a(n_40231), .b(n_39914), .o(n_40298) );
in01s01 g739912 ( .a(n_40124), .o(n_40199) );
oa22s01 g739914 ( .a(n_40049), .b(n_39919), .c(n_40087), .d(n_39920), .o(n_40198) );
in01s01 g739915 ( .a(n_40164), .o(n_40165) );
oa12s02 g739916 ( .a(n_39904), .b(n_40049), .c(n_39820), .o(n_40164) );
in01s01 g739917 ( .a(n_40297), .o(n_40379) );
in01s01 g739918 ( .a(n_40260), .o(n_40297) );
na02f08 g739919 ( .a(n_40231), .b(n_39974), .o(n_40260) );
in01s01 g739920 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_5_), .o(n_40341) );
no02s02 g739922 ( .a(n_40336), .b(n_40116), .o(n_40338) );
no02s02 g739923 ( .a(n_40336), .b(n_40120), .o(n_40337) );
no02f06 g739924 ( .a(n_40436), .b(n_40097), .o(n_40438) );
no02s06 g739925 ( .a(n_40436), .b(n_40332), .o(n_40437) );
in01s01 g739928 ( .a(n_40092), .o(n_40123) );
in01m01 g739929 ( .a(n_40050), .o(n_40092) );
ao12f08 g739930 ( .a(n_39928), .b(n_39959), .c(n_39873), .o(n_40050) );
no02s01 g739931 ( .a(n_40336), .b(n_40195), .o(n_40335) );
in01s01 g739933 ( .a(n_40374), .o(n_40371) );
na02s08 g739934 ( .a(n_40257), .b(n_40156), .o(n_40374) );
oa22s01 g739935 ( .a(n_39961), .b(n_40322), .c(n_39962), .d(n_40323), .o(n_40410) );
in01s01 g739937 ( .a(n_40230), .o(n_40258) );
in01s01 g739938 ( .a(n_40231), .o(n_40230) );
ao12f08 g739939 ( .a(n_39860), .b(n_40086), .c(n_39897), .o(n_40231) );
oa22s01 g739940 ( .a(n_40122), .b(n_40363), .c(n_40159), .d(n_40364), .o(n_40427) );
in01s01 g739941 ( .a(n_40369), .o(n_40370) );
oa12s01 g739942 ( .a(n_40310), .b(n_40122), .c(n_39833), .o(n_40369) );
in01s01 g739943 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_), .o(n_40478) );
no02s01 g739945 ( .a(n_40089), .b(n_39982), .o(n_40091) );
no03s04 TIMEBOOST_cell_3484 ( .a(n_23176), .b(n_23175), .c(delay_add_ln22_unr14_stage6_stallmux_q_7_), .o(n_23251) );
no02s01 g739947 ( .a(n_40228), .b(n_40118), .o(n_40229) );
in01s01 g739949 ( .a(n_40257), .o(n_40336) );
no02s08 g739950 ( .a(n_40228), .b(n_40083), .o(n_40257) );
in01s01 g739952 ( .a(n_40049), .o(n_40087) );
na02m01 g739953 ( .a(n_39960), .b(n_39927), .o(n_40049) );
no02s01 g739954 ( .a(n_40398), .b(n_40131), .o(n_40399) );
in01m08 g739955 ( .a(n_40409), .o(n_40436) );
no02f08 TIMEBOOST_cell_1300 ( .a(n_29301), .b(TIMEBOOST_net_264), .o(n_30192) );
no02m02 TIMEBOOST_cell_1286 ( .a(n_18602), .b(TIMEBOOST_net_257), .o(n_18652) );
no02s01 g739958 ( .a(n_40024), .b(n_40047), .o(n_40048) );
in01s01 g739959 ( .a(n_40089), .o(n_40046) );
na02f08 g739960 ( .a(FE_OCP_RBN3395_FE_RN_1094_0), .b(n_39923), .o(n_40089) );
no02s01 g739961 ( .a(n_40157), .b(n_40041), .o(n_40197) );
in01s01 g739962 ( .a(n_40228), .o(n_40196) );
na02m08 g739963 ( .a(n_40121), .b(n_40044), .o(n_40228) );
in01s01 g739964 ( .a(n_39961), .o(n_39962) );
na02s01 g739965 ( .a(n_39929), .b(n_39796), .o(n_39961) );
in01s01 g739967 ( .a(n_40122), .o(n_40159) );
in01s01 g739968 ( .a(n_40086), .o(n_40122) );
na02f08 g739969 ( .a(n_40022), .b(n_40045), .o(n_40086) );
no02s01 g739970 ( .a(n_40333), .b(n_40133), .o(n_40368) );
in01s01 g739971 ( .a(n_40398), .o(n_40367) );
na02s10 g739972 ( .a(n_40134), .b(n_40295), .o(n_40398) );
na02s01 g739973 ( .a(n_40023), .b(n_40045), .o(n_40085) );
in01s01 g739974 ( .a(n_39959), .o(n_39960) );
no02f08 g739975 ( .a(n_39929), .b(n_39818), .o(n_39959) );
no02m04 TIMEBOOST_cell_1366 ( .a(TIMEBOOST_net_297), .b(n_18871), .o(n_18925) );
oa22s01 g739977 ( .a(n_39875), .b(n_39814), .c(n_39874), .d(n_39815), .o(n_39958) );
in01s01 g739978 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_4_), .o(n_40084) );
in01s01 g739980 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_3_), .o(n_40714) );
na02f06 g739982 ( .a(n_39876), .b(n_39927), .o(n_39928) );
na02f08 g739983 ( .a(n_39849), .b(n_39795), .o(n_39929) );
in01s01 g739985 ( .a(FE_OCP_RBN3394_FE_RN_1094_0), .o(n_40024) );
in01s01 g739988 ( .a(n_40121), .o(n_40157) );
no02m06 g739989 ( .a(n_40020), .b(n_40016), .o(n_40121) );
na02s01 g739990 ( .a(n_40148), .b(n_40072), .o(n_40195) );
no02s06 g739991 ( .a(n_40120), .b(n_40081), .o(n_40156) );
no02m04 TIMEBOOST_cell_1365 ( .a(n_18870), .b(n_18514), .o(TIMEBOOST_net_297) );
in01s01 g739993 ( .a(n_40022), .o(n_40023) );
na02f08 g739994 ( .a(n_39955), .b(n_39857), .o(n_40022) );
no02s02 g739995 ( .a(n_40150), .b(n_40193), .o(n_40194) );
no02s01 g739996 ( .a(n_40255), .b(n_40059), .o(n_40256) );
in01s01 g739998 ( .a(n_40295), .o(n_40333) );
no02m10 g739999 ( .a(n_40255), .b(n_40104), .o(n_40295) );
no02m02 TIMEBOOST_cell_1285 ( .a(n_18317), .b(n_18263), .o(TIMEBOOST_net_257) );
na02s01 g740002 ( .a(n_40141), .b(n_40073), .o(n_40192) );
na02s04 g740003 ( .a(n_40137), .b(n_40188), .o(n_40191) );
no02s01 g740004 ( .a(n_40038), .b(n_40152), .o(n_40153) );
in01s01 g740005 ( .a(n_40150), .o(n_40151) );
na02m01 g740006 ( .a(n_40068), .b(n_40003), .o(n_40150) );
no02s01 g740007 ( .a(n_40189), .b(n_40033), .o(n_40226) );
in01s01 g740008 ( .a(n_40255), .o(n_40225) );
na02m10 g740009 ( .a(n_40136), .b(n_40063), .o(n_40255) );
na02s04 TIMEBOOST_cell_8626 ( .a(FE_RN_1126_0), .b(FE_OCP_RBN4393_n_10682), .o(TIMEBOOST_net_2800) );
in01s01 g740011 ( .a(n_39874), .o(n_39875) );
in01s01 g740012 ( .a(n_39849), .o(n_39874) );
oa12f06 g740013 ( .a(n_39771), .b(n_39824), .c(n_39751), .o(n_39849) );
na02m04 g740015 ( .a(n_39870), .b(n_39816), .o(n_39923) );
no02s02 TIMEBOOST_cell_8547 ( .a(TIMEBOOST_net_2760), .b(FE_RN_1907_0), .o(FE_RN_1908_0) );
no02s01 TIMEBOOST_cell_1244 ( .a(TIMEBOOST_net_236), .b(n_45897), .o(n_38372) );
na02s06 g740018 ( .a(n_39981), .b(FE_OCP_RBN6157_n_39816), .o(n_40044) );
na02s01 TIMEBOOST_cell_1246 ( .a(TIMEBOOST_net_237), .b(n_45897), .o(n_38371) );
in01s01 g740021 ( .a(n_40120), .o(n_40148) );
na02m04 TIMEBOOST_cell_8789 ( .a(TIMEBOOST_net_2881), .b(n_9365), .o(n_9526) );
no02s03 TIMEBOOST_cell_1248 ( .a(TIMEBOOST_net_238), .b(n_19026), .o(n_19272) );
no02s02 g740025 ( .a(n_40006), .b(FE_OCP_RBN6159_n_39816), .o(n_40154) );
oa22s01 g740026 ( .a(n_39784), .b(n_39782), .c(n_39824), .d(n_39783), .o(n_39848) );
in01s01 g740027 ( .a(n_39955), .o(n_39956) );
ao12f06 g740028 ( .a(n_39776), .b(n_39861), .c(n_39806), .o(n_39955) );
no02f08 g740029 ( .a(n_40038), .b(n_40004), .o(n_40080) );
no02f08 TIMEBOOST_cell_1302 ( .a(TIMEBOOST_net_265), .b(FE_RN_1289_0), .o(n_29143) );
oa22s01 g740031 ( .a(n_39899), .b(n_39829), .c(n_39898), .d(n_39830), .o(n_39986) );
in01s01 g740033 ( .a(n_39984), .o(n_39985) );
na02s01 g740034 ( .a(n_39866), .b(n_39846), .o(n_39984) );
no02s04 TIMEBOOST_cell_8563 ( .a(TIMEBOOST_net_2768), .b(n_38042), .o(n_38090) );
no02m08 g740036 ( .a(n_39845), .b(n_39872), .o(n_39873) );
no02s01 g740037 ( .a(n_39907), .b(n_39867), .o(n_39908) );
na02m08 TIMEBOOST_cell_5984 ( .a(TIMEBOOST_net_1843), .b(n_12376), .o(n_12464) );
in01s01 g740039 ( .a(n_40293), .o(n_40294) );
no02s02 g740040 ( .a(n_40254), .b(n_40047), .o(n_40293) );
in01s01 g740041 ( .a(n_40018), .o(n_40019) );
no02s01 g740042 ( .a(n_39983), .b(n_39982), .o(n_40018) );
na02s04 g740043 ( .a(n_39843), .b(n_39869), .o(n_39870) );
no02s02 g740044 ( .a(n_39865), .b(n_39921), .o(n_39922) );
in01s01 g740045 ( .a(n_40330), .o(n_40331) );
na02s01 g740046 ( .a(n_40292), .b(n_40219), .o(n_40330) );
no03m04 TIMEBOOST_cell_8292 ( .a(n_34625), .b(n_34624), .c(n_34971), .o(TIMEBOOST_net_2490) );
na02s03 g740048 ( .a(n_39918), .b(n_39953), .o(n_39954) );
in01s01 g740049 ( .a(n_40078), .o(n_40079) );
no02s01 g740050 ( .a(n_40043), .b(n_40015), .o(n_40078) );
no02s01 g740051 ( .a(n_40016), .b(n_40015), .o(n_40017) );
no03s20 TIMEBOOST_cell_5695 ( .a(n_32568), .b(n_32543), .c(FE_OCP_RBN7008_n_44962), .o(n_32630) );
in01s01 g740054 ( .a(n_40076), .o(n_40077) );
no02s01 g740055 ( .a(n_40042), .b(n_40041), .o(n_40076) );
na02s02 g740056 ( .a(n_39950), .b(n_39561), .o(n_39981) );
in01s01 g740058 ( .a(n_40145), .o(n_40146) );
no02s01 g740059 ( .a(n_40119), .b(n_40118), .o(n_40145) );
na02s01 TIMEBOOST_cell_1245 ( .a(n_37542), .b(n_37308), .o(TIMEBOOST_net_237) );
in01s01 g740062 ( .a(n_40143), .o(n_40144) );
no02s01 g740063 ( .a(n_40117), .b(n_40116), .o(n_40143) );
in01s01 g740064 ( .a(n_40114), .o(n_40115) );
na02s01 g740065 ( .a(n_40073), .b(n_40072), .o(n_40114) );
no03m06 TIMEBOOST_cell_8208 ( .a(n_18115), .b(n_18023), .c(TIMEBOOST_net_1422), .o(n_18164) );
in01s01 g740068 ( .a(n_40113), .o(n_40141) );
na02s06 g740069 ( .a(n_40071), .b(n_40036), .o(n_40113) );
in01s01 g740070 ( .a(n_40139), .o(n_40140) );
no02s01 g740071 ( .a(n_40112), .b(n_40111), .o(n_40139) );
no02s01 TIMEBOOST_cell_1247 ( .a(n_18866), .b(FE_OCPN1709_FE_OFN739_n_17093), .o(TIMEBOOST_net_238) );
no02s02 g740074 ( .a(n_40111), .b(n_40005), .o(n_40006) );
in01m01 g740075 ( .a(n_40137), .o(n_40138) );
no02s01 g740076 ( .a(n_40110), .b(n_40112), .o(n_40137) );
in01s01 g740077 ( .a(n_39919), .o(n_39920) );
na02s01 g740078 ( .a(n_39904), .b(n_39802), .o(n_39919) );
in01s01 g740079 ( .a(n_40328), .o(n_40329) );
na02s02 g740080 ( .a(n_40291), .b(n_40215), .o(n_40328) );
no02s01 g740081 ( .a(n_39998), .b(n_39940), .o(n_40039) );
in01s01 g740084 ( .a(n_40038), .o(n_40068) );
no03f08 TIMEBOOST_cell_7181 ( .a(n_41896), .b(n_41675), .c(n_41754), .o(n_41939) );
na02f06 g740086 ( .a(n_40003), .b(n_39941), .o(n_40004) );
no02s01 g740087 ( .a(n_40107), .b(n_40206), .o(n_40253) );
in01s01 g740089 ( .a(n_40136), .o(n_40189) );
no02m10 g740090 ( .a(n_40034), .b(n_40107), .o(n_40136) );
no02m10 g740091 ( .a(n_40066), .b(n_40032), .o(n_40067) );
no02m04 TIMEBOOST_cell_1301 ( .a(n_29034), .b(FE_RN_469_0), .o(TIMEBOOST_net_265) );
no02f04 g740093 ( .a(n_39801), .b(n_39773), .o(n_39927) );
in01s01 g740094 ( .a(n_40289), .o(n_40290) );
na02m01 g740095 ( .a(n_40187), .b(n_39924), .o(n_40289) );
in01s01 g740096 ( .a(n_40326), .o(n_40327) );
no02s01 g740097 ( .a(n_40220), .b(n_39921), .o(n_40326) );
in01s01 g740098 ( .a(n_40287), .o(n_40288) );
na02s01 g740099 ( .a(n_40186), .b(n_39953), .o(n_40287) );
in01s01 g740100 ( .a(n_40324), .o(n_40325) );
oa22s01 g740101 ( .a(FE_OCP_RBN6155_n_39816), .b(n_39508), .c(FE_OCP_RBN6161_n_39816), .d(n_39535), .o(n_40324) );
in01s01 g740102 ( .a(n_40285), .o(n_40286) );
na02s01 g740103 ( .a(n_40182), .b(n_40013), .o(n_40285) );
in01s01 g740104 ( .a(n_40283), .o(n_40284) );
na02s01 g740105 ( .a(n_40002), .b(n_40181), .o(n_40283) );
in01s01 g740106 ( .a(n_40281), .o(n_40282) );
na02s01 g740107 ( .a(n_40074), .b(n_40180), .o(n_40281) );
in01s01 g740108 ( .a(n_40279), .o(n_40280) );
na02s01 g740109 ( .a(n_40071), .b(n_40179), .o(n_40279) );
in01s01 g740110 ( .a(n_40277), .o(n_40278) );
na02s01 g740111 ( .a(n_40069), .b(n_40178), .o(n_40277) );
in01s01 g740112 ( .a(n_40249), .o(n_40250) );
na02m08 TIMEBOOST_cell_1250 ( .a(n_33622), .b(TIMEBOOST_net_239), .o(n_33677) );
oa12s01 g740114 ( .a(n_39799), .b(n_39798), .c(n_39797), .o(n_39847) );
in01s01 g740115 ( .a(n_40223), .o(n_40224) );
na02s01 g740116 ( .a(n_40188), .b(n_40106), .o(n_40223) );
in01s01 g740117 ( .a(n_40221), .o(n_40222) );
oa22s01 g740118 ( .a(FE_OCP_RBN6158_n_39816), .b(FE_OCP_RBN6811_n_39551), .c(FE_OCP_RBN6157_n_39816), .d(n_39551), .o(n_40221) );
in01s01 g740119 ( .a(n_40322), .o(n_40323) );
oa22s02 g740120 ( .a(FE_OCP_RBN6154_n_39816), .b(n_39800), .c(FE_OCP_RBN6157_n_39816), .d(n_39817), .o(n_40322) );
in01s01 g740121 ( .a(n_40320), .o(n_40321) );
no02s01 g740122 ( .a(n_40217), .b(n_39872), .o(n_40320) );
in01s01 g740123 ( .a(n_40318), .o(n_40319) );
oa22s01 g740124 ( .a(FE_OCP_RBN6152_n_39816), .b(n_39840), .c(FE_OCP_RBN6161_n_39816), .d(n_39460), .o(n_40318) );
in01s01 g740125 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_1_), .o(n_40684) );
in01s01 g740127 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_2_), .o(n_40667) );
in01s01 g740130 ( .a(n_39846), .o(n_39867) );
na02s06 g740131 ( .a(n_39816), .b(FE_OCPN1671_n_39371), .o(n_39846) );
in01s01 g740133 ( .a(n_39866), .o(n_39902) );
in01s01 g740136 ( .a(n_39802), .o(n_39820) );
na02m02 g740137 ( .a(n_39770), .b(n_39785), .o(n_39802) );
no02m02 g740138 ( .a(n_39781), .b(n_39800), .o(n_39801) );
in01s01 g740139 ( .a(n_39845), .o(n_39904) );
no02m08 g740140 ( .a(n_39816), .b(FE_OCP_DRV_N3518_n_39785), .o(n_39845) );
no02m06 g740141 ( .a(n_39816), .b(n_39334), .o(n_39872) );
no02s06 g740142 ( .a(n_39816), .b(n_39817), .o(n_39818) );
na02m04 g740143 ( .a(n_39781), .b(n_39844), .o(n_39924) );
na02s01 g740144 ( .a(FE_OCP_RBN6161_n_39816), .b(n_39459), .o(n_40187) );
in01s01 g740145 ( .a(n_39843), .o(n_40047) );
na02s04 g740146 ( .a(n_39816), .b(n_39864), .o(n_39843) );
no02s02 g740147 ( .a(n_39816), .b(n_39864), .o(n_39865) );
no02s02 g740148 ( .a(FE_OCP_RBN6161_n_39816), .b(n_39864), .o(n_40254) );
no02s02 g740149 ( .a(n_39816), .b(n_39506), .o(n_39921) );
no02s01 g740150 ( .a(FE_OCP_RBN6155_n_39816), .b(n_39869), .o(n_40220) );
no02s02 g740151 ( .a(n_39781), .b(n_39841), .o(n_39982) );
in01s01 g740152 ( .a(n_39918), .o(n_39983) );
na02s01 g740153 ( .a(n_39781), .b(n_39841), .o(n_39918) );
na02s01 g740154 ( .a(n_39781), .b(n_39562), .o(n_39953) );
na02s01 g740155 ( .a(FE_OCP_RBN6161_n_39816), .b(n_39905), .o(n_40186) );
in01s01 g740156 ( .a(n_40218), .o(n_40219) );
no02s01 g740157 ( .a(FE_OCP_RBN6161_n_39816), .b(n_40183), .o(n_40218) );
na02s01 g740158 ( .a(FE_OCP_RBN6161_n_39816), .b(n_40183), .o(n_40292) );
no02s02 g740159 ( .a(n_39812), .b(n_39900), .o(n_40015) );
in01s01 g740160 ( .a(n_39980), .o(n_40043) );
na02s06 g740161 ( .a(FE_OCP_RBN6155_n_39816), .b(n_39900), .o(n_39980) );
na02s01 g740162 ( .a(FE_OCP_RBN6161_n_39816), .b(n_46950), .o(n_40182) );
na02s01 g740163 ( .a(n_39812), .b(n_39548), .o(n_40013) );
in01s01 g740164 ( .a(n_39950), .o(n_40041) );
na02s01 g740165 ( .a(n_39816), .b(n_39917), .o(n_39950) );
no02m01 g740166 ( .a(n_39816), .b(n_39917), .o(n_40042) );
in01s01 g740167 ( .a(n_40001), .o(n_40002) );
no02s01 g740168 ( .a(n_39816), .b(n_39978), .o(n_40001) );
na02s01 g740169 ( .a(FE_OCP_RBN6161_n_39816), .b(n_39978), .o(n_40181) );
no02s01 g740170 ( .a(n_39812), .b(n_46948), .o(n_40118) );
in01s01 g740171 ( .a(n_40037), .o(n_40119) );
na02s02 g740172 ( .a(FE_OCP_RBN6154_n_39816), .b(n_46948), .o(n_40037) );
na02s02 g740173 ( .a(FE_OCP_RBN6154_n_39816), .b(n_39627), .o(n_40074) );
na02s01 g740174 ( .a(FE_OCP_RBN6157_n_39816), .b(n_40011), .o(n_40180) );
no02s03 g740175 ( .a(FE_OCP_RBN6154_n_39816), .b(n_39947), .o(n_40116) );
in01s01 g740176 ( .a(n_40036), .o(n_40117) );
na02s02 g740177 ( .a(FE_OCP_RBN6154_n_39816), .b(n_39947), .o(n_40036) );
na02s02 g740178 ( .a(FE_OCP_RBN6154_n_39816), .b(n_39580), .o(n_40071) );
na02s01 g740179 ( .a(FE_OCP_RBN6157_n_39816), .b(n_40009), .o(n_40179) );
in01s01 g740180 ( .a(n_39977), .o(n_40072) );
no02s01 g740181 ( .a(n_39812), .b(n_39945), .o(n_39977) );
na02s02 g740182 ( .a(FE_OCP_RBN6154_n_39816), .b(n_39945), .o(n_40073) );
na02s01 g740183 ( .a(FE_OCP_RBN6157_n_39816), .b(n_40007), .o(n_40178) );
na02s01 g740184 ( .a(FE_OCP_RBN6154_n_39816), .b(n_39553), .o(n_40069) );
no02m01 g740185 ( .a(FE_OCP_RBN6157_n_39816), .b(n_39531), .o(n_40112) );
no02s01 g740186 ( .a(n_39812), .b(FE_OCP_RBN3108_n_39531), .o(n_40111) );
na02s01 TIMEBOOST_cell_1249 ( .a(n_33184), .b(FE_OCPN1725_n_33136), .o(TIMEBOOST_net_239) );
no02s01 g740188 ( .a(FE_OCP_RBN6157_n_39816), .b(n_40005), .o(n_40110) );
na02s01 g740189 ( .a(n_39798), .b(n_39797), .o(n_39799) );
na02s01 g740190 ( .a(FE_OCP_RBN6157_n_39816), .b(n_39600), .o(n_40106) );
na02s01 g740191 ( .a(FE_OCP_RBN6159_n_39816), .b(n_39586), .o(n_40188) );
in01s01 g740192 ( .a(n_39814), .o(n_39815) );
na02s01 g740193 ( .a(n_39796), .b(n_39795), .o(n_39814) );
no02s01 g740194 ( .a(FE_OCP_RBN6152_n_39816), .b(n_39822), .o(n_40217) );
in01s01 g740195 ( .a(n_40214), .o(n_40215) );
no02s02 g740196 ( .a(FE_OCP_RBN6161_n_39816), .b(n_40177), .o(n_40214) );
na02s02 g740197 ( .a(FE_OCP_RBN6161_n_39816), .b(n_40177), .o(n_40291) );
no02m01 g740198 ( .a(n_40210), .b(n_40247), .o(n_40248) );
in01s01 g740199 ( .a(n_39907), .o(n_39862) );
in01s01 g740201 ( .a(n_39824), .o(n_39784) );
ao12f06 g740202 ( .a(n_39772), .b(n_39750), .c(n_39753), .o(n_39824) );
na02f08 g740203 ( .a(n_39812), .b(n_39461), .o(n_39925) );
in01s01 g740204 ( .a(n_40016), .o(n_39976) );
no02m01 g740205 ( .a(n_39812), .b(n_39536), .o(n_40016) );
na02s01 g740206 ( .a(n_39812), .b(n_39534), .o(n_39944) );
in01s01 g740208 ( .a(n_39975), .o(n_39998) );
na02f04 g740209 ( .a(n_39895), .b(n_39803), .o(n_39975) );
in01s01 g740210 ( .a(n_39898), .o(n_39899) );
in01s01 g740211 ( .a(n_39861), .o(n_39898) );
oa12f08 g740212 ( .a(n_39774), .b(n_39792), .c(n_39758), .o(n_39861) );
na02m06 g740213 ( .a(n_39838), .b(n_39803), .o(n_39897) );
na02s01 TIMEBOOST_cell_8681 ( .a(TIMEBOOST_net_2827), .b(FE_OCP_RBN4468_n_44267), .o(n_22338) );
no02m06 g740215 ( .a(n_39916), .b(n_39973), .o(n_39974) );
na02f06 g740216 ( .a(n_39892), .b(FE_OCP_RBN4430_n_39942), .o(n_40003) );
na02f06 g740217 ( .a(n_39890), .b(FE_OCP_RBN4430_n_39942), .o(n_39941) );
na02m08 g740218 ( .a(n_39996), .b(n_39938), .o(n_39997) );
in01s01 g740219 ( .a(n_40107), .o(n_40064) );
na02s01 TIMEBOOST_cell_3392 ( .a(n_36246), .b(n_36193), .o(TIMEBOOST_net_987) );
no02s06 g740221 ( .a(FE_OCP_RBN6853_n_39793), .b(n_39966), .o(n_40034) );
na03m10 g740222 ( .a(n_39967), .b(n_39995), .c(n_39994), .o(n_40066) );
no02m10 TIMEBOOST_cell_8504 ( .a(n_28385), .b(n_28006), .o(TIMEBOOST_net_2739) );
no02s06 TIMEBOOST_cell_1284 ( .a(TIMEBOOST_net_256), .b(n_7627), .o(n_7693) );
no02m02 TIMEBOOST_cell_8749 ( .a(TIMEBOOST_net_2861), .b(n_13943), .o(n_13940) );
no02f06 TIMEBOOST_cell_1299 ( .a(n_29232), .b(n_28739), .o(TIMEBOOST_net_264) );
no02s06 g740227 ( .a(n_40098), .b(FE_OCP_RBN3342_n_39942), .o(n_40251) );
oa22s01 g740228 ( .a(n_39788), .b(n_39804), .c(n_39789), .d(n_39805), .o(n_39896) );
in01s01 g740229 ( .a(n_39773), .o(n_39796) );
no02m02 g740230 ( .a(n_39764), .b(n_39763), .o(n_39773) );
na02m04 g740231 ( .a(n_39764), .b(n_39763), .o(n_39795) );
no02s01 g740232 ( .a(n_39772), .b(n_39754), .o(n_39798) );
in01s01 g740233 ( .a(n_39782), .o(n_39783) );
na02s01 g740234 ( .a(n_39771), .b(n_39752), .o(n_39782) );
no03s02 TIMEBOOST_cell_8634 ( .a(n_4352), .b(n_4148), .c(n_4147), .o(TIMEBOOST_net_2804) );
na02s06 g740236 ( .a(n_39811), .b(n_39859), .o(n_39860) );
na02m04 g740237 ( .a(n_39807), .b(n_39808), .o(n_39838) );
in01s01 g740238 ( .a(n_39971), .o(n_39972) );
no02s01 g740239 ( .a(n_39973), .b(n_39940), .o(n_39971) );
in01s01 g740240 ( .a(n_40316), .o(n_40317) );
no02s01 g740241 ( .a(n_40274), .b(n_40152), .o(n_40316) );
na02m08 g740242 ( .a(n_39854), .b(n_39853), .o(n_39893) );
na02s02 g740243 ( .a(n_39915), .b(n_39914), .o(n_39916) );
na02f04 g740244 ( .a(n_39852), .b(n_39891), .o(n_39892) );
no02s06 g740245 ( .a(n_39882), .b(n_39939), .o(n_39996) );
in01s01 g740246 ( .a(n_40314), .o(n_40315) );
no02s01 g740247 ( .a(n_40273), .b(n_40193), .o(n_40314) );
na02f06 g740248 ( .a(n_39851), .b(n_39889), .o(n_39890) );
na02s01 TIMEBOOST_cell_1270 ( .a(TIMEBOOST_net_249), .b(n_2144), .o(n_2177) );
in01s01 g740250 ( .a(n_40365), .o(n_40366) );
na02s01 g740251 ( .a(n_40243), .b(n_40313), .o(n_40365) );
no02f10 TIMEBOOST_cell_3391 ( .a(n_36416), .b(TIMEBOOST_net_986), .o(n_36474) );
in01s01 g740253 ( .a(n_40311), .o(n_40312) );
na02s01 g740254 ( .a(n_40207), .b(n_39994), .o(n_40311) );
na02s01 g740255 ( .a(n_39994), .b(n_39967), .o(n_39968) );
no02f06 TIMEBOOST_cell_6326 ( .a(TIMEBOOST_net_2014), .b(FE_RN_1274_0), .o(n_26753) );
in01s01 g740257 ( .a(n_40061), .o(n_40062) );
no02s01 g740258 ( .a(n_40032), .b(n_40033), .o(n_40061) );
no03m06 TIMEBOOST_cell_8439 ( .a(n_25793), .b(n_25762), .c(n_25829), .o(n_25898) );
in01s01 g740260 ( .a(n_40102), .o(n_40103) );
no02s01 g740261 ( .a(n_40060), .b(n_40059), .o(n_40102) );
no02s02 TIMEBOOST_cell_1283 ( .a(n_7612), .b(n_7611), .o(TIMEBOOST_net_256) );
no02s06 g740263 ( .a(n_40057), .b(n_40060), .o(n_40058) );
in01s01 g740264 ( .a(n_40173), .o(n_40174) );
no02s01 g740265 ( .a(n_40133), .b(n_40132), .o(n_40173) );
in01s01 g740266 ( .a(n_40171), .o(n_40172) );
no02s01 g740267 ( .a(n_40131), .b(n_40130), .o(n_40171) );
na02m01 g740268 ( .a(n_40100), .b(n_40054), .o(n_40101) );
no02m02 TIMEBOOST_cell_8748 ( .a(n_13939), .b(n_13821), .o(TIMEBOOST_net_2861) );
in01s01 TIMEBOOST_cell_4568 ( .a(TIMEBOOST_net_1375), .o(TIMEBOOST_net_1374) );
in01s01 g740272 ( .a(n_40212), .o(n_40213) );
na02m01 g740273 ( .a(n_40051), .b(n_40170), .o(n_40212) );
in01s01 g740274 ( .a(n_40210), .o(n_40211) );
na02s02 g740275 ( .a(n_40169), .b(n_40170), .o(n_40210) );
no02s06 g740276 ( .a(n_40097), .b(FE_OCP_RBN6835_n_39577), .o(n_40098) );
na02s01 g740277 ( .a(n_39857), .b(n_40045), .o(n_39858) );
in01s01 g740278 ( .a(n_40363), .o(n_40364) );
na02s01 g740279 ( .a(n_40310), .b(n_39807), .o(n_40363) );
in01s01 g740280 ( .a(n_40361), .o(n_40362) );
na02s01 g740281 ( .a(n_40239), .b(n_40309), .o(n_40361) );
in01f10 g740317 ( .a(n_39816), .o(n_39812) );
in01f10 g740318 ( .a(n_39781), .o(n_39816) );
in01f08 g740321 ( .a(n_39770), .o(n_39781) );
no02f06 g740322 ( .a(n_39733), .b(n_39742), .o(n_39770) );
oa12s01 g740323 ( .a(n_39762), .b(n_39761), .c(n_39760), .o(n_39779) );
in01s01 g740324 ( .a(n_40396), .o(n_40397) );
na02s01 g740325 ( .a(n_40270), .b(n_39915), .o(n_40396) );
in01s01 g740326 ( .a(n_40359), .o(n_40360) );
no02s01 g740327 ( .a(n_40246), .b(n_39939), .o(n_40359) );
in01s01 g740328 ( .a(n_40357), .o(n_40358) );
no02s01 g740329 ( .a(n_40245), .b(n_39937), .o(n_40357) );
in01s01 g740330 ( .a(n_40394), .o(n_40395) );
oa22s01 g740331 ( .a(FE_OCP_RBN3344_n_39942), .b(n_39969), .c(FE_OCP_RBN6853_n_39793), .d(n_39519), .o(n_40394) );
in01s01 g740332 ( .a(n_40392), .o(n_40393) );
na02s01 g740333 ( .a(n_39995), .b(n_40269), .o(n_40392) );
in01s01 g740334 ( .a(n_40355), .o(n_40356) );
no02s01 g740335 ( .a(n_40308), .b(n_40241), .o(n_40355) );
in01s01 g740336 ( .a(n_40407), .o(n_40408) );
no02s01 g740337 ( .a(n_40057), .b(n_40303), .o(n_40407) );
in01s01 g740338 ( .a(n_40390), .o(n_40391) );
na02s01 g740339 ( .a(n_40100), .b(n_40267), .o(n_40390) );
in01s01 g740340 ( .a(n_40353), .o(n_40354) );
no02s01 g740341 ( .a(n_40240), .b(n_40128), .o(n_40353) );
na02s01 g740343 ( .a(n_40169), .b(n_40205), .o(n_40306) );
oa22s01 g740344 ( .a(n_39790), .b(n_39778), .c(n_39791), .d(n_39755), .o(n_39855) );
in01s01 g740345 ( .a(n_40271), .o(n_40272) );
na02s04 TIMEBOOST_cell_1292 ( .a(TIMEBOOST_net_260), .b(FE_RN_519_0), .o(FE_RN_1032_0) );
in01s01 g740347 ( .a(n_40304), .o(n_40305) );
na02s02 g740348 ( .a(n_40204), .b(n_40166), .o(n_40304) );
in01s01 g740349 ( .a(n_40388), .o(n_40389) );
na02s01 g740350 ( .a(n_40266), .b(n_39859), .o(n_40388) );
in01s01 g740351 ( .a(n_40386), .o(n_40387) );
oa22s01 g740352 ( .a(FE_OCP_RBN3345_n_39942), .b(n_39470), .c(FE_OCP_RBN3340_n_39942), .d(n_39894), .o(n_40386) );
no02f06 g740354 ( .a(n_39729), .b(FE_OCP_RBN3284_n_39674), .o(n_39742) );
na02s01 TIMEBOOST_cell_4071 ( .a(n_45072), .b(FE_OCPN6925_n_45081), .o(TIMEBOOST_net_1126) );
na02s04 g740356 ( .a(n_39739), .b(n_39738), .o(n_39771) );
in01s01 g740357 ( .a(n_39753), .o(n_39754) );
na02f04 g740358 ( .a(n_39741), .b(n_39740), .o(n_39753) );
no02f04 g740359 ( .a(n_39741), .b(n_39740), .o(n_39772) );
in01s01 g740360 ( .a(n_39751), .o(n_39752) );
no02f04 g740361 ( .a(n_39739), .b(n_39738), .o(n_39751) );
na02s02 g740362 ( .a(n_39761), .b(n_39760), .o(n_39762) );
no02f10 TIMEBOOST_cell_3379 ( .a(n_31813), .b(TIMEBOOST_net_980), .o(n_31908) );
na02s01 g740364 ( .a(FE_OCP_RBN3344_n_39942), .b(n_40202), .o(n_40309) );
na02s02 g740365 ( .a(FE_OCP_RBN6106_n_39793), .b(n_39810), .o(n_39811) );
na02s01 g740366 ( .a(FE_OCP_RBN3339_n_39942), .b(n_39810), .o(n_40310) );
na02m02 g740367 ( .a(FE_OCP_RBN6106_n_39793), .b(n_39808), .o(n_39859) );
na02s03 g740368 ( .a(n_39793), .b(n_39084), .o(n_39857) );
na02s06 g740369 ( .a(FE_OCP_RBN6105_n_39793), .b(n_39085), .o(n_40045) );
in01s01 g740371 ( .a(n_39807), .o(n_39833) );
na02s02 g740372 ( .a(n_39793), .b(n_39112), .o(n_39807) );
in01s01 g740373 ( .a(n_39854), .o(n_39940) );
na02s06 g740374 ( .a(n_39803), .b(n_39832), .o(n_39854) );
no02s08 g740375 ( .a(FE_OCP_RBN4430_n_39942), .b(n_39832), .o(n_39973) );
na02s01 g740376 ( .a(FE_OCP_RBN3345_n_39942), .b(n_39465), .o(n_40270) );
na02s02 g740377 ( .a(FE_OCP_RBN6106_n_39793), .b(n_39853), .o(n_39915) );
in01s01 g740378 ( .a(n_39852), .o(n_40152) );
na02f04 g740379 ( .a(n_39803), .b(n_39881), .o(n_39852) );
no02s02 g740380 ( .a(n_39803), .b(n_39881), .o(n_39882) );
no02s01 g740381 ( .a(FE_OCP_RBN3344_n_39942), .b(n_39881), .o(n_40274) );
no02s01 g740382 ( .a(FE_OCP_RBN3340_n_39942), .b(n_39891), .o(n_40246) );
no02s03 g740383 ( .a(n_39803), .b(n_39513), .o(n_39939) );
in01s01 g740384 ( .a(n_39851), .o(n_40193) );
na02m04 g740385 ( .a(n_39803), .b(n_39878), .o(n_39851) );
na02m04 TIMEBOOST_cell_8532 ( .a(TIMEBOOST_net_1464), .b(n_41740), .o(TIMEBOOST_net_2753) );
no02s01 g740387 ( .a(FE_OCP_RBN3344_n_39942), .b(n_39878), .o(n_40273) );
no02s01 g740388 ( .a(FE_OCP_RBN3340_n_39942), .b(n_39889), .o(n_40245) );
no02s02 g740389 ( .a(n_39803), .b(n_39520), .o(n_39937) );
in01s01 g740390 ( .a(n_39934), .o(n_40313) );
no02s06 g740391 ( .a(FE_OCP_RBN6853_n_39793), .b(n_39488), .o(n_39934) );
in01s01 g740392 ( .a(n_40242), .o(n_40243) );
no02s01 g740393 ( .a(FE_OCP_RBN3344_n_39942), .b(n_39538), .o(n_40242) );
in01s01 g740394 ( .a(n_40206), .o(n_40207) );
no02s01 g740396 ( .a(FE_OCP_RBN6853_n_39793), .b(n_39910), .o(n_40206) );
na02s06 g740397 ( .a(FE_OCP_RBN6108_n_39793), .b(n_39910), .o(n_39994) );
na02s01 g740398 ( .a(FE_OCP_RBN4429_n_39942), .b(n_39965), .o(n_40269) );
na02s06 g740399 ( .a(FE_OCP_RBN6853_n_39793), .b(n_46949), .o(n_39995) );
in01s01 g740400 ( .a(n_39964), .o(n_40033) );
na02s06 g740401 ( .a(FE_OCP_RBN4429_n_39942), .b(n_39932), .o(n_39964) );
no02s03 g740402 ( .a(FE_OCP_RBN4431_n_39942), .b(n_39932), .o(n_40032) );
no02s01 g740403 ( .a(FE_OCP_RBN3333_n_39942), .b(n_39992), .o(n_40241) );
no02s02 g740404 ( .a(FE_OCP_RBN4431_n_39942), .b(n_39602), .o(n_40308) );
no02s06 g740405 ( .a(FE_OCP_RBN3333_n_39942), .b(n_39543), .o(n_40059) );
no02s02 g740406 ( .a(FE_OCP_RBN4431_n_39942), .b(n_39544), .o(n_40060) );
no02s01 g740407 ( .a(FE_OCP_RBN3333_n_39942), .b(n_39605), .o(n_40303) );
no02s02 g740408 ( .a(FE_OCP_RBN4431_n_39942), .b(n_39989), .o(n_40057) );
in01s01 g740409 ( .a(n_40030), .o(n_40133) );
na02s02 g740410 ( .a(FE_OCP_RBN4431_n_39942), .b(n_39581), .o(n_40030) );
in01s01 g740411 ( .a(n_40054), .o(n_40132) );
na02s01 g740412 ( .a(FE_OCP_RBN3333_n_39942), .b(n_39582), .o(n_40054) );
na02s01 g740413 ( .a(FE_OCP_RBN4431_n_39942), .b(n_39612), .o(n_40267) );
na02s01 g740414 ( .a(FE_OCP_RBN3333_n_39942), .b(n_40028), .o(n_40100) );
no02s06 g740415 ( .a(FE_OCP_RBN3333_n_39942), .b(n_39495), .o(n_40131) );
no02s01 g740416 ( .a(FE_OCP_RBN4431_n_39942), .b(n_39496), .o(n_40130) );
no02s01 g740417 ( .a(FE_OCP_RBN3333_n_39942), .b(n_39555), .o(n_40240) );
no02s01 g740418 ( .a(FE_OCP_RBN3337_n_39942), .b(FE_OCP_RBN6824_n_39542), .o(n_40128) );
in01s01 g740419 ( .a(n_40097), .o(n_40051) );
no02s03 g740420 ( .a(FE_OCP_RBN3333_n_39942), .b(FE_OCP_RBN4382_n_39523), .o(n_40097) );
na02s02 g740421 ( .a(FE_OCP_RBN3333_n_39942), .b(FE_OCP_RBN4382_n_39523), .o(n_40170) );
na02s01 g740422 ( .a(FE_OCP_RBN3337_n_39942), .b(FE_OCP_RBN6835_n_39577), .o(n_40205) );
na02s01 g740423 ( .a(FE_OCP_RBN3341_n_39942), .b(n_39577), .o(n_40169) );
na02m02 TIMEBOOST_cell_1291 ( .a(n_18947), .b(n_17815), .o(TIMEBOOST_net_260) );
no02s02 g740425 ( .a(FE_OCP_RBN3337_n_39942), .b(FE_OCP_RBN3226_n_39575), .o(n_40247) );
na02s01 g740426 ( .a(FE_OCP_RBN3337_n_39942), .b(n_39559), .o(n_40204) );
na02s01 g740427 ( .a(FE_OCP_RBN3341_n_39942), .b(n_39558), .o(n_40166) );
in01s01 g740428 ( .a(n_39829), .o(n_39830) );
na02s01 g740429 ( .a(n_39777), .b(n_39806), .o(n_39829) );
na02s01 g740430 ( .a(FE_OCP_RBN3345_n_39942), .b(n_39427), .o(n_40266) );
in01s01 g740431 ( .a(n_40238), .o(n_40239) );
no02s01 g740432 ( .a(FE_OCP_RBN3344_n_39942), .b(n_40202), .o(n_40238) );
in01s01 g740434 ( .a(n_39750), .o(n_39797) );
na02s02 g740436 ( .a(FE_OCP_RBN6106_n_39793), .b(n_39471), .o(n_39914) );
in01s01 g740437 ( .a(n_39804), .o(n_39805) );
in01s01 g740438 ( .a(n_39792), .o(n_39804) );
ao12f08 g740439 ( .a(n_39756), .b(n_39778), .c(n_39775), .o(n_39792) );
in01s01 g740440 ( .a(n_39967), .o(n_39931) );
na02s08 g740441 ( .a(FE_OCP_RBN6108_n_39793), .b(n_39539), .o(n_39967) );
in01s01 g740442 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_0_), .o(n_39737) );
na02f06 g740444 ( .a(n_39727), .b(n_39668), .o(n_39729) );
no02f02 TIMEBOOST_cell_8604 ( .a(n_20418), .b(n_45060), .o(TIMEBOOST_net_2789) );
na02s03 g740446 ( .a(n_39727), .b(n_39674), .o(n_39728) );
no02s01 TIMEBOOST_cell_5539 ( .a(TIMEBOOST_net_1717), .b(n_43383), .o(n_43467) );
no02s01 g740449 ( .a(n_39718), .b(n_39725), .o(n_39761) );
na02m03 g740450 ( .a(n_39769), .b(n_39768), .o(n_39806) );
in01s01 g740451 ( .a(n_39776), .o(n_39777) );
no02s03 g740452 ( .a(n_39769), .b(n_39768), .o(n_39776) );
in01s01 g740453 ( .a(n_39790), .o(n_39791) );
na02s01 g740454 ( .a(n_39757), .b(n_39775), .o(n_39790) );
in01s01 g740455 ( .a(n_39788), .o(n_39789) );
na02s01 g740456 ( .a(n_39774), .b(n_39759), .o(n_39788) );
no02s03 TIMEBOOST_cell_5607 ( .a(TIMEBOOST_net_1751), .b(n_31764), .o(n_31833) );
na02f04 g740458 ( .a(n_39701), .b(n_39710), .o(n_39741) );
in01f08 g740493 ( .a(FE_OCP_RBN6106_n_39793), .o(n_39803) );
na02f08 g740496 ( .a(n_39749), .b(n_39736), .o(n_39793) );
oa12s01 g740497 ( .a(n_39767), .b(n_39766), .c(n_39765), .o(n_39786) );
no02f02 g740498 ( .a(n_39711), .b(FE_OCP_RBN3329_n_39685), .o(n_39712) );
na02s06 TIMEBOOST_cell_8622 ( .a(FE_OFN4799_n_44498), .b(n_10978), .o(TIMEBOOST_net_2798) );
oa12s06 g740501 ( .a(n_39735), .b(n_39734), .c(FE_OCP_RBN3177_n_39640), .o(n_39736) );
na02m06 g740502 ( .a(n_39672), .b(n_39702), .o(n_39719) );
no02m08 g740503 ( .a(n_39711), .b(n_39655), .o(n_39727) );
na02m02 g740504 ( .a(n_39683), .b(n_39690), .o(n_39701) );
na02f02 g740505 ( .a(n_39684), .b(n_39677), .o(n_39710) );
in01s01 g740506 ( .a(n_39717), .o(n_39718) );
na02f04 g740507 ( .a(n_39698), .b(n_38786), .o(n_39717) );
in01s01 g740508 ( .a(n_39724), .o(n_39725) );
na02m06 g740509 ( .a(n_39699), .b(n_38787), .o(n_39724) );
in01s01 g740510 ( .a(n_39758), .o(n_39759) );
no02m06 g740511 ( .a(n_39746), .b(n_39745), .o(n_39758) );
na02m08 g740512 ( .a(n_39748), .b(FE_OCPN3582_n_39747), .o(n_39775) );
in01s01 g740513 ( .a(n_39756), .o(n_39757) );
no02f06 g740514 ( .a(n_39748), .b(FE_OCPN3582_n_39747), .o(n_39756) );
na02f04 g740515 ( .a(n_39746), .b(n_39745), .o(n_39774) );
na02s01 g740516 ( .a(n_39766), .b(n_39765), .o(n_39767) );
oa12s01 g740517 ( .a(n_39689), .b(n_39676), .c(n_39675), .o(n_39716) );
in01s01 g740518 ( .a(n_39778), .o(n_39755) );
na02f08 g740519 ( .a(n_39732), .b(n_39730), .o(n_39778) );
ao22m04 g740520 ( .a(n_39734), .b(n_39735), .c(n_39744), .d(n_39743), .o(n_39769) );
na02m08 g740522 ( .a(n_39690), .b(n_39656), .o(n_39711) );
no02s06 g740523 ( .a(n_39665), .b(n_39677), .o(n_39702) );
in01s01 g740525 ( .a(n_39689), .o(n_39760) );
na02m04 g740526 ( .a(n_39676), .b(n_39675), .o(n_39689) );
na02f06 g740527 ( .a(n_39722), .b(n_39695), .o(n_39732) );
no02s01 g740528 ( .a(n_39731), .b(n_39723), .o(n_39766) );
na02f08 g740532 ( .a(n_39668), .b(n_45530), .o(n_39674) );
na02f04 g740534 ( .a(n_39672), .b(n_39654), .o(n_39685) );
in01f02 g740535 ( .a(n_39683), .o(n_39684) );
na02f04 g740536 ( .a(n_39656), .b(n_45514), .o(n_39683) );
in01m02 g740537 ( .a(n_39698), .o(n_39699) );
na02m08 TIMEBOOST_cell_7987 ( .a(TIMEBOOST_net_2624), .b(n_30904), .o(n_31018) );
no02s02 TIMEBOOST_cell_6966 ( .a(TIMEBOOST_net_2241), .b(n_3738), .o(TIMEBOOST_net_1909) );
no02s02 TIMEBOOST_cell_4477 ( .a(n_10711), .b(n_10391), .o(TIMEBOOST_net_1329) );
no02s06 TIMEBOOST_cell_3387 ( .a(TIMEBOOST_net_984), .b(n_40374), .o(n_40373) );
na02f04 g740542 ( .a(n_39644), .b(n_39647), .o(n_39667) );
no02s02 TIMEBOOST_cell_6965 ( .a(n_2989), .b(n_3857), .o(TIMEBOOST_net_2241) );
na02f04 g740544 ( .a(FE_OCP_RBN3248_n_39697), .b(n_39693), .o(n_39714) );
na02m06 g740545 ( .a(n_39657), .b(n_39616), .o(n_39677) );
no02m08 g740546 ( .a(n_39621), .b(n_39647), .o(n_39690) );
na02m10 g740547 ( .a(n_39662), .b(FE_OCP_RBN3249_n_39697), .o(n_39734) );
no02s06 g740548 ( .a(n_39697), .b(FE_OCP_RBN3207_n_39662), .o(n_39744) );
no02f06 g740549 ( .a(n_39691), .b(n_45738), .o(n_39709) );
no02m02 TIMEBOOST_cell_5482 ( .a(n_15987), .b(n_15845), .o(TIMEBOOST_net_1689) );
in01s04 g740552 ( .a(n_39656), .o(n_39665) );
in01s06 g740554 ( .a(n_39672), .o(n_39655) );
na02m08 g740555 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n_39629), .o(n_39672) );
in01s02 g740557 ( .a(n_39668), .o(n_39645) );
na02f04 g740559 ( .a(FE_OCP_RBN4398_n_39629), .b(FE_RN_1873_0), .o(n_39654) );
in01s01 g740561 ( .a(n_39722), .o(n_39723) );
na02f04 g740562 ( .a(n_39704), .b(n_38794), .o(n_39722) );
in01s01 g740563 ( .a(n_39730), .o(n_39731) );
na02m06 g740564 ( .a(n_38795), .b(n_39705), .o(n_39730) );
ao22s02 g740565 ( .a(n_39619), .b(n_45840), .c(n_39614), .d(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39676) );
oa12s01 g740566 ( .a(n_39681), .b(n_39680), .c(n_39679), .o(n_39708) );
na02m10 g740570 ( .a(n_39678), .b(n_45740), .o(n_39697) );
na02f08 g740571 ( .a(n_39619), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39657) );
no02m06 g740572 ( .a(n_39614), .b(n_45840), .o(n_39647) );
na02s01 g740573 ( .a(n_39680), .b(n_39679), .o(n_39681) );
in01s01 g740574 ( .a(n_39695), .o(n_39765) );
no02m04 g740575 ( .a(n_39680), .b(n_38712), .o(n_39695) );
in01f02 g740576 ( .a(n_39643), .o(n_39644) );
na02s04 TIMEBOOST_cell_5637 ( .a(TIMEBOOST_net_1766), .b(n_27621), .o(n_27693) );
in01s02 g740578 ( .a(n_39693), .o(n_39694) );
na02f06 g740579 ( .a(n_39662), .b(n_39661), .o(n_39693) );
in01f04 g740580 ( .a(n_39691), .o(n_39692) );
no02s01 TIMEBOOST_cell_4429 ( .a(FE_OCPN1763_n_30708), .b(FE_OCP_DRV_N7081_n_27130), .o(TIMEBOOST_net_1305) );
na02s08 TIMEBOOST_cell_1006 ( .a(n_37270), .b(TIMEBOOST_net_117), .o(n_37277) );
in01m02 g740588 ( .a(n_39704), .o(n_39705) );
no02s01 TIMEBOOST_cell_4449 ( .a(n_4556), .b(n_4606), .o(TIMEBOOST_net_1315) );
no02s04 TIMEBOOST_cell_4448 ( .a(TIMEBOOST_net_1314), .b(FE_OCP_RBN3156_n_4925), .o(n_5163) );
no02m02 g740591 ( .a(n_39648), .b(n_39652), .o(n_39664) );
no02m08 g740594 ( .a(FE_OCP_RBN6836_n_39577), .b(n_45840), .o(n_39607) );
no02f06 g740595 ( .a(n_39577), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39596) );
in01s04 g740597 ( .a(n_39616), .o(n_39621) );
na02m08 g740598 ( .a(n_39592), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39616) );
na03s08 TIMEBOOST_cell_1005 ( .a(n_37271), .b(n_37252), .c(n_37112), .o(TIMEBOOST_net_117) );
na02s02 TIMEBOOST_cell_3343 ( .a(TIMEBOOST_net_962), .b(n_5880), .o(n_5971) );
no02m08 g740601 ( .a(n_39558), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39594) );
no02m06 g740602 ( .a(n_39559), .b(n_45840), .o(n_39579) );
na02s04 TIMEBOOST_cell_5553 ( .a(TIMEBOOST_net_1724), .b(n_6207), .o(n_6301) );
na02f08 g740606 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n_39635), .o(n_39662) );
na02m08 g740607 ( .a(n_39633), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39678) );
na02f04 g740608 ( .a(n_39636), .b(FE_RN_1873_0), .o(n_39661) );
na02s02 TIMEBOOST_cell_4428 ( .a(TIMEBOOST_net_1304), .b(n_36125), .o(n_36228) );
na02s04 g740610 ( .a(n_39640), .b(n_39639), .o(n_39743) );
no02m02 g740611 ( .a(n_39638), .b(FE_OCP_RBN3176_n_39640), .o(n_39735) );
in01f04 g740613 ( .a(n_39614), .o(n_39619) );
na02f08 g740615 ( .a(n_39578), .b(n_39560), .o(n_39614) );
oa22s02 g740616 ( .a(n_39625), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .c(n_39617), .d(FE_RN_1873_0), .o(n_39680) );
na02f06 g740617 ( .a(FE_OCP_RBN6825_n_39542), .b(n_45840), .o(n_39578) );
na02m04 g740618 ( .a(n_39542), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39560) );
in01s02 g740619 ( .a(n_39652), .o(n_39642) );
na02f08 g740620 ( .a(n_39617), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39652) );
na02f08 g740624 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n_39628), .o(n_39640) );
in01m02 g740625 ( .a(n_39638), .o(n_39639) );
no02s04 g740626 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n_39628), .o(n_39638) );
no02s06 TIMEBOOST_cell_6299 ( .a(n_35659), .b(FE_OCPN950_n_44180), .o(TIMEBOOST_net_2001) );
in01f02 g740629 ( .a(n_39592), .o(n_39593) );
in01f02 g740631 ( .a(n_39635), .o(n_39636) );
no02f10 TIMEBOOST_cell_822 ( .a(TIMEBOOST_net_25), .b(n_32595), .o(n_32641) );
in01f02 g740633 ( .a(n_39633), .o(n_39634) );
na02s06 TIMEBOOST_cell_7454 ( .a(FE_OCP_RBN5016_n_12026), .b(FE_RN_231_0), .o(TIMEBOOST_net_2358) );
in01s01 g740635 ( .a(n_39989), .o(n_39605) );
na02s02 g740636 ( .a(n_39556), .b(n_39545), .o(n_39989) );
in01s01 g740637 ( .a(n_40028), .o(n_39612) );
no02s02 g740638 ( .a(n_39557), .b(n_39571), .o(n_40028) );
no02s02 TIMEBOOST_cell_992 ( .a(TIMEBOOST_net_110), .b(n_37389), .o(n_37480) );
in01s01 g740643 ( .a(FE_OCP_RBN3226_n_39575), .o(n_39590) );
no02f06 TIMEBOOST_cell_7094 ( .a(TIMEBOOST_net_2305), .b(TIMEBOOST_net_474), .o(n_20501) );
in01s03 g740649 ( .a(n_39559), .o(n_39558) );
no02s06 TIMEBOOST_cell_3361 ( .a(TIMEBOOST_net_971), .b(n_32280), .o(n_32364) );
na02f02 TIMEBOOST_cell_6251 ( .a(n_4447), .b(n_4488), .o(TIMEBOOST_net_1977) );
na03m08 TIMEBOOST_cell_8307 ( .a(n_24476), .b(FE_OCP_RBN5706_n_24451), .c(FE_OCPN1916_n_22111), .o(n_24623) );
no02s02 TIMEBOOST_cell_4385 ( .a(n_4838), .b(n_4423), .o(TIMEBOOST_net_1283) );
na02f08 g740655 ( .a(n_39597), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39637) );
no02f08 TIMEBOOST_cell_5383 ( .a(TIMEBOOST_net_1639), .b(n_16125), .o(n_16328) );
no02s01 g740657 ( .a(n_39524), .b(n_39529), .o(n_39571) );
no02s01 g740658 ( .a(n_39525), .b(n_39528), .o(n_39557) );
no02m04 g740659 ( .a(n_39480), .b(n_39249), .o(n_39527) );
no02f08 TIMEBOOST_cell_8830 ( .a(n_25730), .b(FE_OFN747_n_22641), .o(TIMEBOOST_net_2902) );
no02f08 g740661 ( .a(n_39482), .b(n_39208), .o(n_39526) );
no02s01 TIMEBOOST_cell_991 ( .a(n_37205), .b(n_37254), .o(TIMEBOOST_net_110) );
na02s01 g740663 ( .a(n_39475), .b(n_39502), .o(n_39545) );
na02s01 g740664 ( .a(n_39476), .b(n_39503), .o(n_39556) );
in01s01 g740665 ( .a(n_40011), .o(n_39627) );
na02s01 g740666 ( .a(n_39587), .b(n_39601), .o(n_40011) );
in01m01 g740668 ( .a(n_39617), .o(n_39625) );
no02m08 TIMEBOOST_cell_998 ( .a(TIMEBOOST_net_113), .b(n_40834), .o(n_40896) );
no02s04 TIMEBOOST_cell_5092 ( .a(n_19270), .b(n_18032), .o(TIMEBOOST_net_1494) );
in01s01 g740671 ( .a(n_39992), .o(n_39602) );
no02m01 g740672 ( .a(n_39554), .b(n_39540), .o(n_39992) );
in01s01 g740673 ( .a(n_39543), .o(n_39544) );
ao12s01 g740674 ( .a(n_39485), .b(n_39484), .c(n_39483), .o(n_39543) );
in01s01 g740675 ( .a(FE_OCP_RBN6824_n_39542), .o(n_39555) );
na02s01 TIMEBOOST_cell_5157 ( .a(TIMEBOOST_net_1526), .b(n_15578), .o(n_15639) );
no02f08 g740680 ( .a(n_39552), .b(FE_RN_1873_0), .o(n_39589) );
no02s06 TIMEBOOST_cell_8686 ( .a(FE_OCPN1711_n_45073), .b(n_21345), .o(TIMEBOOST_net_2830) );
na02s01 TIMEBOOST_cell_7807 ( .a(TIMEBOOST_net_2534), .b(n_16384), .o(n_16262) );
na02s01 g740683 ( .a(n_39566), .b(n_39454), .o(n_39587) );
na02s01 g740684 ( .a(n_39567), .b(n_39453), .o(n_39601) );
no02s01 g740685 ( .a(n_39473), .b(n_39501), .o(n_39554) );
no02s02 g740686 ( .a(n_39474), .b(n_39500), .o(n_39540) );
no02s01 g740687 ( .a(n_39484), .b(n_39483), .o(n_39485) );
na02s01 g740688 ( .a(n_39969), .b(n_39538), .o(n_39539) );
in01s01 g740689 ( .a(n_39524), .o(n_39525) );
ao12s01 g740690 ( .a(n_39421), .b(n_39497), .c(n_39487), .o(n_39524) );
in01m04 g740691 ( .a(n_39481), .o(n_39482) );
ao12f06 g740692 ( .a(FE_OCP_RBN5966_n_39098), .b(n_39450), .c(FE_OCP_RBN5965_n_39097), .o(n_39481) );
in01m02 g740693 ( .a(n_39479), .o(n_39480) );
oa12m04 g740694 ( .a(n_39210), .b(n_39450), .c(n_39155), .o(n_39479) );
in01m04 g740695 ( .a(n_39477), .o(n_39478) );
oa12m08 g740696 ( .a(n_39335), .b(n_39386), .c(n_39211), .o(n_39477) );
in01s01 g740697 ( .a(n_39475), .o(n_39476) );
oa12s01 g740698 ( .a(n_39079), .b(n_39414), .c(n_38987), .o(n_39475) );
in01f04 g740701 ( .a(n_39586), .o(n_39600) );
in01s01 g740704 ( .a(n_40005), .o(n_39599) );
in01s01 g740705 ( .a(n_39584), .o(n_40005) );
in01m02 g740708 ( .a(n_39597), .o(n_39598) );
ao22f06 g740709 ( .a(FE_OCP_RBN3107_n_39531), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .c(n_39531), .d(n_45840), .o(n_39597) );
in01s01 g740710 ( .a(n_46949), .o(n_39965) );
in01s01 g740712 ( .a(n_39581), .o(n_39582) );
oa22s01 g740713 ( .a(n_39497), .b(n_39504), .c(n_39386), .d(n_39505), .o(n_39581) );
in01s01 g740714 ( .a(n_39495), .o(n_39496) );
ao12s01 g740715 ( .a(n_39417), .b(n_39416), .c(n_39415), .o(n_39495) );
no02s01 g740721 ( .a(n_39416), .b(n_39415), .o(n_39417) );
no02s01 g740723 ( .a(n_39408), .b(n_39455), .o(n_39494) );
na02s01 g740724 ( .a(n_39414), .b(n_38983), .o(n_39484) );
in01s01 g740725 ( .a(n_39566), .o(n_39567) );
ao12s01 g740726 ( .a(n_39043), .b(n_39532), .c(n_38988), .o(n_39566) );
in01s01 g740727 ( .a(n_39473), .o(n_39474) );
ao12s02 g740728 ( .a(n_39358), .b(n_39448), .c(n_39425), .o(n_39473) );
na02s10 TIMEBOOST_cell_792 ( .a(n_6642), .b(TIMEBOOST_net_10), .o(n_6745) );
in01s01 g740732 ( .a(n_40009), .o(n_39580) );
na02s01 g740733 ( .a(n_39537), .b(n_39518), .o(n_40009) );
in01s01 g740735 ( .a(n_39553), .o(n_40007) );
in01f06 g740736 ( .a(n_39553), .o(n_39552) );
in01s01 g740742 ( .a(n_39889), .o(n_39520) );
no02s02 g740743 ( .a(n_39413), .b(n_39445), .o(n_39889) );
in01s01 g740744 ( .a(n_39969), .o(n_39519) );
na02s02 g740745 ( .a(n_39412), .b(n_39444), .o(n_39969) );
no02m01 g740746 ( .a(n_39443), .b(n_39411), .o(n_39910) );
oa22s02 g740747 ( .a(n_39448), .b(n_39457), .c(n_39355), .d(n_39458), .o(n_39932) );
na02s01 g740748 ( .a(n_39489), .b(n_39451), .o(n_39518) );
na02s01 g740749 ( .a(n_39490), .b(n_39452), .o(n_39537) );
na02s08 TIMEBOOST_cell_791 ( .a(n_6607), .b(n_6577), .o(TIMEBOOST_net_10) );
no02s01 g740751 ( .a(n_39356), .b(n_39258), .o(n_39416) );
no02s01 g740752 ( .a(n_39311), .b(n_39366), .o(n_39413) );
no02s01 g740753 ( .a(n_39312), .b(n_39367), .o(n_39445) );
na02s01 g740754 ( .a(n_39353), .b(n_39362), .o(n_39412) );
na02s01 g740755 ( .a(n_39352), .b(n_39363), .o(n_39444) );
no02s01 g740756 ( .a(n_39385), .b(n_39077), .o(n_39443) );
no02s01 g740757 ( .a(n_39384), .b(n_39078), .o(n_39411) );
no02s01 g740758 ( .a(n_39535), .b(n_40183), .o(n_39536) );
na02s01 g740759 ( .a(n_39535), .b(n_40183), .o(n_39534) );
no02s01 g740760 ( .a(n_39532), .b(n_39072), .o(n_39533) );
in01m04 g740762 ( .a(n_39516), .o(n_39517) );
oa12m08 g740763 ( .a(n_39183), .b(n_39493), .c(n_39206), .o(n_39516) );
ao12m10 g740765 ( .a(n_39125), .b(n_39493), .c(n_39121), .o(n_39514) );
no03f06 TIMEBOOST_cell_4836 ( .a(n_26174), .b(n_23466), .c(n_26191), .o(n_26373) );
in01s01 g740769 ( .a(n_39386), .o(n_39497) );
na02m40 TIMEBOOST_cell_784 ( .a(n_22816), .b(TIMEBOOST_net_6), .o(n_22990) );
ao12s01 g740771 ( .a(n_39313), .b(n_39314), .c(n_39010), .o(n_39414) );
in01s01 g740772 ( .a(n_39905), .o(n_39562) );
na02s06 g740773 ( .a(n_39512), .b(n_39492), .o(n_39905) );
in01s01 g740774 ( .a(n_46950), .o(n_39548) );
in01s01 g740776 ( .a(n_39561), .o(n_39978) );
ao12s01 g740777 ( .a(n_39511), .b(n_39510), .c(n_39509), .o(n_39561) );
oa22f08 g740781 ( .a(n_39430), .b(FE_OCPN6923_n_39185), .c(n_39493), .d(n_39186), .o(n_39531) );
in01s01 g740782 ( .a(n_39891), .o(n_39513) );
no02s01 g740783 ( .a(n_39442), .b(n_39407), .o(n_39891) );
oa12s01 g740785 ( .a(n_39080), .b(n_39354), .c(n_39081), .o(n_39408) );
na02s02 g740786 ( .a(n_39463), .b(n_39322), .o(n_39512) );
na02s01 g740787 ( .a(n_39462), .b(n_39323), .o(n_39492) );
na02s01 g740789 ( .a(n_39431), .b(n_39391), .o(n_39472) );
no02s01 g740790 ( .a(n_39510), .b(n_39509), .o(n_39511) );
na02m20 TIMEBOOST_cell_783 ( .a(n_22820), .b(n_22708), .o(TIMEBOOST_net_6) );
no02s01 g740792 ( .a(n_39349), .b(n_39365), .o(n_39442) );
no02s01 g740793 ( .a(n_39350), .b(n_39364), .o(n_39407) );
in01s01 g740794 ( .a(n_39355), .o(n_39448) );
no02s01 g740795 ( .a(n_39314), .b(n_39313), .o(n_39355) );
in01s01 g740796 ( .a(n_39384), .o(n_39385) );
na02s01 g740797 ( .a(n_39354), .b(n_38984), .o(n_39384) );
na02s01 g740798 ( .a(n_39470), .b(n_40202), .o(n_39471) );
oa12m08 g740799 ( .a(n_39131), .b(n_39440), .c(n_38981), .o(n_39441) );
no02f08 g740800 ( .a(n_39406), .b(n_39129), .o(n_39469) );
in01s01 g740801 ( .a(n_39489), .o(n_39490) );
oa12s01 g740802 ( .a(n_38980), .b(n_39468), .c(n_39395), .o(n_39489) );
na02s01 TIMEBOOST_cell_5618 ( .a(n_6237), .b(n_6140), .o(TIMEBOOST_net_1757) );
in01m04 g740804 ( .a(n_39466), .o(n_39467) );
ao12f08 g740805 ( .a(n_39280), .b(n_39381), .c(n_39279), .o(n_39466) );
no02f06 g740806 ( .a(n_39293), .b(n_39140), .o(n_39356) );
in01s01 g740807 ( .a(n_39311), .o(n_39312) );
oa12s01 g740808 ( .a(n_39061), .b(n_39264), .c(n_38885), .o(n_39311) );
in01s01 g740809 ( .a(n_39352), .o(n_39353) );
ao12s01 g740810 ( .a(n_39242), .b(n_39291), .c(n_39303), .o(n_39352) );
in01s01 g740811 ( .a(n_39535), .o(n_39508) );
na02s01 g740812 ( .a(n_39438), .b(n_39405), .o(n_39535) );
no02s01 g740813 ( .a(n_39464), .b(n_39439), .o(n_39900) );
oa12s01 g740814 ( .a(n_39435), .b(n_39434), .c(n_39433), .o(n_39917) );
no02s01 g740816 ( .a(n_39437), .b(n_39164), .o(n_39532) );
ao22s01 g740817 ( .a(n_39468), .b(n_39423), .c(n_39381), .d(n_39424), .o(n_39947) );
ao22s01 g740818 ( .a(n_39376), .b(n_39151), .c(n_39440), .d(n_39152), .o(n_39945) );
in01s01 g740819 ( .a(n_39853), .o(n_39465) );
no02s02 g740820 ( .a(n_39383), .b(n_39351), .o(n_39853) );
na02s02 g740821 ( .a(n_39265), .b(n_39292), .o(n_39878) );
in01s01 g740822 ( .a(n_39538), .o(n_39488) );
na02s01 g740823 ( .a(n_39382), .b(n_39404), .o(n_39538) );
no02f08 g740824 ( .a(n_39440), .b(n_38981), .o(n_39406) );
no02s01 g740825 ( .a(n_39401), .b(n_39075), .o(n_39439) );
no02s01 g740826 ( .a(n_39402), .b(n_39074), .o(n_39464) );
na02s01 g740827 ( .a(n_39374), .b(n_39321), .o(n_39405) );
na02s01 g740828 ( .a(n_39375), .b(n_39320), .o(n_39438) );
no02s01 g740829 ( .a(n_39436), .b(n_38998), .o(n_39437) );
no02s01 g740830 ( .a(n_39218), .b(n_39301), .o(n_39351) );
no02s01 g740831 ( .a(n_39219), .b(n_39302), .o(n_39383) );
na02s01 g740832 ( .a(n_39264), .b(n_39057), .o(n_39265) );
na02s01 g740833 ( .a(n_39239), .b(n_39058), .o(n_39292) );
na02s01 g740834 ( .a(n_39291), .b(n_39012), .o(n_39354) );
na02s01 g740835 ( .a(n_39291), .b(n_39329), .o(n_39382) );
na02s01 g740836 ( .a(n_39237), .b(n_39330), .o(n_39404) );
na02s01 g740837 ( .a(n_39434), .b(n_39433), .o(n_39435) );
ao12s01 g740839 ( .a(n_39076), .b(n_39380), .c(n_39045), .o(n_39431) );
in01s01 g740840 ( .a(n_39462), .o(n_39463) );
ao12s02 g740841 ( .a(n_38905), .b(n_39399), .c(n_38990), .o(n_39462) );
no03s08 TIMEBOOST_cell_2771 ( .a(n_46950), .b(FE_OCP_RBN6154_n_39816), .c(n_40015), .o(n_40020) );
in01s01 g740843 ( .a(n_39349), .o(n_39350) );
ao12s01 g740844 ( .a(n_39244), .b(n_39310), .c(n_39304), .o(n_39349) );
in01s01 g740845 ( .a(n_39293), .o(n_39314) );
no02s01 g740847 ( .a(n_39379), .b(n_39400), .o(n_39841) );
in01s01 g740848 ( .a(n_39470), .o(n_39894) );
na02s01 g740849 ( .a(n_39346), .b(n_39345), .o(n_39470) );
in01m08 g740850 ( .a(n_39493), .o(n_39430) );
oa12s02 g740852 ( .a(n_39223), .b(n_39222), .c(n_39221), .o(n_39832) );
na02s01 g740853 ( .a(n_39378), .b(n_39398), .o(n_39881) );
in01s01 g740856 ( .a(n_39381), .o(n_39468) );
na02m06 g740857 ( .a(n_39347), .b(n_39254), .o(n_39381) );
in01s01 g740858 ( .a(n_39401), .o(n_39402) );
no02s01 g740859 ( .a(n_39380), .b(n_38973), .o(n_39401) );
no02s01 g740860 ( .a(n_39399), .b(n_39047), .o(n_39400) );
no02s01 g740861 ( .a(n_39342), .b(n_39046), .o(n_39379) );
na02s01 g740862 ( .a(n_39377), .b(n_38978), .o(n_39436) );
na02s01 g740863 ( .a(n_39310), .b(n_39331), .o(n_39378) );
na02s01 g740864 ( .a(n_39217), .b(n_39332), .o(n_39398) );
na02s01 g740865 ( .a(n_39289), .b(n_39274), .o(n_39346) );
na02s01 g740866 ( .a(n_39288), .b(n_39275), .o(n_39345) );
na02s01 g740867 ( .a(n_39222), .b(n_39221), .o(n_39223) );
na02s01 g740868 ( .a(n_39460), .b(n_40177), .o(n_39461) );
no02s01 g740869 ( .a(n_39377), .b(n_39158), .o(n_39434) );
in01s01 g740870 ( .a(n_39440), .o(n_39376) );
oa12f10 g740871 ( .a(n_39236), .b(n_44312), .c(n_39192), .o(n_39440) );
in01s01 g740872 ( .a(n_39374), .o(n_39375) );
oa12s01 g740873 ( .a(n_39326), .b(n_44309), .c(n_38940), .o(n_39374) );
in01s01 g740874 ( .a(n_39264), .o(n_39239) );
na02s01 g740875 ( .a(n_39168), .b(n_39111), .o(n_39264) );
in01s01 g740877 ( .a(n_39237), .o(n_39291) );
in01s01 g740879 ( .a(n_39220), .o(n_39237) );
oa12f08 g740880 ( .a(n_39145), .b(n_39113), .c(n_39062), .o(n_39220) );
in01s01 g740881 ( .a(n_39218), .o(n_39219) );
ao12s01 g740882 ( .a(n_38967), .b(n_39167), .c(n_38924), .o(n_39218) );
in01s01 g740883 ( .a(n_39844), .o(n_39459) );
no02s02 g740884 ( .a(n_39373), .b(n_39343), .o(n_39844) );
in01s01 g740885 ( .a(n_39869), .o(n_39506) );
no02s01 g740886 ( .a(n_39397), .b(n_39429), .o(n_39869) );
na02s01 g740887 ( .a(n_39428), .b(n_39396), .o(n_40183) );
na02f10 g740888 ( .a(n_39290), .b(n_39191), .o(n_39347) );
no02s01 g740889 ( .a(n_39368), .b(n_39298), .o(n_39397) );
no02s01 g740890 ( .a(n_39369), .b(n_39297), .o(n_39429) );
no02s01 g740891 ( .a(n_39307), .b(n_39269), .o(n_39373) );
no02s01 g740892 ( .a(n_39306), .b(n_39270), .o(n_39343) );
no02s01 g740893 ( .a(n_44309), .b(n_39049), .o(n_39380) );
in01s01 g740894 ( .a(n_39310), .o(n_39217) );
na02s01 g740895 ( .a(n_39147), .b(n_39086), .o(n_39310) );
na02s01 g740896 ( .a(n_39146), .b(n_39060), .o(n_39168) );
no02s01 g740897 ( .a(n_39167), .b(n_38916), .o(n_39222) );
na02s01 g740898 ( .a(n_44311), .b(n_39360), .o(n_39396) );
na02s01 g740899 ( .a(n_44309), .b(n_39361), .o(n_39428) );
no02s01 g740900 ( .a(n_44312), .b(n_39134), .o(n_39377) );
in01s01 g740901 ( .a(n_39342), .o(n_39399) );
na02s01 TIMEBOOST_cell_4129 ( .a(n_35897), .b(FE_OCP_RBN3171_n_44211), .o(TIMEBOOST_net_1155) );
in01s01 g740903 ( .a(n_39288), .o(n_39289) );
ao12s01 g740904 ( .a(n_39203), .b(n_39088), .c(n_39251), .o(n_39288) );
oa12s01 g740906 ( .a(n_39287), .b(n_39286), .c(n_39285), .o(n_39371) );
in01s01 g740907 ( .a(n_39460), .o(n_39840) );
na02s01 g740908 ( .a(n_39309), .b(n_39341), .o(n_39460) );
na02s01 g740909 ( .a(n_39340), .b(n_39370), .o(n_39864) );
na02s01 g740910 ( .a(n_39308), .b(n_39336), .o(n_40202) );
in01s01 g740911 ( .a(n_39808), .o(n_39427) );
ao12s01 g740912 ( .a(n_39339), .b(n_39338), .c(n_39337), .o(n_39808) );
no02f08 TIMEBOOST_cell_3117 ( .a(TIMEBOOST_net_849), .b(n_42738), .o(n_42790) );
na02s01 g740914 ( .a(n_39283), .b(n_39267), .o(n_39309) );
na02s01 g740915 ( .a(n_39284), .b(n_39268), .o(n_39341) );
na02s01 g740916 ( .a(n_39257), .b(n_39299), .o(n_39340) );
na02s01 g740917 ( .a(n_39256), .b(n_39300), .o(n_39370) );
na02s01 g740918 ( .a(n_39286), .b(n_39285), .o(n_39287) );
no02s01 g740919 ( .a(n_39338), .b(n_39337), .o(n_39339) );
no02s01 g740920 ( .a(n_39114), .b(n_38881), .o(n_39167) );
no02f04 g740921 ( .a(n_39258), .b(n_39103), .o(n_39259) );
na02s01 g740922 ( .a(n_39114), .b(n_39277), .o(n_39336) );
na02s01 g740923 ( .a(n_39087), .b(n_39276), .o(n_39308) );
in01s01 g740924 ( .a(n_39368), .o(n_39369) );
no02s01 g740925 ( .a(n_39261), .b(n_39281), .o(n_39368) );
na02s10 TIMEBOOST_cell_776 ( .a(TIMEBOOST_net_2), .b(n_6656), .o(n_6734) );
in01s01 g740928 ( .a(n_39306), .o(n_39307) );
oa12s01 g740929 ( .a(n_39064), .b(n_39214), .c(n_38994), .o(n_39306) );
in01s01 g740930 ( .a(n_39146), .o(n_39147) );
in01s01 g740931 ( .a(n_39113), .o(n_39146) );
na02f08 g740932 ( .a(n_39088), .b(n_39016), .o(n_39113) );
na02m04 TIMEBOOST_cell_8640 ( .a(FE_OCP_RBN6381_n_30824), .b(FE_OCPN5300_n_27130), .o(TIMEBOOST_net_2807) );
in01s01 g740934 ( .a(n_39256), .o(n_39257) );
no02s01 g740935 ( .a(n_39195), .b(n_39083), .o(n_39256) );
no02s01 g740936 ( .a(n_39194), .b(n_38937), .o(n_39261) );
no02s01 g740938 ( .a(n_39213), .b(n_39063), .o(n_39286) );
na02m04 g740939 ( .a(n_39215), .b(n_39027), .o(n_39258) );
na02f06 g740940 ( .a(n_39215), .b(n_39161), .o(n_39216) );
no02f08 g740941 ( .a(n_39212), .b(n_39157), .o(n_39236) );
na02m04 TIMEBOOST_cell_7749 ( .a(TIMEBOOST_net_2505), .b(n_24604), .o(n_24765) );
no02s01 TIMEBOOST_cell_8826 ( .a(FE_OCP_RBN2961_n_4046), .b(FE_OCP_RBN2921_n_3878), .o(TIMEBOOST_net_2900) );
in01s01 g740944 ( .a(n_39283), .o(n_39284) );
oa12s01 g740945 ( .a(n_39246), .b(n_39252), .c(n_39199), .o(n_39283) );
ao12s01 g740946 ( .a(n_38821), .b(n_39065), .c(n_38864), .o(n_39338) );
in01s01 g740947 ( .a(n_39114), .o(n_39087) );
in01s01 g740948 ( .a(n_39088), .o(n_39114) );
ao12f06 g740949 ( .a(n_38865), .b(n_38934), .c(n_38897), .o(n_39088) );
in01s01 g740950 ( .a(n_40177), .o(n_39426) );
na02s01 g740951 ( .a(n_39333), .b(n_39305), .o(n_40177) );
in01s01 g740952 ( .a(n_39822), .o(n_39334) );
ao22s01 g740953 ( .a(n_39138), .b(n_39228), .c(n_39137), .d(n_39229), .o(n_39822) );
in01s01 g740954 ( .a(n_39112), .o(n_39810) );
oa22s01 g740955 ( .a(n_39065), .b(n_38895), .c(n_38971), .d(n_38896), .o(n_39112) );
in01s01 g740956 ( .a(n_39213), .o(n_39214) );
no02s01 g740957 ( .a(n_39252), .b(n_38928), .o(n_39213) );
no02f08 g740958 ( .a(n_39143), .b(n_39053), .o(n_39166) );
na02s01 g740959 ( .a(n_39252), .b(n_39273), .o(n_39333) );
na02s01 g740960 ( .a(n_39135), .b(n_39272), .o(n_39305) );
in01s01 g740961 ( .a(n_39110), .o(n_39111) );
na02f06 g740962 ( .a(n_39086), .b(n_38879), .o(n_39110) );
in01s01 g740963 ( .a(n_39194), .o(n_39195) );
in01s01 g740964 ( .a(n_39165), .o(n_39194) );
no02f10 g740965 ( .a(n_39106), .b(n_39003), .o(n_39165) );
in01s02 g740966 ( .a(n_39215), .o(n_39193) );
no02f08 g740967 ( .a(n_39313), .b(n_39108), .o(n_39215) );
no02m08 TIMEBOOST_cell_8525 ( .a(TIMEBOOST_net_2749), .b(n_33782), .o(TIMEBOOST_net_337) );
in01m06 g740969 ( .a(n_39212), .o(n_39254) );
oa12f08 g740970 ( .a(n_39105), .b(n_39163), .c(n_39133), .o(n_39212) );
na02m08 g740971 ( .a(n_39191), .b(n_39130), .o(n_39192) );
na02s01 g740972 ( .a(n_39109), .b(n_39271), .o(n_39281) );
na02s01 g740973 ( .a(n_39163), .b(n_38975), .o(n_39164) );
in01s01 g740974 ( .a(n_39143), .o(n_39144) );
na02f08 g740975 ( .a(n_39109), .b(n_38900), .o(n_39143) );
na02s06 g740976 ( .a(n_39139), .b(n_39141), .o(n_39142) );
na02s02 g740977 ( .a(n_39139), .b(n_39007), .o(n_39140) );
na02m04 g740978 ( .a(n_39253), .b(n_39233), .o(n_39280) );
no03s04 TIMEBOOST_cell_8226 ( .a(n_23551), .b(delay_add_ln22_unr14_stage6_stallmux_q_18_), .c(n_23664), .o(n_23689) );
na02f08 g740980 ( .a(n_39059), .b(n_38984), .o(n_39313) );
oa12m08 g740981 ( .a(n_38983), .b(n_39005), .c(FE_OCP_RBN4328_n_38878), .o(n_39108) );
in01s01 g740982 ( .a(n_39161), .o(n_39162) );
ao12m04 g740983 ( .a(n_39026), .b(n_39055), .c(FE_OCP_RBN5895_n_38806), .o(n_39161) );
in01s01 TIMEBOOST_cell_8902 ( .a(n_45898), .o(TIMEBOOST_net_2946) );
in01s01 g740985 ( .a(n_39137), .o(n_39138) );
oa12s01 g740986 ( .a(n_38876), .b(n_39107), .c(n_38957), .o(n_39137) );
in01s01 g740988 ( .a(n_39135), .o(n_39252) );
in01s01 g740990 ( .a(n_39106), .o(n_39135) );
oa12f08 g740991 ( .a(n_38926), .b(n_39002), .c(n_38963), .o(n_39106) );
na02m02 g740992 ( .a(n_39141), .b(n_39156), .o(n_39211) );
oa22s01 g740993 ( .a(n_38992), .b(n_39051), .c(n_38991), .d(n_39107), .o(n_39785) );
in01s01 g740994 ( .a(n_39065), .o(n_38971) );
in01s01 g740995 ( .a(n_38934), .o(n_39065) );
ao12f06 g740996 ( .a(n_38831), .b(n_38968), .c(n_38894), .o(n_38934) );
in01s01 g740997 ( .a(n_39084), .o(n_39085) );
oa12s01 g740998 ( .a(n_38970), .b(n_38969), .c(n_38968), .o(n_39084) );
no02m10 g740999 ( .a(n_39134), .b(n_39133), .o(n_39191) );
no02s01 g741000 ( .a(n_38993), .b(n_39063), .o(n_39064) );
ao12m08 g741001 ( .a(n_38974), .b(n_38989), .c(n_44926), .o(n_39105) );
in01s01 g741003 ( .a(n_39163), .o(n_39158) );
no03f04 TIMEBOOST_cell_3810 ( .a(FE_OCP_RBN6102_n_26358), .b(FE_RN_1641_0), .c(n_26406), .o(n_26516) );
in01s01 g741005 ( .a(n_39109), .o(n_39083) );
no02m08 TIMEBOOST_cell_3076 ( .a(n_38601), .b(n_38778), .o(TIMEBOOST_net_829) );
na02s02 TIMEBOOST_cell_2121 ( .a(n_26645), .b(n_26552), .o(TIMEBOOST_net_675) );
na02s01 g741008 ( .a(n_38969), .b(n_38968), .o(n_38970) );
no02m04 g741009 ( .a(n_39234), .b(n_39278), .o(n_39279) );
no02m04 g741010 ( .a(n_38966), .b(n_38932), .o(n_39016) );
in01s02 g741013 ( .a(n_39139), .o(n_39104) );
no02m04 g741015 ( .a(n_39008), .b(n_38986), .o(n_39141) );
na02f04 g741016 ( .a(n_38837), .b(FE_OCP_RBN6756_n_38806), .o(n_38897) );
no02s02 TIMEBOOST_cell_5977 ( .a(n_23237), .b(n_23108), .o(TIMEBOOST_net_1840) );
no02m03 TIMEBOOST_cell_8477 ( .a(FE_OCPN1717_n_12311), .b(TIMEBOOST_net_2725), .o(TIMEBOOST_net_116) );
no02m08 TIMEBOOST_cell_4118 ( .a(TIMEBOOST_net_1149), .b(n_25786), .o(TIMEBOOST_net_495) );
in01s01 g741020 ( .a(n_39209), .o(n_39210) );
na02f08 TIMEBOOST_cell_4138 ( .a(TIMEBOOST_net_1159), .b(n_25911), .o(n_26037) );
na02m04 g741022 ( .a(n_39205), .b(n_39175), .o(n_39234) );
na02m06 g741023 ( .a(n_38864), .b(n_38834), .o(n_38865) );
na02s01 g741024 ( .a(n_38915), .b(n_38860), .o(n_38967) );
na02m02 g741025 ( .a(n_38880), .b(n_38886), .o(n_38932) );
no02s01 g741026 ( .a(n_39030), .b(n_39056), .o(n_39080) );
no02s01 g741028 ( .a(n_39028), .b(n_39004), .o(n_39079) );
na02m02 g741030 ( .a(n_39007), .b(n_39006), .o(n_39008) );
no02s02 g741031 ( .a(n_39155), .b(n_39154), .o(n_39156) );
na02f02 g741032 ( .a(n_38836), .b(n_38820), .o(n_38837) );
in01s01 g741033 ( .a(n_39276), .o(n_39277) );
na02s01 g741034 ( .a(n_39204), .b(n_39251), .o(n_39276) );
in01s01 g741035 ( .a(n_38895), .o(n_38896) );
na02s01 g741036 ( .a(n_38864), .b(n_38836), .o(n_38895) );
no02s01 g741037 ( .a(n_38966), .b(n_38833), .o(n_39221) );
in01s01 g741038 ( .a(n_39331), .o(n_39332) );
na02s01 g741039 ( .a(n_39245), .b(n_39304), .o(n_39331) );
no02m04 g741040 ( .a(n_38833), .b(n_38862), .o(n_38863) );
in01s01 g741041 ( .a(n_39057), .o(n_39058) );
na02s01 g741042 ( .a(n_39061), .b(n_38922), .o(n_39057) );
no02m04 TIMEBOOST_cell_4404 ( .a(TIMEBOOST_net_1292), .b(FE_OCP_RBN5978_n_9682), .o(n_9944) );
in01s01 g741044 ( .a(n_39329), .o(n_39330) );
na02s01 g741045 ( .a(n_39243), .b(n_39303), .o(n_39329) );
in01s01 g741046 ( .a(n_39077), .o(n_39078) );
no02s01 g741047 ( .a(n_39081), .b(n_39056), .o(n_39077) );
in01s01 g741048 ( .a(n_39457), .o(n_39458) );
na02s01 g741049 ( .a(n_39359), .b(n_39425), .o(n_39457) );
na02f08 TIMEBOOST_cell_4137 ( .a(FE_OCP_RBN4368_n_25889), .b(n_26054), .o(TIMEBOOST_net_1159) );
na02s01 g741051 ( .a(n_39037), .b(n_38950), .o(n_39483) );
in01s01 g741052 ( .a(n_39504), .o(n_39505) );
na02s01 g741053 ( .a(n_39422), .b(n_39487), .o(n_39504) );
no02m08 g741054 ( .a(n_39004), .b(n_38548), .o(n_39005) );
no02s01 g741055 ( .a(n_38986), .b(n_39103), .o(n_39415) );
na02s02 g741056 ( .a(n_38985), .b(n_38917), .o(n_39055) );
na02s02 g741058 ( .a(FE_OCP_RBN5963_n_39097), .b(n_39098), .o(n_39189) );
no03s02 TIMEBOOST_cell_8370 ( .a(n_4062), .b(n_3966), .c(n_4110), .o(n_4340) );
na02s01 g741060 ( .a(n_38832), .b(n_38894), .o(n_38969) );
na02s08 g741061 ( .a(n_38929), .b(n_38906), .o(n_39003) );
na02s02 TIMEBOOST_cell_8882 ( .a(n_21075), .b(FE_OCP_RBN4466_n_44267), .o(TIMEBOOST_net_2928) );
na02m06 g741063 ( .a(n_38996), .b(n_39048), .o(n_39134) );
no02s06 g741064 ( .a(n_39042), .b(n_44925), .o(n_39157) );
na02f04 TIMEBOOST_cell_5536 ( .a(n_36534), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_1716) );
no02m06 g741066 ( .a(n_38893), .b(n_44946), .o(n_38963) );
no02s01 TIMEBOOST_cell_6096 ( .a(TIMEBOOST_net_1899), .b(n_34278), .o(n_34366) );
no02f08 g741068 ( .a(n_44954), .b(n_38889), .o(n_39063) );
na03m08 TIMEBOOST_cell_4814 ( .a(n_10475), .b(n_10434), .c(n_10421), .o(n_10607) );
no02f08 TIMEBOOST_cell_8611 ( .a(TIMEBOOST_net_2792), .b(n_25968), .o(n_26118) );
na02s02 g741071 ( .a(n_39184), .b(n_44926), .o(n_39233) );
ao12s01 g741072 ( .a(n_38835), .b(FE_OCPN941_n_39096), .c(n_38144), .o(n_39337) );
in01s01 g741073 ( .a(n_39301), .o(n_39302) );
ao12s01 g741074 ( .a(n_38887), .b(FE_OCPN941_n_39096), .c(n_38862), .o(n_39301) );
in01s01 g741075 ( .a(n_39366), .o(n_39367) );
ao12s01 g741076 ( .a(n_38952), .b(FE_OCPN941_n_39096), .c(n_38930), .o(n_39366) );
oa12s01 g741078 ( .a(n_39013), .b(FE_OCPN1090_n_39089), .c(n_38964), .o(n_39455) );
in01s01 g741079 ( .a(n_39502), .o(n_39503) );
oa12s01 g741080 ( .a(n_39009), .b(FE_OCPN1090_n_39089), .c(n_38919), .o(n_39502) );
na02s02 g741082 ( .a(n_39006), .b(n_39100), .o(n_39187) );
in01s01 g741083 ( .a(n_39249), .o(n_39250) );
no02s06 TIMEBOOST_cell_778 ( .a(TIMEBOOST_net_3), .b(n_17354), .o(n_17499) );
in01s01 g741085 ( .a(n_39800), .o(n_39817) );
ao12s01 g741086 ( .a(n_39034), .b(n_39033), .c(n_39032), .o(n_39800) );
in01s01 g741087 ( .a(n_39107), .o(n_39051) );
in01s01 g741088 ( .a(n_39002), .o(n_39107) );
na02f08 g741089 ( .a(n_38883), .b(n_38868), .o(n_39002) );
oa12f06 g741090 ( .a(n_38804), .b(n_38816), .c(n_38856), .o(n_38968) );
in01s01 g741091 ( .a(n_39274), .o(n_39275) );
oa22s01 g741092 ( .a(FE_OCPN1090_n_39089), .b(n_38404), .c(FE_OCPN941_n_39096), .d(n_38434), .o(n_39274) );
ao12s01 g741093 ( .a(n_38858), .b(n_38857), .c(n_38856), .o(n_39768) );
in01s01 g741094 ( .a(n_39364), .o(n_39365) );
oa22s01 g741095 ( .a(FE_OCPN1090_n_39089), .b(n_38484), .c(FE_OCPN941_n_39096), .d(n_38508), .o(n_39364) );
in01s01 g741096 ( .a(n_39362), .o(n_39363) );
oa22s01 g741097 ( .a(FE_OCPN1090_n_39089), .b(n_38526), .c(FE_OCPN941_n_39096), .d(n_38510), .o(n_39362) );
in01s01 g741098 ( .a(n_39500), .o(n_39501) );
oa22s01 g741099 ( .a(FE_OCPN1090_n_39089), .b(n_38493), .c(FE_OCPN941_n_39096), .d(n_38516), .o(n_39500) );
in01s01 g741100 ( .a(n_39528), .o(n_39529) );
oa22s01 g741101 ( .a(FE_OCPN1090_n_39089), .b(n_38543), .c(FE_OCPN941_n_39096), .d(FE_RN_1859_0), .o(n_39528) );
in01s02 g741102 ( .a(n_39247), .o(n_39248) );
na02s03 g741103 ( .a(n_39150), .b(n_39179), .o(n_39247) );
in01s01 g741104 ( .a(n_39207), .o(n_39208) );
oa22s02 g741105 ( .a(n_39089), .b(FE_OCP_RBN4178_n_38586), .c(FE_OCP_RBN4329_n_38878), .d(n_38608), .o(n_39207) );
na02m08 g741106 ( .a(n_39001), .b(n_38999), .o(n_39133) );
no02s08 g741107 ( .a(n_38958), .b(n_38960), .o(n_39050) );
na02s01 g741108 ( .a(n_39021), .b(n_39044), .o(n_39076) );
no02m06 g741109 ( .a(n_39043), .b(n_39000), .o(n_39001) );
no02m06 g741110 ( .a(n_38998), .b(n_38942), .o(n_38999) );
in01s01 g741111 ( .a(n_39048), .o(n_39049) );
no02m04 g741112 ( .a(n_38940), .b(n_38997), .o(n_39048) );
no02m04 g741113 ( .a(n_38995), .b(n_38939), .o(n_38996) );
no02s06 g741114 ( .a(n_38928), .b(n_38927), .o(n_38929) );
no02s06 g741115 ( .a(n_38957), .b(n_38925), .o(n_38926) );
na02s06 g741116 ( .a(n_38959), .b(n_38904), .o(n_38960) );
na02s08 g741117 ( .a(n_39260), .b(n_38902), .o(n_38958) );
in01s01 g741118 ( .a(n_39205), .o(n_39206) );
no02s06 g741119 ( .a(n_39149), .b(n_39125), .o(n_39205) );
no02s01 g741120 ( .a(n_38993), .b(n_38994), .o(n_39285) );
in01s01 g741121 ( .a(n_39272), .o(n_39273) );
na02s01 g741122 ( .a(n_39200), .b(n_39246), .o(n_39272) );
in01s01 g741123 ( .a(n_38991), .o(n_38992) );
no02s01 g741124 ( .a(n_38957), .b(n_38877), .o(n_38991) );
in01s01 g741125 ( .a(n_39299), .o(n_39300) );
na02s01 g741126 ( .a(n_39271), .b(n_38904), .o(n_39299) );
in01s01 g741127 ( .a(n_39046), .o(n_39047) );
na02s01 g741128 ( .a(n_38990), .b(n_38959), .o(n_39046) );
in01s01 g741129 ( .a(n_39360), .o(n_39361) );
na02s01 g741130 ( .a(n_39326), .b(n_38976), .o(n_39360) );
in01s01 g741131 ( .a(n_39074), .o(n_39075) );
na02s01 g741132 ( .a(n_39045), .b(n_39044), .o(n_39074) );
no02s01 g741133 ( .a(n_39318), .b(n_38942), .o(n_39433) );
no02s01 g741135 ( .a(n_38943), .b(n_39043), .o(n_39072) );
in01s01 g741136 ( .a(n_39423), .o(n_39424) );
no02s01 g741137 ( .a(n_39395), .b(n_39041), .o(n_39423) );
in01s01 g741138 ( .a(n_39151), .o(n_39152) );
no02s01 g741139 ( .a(n_39129), .b(n_38981), .o(n_39151) );
no02s06 g741140 ( .a(n_39041), .b(n_39040), .o(n_39042) );
na02s06 g741141 ( .a(n_38988), .b(n_38588), .o(n_38989) );
no02m06 g741142 ( .a(n_38909), .b(n_38955), .o(n_38956) );
no02m04 g741143 ( .a(n_38853), .b(n_38892), .o(n_38893) );
na02f02 TIMEBOOST_cell_8772 ( .a(n_14254), .b(FE_OCP_RBN2557_n_13141), .o(TIMEBOOST_net_2873) );
no02f06 g741145 ( .a(n_38852), .b(n_38888), .o(n_38889) );
no02s06 TIMEBOOST_cell_5009 ( .a(TIMEBOOST_net_1452), .b(n_28771), .o(n_28805) );
na02s01 TIMEBOOST_cell_6231 ( .a(n_27131), .b(FE_OCPN1340_n_27246), .o(TIMEBOOST_net_1967) );
no02s02 g741148 ( .a(n_39120), .b(n_39125), .o(n_39186) );
na02m02 g741149 ( .a(n_39126), .b(n_39121), .o(n_39185) );
na02s02 g741150 ( .a(n_39183), .b(n_39092), .o(n_39184) );
in01s01 g741151 ( .a(n_39203), .o(n_39204) );
no02s01 g741152 ( .a(FE_OCPN1090_n_39089), .b(n_39181), .o(n_39203) );
in01s01 g741153 ( .a(n_38836), .o(n_38821) );
na02f02 g741154 ( .a(n_38806), .b(n_38060), .o(n_38836) );
in01s01 g741155 ( .a(n_38834), .o(n_38835) );
na02s03 g741156 ( .a(FE_OCP_RBN6754_n_38806), .b(n_38820), .o(n_38834) );
na02s01 g741157 ( .a(FE_OCPN1090_n_39089), .b(n_39181), .o(n_39251) );
in01s01 g741159 ( .a(n_38966), .o(n_38924) );
no02s04 g741160 ( .a(FE_OCP_RBN6756_n_38806), .b(n_38431), .o(n_38966) );
in01s01 g741162 ( .a(n_38833), .o(n_38860) );
no02m04 g741163 ( .a(FE_OCP_RBN6754_n_38806), .b(n_38430), .o(n_38833) );
in01s01 g741164 ( .a(n_38886), .o(n_38887) );
na02s02 g741165 ( .a(FE_OCP_RBN6754_n_38806), .b(n_38466), .o(n_38886) );
na02s01 g741166 ( .a(FE_OCPN1090_n_39089), .b(n_39232), .o(n_39304) );
in01s01 g741167 ( .a(n_39244), .o(n_39245) );
no02s01 g741168 ( .a(FE_OCPN1090_n_39089), .b(n_39232), .o(n_39244) );
na02s06 g741169 ( .a(n_38847), .b(n_38859), .o(n_39061) );
in01s01 g741171 ( .a(n_38885), .o(n_38922) );
in01s01 g741173 ( .a(n_38951), .o(n_38952) );
na02s01 g741175 ( .a(FE_OCPN1090_n_39089), .b(n_39230), .o(n_39303) );
in01s01 g741176 ( .a(n_39242), .o(n_39243) );
no02s01 g741177 ( .a(FE_OCPN1090_n_39089), .b(n_39230), .o(n_39242) );
no02s04 g741178 ( .a(FE_OCP_RBN5897_n_38806), .b(n_38884), .o(n_39081) );
in01s01 g741179 ( .a(n_38921), .o(n_39056) );
na02f08 g741180 ( .a(FE_OCP_RBN5895_n_38806), .b(n_38884), .o(n_38921) );
na02s04 g741181 ( .a(FE_OCP_RBN5893_n_38806), .b(n_38964), .o(n_39013) );
na02s01 g741182 ( .a(FE_OCPN1090_n_39089), .b(n_39324), .o(n_39425) );
in01s01 g741183 ( .a(n_39358), .o(n_39359) );
no02s01 g741184 ( .a(FE_OCPN1090_n_39089), .b(n_39324), .o(n_39358) );
in01s01 g741186 ( .a(n_38987), .o(n_39037) );
in01s01 g741188 ( .a(n_39004), .o(n_38950) );
no02m08 g741189 ( .a(n_38847), .b(n_38512), .o(n_39004) );
na02s04 g741190 ( .a(FE_OCP_RBN5894_n_38806), .b(n_38919), .o(n_39009) );
na02s01 g741191 ( .a(FE_OCPN1090_n_39089), .b(n_39393), .o(n_39487) );
in01s01 g741192 ( .a(n_39421), .o(n_39422) );
no02s01 g741193 ( .a(FE_OCPN1090_n_39089), .b(n_39393), .o(n_39421) );
in01s01 g741195 ( .a(n_38986), .o(n_39035) );
no02s06 g741196 ( .a(FE_OCP_RBN5897_n_38806), .b(FE_OCP_RBN2672_n_38534), .o(n_38986) );
in01s01 g741197 ( .a(n_38985), .o(n_39103) );
na02s02 g741198 ( .a(FE_OCP_RBN6757_n_38806), .b(FE_OCP_RBN2672_n_38534), .o(n_38985) );
na02s02 g741199 ( .a(FE_OCP_RBN5894_n_38806), .b(n_38917), .o(n_39006) );
na02s02 g741200 ( .a(FE_OCP_RBN4329_n_38878), .b(FE_OCP_RBN2682_n_38515), .o(n_39100) );
na02s02 g741202 ( .a(FE_OCP_RBN4328_n_38878), .b(FE_OCP_RBN4173_n_38545), .o(n_39098) );
no02s03 g741204 ( .a(FE_OCP_RBN4328_n_38878), .b(FE_OCP_RBN4173_n_38545), .o(n_39097) );
no02s04 g741205 ( .a(FE_OCP_RBN4329_n_38878), .b(n_39095), .o(n_39154) );
no02s02 TIMEBOOST_cell_777 ( .a(n_17426), .b(n_17425), .o(TIMEBOOST_net_3) );
na02s01 g741207 ( .a(n_39089), .b(n_38622), .o(n_39179) );
na02s01 g741208 ( .a(FE_OCP_RBN4329_n_38878), .b(n_38633), .o(n_39150) );
no02s01 g741209 ( .a(n_39033), .b(n_39032), .o(n_39034) );
na02f06 g741210 ( .a(n_38828), .b(n_38841), .o(n_38883) );
in01s01 g741211 ( .a(n_38831), .o(n_38832) );
no02f04 g741212 ( .a(n_38818), .b(n_38817), .o(n_38831) );
na02m04 g741213 ( .a(n_38818), .b(n_38817), .o(n_38894) );
no02s01 g741214 ( .a(n_38857), .b(n_38856), .o(n_38858) );
in01s01 g741215 ( .a(n_39228), .o(n_39229) );
ao12s01 g741216 ( .a(n_38925), .b(n_44926), .c(n_38892), .o(n_39228) );
in01s01 g741217 ( .a(n_39269), .o(n_39270) );
ao12s01 g741218 ( .a(n_38927), .b(n_44926), .c(n_38890), .o(n_39269) );
in01s01 g741219 ( .a(n_39297), .o(n_39298) );
oa12s01 g741220 ( .a(n_39260), .b(n_44925), .c(n_38873), .o(n_39297) );
in01s01 g741221 ( .a(n_39322), .o(n_39323) );
ao12s01 g741222 ( .a(n_38903), .b(n_44926), .c(n_38953), .o(n_39322) );
in01s01 g741223 ( .a(n_39320), .o(n_39321) );
ao12s01 g741224 ( .a(n_38997), .b(n_44926), .c(n_38907), .o(n_39320) );
ao12s01 g741226 ( .a(n_38995), .b(n_44926), .c(n_38955), .o(n_39391) );
oa12s01 g741227 ( .a(n_38941), .b(n_44925), .c(n_38550), .o(n_39509) );
in01s01 g741228 ( .a(n_39453), .o(n_39454) );
ao12s01 g741229 ( .a(n_39000), .b(n_44926), .c(n_38912), .o(n_39453) );
in01s01 g741230 ( .a(n_39176), .o(n_39177) );
no02s02 g741231 ( .a(n_39069), .b(n_39094), .o(n_39176) );
in01s01 g741232 ( .a(n_39201), .o(n_39202) );
na02s02 g741233 ( .a(n_39175), .b(n_39123), .o(n_39201) );
no02m08 TIMEBOOST_cell_4090 ( .a(TIMEBOOST_net_1135), .b(n_39293), .o(n_39386) );
in01s01 g741236 ( .a(n_38915), .o(n_38916) );
in01s01 g741237 ( .a(n_38882), .o(n_38915) );
no02m02 g741238 ( .a(FE_OCP_RBN6754_n_38806), .b(n_38435), .o(n_38882) );
in01s01 g741239 ( .a(n_38880), .o(n_38881) );
na02s02 g741240 ( .a(FE_OCP_RBN6754_n_38806), .b(n_38433), .o(n_38880) );
na02m04 g741241 ( .a(FE_OCP_RBN5896_n_38806), .b(n_38485), .o(n_38879) );
na02s04 g741242 ( .a(n_38847), .b(n_38509), .o(n_39060) );
in01s01 g741244 ( .a(n_38984), .o(n_39030) );
na02s08 g741245 ( .a(FE_OCP_RBN5897_n_38806), .b(n_38527), .o(n_38984) );
na02s02 g741246 ( .a(FE_OCP_RBN5892_n_38806), .b(n_38511), .o(n_39012) );
na02s04 g741247 ( .a(FE_OCP_RBN5894_n_38806), .b(n_38517), .o(n_39010) );
in01s01 g741249 ( .a(n_38983), .o(n_39028) );
na02s08 g741250 ( .a(FE_OCP_RBN5895_n_38806), .b(n_38494), .o(n_38983) );
in01s01 g741251 ( .a(n_39026), .o(n_39027) );
na02s02 g741253 ( .a(FE_OCP_RBN5894_n_38806), .b(n_38563), .o(n_39007) );
no02s04 g741254 ( .a(FE_OCP_RBN4329_n_38878), .b(n_38612), .o(n_39155) );
in01s01 g741255 ( .a(n_39267), .o(n_39268) );
oa22s01 g741256 ( .a(n_44926), .b(n_38888), .c(n_44925), .d(n_38469), .o(n_39267) );
in01s01 g741257 ( .a(n_39451), .o(n_39452) );
oa22s01 g741258 ( .a(n_44926), .b(n_39040), .c(n_44925), .d(n_38538), .o(n_39451) );
in01s02 g741259 ( .a(n_39226), .o(n_39227) );
na02s02 g741260 ( .a(n_39148), .b(n_39118), .o(n_39226) );
in01s01 g741261 ( .a(n_39199), .o(n_39200) );
no02s01 g741262 ( .a(n_44926), .b(n_38405), .o(n_39199) );
na02s01 g741263 ( .a(n_44926), .b(n_38436), .o(n_39271) );
na02s01 g741264 ( .a(n_44926), .b(n_38908), .o(n_39326) );
in01s01 g741265 ( .a(n_39318), .o(n_39319) );
no02s01 g741266 ( .a(n_44925), .b(n_38473), .o(n_39318) );
no02s01 g741267 ( .a(n_44926), .b(n_38553), .o(n_39395) );
no02s01 g741268 ( .a(n_44925), .b(n_39025), .o(n_39094) );
in01s01 g741269 ( .a(n_39068), .o(n_39069) );
na02s02 g741270 ( .a(n_44925), .b(n_39025), .o(n_39068) );
no02s04 g741274 ( .a(n_44946), .b(FE_OCP_RBN2766_n_38530), .o(n_38981) );
in01s01 g741275 ( .a(n_39041), .o(n_38980) );
no02s06 g741276 ( .a(FE_OCP_RBN2861_n_44921), .b(n_38514), .o(n_39041) );
in01s01 g741277 ( .a(n_38988), .o(n_38943) );
na02m03 g741278 ( .a(n_44944), .b(n_46951), .o(n_38988) );
no02m04 g741279 ( .a(n_44921), .b(n_46951), .o(n_39043) );
no02m04 g741280 ( .a(n_44921), .b(n_38912), .o(n_39000) );
in01s01 g741282 ( .a(n_38942), .o(n_38978) );
no02m04 g741283 ( .a(n_44921), .b(n_38572), .o(n_38942) );
in01s01 g741284 ( .a(n_38998), .o(n_38941) );
no02m04 g741285 ( .a(n_44955), .b(n_38573), .o(n_38998) );
in01s01 g741286 ( .a(n_38909), .o(n_39044) );
no02s06 g741287 ( .a(n_44954), .b(n_38471), .o(n_38909) );
in01s01 g741289 ( .a(n_38940), .o(n_38976) );
no02m02 g741290 ( .a(n_44955), .b(n_38908), .o(n_38940) );
no02m02 g741291 ( .a(n_44955), .b(n_38907), .o(n_38997) );
no02s02 g741292 ( .a(n_44955), .b(n_38955), .o(n_38995) );
in01s01 g741293 ( .a(n_38939), .o(n_39045) );
no02s02 g741294 ( .a(n_44944), .b(n_38472), .o(n_38939) );
no02s03 g741295 ( .a(n_44944), .b(n_38890), .o(n_38927) );
in01s01 g741296 ( .a(n_38906), .o(n_38994) );
na02s03 g741297 ( .a(n_44946), .b(n_38829), .o(n_38906) );
no02s06 g741298 ( .a(n_44955), .b(n_38147), .o(n_38957) );
no02s04 g741299 ( .a(n_44955), .b(n_38892), .o(n_38925) );
in01s01 g741300 ( .a(n_38876), .o(n_38877) );
in01s01 g741301 ( .a(n_38853), .o(n_38876) );
no02m02 g741302 ( .a(n_38830), .b(n_38146), .o(n_38853) );
in01s01 g741303 ( .a(n_38959), .o(n_38905) );
na02s06 g741304 ( .a(n_44946), .b(n_38872), .o(n_38959) );
in01s01 g741306 ( .a(n_38904), .o(n_38937) );
na02s06 g741307 ( .a(n_44946), .b(n_38495), .o(n_38904) );
in01s01 g741308 ( .a(n_38902), .o(n_38903) );
na02s08 g741309 ( .a(n_44925), .b(n_38498), .o(n_38902) );
na02s06 g741310 ( .a(n_44946), .b(n_38873), .o(n_39260) );
no02m04 g741311 ( .a(n_38830), .b(n_38829), .o(n_38993) );
in01s01 g741312 ( .a(n_38852), .o(n_39246) );
no02f04 g741313 ( .a(n_38830), .b(n_38468), .o(n_38852) );
in01s01 g741314 ( .a(n_38901), .o(n_38990) );
no02s06 g741315 ( .a(n_44925), .b(n_38872), .o(n_38901) );
in01s01 g741316 ( .a(n_39131), .o(n_39129) );
na02s03 g741317 ( .a(n_44925), .b(FE_OCP_RBN2766_n_38530), .o(n_39131) );
in01s04 g741319 ( .a(n_39126), .o(n_39125) );
na02s02 g741321 ( .a(n_44925), .b(FE_OCP_RBN4193_n_38537), .o(n_39126) );
no02s02 g741322 ( .a(n_44926), .b(n_38598), .o(n_39149) );
na02s01 g741323 ( .a(n_44926), .b(n_38601), .o(n_39123) );
na02s01 g741324 ( .a(n_44925), .b(n_39092), .o(n_39175) );
in01m04 g741325 ( .a(n_39120), .o(n_39121) );
no02s01 g741327 ( .a(n_44925), .b(FE_OCP_RBN4193_n_38537), .o(n_39120) );
na02s06 TIMEBOOST_cell_4227 ( .a(FE_RN_931_0), .b(FE_RN_930_0), .o(TIMEBOOST_net_1204) );
na02s01 g741329 ( .a(n_44926), .b(n_38641), .o(n_39118) );
na02s01 g741330 ( .a(n_44925), .b(n_38627), .o(n_39148) );
no02s01 g741331 ( .a(n_38869), .b(n_38842), .o(n_39033) );
no02s01 g741332 ( .a(n_38805), .b(n_38816), .o(n_38857) );
in01s01 g741333 ( .a(n_38974), .o(n_38975) );
no02m06 g741334 ( .a(FE_OCP_RBN2861_n_44921), .b(n_38574), .o(n_38974) );
in01s01 g741336 ( .a(n_38973), .o(n_39021) );
no02m06 g741337 ( .a(FE_OCP_RBN2861_n_44921), .b(n_38518), .o(n_38973) );
na02s03 g741338 ( .a(n_44925), .b(n_38554), .o(n_39130) );
no02s03 g741339 ( .a(n_44944), .b(n_38470), .o(n_38928) );
na02s02 g741340 ( .a(n_44944), .b(n_38496), .o(n_38900) );
na02s03 g741341 ( .a(n_44926), .b(n_38603), .o(n_39183) );
ao12s01 g741342 ( .a(n_38845), .b(n_38844), .c(n_38843), .o(n_39763) );
in01s01 g741343 ( .a(n_38828), .o(n_39032) );
oa12f04 g741344 ( .a(n_38802), .b(n_38843), .c(n_38813), .o(n_38828) );
ao12f06 g741346 ( .a(n_38761), .b(n_38801), .c(n_38783), .o(n_38856) );
oa12f01 g741347 ( .a(n_38798), .b(n_38801), .c(n_38797), .o(n_39745) );
in01s06 g741381 ( .a(FE_OCP_RBN4329_n_38878), .o(n_39089) );
in01m08 g741394 ( .a(FE_OCP_RBN6757_n_38806), .o(n_38847) );
no02m08 TIMEBOOST_cell_3000 ( .a(n_29062), .b(n_25738), .o(TIMEBOOST_net_791) );
no02s01 g741401 ( .a(n_38843), .b(n_38844), .o(n_38845) );
in01s01 g741402 ( .a(n_38841), .o(n_38842) );
na02m04 g741403 ( .a(n_38811), .b(n_38067), .o(n_38841) );
in01s01 g741404 ( .a(n_38868), .o(n_38869) );
na02s06 g741405 ( .a(n_38812), .b(n_38068), .o(n_38868) );
ao12f06 g741406 ( .a(n_38677), .b(n_38770), .c(n_38708), .o(n_38785) );
no02f04 g741407 ( .a(n_38800), .b(n_38799), .o(n_38816) );
in01s01 g741408 ( .a(n_38804), .o(n_38805) );
na02f04 g741409 ( .a(n_38800), .b(n_38799), .o(n_38804) );
na02s01 g741410 ( .a(n_38801), .b(n_38797), .o(n_38798) );
no02f10 g741448 ( .a(n_38796), .b(n_38779), .o(n_38830) );
na02f08 TIMEBOOST_cell_2999 ( .a(n_34276), .b(TIMEBOOST_net_790), .o(n_34390) );
no02m04 g741450 ( .a(n_38763), .b(n_38707), .o(n_38784) );
na02m02 g741451 ( .a(n_38770), .b(n_38691), .o(n_38769) );
no02s01 g741452 ( .a(n_38803), .b(n_38813), .o(n_38844) );
ao12f08 g741453 ( .a(FE_OCP_RBN4194_n_38683), .b(n_38788), .c(n_38778), .o(n_38796) );
oa12s01 g741454 ( .a(n_38809), .b(n_38808), .c(n_38807), .o(n_39738) );
ao12f04 g741455 ( .a(n_38772), .b(n_38807), .c(n_38790), .o(n_38843) );
in01s02 g741456 ( .a(n_38811), .o(n_38812) );
in01s01 TIMEBOOST_cell_7387 ( .a(TIMEBOOST_net_2323), .o(TIMEBOOST_net_2322) );
oa12f04 g741459 ( .a(n_38744), .b(n_38780), .c(n_38760), .o(n_38801) );
ao12s01 g741460 ( .a(n_38782), .b(n_38781), .c(n_38780), .o(n_39747) );
in01s01 g741461 ( .a(n_38794), .o(n_38795) );
ao12s01 g741462 ( .a(n_38768), .b(n_38767), .c(n_38766), .o(n_38794) );
na02m04 g741463 ( .a(n_44166), .b(n_38729), .o(n_38793) );
no02s03 TIMEBOOST_cell_6922 ( .a(TIMEBOOST_net_2219), .b(TIMEBOOST_net_315), .o(n_8051) );
in01m02 g741465 ( .a(n_38770), .o(n_38763) );
na02f08 g741466 ( .a(n_38746), .b(n_38721), .o(n_38770) );
na02s01 g741467 ( .a(n_38807), .b(n_38808), .o(n_38809) );
in01s01 g741468 ( .a(n_38802), .o(n_38803) );
na02m02 g741469 ( .a(n_38792), .b(n_38791), .o(n_38802) );
no02m02 g741470 ( .a(n_38792), .b(n_38791), .o(n_38813) );
na02s01 g741471 ( .a(n_38762), .b(n_38783), .o(n_38797) );
no02s01 g741472 ( .a(n_38781), .b(n_38780), .o(n_38782) );
no02s01 g741473 ( .a(n_38767), .b(n_38766), .o(n_38768) );
no02s08 g741474 ( .a(n_38759), .b(n_38778), .o(n_38779) );
no02f08 g741476 ( .a(n_38758), .b(n_38716), .o(n_38788) );
na02s01 g741477 ( .a(n_38790), .b(n_38773), .o(n_38808) );
in01s01 g741478 ( .a(n_38761), .o(n_38762) );
no02f04 g741479 ( .a(n_38753), .b(n_38752), .o(n_38761) );
na02f04 g741480 ( .a(n_38753), .b(n_38752), .o(n_38783) );
no02s01 g741481 ( .a(n_38745), .b(n_38760), .o(n_38781) );
ao12s01 g741482 ( .a(n_38776), .b(n_38775), .c(n_38774), .o(n_39740) );
ao22m02 g741483 ( .a(n_38749), .b(n_38726), .c(n_38748), .d(n_38727), .o(n_38792) );
oa12f06 g741484 ( .a(n_38740), .b(n_38774), .c(n_38754), .o(n_38807) );
ao12s01 g741486 ( .a(n_38737), .b(n_38747), .c(n_38736), .o(n_38767) );
in01f02 g741488 ( .a(n_38746), .o(n_38750) );
oa12f06 g741489 ( .a(n_38711), .b(n_38710), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38746) );
in01s04 g741490 ( .a(n_38758), .o(n_38759) );
no02f08 g741491 ( .a(n_38743), .b(n_38715), .o(n_38758) );
no02s01 g741492 ( .a(n_38774), .b(n_38775), .o(n_38776) );
na02f03 g741493 ( .a(n_38765), .b(n_38764), .o(n_38790) );
in01s01 g741494 ( .a(n_38772), .o(n_38773) );
no02m02 g741495 ( .a(n_38765), .b(n_38764), .o(n_38772) );
no02f02 g741496 ( .a(n_38739), .b(n_38738), .o(n_38760) );
in01s01 g741497 ( .a(n_38744), .o(n_38745) );
na02m02 g741498 ( .a(n_38739), .b(n_38738), .o(n_38744) );
no02s01 g741499 ( .a(n_38747), .b(n_38736), .o(n_38737) );
in01s01 g741500 ( .a(n_38786), .o(n_38787) );
ao12s01 g741501 ( .a(n_38757), .b(n_38756), .c(n_38755), .o(n_38786) );
na02m06 g741503 ( .a(n_38709), .b(FE_OCP_RBN6689_n_38655), .o(n_38711) );
no02s01 g741504 ( .a(n_38756), .b(n_38755), .o(n_38757) );
no02s01 g741505 ( .a(n_38754), .b(n_38741), .o(n_38775) );
in01m02 g741506 ( .a(n_38748), .o(n_38749) );
in01m01 g741507 ( .a(n_38743), .o(n_38748) );
na03f10 TIMEBOOST_cell_5885 ( .a(n_39893), .b(FE_OCP_RBN4430_n_39942), .c(n_39975), .o(n_40038) );
no02f06 g741509 ( .a(n_38709), .b(n_38656), .o(n_38710) );
ao12f06 g741510 ( .a(n_38724), .b(n_38742), .c(n_38755), .o(n_38774) );
na02s04 TIMEBOOST_cell_7610 ( .a(FE_OCP_RBN2857_n_9082), .b(FE_OCPN4535_n_9012), .o(TIMEBOOST_net_2436) );
in01m02 g741512 ( .a(n_38734), .o(n_38735) );
na02m04 g741513 ( .a(n_38704), .b(n_38695), .o(n_38734) );
no03s20 TIMEBOOST_cell_2208 ( .a(n_23378), .b(FE_RN_1256_0), .c(FE_RN_1255_0), .o(n_23178) );
na02m02 g741517 ( .a(n_38717), .b(n_38696), .o(n_38728) );
no02s02 TIMEBOOST_cell_7609 ( .a(TIMEBOOST_net_2435), .b(n_29279), .o(TIMEBOOST_net_2230) );
no02s06 g741519 ( .a(n_38707), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38708) );
in01f02 g741520 ( .a(n_38705), .o(n_38706) );
in01m01 g741521 ( .a(n_38709), .o(n_38705) );
no02f08 g741522 ( .a(n_38667), .b(n_38629), .o(n_38709) );
na02s02 g741523 ( .a(n_38676), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38695) );
na02m04 g741524 ( .a(n_38677), .b(n_38778), .o(n_38704) );
na02m02 g741525 ( .a(n_38721), .b(n_38691), .o(n_38722) );
no02m02 g741526 ( .a(n_38707), .b(n_38692), .o(n_38720) );
na02s01 g741527 ( .a(n_38725), .b(n_38742), .o(n_38756) );
no02m06 g741528 ( .a(n_38732), .b(FE_OCPN3564_n_38731), .o(n_38754) );
in01s01 g741529 ( .a(n_38740), .o(n_38741) );
na02f04 g741530 ( .a(n_38732), .b(FE_OCPN3564_n_38731), .o(n_38740) );
ao12f06 g741531 ( .a(n_38690), .b(n_45623), .c(FE_OFN5092_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38719) );
in01s02 g741532 ( .a(n_38729), .o(n_38730) );
oa22s04 g741533 ( .a(FE_OCP_RBN4195_n_38683), .b(n_38778), .c(n_38683), .d(FE_OFN5092_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38729) );
in01m02 g741534 ( .a(n_38693), .o(n_38694) );
oa22f02 g741535 ( .a(FE_OCP_RBN6690_n_38655), .b(n_38778), .c(n_38655), .d(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38693) );
in01s01 g741537 ( .a(n_38703), .o(n_38717) );
no02m08 g741538 ( .a(n_38671), .b(n_38649), .o(n_38703) );
in01m02 g741539 ( .a(n_38726), .o(n_38727) );
no02m02 g741540 ( .a(n_38716), .b(n_38715), .o(n_38726) );
in01m01 g741541 ( .a(n_38721), .o(n_38692) );
na02m08 g741542 ( .a(n_38680), .b(FE_OFN5090_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38721) );
na02f04 g741543 ( .a(n_38655), .b(n_38652), .o(n_38656) );
in01s02 g741544 ( .a(n_38707), .o(n_38691) );
no02m08 g741547 ( .a(n_38680), .b(FE_OFN5091_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38707) );
na02f04 g741548 ( .a(n_38714), .b(n_38713), .o(n_38742) );
in01s01 g741549 ( .a(n_38724), .o(n_38725) );
no02f04 g741550 ( .a(n_38714), .b(n_38713), .o(n_38724) );
in01m02 g741554 ( .a(n_38667), .o(n_38678) );
ao12f08 g741555 ( .a(n_38778), .b(n_38654), .c(n_38624), .o(n_38667) );
oa12s01 g741556 ( .a(n_38687), .b(n_38686), .c(n_38685), .o(n_39675) );
no02s01 TIMEBOOST_cell_5292 ( .a(FE_OCP_RBN5935_n_44563), .b(FE_OCP_RBN5906_n_44563), .o(TIMEBOOST_net_1594) );
in01s02 g741558 ( .a(n_38696), .o(n_38697) );
oa22f02 g741559 ( .a(n_38690), .b(FE_OFN5092_delay_sub_ln23_0_unr25_stage9_stallmux_q), .c(n_38647), .d(n_38778), .o(n_38696) );
in01s01 g741560 ( .a(n_38712), .o(n_39679) );
ao12s01 g741561 ( .a(n_38670), .b(n_38669), .c(n_38668), .o(n_38712) );
in01s04 g741562 ( .a(n_38676), .o(n_38677) );
na02m04 TIMEBOOST_cell_6009 ( .a(n_41208), .b(n_41046), .o(TIMEBOOST_net_1856) );
in01f02 g741565 ( .a(n_38673), .o(n_38674) );
no02f08 g741568 ( .a(n_38651), .b(n_38648), .o(n_38671) );
no02s04 g741569 ( .a(n_38660), .b(n_38663), .o(n_38689) );
no02s06 g741571 ( .a(n_38658), .b(n_38778), .o(n_38715) );
no02m06 g741572 ( .a(n_38659), .b(FE_OFN5092_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38716) );
no02s06 TIMEBOOST_cell_5239 ( .a(TIMEBOOST_net_1567), .b(FE_OCP_RBN2664_n_24372), .o(n_24534) );
no02s01 TIMEBOOST_cell_3824 ( .a(TIMEBOOST_net_1002), .b(n_6600), .o(n_6652) );
na02f02 g741575 ( .a(n_38643), .b(n_38652), .o(n_38653) );
no02f02 g741576 ( .a(n_38629), .b(n_38630), .o(n_38666) );
na02s01 g741577 ( .a(n_38686), .b(n_38685), .o(n_38687) );
na02s04 g741578 ( .a(n_38657), .b(n_38685), .o(n_38755) );
no02s01 g741579 ( .a(n_38669), .b(n_38668), .o(n_38670) );
na02m06 g741580 ( .a(n_38669), .b(n_37636), .o(n_38766) );
no02m08 TIMEBOOST_cell_2094 ( .a(n_26537), .b(TIMEBOOST_net_661), .o(n_26985) );
na02f04 g741584 ( .a(n_38664), .b(n_38665), .o(n_38714) );
no02m04 TIMEBOOST_cell_6780 ( .a(TIMEBOOST_net_2147), .b(n_9742), .o(TIMEBOOST_net_1630) );
na02s01 TIMEBOOST_cell_8860 ( .a(n_6368), .b(n_6268), .o(TIMEBOOST_net_2917) );
na02m02 g741588 ( .a(n_38635), .b(n_38640), .o(n_38665) );
na02f02 g741589 ( .a(n_38636), .b(n_38639), .o(n_38664) );
in01s02 g741590 ( .a(n_38662), .o(n_38663) );
in01s01 g741591 ( .a(n_38651), .o(n_38662) );
na02f06 g741592 ( .a(n_38626), .b(n_38623), .o(n_38651) );
na02f06 TIMEBOOST_cell_5525 ( .a(TIMEBOOST_net_1710), .b(n_36458), .o(n_36549) );
no02s06 g741594 ( .a(n_38633), .b(n_38778), .o(n_38650) );
no02m02 g741596 ( .a(n_38649), .b(n_38648), .o(n_38660) );
no02m06 TIMEBOOST_cell_4226 ( .a(TIMEBOOST_net_1203), .b(n_37516), .o(n_37649) );
no02s01 TIMEBOOST_cell_8541 ( .a(TIMEBOOST_net_2757), .b(n_14352), .o(n_14489) );
in01m01 g741599 ( .a(n_38652), .o(n_38630) );
na02f04 g741600 ( .a(n_38616), .b(n_38778), .o(n_38652) );
no02f08 g741601 ( .a(n_38587), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38604) );
no02m08 TIMEBOOST_cell_5005 ( .a(TIMEBOOST_net_1450), .b(n_37763), .o(n_37794) );
in01m01 g741604 ( .a(n_38629), .o(n_38643) );
no02m08 g741605 ( .a(n_38616), .b(n_38778), .o(n_38629) );
na02s01 g741606 ( .a(n_38587), .b(FE_OCP_RBN4193_n_38537), .o(n_38603) );
in01m02 g741607 ( .a(n_38658), .o(n_38659) );
no02s02 TIMEBOOST_cell_6666 ( .a(TIMEBOOST_net_2090), .b(n_3238), .o(n_3338) );
in01s01 g741609 ( .a(n_38657), .o(n_38686) );
ao22s02 g741610 ( .a(n_38610), .b(n_38778), .c(n_38609), .d(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38657) );
in01f02 g741612 ( .a(n_38654), .o(n_38628) );
na02f08 g741613 ( .a(n_38589), .b(n_38584), .o(n_38654) );
in01s01 g741615 ( .a(n_38627), .o(n_38641) );
in01s02 g741616 ( .a(n_38615), .o(n_38627) );
oa22m02 g741617 ( .a(n_38571), .b(n_38258), .c(n_38570), .d(n_38259), .o(n_38615) );
in01m02 g741618 ( .a(n_38690), .o(n_38647) );
na03f06 TIMEBOOST_cell_8410 ( .a(n_16624), .b(n_16599), .c(TIMEBOOST_net_1755), .o(n_16757) );
in01s02 g741620 ( .a(n_38639), .o(n_38640) );
in01s01 g741621 ( .a(n_38626), .o(n_38639) );
na02f06 g741622 ( .a(n_38596), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38626) );
no02f06 g741623 ( .a(n_38594), .b(n_38778), .o(n_38648) );
na02m08 TIMEBOOST_cell_4240 ( .a(n_12761), .b(TIMEBOOST_net_1210), .o(n_12921) );
no02s04 g741625 ( .a(n_38586), .b(n_38778), .o(n_38602) );
no02m06 g741626 ( .a(n_38595), .b(FE_OFN5092_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38649) );
no02s02 TIMEBOOST_cell_2091 ( .a(n_30558), .b(n_45744), .o(TIMEBOOST_net_660) );
no02m10 TIMEBOOST_cell_2909 ( .a(TIMEBOOST_net_745), .b(n_33550), .o(n_33664) );
na02f06 g741629 ( .a(FE_OCP_RBN5735_n_38569), .b(n_38778), .o(n_38589) );
in01s01 g741631 ( .a(n_38624), .o(n_38637) );
na02m08 g741632 ( .a(n_38591), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38624) );
na02m04 g741633 ( .a(n_38569), .b(FE_OFN5093_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38584) );
no02s01 g741634 ( .a(FE_OCP_RBN4178_n_38586), .b(FE_OCP_RBN4173_n_38545), .o(n_38612) );
in01m02 g741635 ( .a(n_38635), .o(n_38636) );
na02m02 g741636 ( .a(n_38597), .b(n_38623), .o(n_38635) );
in01s02 g741638 ( .a(n_38622), .o(n_38633) );
ao22s04 g741640 ( .a(n_38577), .b(n_38212), .c(FE_OCP_RBN5698_n_38577), .d(n_38211), .o(n_38622) );
in01s01 g741641 ( .a(n_38912), .o(n_38588) );
na02s02 g741642 ( .a(n_38541), .b(n_38555), .o(n_38912) );
in01s06 g741644 ( .a(n_38601), .o(n_39092) );
na02m08 g741646 ( .a(n_38556), .b(n_38575), .o(n_38601) );
in01s01 g741649 ( .a(n_38587), .o(n_38598) );
in01f04 g741650 ( .a(n_38583), .o(n_38587) );
na02f04 g741653 ( .a(n_38579), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38623) );
na02m02 g741654 ( .a(n_38580), .b(n_38778), .o(n_38597) );
na02m04 g741657 ( .a(n_38539), .b(n_38239), .o(n_38556) );
na02m08 g741658 ( .a(n_38540), .b(n_38240), .o(n_38575) );
na02s01 g741659 ( .a(n_38522), .b(n_38374), .o(n_38555) );
na02s01 g741660 ( .a(n_38521), .b(n_38375), .o(n_38541) );
no02s01 g741661 ( .a(n_38573), .b(n_38572), .o(n_38574) );
na02s01 g741662 ( .a(n_39040), .b(n_38553), .o(n_38554) );
in01s01 g741663 ( .a(n_38570), .o(n_38571) );
no02s01 TIMEBOOST_cell_6854 ( .a(TIMEBOOST_net_2184), .b(FE_OCPN5113_n_22249), .o(n_22501) );
in01s02 g741665 ( .a(n_38609), .o(n_38610) );
in01s01 g741666 ( .a(n_38596), .o(n_38609) );
na02s06 TIMEBOOST_cell_2894 ( .a(n_2007), .b(n_2006), .o(TIMEBOOST_net_738) );
in01m02 g741668 ( .a(n_38594), .o(n_38595) );
in01s01 g741672 ( .a(FE_OCP_RBN4178_n_38586), .o(n_38608) );
in01s01 g741677 ( .a(FE_OCP_RBN4180_n_38592), .o(n_39095) );
oa22m06 g741679 ( .a(n_38546), .b(n_38234), .c(n_38547), .d(n_38233), .o(n_38592) );
in01s01 g741680 ( .a(FE_OCP_RBN5736_n_38569), .o(n_39025) );
in01m02 g741684 ( .a(n_38605), .o(n_38606) );
in01m02 g741685 ( .a(n_38591), .o(n_38605) );
na02s01 TIMEBOOST_cell_6054 ( .a(TIMEBOOST_net_1878), .b(n_784), .o(n_848) );
no02f10 TIMEBOOST_cell_2893 ( .a(n_33273), .b(TIMEBOOST_net_737), .o(n_33331) );
no02f04 TIMEBOOST_cell_8636 ( .a(FE_RN_1964_0), .b(FE_RN_1963_0), .o(TIMEBOOST_net_2805) );
no02m08 TIMEBOOST_cell_5084 ( .a(n_17732), .b(n_18950), .o(TIMEBOOST_net_1490) );
na02m02 TIMEBOOST_cell_8599 ( .a(TIMEBOOST_net_2786), .b(n_26175), .o(n_26202) );
in01m04 g741691 ( .a(n_38539), .o(n_38540) );
na02m06 g741692 ( .a(n_38523), .b(n_38217), .o(n_38539) );
no02s01 TIMEBOOST_cell_5955 ( .a(n_32603), .b(n_32443), .o(TIMEBOOST_net_1829) );
na02s01 g741695 ( .a(n_38564), .b(n_38562), .o(n_38563) );
in01s01 g741696 ( .a(n_38521), .o(n_38522) );
oa12s01 g741697 ( .a(n_38089), .b(n_38478), .c(n_37949), .o(n_38521) );
ao12f04 g741699 ( .a(n_38102), .b(n_38506), .c(n_46416), .o(n_38519) );
in01m01 g741700 ( .a(n_38579), .o(n_38580) );
no02f08 TIMEBOOST_cell_2048 ( .a(TIMEBOOST_net_638), .b(FE_OCP_RBN2733_n_29657), .o(n_29696) );
in01s01 g741704 ( .a(n_39040), .o(n_38538) );
oa12s02 g741705 ( .a(n_38482), .b(n_38481), .c(n_38480), .o(n_39040) );
in01s01 g741707 ( .a(n_38573), .o(n_38550) );
na02s01 g741708 ( .a(n_38477), .b(n_38504), .o(n_38573) );
in01s01 g741715 ( .a(n_38919), .o(n_38548) );
ao12s01 g741716 ( .a(n_38503), .b(n_38502), .c(n_38501), .o(n_38919) );
na02s01 g741717 ( .a(n_38481), .b(n_38480), .o(n_38482) );
na02s04 g741718 ( .a(n_38506), .b(n_38156), .o(n_38523) );
na02s01 g741719 ( .a(n_38478), .b(n_38085), .o(n_38479) );
na02s01 g741721 ( .a(n_38457), .b(n_38349), .o(n_38477) );
na02s01 g741722 ( .a(n_38458), .b(n_38350), .o(n_38504) );
in01m04 g741723 ( .a(n_38546), .o(n_38547) );
na02m08 g741724 ( .a(n_46417), .b(n_38199), .o(n_38546) );
na02f06 TIMEBOOST_cell_6722 ( .a(TIMEBOOST_net_2118), .b(n_24071), .o(n_24181) );
no02s01 g741726 ( .a(n_38907), .b(n_38908), .o(n_38518) );
no02s01 g741727 ( .a(n_38502), .b(n_38501), .o(n_38503) );
in01f02 g741728 ( .a(n_38499), .o(n_38500) );
oa12f06 g741729 ( .a(n_38051), .b(n_38421), .c(FE_OCPN1056_n_38087), .o(n_38499) );
na02f06 g741735 ( .a(n_38497), .b(n_38476), .o(n_38545) );
na02m06 g741737 ( .a(n_38475), .b(n_38134), .o(n_38531) );
oa12s02 g741741 ( .a(n_38463), .b(n_38462), .c(n_38461), .o(n_38955) );
in01s01 g741742 ( .a(n_38498), .o(n_38953) );
ao12s02 g741743 ( .a(n_38428), .b(n_38427), .c(n_38426), .o(n_38498) );
in01s01 g741744 ( .a(FE_RN_1859_0), .o(n_38543) );
oa12s01 g741745 ( .a(n_38492), .b(n_38491), .c(n_38490), .o(n_38564) );
no02s01 g741746 ( .a(n_38427), .b(n_38426), .o(n_38428) );
na02s01 g741747 ( .a(n_38462), .b(n_38461), .o(n_38463) );
na02f06 g741748 ( .a(FE_OCP_RBN5683_n_38474), .b(n_38158), .o(n_38497) );
na02s04 g741749 ( .a(n_38474), .b(n_38159), .o(n_38476) );
na02m04 g741750 ( .a(n_38474), .b(FE_OCPN1626_n_38135), .o(n_38475) );
na02s01 g741751 ( .a(n_38873), .b(n_38495), .o(n_38496) );
na02s01 g741752 ( .a(n_38516), .b(n_38467), .o(n_38517) );
na02s01 g741753 ( .a(n_38493), .b(n_39324), .o(n_38494) );
na02s01 g741754 ( .a(n_38491), .b(n_38490), .o(n_38492) );
oa12s01 g741755 ( .a(n_38328), .b(n_38455), .c(n_38378), .o(n_38481) );
in01m02 g741756 ( .a(n_38506), .o(n_38460) );
na02f08 g741757 ( .a(n_38369), .b(n_38168), .o(n_38506) );
oa22s01 g741759 ( .a(n_38425), .b(n_38036), .c(n_38236), .d(n_37639), .o(n_38478) );
in01s01 g741760 ( .a(n_38457), .o(n_38458) );
oa12s01 g741761 ( .a(n_38314), .b(n_38425), .c(n_38333), .o(n_38457) );
in01s01 g741763 ( .a(FE_OCP_RBN2681_n_38515), .o(n_38917) );
in01s01 g741768 ( .a(n_38553), .o(n_38514) );
oa12s01 g741769 ( .a(n_38456), .b(n_38455), .c(n_38454), .o(n_38553) );
in01s01 g741770 ( .a(n_38572), .o(n_38473) );
oa12s01 g741771 ( .a(n_38403), .b(n_38425), .c(n_38402), .o(n_38572) );
oa12s01 g741772 ( .a(n_38424), .b(n_38423), .c(n_38422), .o(n_38907) );
in01s01 g741773 ( .a(n_38471), .o(n_38472) );
ao12s01 g741774 ( .a(n_38401), .b(n_38400), .c(n_38399), .o(n_38471) );
ao12s02 g741776 ( .a(n_38452), .b(n_38451), .c(n_38450), .o(n_38512) );
oa12s01 g741777 ( .a(n_38323), .b(n_38389), .c(n_38373), .o(n_38502) );
na02s01 g741778 ( .a(n_38455), .b(n_38454), .o(n_38456) );
na02s01 g741779 ( .a(n_38425), .b(n_38402), .o(n_38403) );
na02s01 g741780 ( .a(n_38423), .b(n_38422), .o(n_38424) );
no02s01 g741781 ( .a(n_38400), .b(n_38399), .o(n_38401) );
na02s01 g741785 ( .a(n_38526), .b(n_39230), .o(n_38527) );
na02s01 g741786 ( .a(n_38510), .b(n_38483), .o(n_38511) );
no02s01 g741787 ( .a(n_38451), .b(n_38450), .o(n_38452) );
na02f06 g741788 ( .a(n_38344), .b(n_38113), .o(n_38369) );
ao12s01 g741789 ( .a(n_38332), .b(n_38397), .c(n_38281), .o(n_38427) );
in01m04 g741790 ( .a(n_38448), .o(n_38449) );
in01m04 g741791 ( .a(n_38421), .o(n_38448) );
na02f08 g741792 ( .a(n_38343), .b(n_38204), .o(n_38421) );
oa12s01 g741793 ( .a(n_38058), .b(n_38322), .c(n_38084), .o(n_38462) );
in01f02 g741794 ( .a(n_38446), .o(n_38447) );
oa12f04 g741795 ( .a(FE_OCP_RBN4062_n_44030), .b(n_38420), .c(n_38139), .o(n_38446) );
ao12s02 g741796 ( .a(n_38398), .b(n_38397), .c(n_38396), .o(n_38872) );
ao12s02 g741797 ( .a(n_38395), .b(n_38394), .c(n_38393), .o(n_38873) );
ao12s02 g741798 ( .a(n_38445), .b(n_38444), .c(n_38443), .o(n_38964) );
in01s01 g741799 ( .a(n_38493), .o(n_38516) );
ao12s01 g741800 ( .a(n_38392), .b(n_38391), .c(n_38390), .o(n_38493) );
in01s01 g741801 ( .a(FE_RN_1858_0), .o(n_39393) );
oa12s01 g741802 ( .a(n_38442), .b(n_38441), .c(n_38440), .o(n_38562) );
ao12s01 g741803 ( .a(n_38307), .b(n_38388), .c(n_38347), .o(n_38491) );
in01s01 g741804 ( .a(n_38344), .o(n_38455) );
oa12f04 g741805 ( .a(n_38188), .b(n_38288), .c(n_38169), .o(n_38344) );
no02s01 g741806 ( .a(n_38397), .b(n_38396), .o(n_38398) );
no02s01 g741807 ( .a(n_38394), .b(n_38393), .o(n_38395) );
no02s01 g741808 ( .a(n_38342), .b(n_38142), .o(n_38425) );
no02s01 g741809 ( .a(n_38321), .b(n_38121), .o(n_38400) );
no02s01 g741810 ( .a(n_38469), .b(n_38468), .o(n_38470) );
na02s01 g741811 ( .a(n_38484), .b(n_39232), .o(n_38485) );
na02s01 g741812 ( .a(n_38508), .b(n_38429), .o(n_38509) );
no02s02 g741813 ( .a(n_38444), .b(n_38443), .o(n_38445) );
no02s01 g741814 ( .a(n_38391), .b(n_38390), .o(n_38392) );
na02s01 g741815 ( .a(n_38441), .b(n_38440), .o(n_38442) );
na02f06 g741816 ( .a(n_38342), .b(n_38143), .o(n_38343) );
ao12s01 g741817 ( .a(n_38311), .b(n_38368), .c(n_38352), .o(n_38423) );
in01m02 g741818 ( .a(n_38418), .o(n_38419) );
na02s06 TIMEBOOST_cell_2890 ( .a(n_1969), .b(n_1968), .o(TIMEBOOST_net_736) );
oa22s01 g741820 ( .a(n_38368), .b(n_38376), .c(n_38285), .d(n_38377), .o(n_38908) );
oa12s02 g741821 ( .a(n_38367), .b(n_38366), .c(n_38365), .o(n_38890) );
oa12s02 g741823 ( .a(n_38439), .b(n_38438), .c(n_38437), .o(n_38930) );
in01s01 g741824 ( .a(n_38510), .o(n_38526) );
oa12s01 g741825 ( .a(n_38417), .b(n_38416), .c(n_38415), .o(n_38510) );
oa12s02 g741826 ( .a(n_38414), .b(n_38413), .c(n_38412), .o(n_38884) );
in01s01 g741827 ( .a(n_39324), .o(n_38467) );
ao12s01 g741828 ( .a(n_38387), .b(n_38386), .c(n_38385), .o(n_39324) );
in01s01 g741829 ( .a(n_38389), .o(n_38451) );
oa12s01 g741830 ( .a(n_38118), .b(n_38386), .c(n_38082), .o(n_38389) );
no02f06 g741831 ( .a(n_38288), .b(n_38116), .o(n_38342) );
na02s01 g741832 ( .a(n_38366), .b(n_38365), .o(n_38367) );
in01s01 g741833 ( .a(n_38321), .o(n_38322) );
no02s01 g741834 ( .a(n_38288), .b(n_38038), .o(n_38321) );
na02m08 TIMEBOOST_cell_2889 ( .a(n_2106), .b(TIMEBOOST_net_735), .o(n_2158) );
in01s01 g741836 ( .a(n_38388), .o(n_38441) );
in01s01 g741837 ( .a(n_38420), .o(n_38388) );
na02f08 g741838 ( .a(n_38340), .b(n_38219), .o(n_38420) );
na02s01 g741839 ( .a(n_38438), .b(n_38437), .o(n_38439) );
na02s01 g741840 ( .a(n_38416), .b(n_38415), .o(n_38417) );
na02s01 g741841 ( .a(n_38413), .b(n_38412), .o(n_38414) );
no02s01 g741842 ( .a(n_38386), .b(n_38385), .o(n_38387) );
ao12s01 g741843 ( .a(n_38063), .b(n_38363), .c(n_37940), .o(n_38397) );
ao12s01 g741844 ( .a(n_38255), .b(n_38363), .c(n_38316), .o(n_38394) );
in01s01 g741845 ( .a(n_38469), .o(n_38888) );
ao12s01 g741846 ( .a(n_38361), .b(n_38360), .c(n_38359), .o(n_38469) );
ao12s01 g741847 ( .a(n_38263), .b(n_38262), .c(n_38261), .o(n_38829) );
in01s01 g741848 ( .a(n_38495), .o(n_38436) );
ao12s02 g741849 ( .a(n_38364), .b(n_38363), .c(n_38362), .o(n_38495) );
in01s01 g741850 ( .a(n_38484), .o(n_38508) );
ao12s01 g741851 ( .a(n_38384), .b(n_38383), .c(n_38382), .o(n_38484) );
ao12s01 g741852 ( .a(n_38411), .b(n_38410), .c(n_38409), .o(n_38859) );
ao12s02 g741853 ( .a(n_38327), .b(n_38287), .c(n_38304), .o(n_38444) );
ao12s01 g741854 ( .a(n_38284), .b(n_38286), .c(n_38271), .o(n_38391) );
no02s01 g741855 ( .a(n_38363), .b(n_38362), .o(n_38364) );
no02s01 g741856 ( .a(n_38360), .b(n_38359), .o(n_38361) );
no02s01 g741857 ( .a(n_38262), .b(n_38261), .o(n_38263) );
no02s01 g741858 ( .a(n_38434), .b(n_38432), .o(n_38435) );
na02s01 g741859 ( .a(n_38434), .b(n_38432), .o(n_38433) );
no02s01 g741860 ( .a(n_38383), .b(n_38382), .o(n_38384) );
no02s01 g741861 ( .a(n_38410), .b(n_38409), .o(n_38411) );
ao12s01 g741862 ( .a(n_38296), .b(n_38243), .c(n_38309), .o(n_38438) );
no02s01 g741863 ( .a(n_38287), .b(n_38026), .o(n_38413) );
no02s01 g741864 ( .a(n_38286), .b(n_38166), .o(n_38386) );
in01s01 g741865 ( .a(n_38368), .o(n_38285) );
in01s01 g741866 ( .a(n_38288), .o(n_38368) );
oa12s01 g741868 ( .a(n_38014), .b(n_38190), .c(n_38016), .o(n_38366) );
na02f08 g741869 ( .a(n_38286), .b(n_38083), .o(n_38340) );
in01s01 g741870 ( .a(n_38862), .o(n_38466) );
oa12s01 g741871 ( .a(n_38381), .b(n_38380), .c(n_38379), .o(n_38862) );
in01s01 g741872 ( .a(n_38483), .o(n_39230) );
oa12s01 g741873 ( .a(n_38408), .b(n_38407), .c(n_38406), .o(n_38483) );
oa12s01 g741874 ( .a(n_38348), .b(n_38244), .c(n_38301), .o(n_38416) );
na02s01 g741875 ( .a(n_38205), .b(n_38122), .o(n_38363) );
no02s01 g741876 ( .a(n_38191), .b(n_38062), .o(n_38262) );
na02s01 g741877 ( .a(n_38380), .b(n_38379), .o(n_38381) );
na02s01 g741878 ( .a(n_38407), .b(n_38406), .o(n_38408) );
no02s01 g741879 ( .a(n_38244), .b(n_44034), .o(n_38287) );
ao12s01 g741881 ( .a(n_38238), .b(n_38338), .c(n_38283), .o(n_38360) );
no02f08 g741882 ( .a(n_38244), .b(n_38055), .o(n_38286) );
in01s01 g741883 ( .a(n_38468), .o(n_38405) );
ao12s01 g741884 ( .a(n_38339), .b(n_38338), .c(n_38337), .o(n_38468) );
in01s01 g741885 ( .a(n_38434), .o(n_38404) );
oa12s01 g741886 ( .a(n_38336), .b(n_38335), .c(n_38334), .o(n_38434) );
in01s01 g741887 ( .a(n_38430), .o(n_38431) );
ao12s01 g741888 ( .a(n_38357), .b(n_38356), .c(n_38355), .o(n_38430) );
in01s01 g741889 ( .a(n_39232), .o(n_38429) );
ao12s01 g741890 ( .a(n_38354), .b(n_38358), .c(n_38353), .o(n_39232) );
oa12s01 g741891 ( .a(n_38250), .b(n_38242), .c(n_38310), .o(n_38383) );
ao12s01 g741892 ( .a(n_37907), .b(n_38358), .c(n_38267), .o(n_38410) );
in01s01 g741893 ( .a(n_38190), .o(n_38191) );
na02s01 g741894 ( .a(n_38338), .b(n_37956), .o(n_38190) );
no02s01 g741895 ( .a(n_38338), .b(n_38337), .o(n_38339) );
na02s01 g741896 ( .a(n_38335), .b(n_38334), .o(n_38336) );
no02s01 g741897 ( .a(n_38356), .b(n_38355), .o(n_38357) );
no02s01 g741898 ( .a(n_38358), .b(n_38353), .o(n_38354) );
na02s01 g741899 ( .a(n_38242), .b(n_38010), .o(n_38243) );
in01s01 g741901 ( .a(n_38244), .o(n_38407) );
no02f06 g741902 ( .a(n_38172), .b(n_38091), .o(n_38244) );
oa12s02 g741903 ( .a(n_38127), .b(n_38126), .c(n_38125), .o(n_38892) );
oa12s01 g741904 ( .a(n_38260), .b(n_38320), .c(n_38228), .o(n_38380) );
no02f08 g741905 ( .a(n_38075), .b(n_37979), .o(n_38338) );
na02s01 g741906 ( .a(n_38126), .b(n_38125), .o(n_38127) );
na02s01 g741907 ( .a(n_38320), .b(n_38012), .o(n_38356) );
in01s01 g741908 ( .a(n_38242), .o(n_38358) );
na02s01 g741909 ( .a(n_38171), .b(n_38090), .o(n_38242) );
in01s01 g741911 ( .a(n_38432), .o(n_39181) );
oa12s01 g741912 ( .a(n_38319), .b(n_38170), .c(n_38317), .o(n_38432) );
oa12s01 g741913 ( .a(n_38232), .b(n_38170), .c(n_38254), .o(n_38335) );
na02s01 g741914 ( .a(n_38170), .b(n_38317), .o(n_38319) );
na02s01 g741915 ( .a(n_38145), .b(n_38208), .o(n_38320) );
na02s01 g741916 ( .a(n_38145), .b(n_38035), .o(n_38171) );
ao12f06 g741917 ( .a(n_37954), .b(n_38074), .c(n_38073), .o(n_38075) );
in01s01 g741918 ( .a(n_38146), .o(n_38147) );
ao12s01 g741919 ( .a(n_38072), .b(n_38074), .c(n_38071), .o(n_38146) );
oa12s01 g741920 ( .a(n_38073), .b(n_38074), .c(n_37941), .o(n_38126) );
no02m04 g741921 ( .a(n_38187), .b(n_38167), .o(n_38204) );
no02s01 g741922 ( .a(n_38074), .b(n_38071), .o(n_38072) );
in01s01 g741925 ( .a(n_38145), .o(n_38170) );
in01s01 g741926 ( .a(n_38124), .o(n_38145) );
oa12f04 g741927 ( .a(n_37972), .b(n_38092), .c(n_37887), .o(n_38124) );
in01s01 g741928 ( .a(n_38820), .o(n_38144) );
ao12s01 g741929 ( .a(n_38070), .b(n_38092), .c(n_38069), .o(n_38820) );
na02m02 g741930 ( .a(n_38186), .b(n_38219), .o(n_38220) );
no02s01 g741931 ( .a(n_38092), .b(n_38069), .o(n_38070) );
in01m04 g741932 ( .a(n_38187), .o(n_38188) );
na02f06 g741933 ( .a(n_38141), .b(n_44029), .o(n_38187) );
ao12f08 g741936 ( .a(n_37905), .b(n_37991), .c(n_37867), .o(n_38074) );
in01s01 g741937 ( .a(n_38067), .o(n_38068) );
ao12s01 g741938 ( .a(n_37990), .b(n_37991), .c(n_37989), .o(n_38067) );
na02m06 g741939 ( .a(n_38117), .b(n_38115), .o(n_38169) );
no02s03 g741940 ( .a(n_38114), .b(n_38111), .o(n_38143) );
in01s01 g741943 ( .a(n_38141), .o(n_38142) );
no02s02 TIMEBOOST_cell_7390 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_9_), .b(delay_xor_ln22_unr18_stage7_stallmux_q_10_), .o(TIMEBOOST_net_2326) );
no02s01 g741947 ( .a(n_37991), .b(n_37989), .o(n_37990) );
no02s02 g741948 ( .a(n_38110), .b(n_38167), .o(n_38168) );
na02s01 g741949 ( .a(n_38140), .b(n_38247), .o(n_38284) );
na02m04 g741950 ( .a(n_38090), .b(n_38041), .o(n_38091) );
oa12f06 g741951 ( .a(n_37842), .b(n_44036), .c(n_37881), .o(n_38092) );
no02m06 g741952 ( .a(n_38119), .b(n_38166), .o(n_38219) );
oa12s01 g741954 ( .a(n_37988), .b(n_44036), .c(n_37987), .o(n_38060) );
na02f04 TIMEBOOST_cell_8169 ( .a(TIMEBOOST_net_2715), .b(n_21148), .o(n_21344) );
na02s04 TIMEBOOST_cell_5647 ( .a(TIMEBOOST_net_1771), .b(n_6277), .o(n_6376) );
in01s02 g741957 ( .a(n_38185), .o(n_38186) );
no02s02 TIMEBOOST_cell_6698 ( .a(TIMEBOOST_net_2106), .b(n_8019), .o(n_8199) );
in01s01 g741959 ( .a(n_38166), .o(n_38140) );
na02m06 g741960 ( .a(n_47336), .b(n_38120), .o(n_38166) );
na02s04 g741961 ( .a(n_38118), .b(n_38053), .o(n_38119) );
na02s01 g741963 ( .a(n_44036), .b(n_37987), .o(n_37988) );
no02s01 g741964 ( .a(n_38042), .b(n_38229), .o(n_38260) );
in01m04 g741967 ( .a(n_38116), .o(n_38117) );
na02m08 g741968 ( .a(n_38039), .b(n_38033), .o(n_38116) );
in01m04 g741969 ( .a(n_38114), .o(n_38115) );
na02m06 g741970 ( .a(n_38089), .b(n_38037), .o(n_38114) );
na02s04 TIMEBOOST_cell_5649 ( .a(TIMEBOOST_net_1772), .b(FE_RN_1944_0), .o(n_46993) );
na02f08 TIMEBOOST_cell_8630 ( .a(n_39166), .b(n_39050), .o(TIMEBOOST_net_2802) );
ao12f08 g741975 ( .a(n_37833), .b(n_37917), .c(n_37866), .o(n_37991) );
oa12s01 g741976 ( .a(n_37919), .b(n_37918), .c(n_37917), .o(n_38791) );
ao12s01 g741977 ( .a(n_37952), .b(n_37951), .c(n_37950), .o(n_38817) );
no02m06 g741980 ( .a(n_38008), .b(n_38038), .o(n_38039) );
no02m04 g741981 ( .a(n_38036), .b(n_38005), .o(n_38037) );
no02s01 g741982 ( .a(n_38121), .b(n_38057), .o(n_38058) );
no02s01 g741983 ( .a(n_38062), .b(n_37980), .o(n_38014) );
na02s01 g741984 ( .a(n_38216), .b(n_38217), .o(n_38218) );
na02m04 g741985 ( .a(n_37984), .b(n_37983), .o(n_37985) );
na02s10 TIMEBOOST_cell_1938 ( .a(n_1398), .b(TIMEBOOST_net_583), .o(n_1533) );
na02m04 g741987 ( .a(n_37895), .b(n_37906), .o(n_37954) );
in01s02 g741990 ( .a(n_38108), .o(n_38109) );
no02s03 g741991 ( .a(n_38088), .b(FE_OCPN1056_n_38087), .o(n_38108) );
no02s01 g741992 ( .a(n_38378), .b(n_38329), .o(n_38454) );
na02s01 g741994 ( .a(n_38089), .b(n_37984), .o(n_38085) );
no02s01 g741995 ( .a(n_38333), .b(n_38313), .o(n_38402) );
in01s01 g741996 ( .a(n_38376), .o(n_38377) );
na02s01 g741997 ( .a(n_38352), .b(n_38312), .o(n_38376) );
no02s01 g741998 ( .a(n_38084), .b(n_38057), .o(n_38399) );
na02s01 g741999 ( .a(n_38283), .b(n_38237), .o(n_38337) );
no02s01 g742000 ( .a(n_38016), .b(n_37980), .o(n_38261) );
no02s01 g742001 ( .a(n_37979), .b(n_37896), .o(n_38125) );
no02s01 g742002 ( .a(n_38332), .b(n_38282), .o(n_38396) );
na02s01 g742003 ( .a(n_38316), .b(n_38256), .o(n_38362) );
in01s01 g742004 ( .a(n_38239), .o(n_38240) );
na02s01 g742005 ( .a(n_38181), .b(n_38216), .o(n_38239) );
na03m08 TIMEBOOST_cell_7138 ( .a(TIMEBOOST_net_1033), .b(n_18190), .c(n_17947), .o(n_18266) );
na02s02 g742007 ( .a(FE_OCP_RBN4061_n_44030), .b(n_47252), .o(n_38164) );
na02s01 g742008 ( .a(n_38073), .b(n_37906), .o(n_38071) );
na02s01 g742009 ( .a(n_37918), .b(n_37917), .o(n_37919) );
no02s01 g742010 ( .a(n_37951), .b(n_37950), .o(n_37952) );
in01s01 g742011 ( .a(n_38183), .o(n_38184) );
na02s02 TIMEBOOST_cell_6643 ( .a(n_33576), .b(n_33579), .o(TIMEBOOST_net_2079) );
in01s01 g742013 ( .a(n_38374), .o(n_38375) );
oa12s01 g742014 ( .a(n_38006), .b(n_38236), .c(n_37983), .o(n_38374) );
oa12s01 g742015 ( .a(n_38009), .b(n_38236), .c(n_37566), .o(n_38461) );
oa12s01 g742016 ( .a(n_37955), .b(n_38236), .c(n_37894), .o(n_38365) );
oa12s01 g742017 ( .a(n_37947), .b(n_38236), .c(n_37981), .o(n_38426) );
na02s06 g742018 ( .a(n_44035), .b(n_38004), .o(n_38055) );
in01s01 g742019 ( .a(n_38042), .o(n_38012) );
no02s04 g742020 ( .a(n_44872), .b(n_37911), .o(n_38042) );
in01s01 TIMEBOOST_cell_5903 ( .a(n_27131), .o(TIMEBOOST_net_1792) );
no02s02 g742022 ( .a(n_37908), .b(n_44866), .o(n_37976) );
in01s01 g742023 ( .a(n_38034), .o(n_38035) );
no03m04 TIMEBOOST_cell_8457 ( .a(FE_OCP_RBN1604_n_20995), .b(n_44158), .c(n_21153), .o(TIMEBOOST_net_2692) );
na02f04 g742026 ( .a(n_38010), .b(n_37943), .o(n_38011) );
no02s06 g742027 ( .a(n_38082), .b(n_44033), .o(n_38083) );
in01s01 g742028 ( .a(n_38138), .o(n_38139) );
na02s06 g742029 ( .a(n_38050), .b(FE_OCP_RBN6571_n_44875), .o(n_38138) );
na02s02 g742031 ( .a(n_38001), .b(n_44875), .o(n_38118) );
na02s02 g742032 ( .a(n_38000), .b(n_44875), .o(n_38053) );
in01s01 g742033 ( .a(n_38349), .o(n_38350) );
oa22s01 g742034 ( .a(n_38196), .b(n_37589), .c(n_38236), .d(n_37619), .o(n_38349) );
ao22s01 g742035 ( .a(n_38236), .b(n_37554), .c(n_38196), .d(n_37569), .o(n_38422) );
ao22s01 g742036 ( .a(n_38236), .b(n_37364), .c(n_38196), .d(n_37393), .o(n_38359) );
ao22s01 g742037 ( .a(n_38236), .b(n_37518), .c(n_38196), .d(n_37545), .o(n_38393) );
in01s01 g742038 ( .a(n_38258), .o(n_38259) );
oa22s01 g742039 ( .a(FE_OCP_RBN4133_n_38028), .b(n_37700), .c(n_37945), .d(n_37701), .o(n_38258) );
oa22s01 g742040 ( .a(n_38196), .b(n_37520), .c(n_38236), .d(n_37499), .o(n_38480) );
in01s01 g742041 ( .a(n_38214), .o(n_38215) );
na02f04 TIMEBOOST_cell_8786 ( .a(FE_OCP_RBN3013_n_14985), .b(FE_OCP_RBN2838_n_13962), .o(TIMEBOOST_net_2880) );
in01s01 g742043 ( .a(n_38201), .o(n_38202) );
no02f06 TIMEBOOST_cell_8072 ( .a(n_20337), .b(FE_OCP_RBN1844_n_20616), .o(TIMEBOOST_net_2667) );
in01s01 g742045 ( .a(n_38088), .o(n_38051) );
no02s02 g742046 ( .a(n_38028), .b(FE_OCP_RBN5556_n_37559), .o(n_38088) );
in01s01 g742047 ( .a(n_37984), .o(n_37949) );
na02s02 g742048 ( .a(n_37913), .b(n_37587), .o(n_37984) );
no02m02 g742049 ( .a(n_37900), .b(n_37948), .o(n_38057) );
in01s01 g742050 ( .a(n_37946), .o(n_37947) );
no02s02 g742051 ( .a(n_37904), .b(n_37544), .o(n_37946) );
in01s01 g742052 ( .a(n_37975), .o(n_38332) );
in01s01 g742054 ( .a(n_37895), .o(n_37896) );
na02s02 g742055 ( .a(n_37844), .b(n_37877), .o(n_37895) );
no02s02 g742056 ( .a(n_37904), .b(n_37877), .o(n_37979) );
na02s02 g742057 ( .a(n_37893), .b(n_37894), .o(n_37955) );
no02s02 g742058 ( .a(n_37904), .b(n_37385), .o(n_38016) );
in01s01 g742059 ( .a(n_38281), .o(n_38282) );
na02s01 g742061 ( .a(n_38196), .b(n_37912), .o(n_38281) );
no02s04 g742062 ( .a(n_37893), .b(n_37384), .o(n_37980) );
in01s01 g742063 ( .a(n_38008), .o(n_38009) );
no02m04 g742064 ( .a(n_37973), .b(n_37974), .o(n_38008) );
in01s01 g742065 ( .a(n_38033), .o(n_38084) );
na02m06 g742066 ( .a(n_38007), .b(n_37948), .o(n_38033) );
in01s01 g742068 ( .a(n_38005), .o(n_38006) );
no02m04 g742069 ( .a(n_37973), .b(n_37637), .o(n_38005) );
no02s01 g742070 ( .a(n_37945), .b(n_37559), .o(n_38087) );
no02f04 TIMEBOOST_cell_6637 ( .a(FE_RN_960_0), .b(n_23329), .o(TIMEBOOST_net_2076) );
no02s01 g742072 ( .a(n_38028), .b(n_38032), .o(n_38112) );
in01s01 g742073 ( .a(n_38328), .o(n_38329) );
na02s01 g742074 ( .a(n_38196), .b(n_38315), .o(n_38328) );
no02s01 g742075 ( .a(n_38196), .b(n_38315), .o(n_38378) );
in01s01 g742076 ( .a(n_38313), .o(n_38314) );
no02s01 g742077 ( .a(n_38236), .b(n_37618), .o(n_38313) );
no02s01 g742078 ( .a(n_38196), .b(n_37548), .o(n_38333) );
na02s01 g742079 ( .a(n_38236), .b(n_38279), .o(n_38352) );
in01s01 g742080 ( .a(n_38311), .o(n_38312) );
no02s01 g742081 ( .a(n_38236), .b(n_38279), .o(n_38311) );
in01s01 g742082 ( .a(n_38237), .o(n_38238) );
na02s01 g742083 ( .a(n_38196), .b(n_37392), .o(n_38237) );
na02s01 g742084 ( .a(n_37945), .b(n_37309), .o(n_38283) );
in01s01 g742085 ( .a(n_38255), .o(n_38256) );
no02s01 g742086 ( .a(n_38236), .b(n_38235), .o(n_38255) );
na02s01 g742087 ( .a(n_38236), .b(n_38235), .o(n_38316) );
na02s01 g742088 ( .a(FE_OCP_RBN4133_n_38028), .b(n_37597), .o(n_38216) );
in01s01 g742089 ( .a(n_38181), .o(n_38182) );
na02s01 g742090 ( .a(n_37945), .b(n_37760), .o(n_38181) );
na02s01 TIMEBOOST_cell_7065 ( .a(FE_OCP_RBN4483_n_11439), .b(FE_OCPN1218_n_11012), .o(TIMEBOOST_net_2291) );
no02s01 g742093 ( .a(n_37945), .b(FE_OCP_RBN5563_n_37551), .o(n_38102) );
in01s01 TIMEBOOST_cell_7376 ( .a(TIMEBOOST_net_2312), .o(rst) );
na02s01 TIMEBOOST_cell_6107 ( .a(n_42160), .b(n_42569), .o(TIMEBOOST_net_1905) );
no02m08 TIMEBOOST_cell_3336 ( .a(n_26985), .b(n_26354), .o(TIMEBOOST_net_959) );
no02s06 TIMEBOOST_cell_8679 ( .a(TIMEBOOST_net_2826), .b(n_36585), .o(n_36690) );
no03s40 TIMEBOOST_cell_2166 ( .a(FE_OCP_RBN7009_n_44962), .b(FE_RN_1646_0), .c(n_32731), .o(n_32659) );
no03s20 TIMEBOOST_cell_2167 ( .a(n_32600), .b(FE_OCP_RBN7006_n_44962), .c(n_32389), .o(n_32551) );
no02s02 TIMEBOOST_cell_1897 ( .a(n_16977), .b(FE_OCP_RBN6073_n_16086), .o(TIMEBOOST_net_563) );
no02f06 TIMEBOOST_cell_1853 ( .a(n_26799), .b(n_26692), .o(TIMEBOOST_net_541) );
in01s01 g742106 ( .a(n_38010), .o(n_37907) );
no02s01 TIMEBOOST_cell_8629 ( .a(TIMEBOOST_net_2801), .b(n_43362), .o(n_43617) );
na02s02 g742108 ( .a(n_37970), .b(n_37968), .o(n_38082) );
na03s01 TIMEBOOST_cell_7174 ( .a(n_14213), .b(n_14212), .c(n_14077), .o(n_14214) );
no03m04 TIMEBOOST_cell_8323 ( .a(n_44594), .b(FE_OCP_RBN2902_n_8902), .c(n_8988), .o(n_9240) );
na03m08 TIMEBOOST_cell_7293 ( .a(n_35334), .b(n_35234), .c(n_35353), .o(n_35428) );
in01m02 g742114 ( .a(n_38160), .o(n_38161) );
no02f08 TIMEBOOST_cell_5144 ( .a(n_14551), .b(n_14635), .o(TIMEBOOST_net_1520) );
in01s02 g742116 ( .a(n_38158), .o(n_38159) );
na02s02 g742117 ( .a(n_38135), .b(n_38134), .o(n_38158) );
in01s01 g742118 ( .a(n_38233), .o(n_38234) );
no02s02 g742119 ( .a(n_38180), .b(n_38213), .o(n_38233) );
no02s02 g742120 ( .a(n_38078), .b(n_38157), .o(n_38486) );
na02s02 g742121 ( .a(n_38179), .b(n_38199), .o(n_38200) );
na02m06 g742122 ( .a(n_37862), .b(n_37275), .o(n_38073) );
in01s01 g742124 ( .a(n_37906), .o(n_37941) );
na02s04 g742125 ( .a(n_37861), .b(n_37274), .o(n_37906) );
no02s01 g742126 ( .a(n_37868), .b(n_37905), .o(n_37989) );
no02s01 g742127 ( .a(n_38254), .b(n_38231), .o(n_38317) );
no02s01 g742128 ( .a(n_37891), .b(n_37809), .o(n_37951) );
na02s01 g742129 ( .a(n_37972), .b(n_37888), .o(n_38069) );
na02s01 g742130 ( .a(n_38227), .b(n_38230), .o(n_38355) );
no02s01 g742131 ( .a(n_38310), .b(n_38249), .o(n_38353) );
na02s01 g742132 ( .a(n_38297), .b(n_38277), .o(n_38409) );
no02s01 g742133 ( .a(n_38266), .b(n_38276), .o(n_38309) );
na02s01 g742134 ( .a(n_38348), .b(n_38302), .o(n_38406) );
no02s01 g742135 ( .a(n_38292), .b(n_38303), .o(n_38412) );
na02s02 g742136 ( .a(n_38120), .b(n_38291), .o(n_38327) );
no02s01 g742137 ( .a(n_38272), .b(n_38248), .o(n_38385) );
no02s01 g742138 ( .a(n_38324), .b(n_38373), .o(n_38450) );
na02s01 g742139 ( .a(n_38347), .b(n_38308), .o(n_38440) );
no02s01 g742141 ( .a(n_37945), .b(n_37590), .o(n_38167) );
in01s01 g742142 ( .a(n_37939), .o(n_37940) );
no02s04 g742143 ( .a(n_37904), .b(n_37519), .o(n_37939) );
no02m06 g742145 ( .a(n_37900), .b(n_37546), .o(n_38063) );
no02s06 g742146 ( .a(n_37900), .b(n_37391), .o(n_38062) );
no02s02 g742147 ( .a(n_37913), .b(n_37555), .o(n_38038) );
no02s02 g742148 ( .a(n_38028), .b(n_37568), .o(n_38111) );
no02s02 g742149 ( .a(n_37913), .b(n_37617), .o(n_38036) );
oa12s01 g742150 ( .a(n_37945), .b(n_37574), .c(FE_OCP_RBN5563_n_37551), .o(n_38156) );
oa12s01 g742151 ( .a(FE_OCP_RBN4133_n_38028), .b(n_37556), .c(n_37551), .o(n_38217) );
in01s01 g742152 ( .a(n_38153), .o(n_38154) );
no02s03 TIMEBOOST_cell_4061 ( .a(n_10517), .b(n_10364), .o(TIMEBOOST_net_1121) );
in01s01 g742154 ( .a(n_38197), .o(n_38198) );
no02s02 g742155 ( .a(n_38157), .b(n_38130), .o(n_38197) );
oa12f08 g742156 ( .a(n_37810), .b(n_37863), .c(n_37832), .o(n_37917) );
ao12s01 g742157 ( .a(n_37865), .b(n_37864), .c(n_37863), .o(n_38764) );
oa12s01 g742158 ( .a(n_37846), .b(n_37853), .c(n_37845), .o(n_38799) );
oa22s01 g742159 ( .a(FE_OCP_RBN2549_n_44881), .b(n_37398), .c(n_44887), .d(n_37910), .o(n_38334) );
oa12s01 g742160 ( .a(n_38253), .b(FE_OCP_RBN2549_n_44881), .c(n_38251), .o(n_38379) );
ao12s01 g742161 ( .a(n_37892), .b(n_44887), .c(n_37852), .o(n_38382) );
oa12s01 g742162 ( .a(n_38295), .b(FE_OCP_RBN2549_n_44881), .c(n_38293), .o(n_38437) );
oa12s01 g742163 ( .a(n_38300), .b(FE_OCP_RBN2549_n_44881), .c(n_38298), .o(n_38415) );
ao12s01 g742164 ( .a(n_38003), .b(n_44887), .c(n_37935), .o(n_38443) );
ao12s01 g742165 ( .a(n_38274), .b(n_44887), .c(n_38273), .o(n_38390) );
ao12s01 g742166 ( .a(n_38326), .b(n_44887), .c(n_38325), .o(n_38501) );
oa12s01 g742167 ( .a(n_38306), .b(FE_OCP_RBN2549_n_44881), .c(FE_OCP_RBN4026_n_37577), .o(n_38490) );
in01s01 g742168 ( .a(n_38211), .o(n_38212) );
oa22s01 g742169 ( .a(FE_OCP_RBN6575_n_44875), .b(n_37838), .c(FE_OCP_RBN6574_n_44875), .d(n_37823), .o(n_38211) );
in01s01 g742172 ( .a(n_38307), .o(n_38308) );
no02s01 g742174 ( .a(n_44887), .b(n_38270), .o(n_38307) );
na02s01 g742176 ( .a(FE_OCP_RBN2549_n_44881), .b(FE_OCP_RBN4026_n_37577), .o(n_38306) );
in01s02 g742177 ( .a(n_38303), .o(n_38304) );
na02s01 TIMEBOOST_cell_3342 ( .a(n_5876), .b(n_5659), .o(TIMEBOOST_net_962) );
no02s01 g742179 ( .a(n_44887), .b(n_38269), .o(n_38303) );
no02s02 g742180 ( .a(n_44867), .b(n_37935), .o(n_38003) );
in01s01 g742181 ( .a(n_38301), .o(n_38302) );
no02s01 g742183 ( .a(n_44887), .b(n_38268), .o(n_38301) );
na02s01 g742185 ( .a(FE_OCP_RBN2549_n_44881), .b(n_38298), .o(n_38300) );
in01s01 g742186 ( .a(n_38231), .o(n_38232) );
na02s01 TIMEBOOST_cell_6631 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_23_), .o(TIMEBOOST_net_2073) );
no02s01 g742188 ( .a(FE_OCP_RBN2549_n_44881), .b(n_37875), .o(n_38231) );
in01s01 g742189 ( .a(n_38229), .o(n_38230) );
no02m02 TIMEBOOST_cell_1822 ( .a(TIMEBOOST_net_525), .b(n_31400), .o(FE_RN_2675_0) );
no02s01 g742191 ( .a(FE_OCP_RBN2549_n_44881), .b(n_38209), .o(n_38229) );
in01s01 g742192 ( .a(n_38276), .o(n_38277) );
na03m08 TIMEBOOST_cell_8312 ( .a(n_16070), .b(FE_OCP_RBN4204_n_13796), .c(TIMEBOOST_net_651), .o(n_14547) );
no02s01 g742194 ( .a(FE_OCP_RBN2549_n_44881), .b(n_37871), .o(n_38276) );
no02f08 TIMEBOOST_cell_5481 ( .a(TIMEBOOST_net_1688), .b(n_35157), .o(n_35293) );
na02s01 g742196 ( .a(FE_OCP_RBN2549_n_44881), .b(n_38251), .o(n_38253) );
in01s01 g742197 ( .a(n_38227), .o(n_38228) );
na02s01 g742199 ( .a(FE_OCP_RBN2549_n_44881), .b(n_38209), .o(n_38227) );
na02s06 g742200 ( .a(n_44877), .b(n_37869), .o(n_37972) );
in01s01 g742201 ( .a(n_37887), .o(n_37888) );
no02s02 g742202 ( .a(n_44869), .b(n_37869), .o(n_37887) );
no02f08 g742203 ( .a(n_37853), .b(n_37808), .o(n_37891) );
in01s01 g742204 ( .a(n_38296), .o(n_38297) );
na02s01 TIMEBOOST_cell_6829 ( .a(n_31476), .b(n_30906), .o(TIMEBOOST_net_2172) );
no02s01 g742206 ( .a(n_44887), .b(n_37884), .o(n_38296) );
no02m04 g742207 ( .a(n_44867), .b(n_37882), .o(n_37883) );
na02s01 g742208 ( .a(FE_OCP_RBN2549_n_44881), .b(n_38293), .o(n_38295) );
no02f06 g742209 ( .a(n_44920), .b(n_37852), .o(n_37892) );
in01s01 g742210 ( .a(n_38249), .o(n_38250) );
no02f10 TIMEBOOST_cell_3331 ( .a(n_31974), .b(TIMEBOOST_net_956), .o(n_32081) );
no02s01 g742212 ( .a(n_44887), .b(n_37849), .o(n_38249) );
na02s02 g742213 ( .a(n_44877), .b(n_37969), .o(n_37970) );
no02s01 g742214 ( .a(n_44887), .b(n_38273), .o(n_38274) );
in01s01 g742215 ( .a(n_38271), .o(n_38272) );
na02s02 g742216 ( .a(n_44877), .b(n_37967), .o(n_37968) );
na02s01 g742217 ( .a(FE_OCP_RBN2549_n_44881), .b(n_37967), .o(n_38271) );
no02s01 g742219 ( .a(n_44887), .b(n_38325), .o(n_38326) );
in01s01 g742220 ( .a(n_38323), .o(n_38324) );
na02s01 g742222 ( .a(FE_OCP_RBN2549_n_44881), .b(n_38290), .o(n_38323) );
in01s01 TIMEBOOST_cell_8900 ( .a(n_1014), .o(TIMEBOOST_net_2944) );
no02f08 TIMEBOOST_cell_5143 ( .a(TIMEBOOST_net_1519), .b(n_38602), .o(n_38690) );
na02f02 TIMEBOOST_cell_4481 ( .a(n_39643), .b(n_39657), .o(TIMEBOOST_net_1331) );
na02s01 g742226 ( .a(n_44887), .b(n_38270), .o(n_38347) );
in01s01 g742227 ( .a(n_38291), .o(n_38292) );
na02s01 g742229 ( .a(n_44887), .b(n_38269), .o(n_38291) );
in01s01 g742230 ( .a(n_38247), .o(n_38248) );
na02f08 TIMEBOOST_cell_8075 ( .a(TIMEBOOST_net_2668), .b(n_20683), .o(n_20846) );
na02s01 g742232 ( .a(n_44887), .b(n_37929), .o(n_38247) );
in01s01 TIMEBOOST_cell_7375 ( .a(TIMEBOOST_net_2310), .o(TIMEBOOST_net_2311) );
no02s01 g742234 ( .a(FE_OCP_RBN2549_n_44881), .b(n_38290), .o(n_38373) );
no02s02 g742235 ( .a(FE_OCP_RBN6571_n_44875), .b(n_37654), .o(n_38131) );
no02f04 TIMEBOOST_cell_4060 ( .a(TIMEBOOST_net_1120), .b(FE_OCP_RBN3277_n_5284), .o(n_5456) );
na02s01 g742237 ( .a(FE_OCP_RBN6572_n_44875), .b(n_38047), .o(n_38135) );
in01s01 g742238 ( .a(n_38078), .o(n_38134) );
no02s02 g742239 ( .a(FE_OCP_RBN6572_n_44875), .b(n_38047), .o(n_38078) );
no02s01 g742240 ( .a(FE_OCP_RBN4059_n_44875), .b(n_37692), .o(n_38130) );
no02s01 g742241 ( .a(FE_OCP_RBN6575_n_44875), .b(n_37697), .o(n_38157) );
no02s02 g742242 ( .a(FE_OCP_RBN6575_n_44875), .b(FE_OCP_RBN4042_n_37707), .o(n_38213) );
in01s01 g742243 ( .a(n_38179), .o(n_38180) );
na02s02 g742244 ( .a(FE_OCP_RBN6575_n_44875), .b(FE_OCP_RBN4042_n_37707), .o(n_38179) );
no02m04 g742245 ( .a(n_37848), .b(n_37847), .o(n_37905) );
in01s01 g742246 ( .a(n_37867), .o(n_37868) );
na02s06 g742247 ( .a(n_37848), .b(n_37847), .o(n_37867) );
na02s01 g742248 ( .a(n_37834), .b(n_37866), .o(n_37918) );
no02s01 g742249 ( .a(n_37864), .b(n_37863), .o(n_37865) );
no02s01 g742250 ( .a(n_44887), .b(n_37334), .o(n_38254) );
na02s01 g742251 ( .a(n_37853), .b(n_37845), .o(n_37846) );
no02s01 g742252 ( .a(n_37843), .b(n_37881), .o(n_37987) );
no02s01 g742253 ( .a(FE_OCP_RBN2549_n_44881), .b(n_37352), .o(n_38310) );
na02s01 g742254 ( .a(n_44887), .b(n_38268), .o(n_38348) );
in01s01 g742255 ( .a(n_38266), .o(n_38267) );
no03s01 TIMEBOOST_cell_7219 ( .a(TIMEBOOST_net_2252), .b(n_15455), .c(n_44051), .o(n_15604) );
no02s01 g742257 ( .a(FE_OCP_RBN2549_n_44881), .b(n_37901), .o(n_38266) );
na02s06 TIMEBOOST_cell_8043 ( .a(TIMEBOOST_net_2652), .b(n_31847), .o(FE_RN_604_0) );
na02s01 g742259 ( .a(FE_OCP_RBN2549_n_44881), .b(n_37415), .o(n_38208) );
in01s01 g742260 ( .a(n_38120), .o(n_38026) );
na02s06 g742261 ( .a(n_44875), .b(n_37511), .o(n_38120) );
oa12s02 g742262 ( .a(FE_OCP_RBN6575_n_44875), .b(n_37697), .c(n_38047), .o(n_38199) );
in01m02 g742263 ( .a(n_37861), .o(n_37862) );
no02f04 TIMEBOOST_cell_7055 ( .a(n_19942), .b(n_19943), .o(TIMEBOOST_net_2286) );
oa12s01 g742265 ( .a(n_37820), .b(n_37819), .c(n_37818), .o(n_38731) );
in01s02 g742280 ( .a(n_38196), .o(n_38236) );
in01s01 g742282 ( .a(n_37945), .o(n_38196) );
in01s04 g742293 ( .a(n_37945), .o(n_38028) );
in01m08 g742294 ( .a(n_37904), .o(n_37945) );
in01m08 g742295 ( .a(n_37893), .o(n_37904) );
in01s08 g742298 ( .a(n_37973), .o(n_38007) );
in01s08 g742299 ( .a(n_37900), .o(n_37973) );
in01m08 g742300 ( .a(n_37913), .o(n_37900) );
in01m08 g742301 ( .a(n_37893), .o(n_37913) );
in01m08 g742302 ( .a(n_37844), .o(n_37893) );
oa12m08 g742303 ( .a(n_37783), .b(n_37838), .c(n_37795), .o(n_37844) );
in01s01 g742304 ( .a(n_37842), .o(n_37843) );
na02s04 g742305 ( .a(n_37837), .b(n_37836), .o(n_37842) );
no02m04 g742306 ( .a(n_37837), .b(n_37836), .o(n_37881) );
na02f06 g742307 ( .a(n_37815), .b(n_37778), .o(n_37835) );
no02s08 TIMEBOOST_cell_6594 ( .a(n_17192), .b(TIMEBOOST_net_2054), .o(n_17401) );
na02s02 TIMEBOOST_cell_4025 ( .a(n_4463), .b(n_4237), .o(TIMEBOOST_net_1103) );
in01s01 g742310 ( .a(n_37833), .o(n_37834) );
no02m04 g742311 ( .a(n_37822), .b(n_37821), .o(n_37833) );
na02m04 g742312 ( .a(n_37822), .b(n_37821), .o(n_37866) );
na02s01 g742313 ( .a(n_37819), .b(n_37818), .o(n_37820) );
no02s01 g742314 ( .a(n_37832), .b(n_37811), .o(n_37864) );
no02s01 g742315 ( .a(n_37831), .b(n_37816), .o(n_37950) );
ao12f08 g742359 ( .a(n_37704), .b(n_37782), .c(n_37701), .o(n_37850) );
oa12f06 g742360 ( .a(n_37777), .b(n_37817), .c(n_37757), .o(n_37853) );
ao12f06 g742362 ( .a(n_37767), .b(n_37818), .c(n_37799), .o(n_37863) );
ao12s01 g742363 ( .a(n_37798), .b(n_37797), .c(n_37796), .o(n_38713) );
ao12s01 g742364 ( .a(n_37807), .b(n_37806), .c(n_37817), .o(n_38752) );
na02m08 g742365 ( .a(n_37838), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37783) );
in01s01 g742366 ( .a(n_37815), .o(n_37816) );
na02f04 g742367 ( .a(n_37791), .b(n_37240), .o(n_37815) );
in01s01 g742368 ( .a(n_37916), .o(n_37831) );
na02m06 g742369 ( .a(n_37792), .b(n_37241), .o(n_37916) );
no02f04 g742370 ( .a(n_37801), .b(n_37800), .o(n_37832) );
in01s01 g742371 ( .a(n_37810), .o(n_37811) );
na02s04 g742372 ( .a(n_37801), .b(n_37800), .o(n_37810) );
na02s01 g742373 ( .a(n_37768), .b(n_37799), .o(n_37819) );
no02s01 g742374 ( .a(n_37797), .b(n_37796), .o(n_37798) );
no02s01 g742375 ( .a(n_37809), .b(n_37808), .o(n_37845) );
no02s01 g742376 ( .a(n_37817), .b(n_37806), .o(n_37807) );
in01m06 g742377 ( .a(n_37794), .o(n_37795) );
no02s08 TIMEBOOST_cell_7416 ( .a(n_17129), .b(TIMEBOOST_net_36), .o(TIMEBOOST_net_2339) );
na02m04 g742380 ( .a(n_37772), .b(n_37781), .o(n_37837) );
na02s04 g742381 ( .a(n_37769), .b(n_37746), .o(n_37822) );
oa12s01 g742382 ( .a(n_37766), .b(n_37765), .c(n_37764), .o(n_38738) );
no02s01 TIMEBOOST_cell_1835 ( .a(FE_OCP_RBN6024_n_30711), .b(n_31835), .o(TIMEBOOST_net_532) );
na02f08 g742384 ( .a(n_37780), .b(n_37753), .o(n_37782) );
na02s01 TIMEBOOST_cell_1741 ( .a(n_39163), .b(n_39319), .o(TIMEBOOST_net_485) );
na02s02 g742386 ( .a(n_37780), .b(n_37701), .o(n_37781) );
in01s01 g742387 ( .a(n_37778), .o(n_37809) );
na02m04 g742388 ( .a(n_37771), .b(n_37770), .o(n_37778) );
no02f04 g742389 ( .a(n_37771), .b(n_37770), .o(n_37808) );
na02s02 g742390 ( .a(n_37721), .b(n_37697), .o(n_37746) );
no02m02 TIMEBOOST_cell_4035 ( .a(n_19921), .b(n_19945), .o(TIMEBOOST_net_1108) );
na02f04 g742392 ( .a(n_37745), .b(n_37744), .o(n_37799) );
in01s01 g742393 ( .a(n_37767), .o(n_37768) );
no02f04 g742394 ( .a(n_37745), .b(n_37744), .o(n_37767) );
na02s01 g742395 ( .a(n_37758), .b(n_37777), .o(n_37806) );
na02s01 g742396 ( .a(n_37764), .b(n_37765), .o(n_37766) );
in01m02 g742397 ( .a(n_37775), .o(n_37776) );
in01m02 g742398 ( .a(n_37763), .o(n_37775) );
no02s02 TIMEBOOST_cell_8752 ( .a(FE_OCP_RBN2634_n_9003), .b(n_8195), .o(TIMEBOOST_net_2863) );
in01s02 g742400 ( .a(n_37791), .o(n_37792) );
na02s01 TIMEBOOST_cell_6032 ( .a(TIMEBOOST_net_1867), .b(n_47252), .o(n_38160) );
na02f06 g742402 ( .a(n_37759), .b(n_37738), .o(n_37817) );
in01s02 g742403 ( .a(n_37838), .o(n_37823) );
na02m10 g742404 ( .a(n_37722), .b(n_37708), .o(n_37838) );
oa12f06 g742405 ( .a(n_37664), .b(n_37762), .c(n_37663), .o(n_37818) );
na03m06 TIMEBOOST_cell_8311 ( .a(n_29616), .b(n_29596), .c(n_29634), .o(n_29672) );
ao12s01 g742407 ( .a(n_37740), .b(n_37762), .c(n_37739), .o(n_37797) );
no02m04 TIMEBOOST_cell_8800 ( .a(n_3602), .b(n_3542), .o(TIMEBOOST_net_2887) );
na03m06 TIMEBOOST_cell_8421 ( .a(n_5648), .b(n_45474), .c(n_6363), .o(n_6463) );
na03f06 TIMEBOOST_cell_8387 ( .a(TIMEBOOST_net_1983), .b(n_5614), .c(FE_OCP_RBN6098_n_5614), .o(n_5810) );
no02f02 g742412 ( .a(n_37720), .b(n_37649), .o(n_37723) );
na02m04 g742413 ( .a(n_37742), .b(n_37741), .o(n_37777) );
na02f04 g742414 ( .a(n_37764), .b(n_37737), .o(n_37759) );
in01s01 g742415 ( .a(n_37757), .o(n_37758) );
no02f04 g742416 ( .a(n_37742), .b(n_37741), .o(n_37757) );
na02m08 g742417 ( .a(n_37695), .b(n_37054), .o(n_37722) );
na02s08 g742418 ( .a(n_37694), .b(n_37055), .o(n_37708) );
no02s01 g742419 ( .a(n_37762), .b(n_37739), .o(n_37740) );
na02s01 g742420 ( .a(n_37737), .b(n_37738), .o(n_37765) );
oa12f04 g742422 ( .a(n_37709), .b(n_37703), .c(n_37667), .o(n_37753) );
no02f08 TIMEBOOST_cell_4034 ( .a(TIMEBOOST_net_1107), .b(FE_OCP_RBN6818_n_25997), .o(n_26190) );
no02s02 g742424 ( .a(n_37720), .b(n_37670), .o(n_37721) );
in01s02 g742427 ( .a(FE_OCP_RBN4040_n_37707), .o(n_37734) );
na02s02 TIMEBOOST_cell_1830 ( .a(TIMEBOOST_net_529), .b(n_31718), .o(n_31807) );
na02f04 g742430 ( .a(n_37668), .b(n_37696), .o(n_37745) );
in01s01 g742431 ( .a(n_38698), .o(n_38736) );
na02s01 TIMEBOOST_cell_1829 ( .a(n_31740), .b(n_31773), .o(TIMEBOOST_net_529) );
no02f06 TIMEBOOST_cell_5595 ( .a(TIMEBOOST_net_1745), .b(n_26019), .o(n_26167) );
na02m08 g742435 ( .a(n_37702), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37756) );
in01s04 g742436 ( .a(n_37670), .o(n_37671) );
no02m06 g742438 ( .a(n_37649), .b(n_37709), .o(n_37670) );
na02s06 g742439 ( .a(n_37658), .b(n_36948), .o(n_37738) );
na02f02 g742440 ( .a(n_37657), .b(FE_OCPN1622_n_36947), .o(n_37737) );
na02f02 g742441 ( .a(n_37693), .b(FE_OCP_RBN2498_n_37624), .o(n_37696) );
oa12m02 g742442 ( .a(n_37624), .b(n_37646), .c(n_37645), .o(n_37668) );
no03s06 TIMEBOOST_cell_8409 ( .a(n_5310), .b(n_5426), .c(FE_RN_1929_0), .o(n_47001) );
no02s02 TIMEBOOST_cell_5379 ( .a(TIMEBOOST_net_1637), .b(n_3472), .o(n_3989) );
in01m06 g742445 ( .a(n_37694), .o(n_37695) );
no02s02 TIMEBOOST_cell_4525 ( .a(n_25697), .b(n_25627), .o(TIMEBOOST_net_1353) );
na02f08 g742450 ( .a(n_37693), .b(n_37628), .o(n_37720) );
no02m06 TIMEBOOST_cell_4021 ( .a(n_34981), .b(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(TIMEBOOST_net_1101) );
oa12f04 g742452 ( .a(n_37715), .b(n_37716), .c(n_37687), .o(n_37764) );
in01s02 g742455 ( .a(n_37697), .o(n_37692) );
na02m08 g742456 ( .a(n_37583), .b(n_37607), .o(n_37697) );
na02f04 g742457 ( .a(n_37665), .b(n_37647), .o(n_37762) );
no02f04 TIMEBOOST_cell_6731 ( .a(TIMEBOOST_net_1922), .b(n_15083), .o(TIMEBOOST_net_2123) );
no03f02 TIMEBOOST_cell_2530 ( .a(n_14051), .b(n_14104), .c(n_14121), .o(n_14122) );
no02s06 g742462 ( .a(n_37686), .b(n_37709), .o(n_37704) );
no02f08 g742465 ( .a(n_37667), .b(n_37709), .o(n_37690) );
no04m20 TIMEBOOST_cell_6406 ( .a(n_32600), .b(n_32599), .c(n_32602), .d(n_32601), .o(n_32617) );
ao12m02 g742467 ( .a(n_37551), .b(n_37644), .c(n_37604), .o(n_37648) );
na02m06 g742468 ( .a(n_37606), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37628) );
na02f02 g742469 ( .a(n_37646), .b(n_37623), .o(n_37647) );
na02f02 g742470 ( .a(n_37626), .b(n_37598), .o(n_37665) );
na02s03 g742471 ( .a(n_37662), .b(FE_OCPN1624_n_37661), .o(n_37664) );
no02s04 g742472 ( .a(n_37662), .b(FE_OCPN1661_n_37661), .o(n_37663) );
in01s01 g742473 ( .a(n_37732), .o(n_37733) );
na02s01 g742474 ( .a(n_37688), .b(n_37715), .o(n_37732) );
in01m02 g742475 ( .a(n_37755), .o(n_37689) );
no02s02 TIMEBOOST_cell_1724 ( .a(TIMEBOOST_net_476), .b(n_20404), .o(n_20466) );
no02f08 g742478 ( .a(n_37646), .b(n_37645), .o(n_37693) );
in01s02 g742479 ( .a(n_37657), .o(n_37658) );
in01s01 g742481 ( .a(n_37649), .o(n_38047) );
no02m02 TIMEBOOST_cell_1821 ( .a(n_31074), .b(FE_OCP_RBN6843_n_31194), .o(TIMEBOOST_net_525) );
oa22s01 g742483 ( .a(FE_OCP_RBN4025_n_37577), .b(n_36686), .c(FE_OCP_RBN4026_n_37577), .d(n_37625), .o(n_38685) );
in01m04 g742484 ( .a(n_37702), .o(n_37703) );
no02m02 TIMEBOOST_cell_1806 ( .a(TIMEBOOST_net_517), .b(n_21713), .o(n_21768) );
no02f08 TIMEBOOST_cell_8831 ( .a(TIMEBOOST_net_2902), .b(TIMEBOOST_net_882), .o(n_25874) );
na02m08 TIMEBOOST_cell_2140 ( .a(TIMEBOOST_net_684), .b(n_44356), .o(n_11914) );
no02s20 TIMEBOOST_cell_8699 ( .a(TIMEBOOST_net_2836), .b(n_28092), .o(n_27964) );
no02f04 TIMEBOOST_cell_4012 ( .a(n_20314), .b(TIMEBOOST_net_1096), .o(n_20412) );
in01f01 g742490 ( .a(n_37646), .o(n_37626) );
no02f08 g742491 ( .a(n_37577), .b(n_37709), .o(n_37646) );
no02f06 g742492 ( .a(n_37578), .b(n_37709), .o(n_37645) );
in01s01 g742493 ( .a(n_37687), .o(n_37688) );
no02f04 g742494 ( .a(n_37656), .b(n_37655), .o(n_37687) );
na02f04 g742495 ( .a(n_37656), .b(n_37655), .o(n_37715) );
in01s01 g742498 ( .a(n_37662), .o(n_37796) );
na02s04 g742499 ( .a(FE_OCP_RBN4023_n_37577), .b(n_37625), .o(n_37662) );
no03f04 TIMEBOOST_cell_6539 ( .a(n_4321), .b(n_4490), .c(n_4894), .o(n_5077) );
in01s06 g742501 ( .a(n_37700), .o(n_37701) );
in01s06 g742504 ( .a(n_37686), .o(n_37700) );
ao22s08 g742505 ( .a(n_37594), .b(n_37087), .c(n_37593), .d(n_37086), .o(n_37686) );
na03m10 TIMEBOOST_cell_7133 ( .a(n_28283), .b(n_28249), .c(n_28089), .o(n_28343) );
in01s01 g742509 ( .a(n_37653), .o(n_37654) );
in01s01 g742510 ( .a(FE_OCP_RBN2498_n_37624), .o(n_37653) );
in01f02 g742512 ( .a(n_37606), .o(n_37624) );
no02m04 g742514 ( .a(n_37515), .b(n_37514), .o(n_37516) );
na02s10 g742515 ( .a(n_37515), .b(n_37069), .o(n_37563) );
in01s02 g742516 ( .a(n_37604), .o(n_37605) );
in01f02 g742518 ( .a(n_37601), .o(n_37602) );
na02m02 g742519 ( .a(n_37581), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37604) );
na02f02 g742520 ( .a(n_37581), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37601) );
na02s01 TIMEBOOST_cell_5410 ( .a(n_43265), .b(n_43187), .o(TIMEBOOST_net_1653) );
na02s04 g742522 ( .a(n_37535), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37560) );
oa12f06 g742526 ( .a(n_37557), .b(n_37559), .c(n_37709), .o(n_37579) );
ao12f04 g742527 ( .a(n_37531), .b(FE_OCP_RBN5558_n_37559), .c(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37644) );
in01m02 g742532 ( .a(n_37598), .o(n_37623) );
in01m02 g742533 ( .a(n_37578), .o(n_37598) );
no02f04 g742534 ( .a(n_37494), .b(n_37512), .o(n_37578) );
in01s02 g742535 ( .a(n_37760), .o(n_37622) );
in01s01 g742537 ( .a(n_37597), .o(n_37760) );
in01s04 g742538 ( .a(n_37597), .o(n_37596) );
na02m08 g742539 ( .a(n_37513), .b(n_37536), .o(n_37597) );
na02f06 g742546 ( .a(n_37576), .b(n_37558), .o(n_37656) );
oa12m06 g742548 ( .a(n_37155), .b(n_37467), .c(n_37350), .o(n_37513) );
na02f06 TIMEBOOST_cell_2142 ( .a(TIMEBOOST_net_685), .b(n_36510), .o(n_36588) );
ao12f02 g742550 ( .a(n_37124), .b(n_37446), .c(n_37258), .o(n_37494) );
no02m06 g742552 ( .a(n_37527), .b(n_37709), .o(n_37659) );
na02f04 g742553 ( .a(FE_OCP_RBN5557_n_37559), .b(n_37557), .o(n_37558) );
na02f04 g742554 ( .a(n_37531), .b(n_37559), .o(n_37576) );
na02s01 g742555 ( .a(n_38298), .b(n_37411), .o(n_37511) );
oa12f08 g742557 ( .a(n_37273), .b(n_37421), .c(FE_OCP_DRV_N6261_n_37471), .o(n_37509) );
in01s01 g742558 ( .a(n_37638), .o(n_37639) );
na02s01 g742559 ( .a(n_37619), .b(n_37618), .o(n_37638) );
no02s01 g742560 ( .a(n_37619), .b(n_37618), .o(n_37617) );
in01s06 g742561 ( .a(n_37593), .o(n_37594) );
no02f08 TIMEBOOST_cell_3385 ( .a(TIMEBOOST_net_983), .b(n_40089), .o(n_40090) );
in01s01 g742564 ( .a(n_37575), .o(n_38032) );
in01f01 g742565 ( .a(n_37581), .o(n_37575) );
in01s02 g742570 ( .a(n_37556), .o(n_37574) );
in01s01 g742571 ( .a(n_37535), .o(n_37556) );
in01f02 g742572 ( .a(n_37535), .o(n_37534) );
oa12s02 g742574 ( .a(n_37508), .b(n_37507), .c(n_37506), .o(n_38270) );
oa12s01 g742576 ( .a(n_37470), .b(n_37469), .c(n_37468), .o(n_37935) );
in01s01 g742577 ( .a(n_37969), .o(n_38273) );
ao12s01 g742578 ( .a(n_37433), .b(n_37432), .c(n_37431), .o(n_37969) );
in01s01 g742579 ( .a(n_37493), .o(n_38290) );
oa12s01 g742580 ( .a(n_37430), .b(n_37429), .c(n_37428), .o(n_37493) );
in01s01 g742581 ( .a(n_37637), .o(n_37983) );
oa12s02 g742582 ( .a(n_37573), .b(n_37572), .c(n_37571), .o(n_37637) );
in01s01 g742583 ( .a(n_37636), .o(n_38668) );
oa22s01 g742584 ( .a(n_37499), .b(n_37504), .c(n_37520), .d(n_36768), .o(n_37636) );
in01s01 g742585 ( .a(n_37965), .o(n_38325) );
ao22s01 g742586 ( .a(n_37460), .b(n_37061), .c(n_37459), .d(n_37062), .o(n_37965) );
no02s03 TIMEBOOST_cell_1803 ( .a(n_11146), .b(n_44511), .o(TIMEBOOST_net_516) );
na02s01 g742588 ( .a(n_37469), .b(n_37468), .o(n_37470) );
no02s01 g742589 ( .a(n_37432), .b(n_37431), .o(n_37433) );
na02s01 g742590 ( .a(n_37572), .b(n_37571), .o(n_37573) );
na02s01 g742591 ( .a(n_37507), .b(n_37506), .o(n_37508) );
in01f04 g742592 ( .a(n_37557), .o(n_37531) );
na02f08 g742594 ( .a(n_37505), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37557) );
na02s01 g742595 ( .a(n_37429), .b(n_37428), .o(n_37430) );
in01s01 g742596 ( .a(n_37716), .o(n_37529) );
na02m01 g742597 ( .a(n_37505), .b(n_37504), .o(n_37716) );
no02s01 g742599 ( .a(n_37520), .b(n_38315), .o(n_37590) );
no02s01 g742600 ( .a(n_37554), .b(n_38279), .o(n_37555) );
no02s01 g742601 ( .a(n_37547), .b(n_37499), .o(n_37568) );
no02f08 g742606 ( .a(n_37451), .b(n_37427), .o(n_37559) );
in01m02 g742610 ( .a(n_37527), .o(n_37551) );
na02s01 TIMEBOOST_cell_6868 ( .a(TIMEBOOST_net_2192), .b(n_32426), .o(n_32557) );
in01m02 g742612 ( .a(n_46952), .o(n_37492) );
oa12s01 g742614 ( .a(n_37466), .b(n_37465), .c(n_37464), .o(n_38269) );
in01s01 g742615 ( .a(n_38298), .o(n_37490) );
ao12s01 g742616 ( .a(n_37425), .b(n_37424), .c(n_37423), .o(n_38298) );
in01s01 g742617 ( .a(n_37929), .o(n_37967) );
oa12s01 g742618 ( .a(n_37404), .b(n_37403), .c(n_37402), .o(n_37929) );
in01s01 g742619 ( .a(n_37619), .o(n_37589) );
ao12s01 g742620 ( .a(n_37526), .b(n_37525), .c(n_37524), .o(n_37619) );
oa12s01 g742622 ( .a(n_37523), .b(n_37522), .c(n_37521), .o(n_37587) );
in01s01 g742623 ( .a(n_37974), .o(n_37566) );
oa12s02 g742624 ( .a(n_37502), .b(n_37501), .c(n_37500), .o(n_37974) );
in01s04 g742625 ( .a(n_37488), .o(n_37489) );
in01m04 g742626 ( .a(n_37467), .o(n_37488) );
ao12m04 g742628 ( .a(n_37153), .b(n_37373), .c(n_37296), .o(n_37427) );
na02f04 TIMEBOOST_cell_7904 ( .a(n_20553), .b(n_20642), .o(TIMEBOOST_net_2583) );
oa12f06 g742631 ( .a(n_37316), .b(n_37399), .c(n_37426), .o(n_37449) );
no02s01 g742632 ( .a(n_37413), .b(n_37233), .o(n_37507) );
no02s01 g742633 ( .a(n_37424), .b(n_37423), .o(n_37425) );
na02s01 g742634 ( .a(n_37403), .b(n_37402), .o(n_37404) );
no02s01 g742635 ( .a(n_37525), .b(n_37524), .o(n_37526) );
na02s02 g742636 ( .a(n_37501), .b(n_37500), .o(n_37502) );
na02s01 g742637 ( .a(n_37522), .b(n_37521), .o(n_37523) );
na02s01 g742639 ( .a(n_37465), .b(n_37464), .o(n_37466) );
na02m06 TIMEBOOST_cell_7771 ( .a(TIMEBOOST_net_2516), .b(n_42173), .o(n_42189) );
no02f02 TIMEBOOST_cell_1814 ( .a(TIMEBOOST_net_521), .b(n_45332), .o(n_16161) );
in01f02 g742642 ( .a(n_37446), .o(n_37447) );
na02m08 g742643 ( .a(FE_OCP_RBN6550_n_37377), .b(n_37419), .o(n_37421) );
na02m04 g742644 ( .a(FE_OCP_RBN6549_n_37377), .b(n_37419), .o(n_37446) );
in01f02 g742645 ( .a(n_37461), .o(n_37462) );
na02m02 TIMEBOOST_cell_8024 ( .a(n_16555), .b(n_16556), .o(TIMEBOOST_net_2643) );
no02s01 g742647 ( .a(n_37852), .b(n_37849), .o(n_37901) );
in01s01 g742648 ( .a(n_37459), .o(n_37460) );
no02s04 TIMEBOOST_cell_1712 ( .a(TIMEBOOST_net_470), .b(FE_OCP_RBN6006_n_15704), .o(n_15858) );
ao12s01 g742650 ( .a(n_37199), .b(n_37380), .c(n_37375), .o(n_37429) );
ao12s01 g742651 ( .a(n_37255), .b(n_37455), .c(n_37095), .o(n_37572) );
ao12s01 g742652 ( .a(n_37011), .b(n_37371), .c(n_37133), .o(n_37469) );
in01s01 g742656 ( .a(n_37499), .o(n_37520) );
in01s01 g742657 ( .a(n_37505), .o(n_37499) );
na02f06 g742658 ( .a(n_37418), .b(n_37401), .o(n_37505) );
ao12s01 g742659 ( .a(n_37196), .b(n_37380), .c(n_36963), .o(n_37432) );
in01s01 g742660 ( .a(n_37618), .o(n_37548) );
ao12s01 g742661 ( .a(n_37484), .b(n_37483), .c(n_37482), .o(n_37618) );
in01s01 g742662 ( .a(n_37554), .o(n_37569) );
ao12s01 g742663 ( .a(n_37458), .b(n_37457), .c(n_37456), .o(n_37554) );
ao12s01 g742664 ( .a(n_37498), .b(n_37497), .c(n_37496), .o(n_37948) );
in01s01 g742665 ( .a(n_37547), .o(n_38315) );
ao12s01 g742666 ( .a(n_37487), .b(n_37486), .c(n_37485), .o(n_37547) );
no02f04 TIMEBOOST_cell_3285 ( .a(TIMEBOOST_net_933), .b(n_26688), .o(n_26795) );
na02s10 TIMEBOOST_cell_8608 ( .a(n_23486), .b(FE_OCP_RBN4392_n_26146), .o(TIMEBOOST_net_2791) );
no02s02 TIMEBOOST_cell_1692 ( .a(TIMEBOOST_net_460), .b(n_3508), .o(n_5447) );
no02s01 g742670 ( .a(n_37380), .b(n_37188), .o(n_37403) );
in01s02 g742671 ( .a(n_37416), .o(n_37417) );
na02s04 g742672 ( .a(n_37399), .b(n_37278), .o(n_37416) );
na02s01 g742673 ( .a(n_37372), .b(n_37135), .o(n_37465) );
no02s01 g742674 ( .a(n_37457), .b(n_37456), .o(n_37458) );
no02s01 g742675 ( .a(n_37486), .b(n_37485), .o(n_37487) );
na02s01 g742676 ( .a(n_37454), .b(n_37270), .o(n_37522) );
no02s01 g742677 ( .a(n_37497), .b(n_37496), .o(n_37498) );
oa12s01 g742678 ( .a(n_37075), .b(n_37379), .c(n_36960), .o(n_37424) );
in01s01 g742679 ( .a(n_37414), .o(n_37415) );
no02s02 g742680 ( .a(n_37398), .b(n_37875), .o(n_37414) );
no02s01 g742681 ( .a(n_37483), .b(n_37482), .o(n_37484) );
no02s02 g742682 ( .a(n_37518), .b(n_38235), .o(n_37519) );
no02s04 g742683 ( .a(n_37545), .b(n_37452), .o(n_37546) );
ao12s02 g742684 ( .a(n_37107), .b(n_37407), .c(n_37148), .o(n_37501) );
in01s01 g742686 ( .a(n_37412), .o(n_37413) );
in01m06 g742687 ( .a(FE_OCP_RBN6550_n_37377), .o(n_37412) );
na02f08 g742689 ( .a(n_37380), .b(n_37185), .o(n_37377) );
no02m04 TIMEBOOST_cell_1678 ( .a(TIMEBOOST_net_453), .b(n_26156), .o(n_26157) );
in01s01 g742691 ( .a(n_37411), .o(n_38268) );
ao22s01 g742692 ( .a(n_37379), .b(n_37123), .c(n_37317), .d(n_37122), .o(n_37411) );
in01s01 g742693 ( .a(n_37889), .o(n_38251) );
oa12s01 g742694 ( .a(n_37356), .b(n_37355), .c(n_37354), .o(n_37889) );
in01s01 g742695 ( .a(n_37871), .o(n_37884) );
ao12s01 g742696 ( .a(n_37324), .b(n_37323), .c(n_37322), .o(n_37871) );
oa12s02 g742697 ( .a(n_37327), .b(n_37326), .c(n_37325), .o(n_37852) );
no02f02 TIMEBOOST_cell_1707 ( .a(n_20186), .b(n_20125), .o(TIMEBOOST_net_468) );
in01s02 g742699 ( .a(n_37544), .o(n_37981) );
oa12s02 g742700 ( .a(n_37481), .b(n_37480), .c(n_37479), .o(n_37544) );
in01s01 g742701 ( .a(n_37882), .o(n_38293) );
oa22s01 g742702 ( .a(n_37348), .b(n_37064), .c(n_37349), .d(n_37063), .o(n_37882) );
in01m02 g742703 ( .a(n_37373), .o(n_37374) );
no02s01 g742705 ( .a(n_37397), .b(n_37098), .o(n_37410) );
no02s01 g742706 ( .a(n_37396), .b(n_37276), .o(n_37486) );
in01s01 g742707 ( .a(n_37371), .o(n_37372) );
no02s01 g742708 ( .a(n_37379), .b(n_37017), .o(n_37371) );
na02s01 g742709 ( .a(n_37355), .b(n_37354), .o(n_37356) );
na02s01 g742710 ( .a(n_37326), .b(n_37325), .o(n_37327) );
no02s01 g742711 ( .a(n_37444), .b(n_37445), .o(n_37483) );
in01s01 g742712 ( .a(n_37454), .o(n_37455) );
na02s01 g742713 ( .a(n_37444), .b(n_44038), .o(n_37454) );
na02s02 g742714 ( .a(n_37480), .b(n_37479), .o(n_37481) );
na02s01 g742715 ( .a(n_37408), .b(FE_OCP_RBN3985_FE_RN_158_0), .o(n_37497) );
no02s01 g742716 ( .a(n_37323), .b(n_37322), .o(n_37324) );
oa12s01 g742718 ( .a(n_37149), .b(n_37409), .c(n_37038), .o(n_37457) );
na02m20 TIMEBOOST_cell_6006 ( .a(TIMEBOOST_net_1854), .b(n_23482), .o(n_23563) );
no02s06 TIMEBOOST_cell_2136 ( .a(TIMEBOOST_net_682), .b(n_22099), .o(n_22235) );
in01s01 g742721 ( .a(n_37398), .o(n_37910) );
ao12s01 g742722 ( .a(n_37321), .b(n_37320), .c(n_37319), .o(n_37398) );
ao12s02 g742723 ( .a(n_37341), .b(n_37340), .c(n_37339), .o(n_38209) );
in01s01 g742724 ( .a(n_37849), .o(n_37352) );
oa12s01 g742725 ( .a(n_37303), .b(n_37302), .c(n_37301), .o(n_37849) );
ao22s01 g742727 ( .a(n_37409), .b(n_37179), .c(n_37365), .d(n_37178), .o(n_38279) );
in01s02 g742728 ( .a(n_37518), .o(n_37545) );
ao12s01 g742729 ( .a(n_37443), .b(n_37442), .c(n_37441), .o(n_37518) );
oa12s02 g742731 ( .a(n_37440), .b(n_37439), .c(n_37438), .o(n_37912) );
in01s01 g742732 ( .a(n_37397), .o(n_37444) );
na02s01 g742733 ( .a(n_37353), .b(n_37207), .o(n_37397) );
no02s06 g742734 ( .a(n_37350), .b(n_37052), .o(n_37351) );
no02s01 g742735 ( .a(n_37320), .b(n_37319), .o(n_37321) );
na02s01 g742736 ( .a(n_37302), .b(n_37301), .o(n_37303) );
no02s02 g742738 ( .a(n_37442), .b(n_37441), .o(n_37443) );
na02s02 g742739 ( .a(n_37439), .b(n_37438), .o(n_37440) );
in01s01 g742740 ( .a(n_37395), .o(n_37396) );
na02m06 g742741 ( .a(n_37353), .b(n_37366), .o(n_37395) );
in01s01 g742742 ( .a(n_37407), .o(n_37408) );
no02s02 g742743 ( .a(n_37409), .b(n_36984), .o(n_37407) );
na02f06 g742744 ( .a(n_37353), .b(n_37265), .o(n_37369) );
no02s02 g742745 ( .a(n_37340), .b(n_37339), .o(n_37341) );
ao12s01 g742746 ( .a(n_37222), .b(n_37291), .c(n_37288), .o(n_37323) );
in01s01 g742747 ( .a(n_37348), .o(n_37349) );
no02m02 TIMEBOOST_cell_8731 ( .a(TIMEBOOST_net_2852), .b(n_12630), .o(n_13889) );
na02s01 TIMEBOOST_cell_5156 ( .a(n_15518), .b(FE_OCP_RBN6801_n_15156), .o(TIMEBOOST_net_1526) );
no02s01 g742751 ( .a(n_37393), .b(n_37392), .o(n_37391) );
in01s01 g742753 ( .a(n_37317), .o(n_37379) );
in01s01 g742755 ( .a(n_37299), .o(n_37317) );
ao12f08 g742756 ( .a(n_37231), .b(n_37291), .c(n_37186), .o(n_37299) );
ao12s01 g742757 ( .a(n_37009), .b(n_37298), .c(n_37131), .o(n_37355) );
ao12s01 g742758 ( .a(n_37221), .b(n_37291), .c(n_36969), .o(n_37326) );
in01s01 g742759 ( .a(n_38235), .o(n_37452) );
ao12s01 g742760 ( .a(n_37388), .b(n_37387), .c(n_37386), .o(n_38235) );
ao12s01 g742762 ( .a(n_37347), .b(n_37346), .c(n_37345), .o(n_37894) );
in01s01 g742763 ( .a(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n_43012) );
no02s01 g742765 ( .a(n_37291), .b(n_37214), .o(n_37302) );
no02f04 TIMEBOOST_cell_1786 ( .a(TIMEBOOST_net_507), .b(n_15500), .o(n_15545) );
na02s01 g742767 ( .a(n_37389), .b(n_37253), .o(n_37439) );
in01m06 g742768 ( .a(n_37350), .o(n_37337) );
na02s10 g742769 ( .a(n_37316), .b(n_37150), .o(n_37350) );
no02s01 g742770 ( .a(n_37298), .b(n_36952), .o(n_37340) );
no02s02 g742771 ( .a(n_37514), .b(n_36957), .o(n_37561) );
no02s01 g742772 ( .a(n_37387), .b(n_37386), .o(n_37388) );
no02s01 g742773 ( .a(n_37346), .b(n_37345), .o(n_37347) );
in01m01 g742774 ( .a(n_37290), .o(n_37608) );
no02m03 g742775 ( .a(n_37514), .b(n_36997), .o(n_37290) );
oa12s01 g742776 ( .a(n_37074), .b(n_37281), .c(n_36958), .o(n_37320) );
in01s01 g742778 ( .a(n_37409), .o(n_37365) );
in01s01 g742779 ( .a(n_37353), .o(n_37409) );
no02s01 TIMEBOOST_cell_4502 ( .a(TIMEBOOST_net_1341), .b(n_31992), .o(n_32128) );
in01s01 g742784 ( .a(n_37875), .o(n_37334) );
no02s01 g742785 ( .a(n_37287), .b(n_37282), .o(n_37875) );
na02s02 TIMEBOOST_cell_2878 ( .a(FE_RN_837_0), .b(n_7134), .o(TIMEBOOST_net_730) );
in01s01 g742787 ( .a(n_37393), .o(n_37364) );
oa12s01 g742788 ( .a(n_37315), .b(n_37314), .c(n_37313), .o(n_37393) );
in01s01 g742789 ( .a(n_37384), .o(n_37385) );
ao12s01 g742790 ( .a(n_37332), .b(n_37331), .c(n_37330), .o(n_37384) );
no02s04 g742791 ( .a(n_37272), .b(n_37126), .o(n_37273) );
na02m01 g742792 ( .a(n_37344), .b(n_37157), .o(n_37389) );
no02s01 g742793 ( .a(n_37344), .b(n_37343), .o(n_37387) );
no02m10 g742794 ( .a(n_37277), .b(n_37099), .o(n_37316) );
no02s02 g742795 ( .a(n_37281), .b(n_37014), .o(n_37298) );
na02s01 g742796 ( .a(n_37314), .b(n_37313), .o(n_37315) );
no02s01 g742797 ( .a(n_37310), .b(n_37147), .o(n_37333) );
na02s10 g742798 ( .a(n_37258), .b(n_37127), .o(n_37514) );
no02s01 g742799 ( .a(n_37331), .b(n_37330), .o(n_37332) );
no02m08 g742800 ( .a(n_37245), .b(n_37132), .o(n_37291) );
no02s01 g742801 ( .a(n_37256), .b(n_37120), .o(n_37287) );
no02s01 g742802 ( .a(n_37281), .b(n_37121), .o(n_37282) );
ao12s01 g742805 ( .a(n_37244), .b(n_37243), .c(n_37242), .o(n_37869) );
ao12s01 g742806 ( .a(n_37105), .b(n_37297), .c(n_37045), .o(n_37346) );
no02s08 g742807 ( .a(n_37311), .b(n_37111), .o(n_37312) );
in01s02 g742808 ( .a(n_37258), .o(n_37272) );
no02s10 g742809 ( .a(n_37083), .b(n_37233), .o(n_37258) );
no02s02 g742810 ( .a(n_37233), .b(n_37067), .o(n_37232) );
no02s01 g742811 ( .a(n_37297), .b(n_37028), .o(n_37331) );
in01s01 g742812 ( .a(n_37277), .o(n_37278) );
no02m04 TIMEBOOST_cell_1660 ( .a(TIMEBOOST_net_444), .b(n_9019), .o(n_9157) );
in01s01 g742815 ( .a(n_37256), .o(n_37281) );
in01s01 g742817 ( .a(n_37245), .o(n_37256) );
oa12m08 g742818 ( .a(n_36967), .b(n_37223), .c(n_37013), .o(n_37245) );
in01s01 g742819 ( .a(n_37310), .o(n_37344) );
na02m01 g742820 ( .a(n_37297), .b(n_37279), .o(n_37310) );
no02s01 g742821 ( .a(n_37243), .b(n_37242), .o(n_37244) );
oa12s01 g742822 ( .a(n_37145), .b(n_37286), .c(n_37036), .o(n_37314) );
oa22s01 g742823 ( .a(n_38173), .b(n_45891), .c(n_45899), .d(n_45895), .o(n_38525) );
in01s01 g742824 ( .a(n_37392), .o(n_37309) );
oa22s01 g742825 ( .a(n_37286), .b(n_37177), .c(n_37266), .d(n_37176), .o(n_37392) );
na02s10 g742826 ( .a(n_37215), .b(n_37130), .o(n_37233) );
na02m08 g742827 ( .a(n_37230), .b(n_37129), .o(n_37231) );
no02s06 g742828 ( .a(n_37276), .b(n_37110), .o(n_37368) );
no02s01 g742829 ( .a(n_37223), .b(n_36990), .o(n_37243) );
no02m01 g742830 ( .a(n_37286), .b(n_37034), .o(n_37297) );
in01m02 g742831 ( .a(n_37311), .o(n_37296) );
na02m10 g742832 ( .a(n_37268), .b(n_37271), .o(n_37311) );
oa12s01 g742833 ( .a(n_37198), .b(n_37200), .c(n_37197), .o(n_37836) );
in01s01 g742834 ( .a(n_37240), .o(n_37241) );
oa12s01 g742835 ( .a(n_37213), .b(n_37212), .c(n_37211), .o(n_37240) );
no02m10 g742836 ( .a(n_37200), .b(n_36989), .o(n_37223) );
na02s01 g742837 ( .a(n_37270), .b(FE_RN_199_0), .o(n_37255) );
na02s01 g742838 ( .a(n_37253), .b(n_37161), .o(n_37254) );
in01s01 g742839 ( .a(n_37215), .o(n_37199) );
no02s10 g742840 ( .a(n_37188), .b(n_37081), .o(n_37215) );
in01s01 g742841 ( .a(n_37230), .o(n_37222) );
no02m08 g742842 ( .a(n_37214), .b(n_37080), .o(n_37230) );
na02s01 g742843 ( .a(n_37195), .b(n_37079), .o(n_37221) );
na02s01 g742844 ( .a(n_37200), .b(n_37197), .o(n_37198) );
na02s01 g742845 ( .a(n_37212), .b(n_37211), .o(n_37213) );
na02s01 g742846 ( .a(n_37165), .b(n_36975), .o(n_37196) );
in01m08 g742847 ( .a(n_37276), .o(n_37268) );
na02m10 g742848 ( .a(n_37252), .b(n_37270), .o(n_37276) );
in01s01 g742850 ( .a(n_37286), .o(n_37266) );
in01m01 g742851 ( .a(n_37251), .o(n_37286) );
ao12f08 g742852 ( .a(n_37089), .b(n_37193), .c(n_37209), .o(n_37251) );
in01s01 g742854 ( .a(n_37274), .o(n_37275) );
oa12s01 g742855 ( .a(n_37238), .b(n_37237), .c(n_37236), .o(n_37274) );
oa12s01 g742856 ( .a(n_37250), .b(n_37249), .c(n_37248), .o(n_37877) );
no02m04 g742857 ( .a(n_37235), .b(n_37109), .o(n_37265) );
in01s01 g742858 ( .a(n_37188), .o(n_37165) );
oa12s10 g742859 ( .a(n_37135), .b(n_44039), .c(FE_OCP_RBN3939_n_46254), .o(n_37188) );
in01s01 g742860 ( .a(n_37214), .o(n_37195) );
na02s08 g742861 ( .a(n_37128), .b(n_37008), .o(n_37214) );
no02m10 g742862 ( .a(n_37445), .b(n_37164), .o(n_37270) );
no02m10 g742864 ( .a(n_37343), .b(n_37163), .o(n_37253) );
ao12m10 g742865 ( .a(n_36937), .b(n_37058), .c(n_36924), .o(n_37200) );
na02s01 g742866 ( .a(n_37237), .b(n_37236), .o(n_37238) );
na02s01 g742867 ( .a(n_37249), .b(n_37248), .o(n_37250) );
oa12s01 g742868 ( .a(n_36936), .b(n_37187), .c(n_36923), .o(n_37212) );
oa22s01 g742869 ( .a(n_37113), .b(n_36919), .c(n_37187), .d(n_36920), .o(n_37770) );
oa12s02 g742870 ( .a(n_37229), .b(n_37228), .c(n_37227), .o(n_37847) );
na02m10 g742871 ( .a(n_37184), .b(FE_OCP_RBN3986_FE_RN_158_0), .o(n_37445) );
na02m10 g742872 ( .a(n_37183), .b(n_37104), .o(n_37343) );
no03s10 g742874 ( .a(n_37077), .b(n_37002), .c(n_37072), .o(n_37186) );
na02s06 g742875 ( .a(n_37015), .b(n_37131), .o(n_37132) );
na03s02 TIMEBOOST_cell_7184 ( .a(FE_RN_1618_0), .b(FE_RN_1617_0), .c(TIMEBOOST_net_2231), .o(n_2495) );
na02s01 g742878 ( .a(n_37228), .b(n_37227), .o(n_37229) );
no02s01 g742879 ( .a(n_37194), .b(n_37203), .o(n_37249) );
in01m02 g742880 ( .a(n_37366), .o(n_37235) );
no02m10 g742881 ( .a(FE_OCP_RBN2428_n_37207), .b(n_37115), .o(n_37366) );
ao12s06 g742882 ( .a(FE_OCP_RBN3939_n_46254), .b(n_36954), .c(n_36563), .o(n_37083) );
no02s02 TIMEBOOST_cell_1779 ( .a(n_43147), .b(FE_OCP_RBN3307_n_43022), .o(TIMEBOOST_net_504) );
no02s03 TIMEBOOST_cell_1780 ( .a(TIMEBOOST_net_504), .b(n_43271), .o(n_43233) );
ao12m03 g742885 ( .a(FE_OCP_RBN3939_n_46254), .b(n_44021), .c(n_36470), .o(n_37081) );
oa12m03 g742886 ( .a(n_46254), .b(n_37071), .c(delay_add_ln22_unr23_stage9_stallmux_q_23_), .o(n_37130) );
oa12s06 g742887 ( .a(n_46254), .b(n_37073), .c(delay_add_ln22_unr23_stage9_stallmux_q_15_), .o(n_37129) );
no02s02 TIMEBOOST_cell_3841 ( .a(n_172), .b(n_156), .o(TIMEBOOST_net_1011) );
ao12s06 g742889 ( .a(FE_OCP_RBN3939_n_46254), .b(n_37079), .c(n_36466), .o(n_37080) );
oa12s03 g742890 ( .a(FE_OCP_RBN3938_n_46254), .b(n_37126), .c(delay_add_ln22_unr23_stage9_stallmux_q_27_), .o(n_37127) );
oa12s01 g742891 ( .a(n_37144), .b(n_37204), .c(n_37030), .o(n_37237) );
in01s06 g742892 ( .a(n_37419), .o(n_37078) );
no02s03 g742893 ( .a(n_37019), .b(n_37005), .o(n_37419) );
in01s06 g742895 ( .a(n_37288), .o(n_37077) );
no02s06 g742896 ( .a(n_37001), .b(n_37016), .o(n_37288) );
no02s06 g742897 ( .a(n_37014), .b(n_37003), .o(n_37015) );
na02s10 g742898 ( .a(n_36964), .b(n_36935), .o(n_37013) );
in01s02 g742899 ( .a(n_37375), .o(n_37076) );
no02s02 g742900 ( .a(n_37012), .b(n_37000), .o(n_37375) );
na02s01 g742901 ( .a(n_37135), .b(n_37010), .o(n_37011) );
na02s01 g742902 ( .a(n_37008), .b(n_37006), .o(n_37009) );
in01s01 g742903 ( .a(n_37124), .o(n_37125) );
no02s01 g742904 ( .a(n_37126), .b(n_37471), .o(n_37124) );
no02m06 TIMEBOOST_cell_3840 ( .a(n_28205), .b(TIMEBOOST_net_1010), .o(n_28298) );
na02s01 g742907 ( .a(n_37133), .b(n_37010), .o(n_37464) );
in01s01 g742908 ( .a(n_37122), .o(n_37123) );
na02s01 g742909 ( .a(n_36961), .b(n_37075), .o(n_37122) );
in01s01 g742910 ( .a(n_37120), .o(n_37121) );
na02s01 g742911 ( .a(n_36959), .b(n_37074), .o(n_37120) );
no02s01 g742912 ( .a(n_36972), .b(n_36968), .o(n_37339) );
no02s01 g742913 ( .a(n_37073), .b(n_37072), .o(n_37322) );
no02s01 g742914 ( .a(n_36971), .b(n_37016), .o(n_37301) );
no02s01 g742915 ( .a(n_36965), .b(n_36966), .o(n_37242) );
no02s01 g742916 ( .a(n_36976), .b(n_37012), .o(n_37402) );
no02s01 g742917 ( .a(n_37071), .b(n_37070), .o(n_37428) );
in01s01 g742918 ( .a(n_37118), .o(n_37119) );
na02s01 g742919 ( .a(n_36996), .b(n_37069), .o(n_37118) );
in01s01 g742920 ( .a(n_37116), .o(n_37117) );
na02s03 g742921 ( .a(n_36956), .b(n_37068), .o(n_37116) );
no02s01 g742922 ( .a(n_37067), .b(n_37019), .o(n_37506) );
in01s02 g742923 ( .a(n_37219), .o(n_37220) );
no02m08 TIMEBOOST_cell_8610 ( .a(FE_OFN748_n_22641), .b(FE_OCP_RBN6033_n_46962), .o(TIMEBOOST_net_2792) );
no02s08 g742926 ( .a(n_37159), .b(n_37048), .o(n_37207) );
na02s06 g742927 ( .a(n_44038), .b(n_44037), .o(n_37115) );
in01s01 g742929 ( .a(n_37065), .o(n_37066) );
ao12s01 g742930 ( .a(n_37005), .b(FE_OCP_RBN3938_n_46254), .c(delay_add_ln22_unr23_stage9_stallmux_q_25_), .o(n_37065) );
ao12s01 g742931 ( .a(n_37004), .b(FE_OCP_RBN3938_n_46254), .c(delay_add_ln22_unr23_stage9_stallmux_q_19_), .o(n_37468) );
ao12s01 g742932 ( .a(n_37003), .b(FE_OCP_RBN3938_n_46254), .c(delay_add_ln22_unr23_stage9_stallmux_q_11_), .o(n_37354) );
in01s01 g742933 ( .a(n_37063), .o(n_37064) );
ao12s01 g742934 ( .a(n_37002), .b(FE_OCP_RBN3938_n_46254), .c(delay_add_ln22_unr23_stage9_stallmux_q_15_), .o(n_37063) );
ao12s01 g742935 ( .a(n_37001), .b(FE_OCP_RBN3938_n_46254), .c(delay_add_ln22_unr23_stage9_stallmux_q_13_), .o(n_37325) );
ao12s01 g742936 ( .a(n_37000), .b(FE_OCP_RBN3938_n_46254), .c(delay_add_ln22_unr23_stage9_stallmux_q_21_), .o(n_37431) );
in01s01 g742937 ( .a(n_37061), .o(n_37062) );
ao12s01 g742938 ( .a(n_36999), .b(FE_OCP_RBN3938_n_46254), .c(delay_add_ln22_unr23_stage9_stallmux_q_23_), .o(n_37061) );
in01s01 g742939 ( .a(n_37059), .o(n_37060) );
ao12s01 g742940 ( .a(n_36998), .b(FE_OCP_RBN3938_n_46254), .c(delay_add_ln22_unr23_stage9_stallmux_q_27_), .o(n_37059) );
oa12m01 g742941 ( .a(n_36996), .b(FE_OCP_RBN3939_n_46254), .c(n_36994), .o(n_36997) );
na02s01 g742942 ( .a(n_37204), .b(n_36944), .o(n_37228) );
in01s01 g742943 ( .a(n_37187), .o(n_37113) );
in01s01 g742944 ( .a(n_37058), .o(n_37187) );
oa12s04 g742946 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_37111), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_27_), .o(n_37112) );
oa12m10 g742947 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_37050), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_19_), .o(n_37184) );
na02f08 TIMEBOOST_cell_1606 ( .a(n_30895), .b(TIMEBOOST_net_417), .o(n_31044) );
oa12s08 g742950 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_37110), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_25_), .o(n_37271) );
na02m10 g742951 ( .a(n_37103), .b(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37183) );
ao12s06 g742952 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_37042), .c(n_36429), .o(n_37163) );
in01s01 g742954 ( .a(n_37193), .o(n_37194) );
na02s01 g742956 ( .a(n_37174), .b(n_37084), .o(n_37203) );
oa22s01 g742957 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_17_), .c(FE_OCP_RBN3939_n_46254), .d(n_36486), .o(n_37423) );
oa22s01 g742958 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_9_), .c(FE_OCP_RBN3939_n_46254), .d(n_36151), .o(n_37319) );
ao22s01 g742959 ( .a(FE_OCP_RBN5525_n_36921), .b(n_36913), .c(n_36921), .d(n_36912), .o(n_37741) );
in01s01 g742960 ( .a(n_37056), .o(n_37057) );
ao22s01 g742961 ( .a(FE_OCP_RBN3939_n_46254), .b(n_36994), .c(FE_OCP_RBN3938_n_46254), .d(delay_add_ln22_unr23_stage9_stallmux_q_29_), .o(n_37056) );
in01s01 g742962 ( .a(n_37054), .o(n_37055) );
oa22m01 g742963 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_31_), .c(FE_OCP_RBN3939_n_46254), .d(n_36650), .o(n_37054) );
no02s02 TIMEBOOST_cell_8635 ( .a(TIMEBOOST_net_2804), .b(n_4353), .o(n_4643) );
no02s06 g742966 ( .a(FE_OCP_RBN3939_n_46254), .b(n_36610), .o(n_37126) );
no02s06 g742967 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_26_), .o(n_37471) );
na02s01 g742968 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_18_), .o(n_37010) );
in01s01 g742969 ( .a(n_36975), .o(n_36976) );
na02s01 g742971 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_20_), .o(n_36975) );
in01m03 g742972 ( .a(n_36974), .o(n_37071) );
na02m03 g742973 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_22_), .o(n_36974) );
no02s06 g742974 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_25_), .o(n_37005) );
no02s01 g742975 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_19_), .o(n_37004) );
na02s06 g742976 ( .a(FE_OCP_RBN3939_n_46254), .b(n_36503), .o(n_37133) );
in01s06 g742977 ( .a(n_36973), .o(n_37073) );
na02s03 g742978 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_14_), .o(n_36973) );
in01s01 g742979 ( .a(n_37006), .o(n_36972) );
na02s10 g742980 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_10_), .o(n_37006) );
in01s01 g742981 ( .a(n_37079), .o(n_36971) );
na02s10 g742982 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_12_), .o(n_37079) );
in01s01 g742983 ( .a(n_37072), .o(n_36970) );
no02s06 g742984 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_14_), .o(n_37072) );
no02s06 g742985 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_15_), .o(n_37002) );
no02s06 g742986 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_13_), .o(n_37001) );
in01s01 g742987 ( .a(n_37016), .o(n_36969) );
no02s06 g742988 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_12_), .o(n_37016) );
in01m01 g742989 ( .a(n_36968), .o(n_37131) );
no02s06 g742990 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_10_), .o(n_36968) );
no02s06 g742991 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_11_), .o(n_37003) );
in01s10 g742992 ( .a(n_36966), .o(n_36967) );
no02s40 g742993 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_7_), .b(delay_add_ln22_unr23_stage9_stallmux_q_7_), .o(n_36966) );
in01s01 g742994 ( .a(n_36964), .o(n_36965) );
na02s20 g742995 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_7_), .b(delay_add_ln22_unr23_stage9_stallmux_q_7_), .o(n_36964) );
in01s01 g742996 ( .a(n_37012), .o(n_36963) );
no02s02 g742997 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_20_), .o(n_37012) );
no02s01 g742998 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_21_), .o(n_37000) );
no02s01 g742999 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_23_), .o(n_36999) );
in01s01 g743000 ( .a(n_37070), .o(n_36962) );
no02s01 g743001 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_22_), .o(n_37070) );
in01s03 g743002 ( .a(n_37357), .o(n_37160) );
no02s10 g743003 ( .a(n_37094), .b(n_37109), .o(n_37357) );
na02s08 g743004 ( .a(n_36983), .b(n_37047), .o(n_37159) );
no02s10 g743007 ( .a(n_37108), .b(n_37088), .o(n_37279) );
no02s10 g743009 ( .a(n_37147), .b(n_37091), .o(n_37157) );
in01s01 g743010 ( .a(n_36960), .o(n_36961) );
no02s01 g743011 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_16_), .o(n_36960) );
na02s01 g743012 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_16_), .o(n_37075) );
na02s01 g743013 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_8_), .o(n_37074) );
in01s01 g743014 ( .a(n_36958), .o(n_36959) );
no02s01 g743015 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_8_), .o(n_36958) );
no02s03 g743016 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_27_), .b(FE_OCP_RBN3938_n_46254), .o(n_36998) );
in01s01 g743017 ( .a(n_36996), .o(n_36957) );
na02s02 g743018 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_28_), .o(n_36996) );
na02s06 g743019 ( .a(FE_OCP_RBN3939_n_46254), .b(n_36625), .o(n_37069) );
na02m01 g743020 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_30_), .o(n_37068) );
in01s03 g743021 ( .a(n_36955), .o(n_36956) );
no02m01 g743022 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_30_), .o(n_36955) );
na02s01 g743024 ( .a(FE_OCP_RBN3985_FE_RN_158_0), .b(n_37106), .o(n_37107) );
na02s01 g743025 ( .a(n_37104), .b(n_37102), .o(n_37105) );
no02s06 TIMEBOOST_cell_1600 ( .a(n_34873), .b(TIMEBOOST_net_414), .o(n_34900) );
na02m10 g743027 ( .a(n_37102), .b(n_36435), .o(n_37103) );
no02s01 g743028 ( .a(n_36990), .b(n_36989), .o(n_37197) );
in01s01 g743029 ( .a(n_37155), .o(n_37156) );
na02s02 g743030 ( .a(n_37051), .b(n_37101), .o(n_37155) );
in01s01 g743031 ( .a(n_37153), .o(n_37154) );
no02s01 g743032 ( .a(n_37100), .b(n_37111), .o(n_37153) );
in01s01 g743033 ( .a(n_37151), .o(n_37152) );
no02m01 g743034 ( .a(n_37426), .b(n_37099), .o(n_37151) );
in01s01 g743035 ( .a(n_37180), .o(n_37181) );
na02s02 g743036 ( .a(n_37150), .b(n_37041), .o(n_37180) );
no02s01 g743037 ( .a(n_37098), .b(n_37097), .o(n_37482) );
na02s01 g743038 ( .a(FE_RN_199_0), .b(n_37095), .o(n_37521) );
in01s01 g743039 ( .a(n_37178), .o(n_37179) );
na02s01 g743040 ( .a(n_37149), .b(n_37039), .o(n_37178) );
na02s01 g743041 ( .a(n_37148), .b(n_37106), .o(n_37496) );
no02s01 g743042 ( .a(n_37109), .b(n_37110), .o(n_37485) );
no02s01 g743043 ( .a(n_37147), .b(n_37146), .o(n_37386) );
na02s01 g743044 ( .a(n_37044), .b(n_37161), .o(n_37438) );
in01s01 g743045 ( .a(n_37176), .o(n_37177) );
na02s01 g743046 ( .a(n_37145), .b(n_37037), .o(n_37176) );
no02s01 g743047 ( .a(n_37043), .b(n_37108), .o(n_37330) );
in01s01 g743048 ( .a(n_36954), .o(n_37067) );
na02s06 g743049 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_24_), .o(n_36954) );
no02s06 g743051 ( .a(FE_OCP_RBN3938_n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_24_), .o(n_37019) );
oa12s10 g743052 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_17_), .c(delay_add_ln22_unr23_stage9_stallmux_q_16_), .o(n_37135) );
ao12s02 g743053 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_17_), .c(delay_add_ln22_unr23_stage9_stallmux_q_16_), .o(n_37017) );
in01s01 g743054 ( .a(n_37008), .o(n_36952) );
oa12s06 g743055 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_8_), .c(delay_add_ln22_unr23_stage9_stallmux_q_9_), .o(n_37008) );
no02s01 TIMEBOOST_cell_7887 ( .a(TIMEBOOST_net_2574), .b(n_35937), .o(TIMEBOOST_net_1568) );
ao12m20 g743057 ( .a(n_36922), .b(n_36936), .c(n_36934), .o(n_36937) );
na02s01 g743058 ( .a(n_37171), .b(n_37175), .o(n_37204) );
in01s01 g743059 ( .a(n_37173), .o(n_37174) );
no02f10 g743060 ( .a(n_37144), .b(n_37029), .o(n_37173) );
in01s01 g743061 ( .a(n_37142), .o(n_37143) );
no02m06 TIMEBOOST_cell_1570 ( .a(TIMEBOOST_net_399), .b(n_8266), .o(n_8364) );
in01s01 g743063 ( .a(n_37140), .o(n_37141) );
ao12s01 g743064 ( .a(n_37093), .b(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_27_), .o(n_37140) );
ao22s01 g743065 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_21_), .c(n_36991), .d(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37524) );
ao22s01 g743066 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_23_), .c(n_36992), .d(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37571) );
ao12s01 g743067 ( .a(n_37046), .b(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_19_), .o(n_37500) );
ao12s01 g743068 ( .a(n_37092), .b(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_15_), .o(n_37479) );
ao12s01 g743069 ( .a(n_37091), .b(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_13_), .o(n_37441) );
no02s01 g743070 ( .a(n_37171), .b(n_36928), .o(n_37172) );
no03m03 TIMEBOOST_cell_6419 ( .a(FE_RN_242_0), .b(n_17929), .c(FE_OCP_RBN5550_n_17914), .o(n_18021) );
no02s01 g743072 ( .a(n_37090), .b(n_37089), .o(n_37248) );
ao12s01 g743073 ( .a(n_37088), .b(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_11_), .o(n_37345) );
oa12s01 g743074 ( .a(n_36987), .b(n_36986), .c(n_36985), .o(n_37800) );
in01s01 g743075 ( .a(n_37086), .o(n_37087) );
oa22s02 g743076 ( .a(n_36590), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .d(delay_sub_ln21_0_unr23_stage9_stallmux_q_31_), .o(n_37086) );
oa22s01 g743077 ( .a(n_36461), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .d(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_), .o(n_37456) );
oa22s01 g743078 ( .a(n_36014), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .d(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_), .o(n_37313) );
in01s01 g743082 ( .a(n_36935), .o(n_36990) );
na02s06 g743083 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_6_), .b(delay_add_ln22_unr23_stage9_stallmux_q_6_), .o(n_36935) );
no02s40 g743084 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_6_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_6_), .o(n_36989) );
no02s20 g743085 ( .a(n_36922), .b(n_36923), .o(n_36924) );
in01s01 g743086 ( .a(n_37051), .o(n_37052) );
na02s01 g743087 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_30_), .o(n_37051) );
no02s06 g743088 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_36591), .o(n_37111) );
in01m10 g743089 ( .a(n_37106), .o(n_37050) );
na02s20 g743090 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_18_), .o(n_37106) );
no02s06 g743091 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(FE_OCP_RBN2337_delay_sub_ln21_0_unr23_stage9_stallmux_q_20_), .o(n_37097) );
no02s06 g743093 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_36950), .o(n_36988) );
no02s08 g743094 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_36537), .o(n_37110) );
no02s06 g743095 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_36564), .o(n_37099) );
na02m02 g743096 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_29_), .o(n_37150) );
no02s03 g743097 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_28_), .o(n_37426) );
no02s06 g743098 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_27_), .o(n_37093) );
in01s01 g743099 ( .a(n_37100), .o(n_37049) );
no02s10 g743100 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_26_), .o(n_37100) );
no02s10 g743101 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_25_), .o(n_37094) );
no02s10 g743102 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_24_), .o(n_37109) );
in01s01 g743103 ( .a(n_37048), .o(n_37148) );
no02s06 g743104 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_18_), .o(n_37048) );
in01s08 g743105 ( .a(n_37046), .o(n_37047) );
no02s10 g743106 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_19_), .o(n_37046) );
na02s01 g743107 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_36950), .o(n_37095) );
no02s01 g743108 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_20_), .o(n_37098) );
no02s20 g743109 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_7_), .b(n_35713), .o(n_37090) );
no02s06 g743110 ( .a(n_36933), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_7_), .o(n_37089) );
no02s10 g743111 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_11_), .o(n_37088) );
in01s01 g743112 ( .a(n_37108), .o(n_37045) );
no02s10 g743113 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_10_), .o(n_37108) );
no02s03 g743114 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_15_), .o(n_37092) );
in01s01 g743115 ( .a(n_37205), .o(n_37044) );
no02s10 g743116 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_14_), .o(n_37205) );
no02s10 g743117 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_12_), .o(n_37147) );
no02s10 g743118 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_13_), .o(n_37091) );
in01s01 g743119 ( .a(n_37102), .o(n_37043) );
na02s20 g743120 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_10_), .o(n_37102) );
in01s01 g743121 ( .a(n_37042), .o(n_37146) );
na02s10 g743122 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_12_), .o(n_37042) );
in01s01 g743123 ( .a(n_37040), .o(n_37041) );
no02s02 g743124 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_29_), .o(n_37040) );
na02s06 g743125 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_14_), .o(n_37161) );
na02s02 g743126 ( .a(n_36636), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37101) );
na02m06 TIMEBOOST_cell_7848 ( .a(n_14805), .b(n_16038), .o(TIMEBOOST_net_2555) );
na02s01 g743128 ( .a(n_36914), .b(n_36934), .o(n_37211) );
na02s01 g743129 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_), .o(n_37149) );
in01s01 g743130 ( .a(n_37038), .o(n_37039) );
no02s01 g743131 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_), .o(n_37038) );
in01s01 g743132 ( .a(n_37036), .o(n_37037) );
no02s01 g743133 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_), .o(n_37036) );
na02s01 g743134 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_), .o(n_37145) );
na02s01 g743135 ( .a(n_36986), .b(n_36985), .o(n_36987) );
in01s01 g743137 ( .a(n_36983), .o(n_36984) );
na02m04 TIMEBOOST_cell_7843 ( .a(TIMEBOOST_net_2552), .b(n_15800), .o(n_15895) );
ao12s06 g743140 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_), .o(n_37034) );
in01s01 g743141 ( .a(n_37085), .o(n_37171) );
na02s01 g743142 ( .a(n_37033), .b(n_37032), .o(n_37085) );
no02m20 g743143 ( .a(n_37029), .b(n_37030), .o(n_37031) );
in01s01 g743144 ( .a(n_37104), .o(n_37028) );
oa12s10 g743145 ( .a(FE_OCP_RBN3964_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_), .o(n_37104) );
na02s01 g743146 ( .a(n_36982), .b(n_37084), .o(n_37236) );
no02s06 TIMEBOOST_cell_5380 ( .a(n_35282), .b(n_35283), .o(TIMEBOOST_net_1638) );
in01s01 g743151 ( .a(n_36947), .o(n_36948) );
ao12s01 g743152 ( .a(n_36911), .b(n_36910), .c(n_36909), .o(n_36947) );
in01s06 g743156 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_7_), .o(n_36933) );
na02m40 g743158 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_5_), .b(delay_add_ln22_unr23_stage9_stallmux_q_5_), .o(n_36934) );
in01s01 g743159 ( .a(n_36922), .o(n_36914) );
no02s80 g743160 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_5_), .b(delay_add_ln22_unr23_stage9_stallmux_q_5_), .o(n_36922) );
in01s01 g743162 ( .a(n_37029), .o(n_36982) );
no02m80 g743163 ( .a(n_36946), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_6_), .o(n_37029) );
in01s03 g743164 ( .a(n_37084), .o(n_36981) );
na02s06 g743165 ( .a(n_36946), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_6_), .o(n_37084) );
in01s01 g743166 ( .a(n_36919), .o(n_36920) );
na02s01 g743167 ( .a(n_36888), .b(n_36936), .o(n_36919) );
in01s01 g743168 ( .a(n_36912), .o(n_36913) );
na02s01 g743169 ( .a(n_36879), .b(n_36897), .o(n_36912) );
no02s01 g743170 ( .a(n_36910), .b(n_36909), .o(n_36911) );
na02s01 g743171 ( .a(n_36932), .b(n_36931), .o(n_36986) );
in01s02 TIMEBOOST_cell_7386 ( .a(TIMEBOOST_net_2322), .o(FE_OFN2_n_43918) );
na02s01 g743173 ( .a(n_36930), .b(n_36943), .o(n_37227) );
ao12s02 g743175 ( .a(n_36709), .b(n_36889), .c(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36891) );
oa12s01 g743177 ( .a(n_36877), .b(n_36876), .c(n_36875), .o(n_37655) );
ao12s01 g743178 ( .a(n_36907), .b(n_36908), .c(n_36906), .o(n_37744) );
in01s01 g743179 ( .a(n_45896), .o(n_38193) );
in01s06 g743181 ( .a(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42196) );
in01m80 g743184 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_6_), .o(n_36946) );
na02s40 g743186 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_4_), .b(delay_add_ln22_unr23_stage9_stallmux_q_4_), .o(n_36936) );
na02s06 g743187 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_3_), .b(delay_add_ln22_unr23_stage9_stallmux_q_3_), .o(n_36897) );
in01s01 g743188 ( .a(n_36878), .o(n_36879) );
no02s40 g743189 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_3_), .b(delay_add_ln22_unr23_stage9_stallmux_q_3_), .o(n_36878) );
in01s01 g743190 ( .a(n_36923), .o(n_36888) );
no02s40 g743191 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_4_), .b(delay_add_ln22_unr23_stage9_stallmux_q_4_), .o(n_36923) );
in01s01 g743192 ( .a(n_37030), .o(n_36930) );
no02m40 g743193 ( .a(n_36918), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_5_), .o(n_37030) );
na02s20 g743194 ( .a(n_36918), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_5_), .o(n_36943) );
na02s01 g743195 ( .a(n_36887), .b(n_36886), .o(n_36909) );
na02s01 g743196 ( .a(n_36876), .b(n_36875), .o(n_36877) );
na02s10 g743197 ( .a(n_36908), .b(n_36884), .o(n_36932) );
no02s01 g743198 ( .a(n_36908), .b(n_36906), .o(n_36907) );
oa12s20 g743200 ( .a(n_36802), .b(n_36847), .c(n_36875), .o(n_36910) );
in01s01 g743201 ( .a(n_36928), .o(n_36929) );
na02s01 g743202 ( .a(n_37175), .b(n_36944), .o(n_36928) );
na02s01 g743203 ( .a(n_37032), .b(n_36917), .o(n_36985) );
ao12f02 g743204 ( .a(n_36751), .b(n_36894), .c(TIMEBOOST_net_2311), .o(n_36896) );
no02s03 TIMEBOOST_cell_1764 ( .a(TIMEBOOST_net_496), .b(n_20973), .o(n_21037) );
no02s01 g743206 ( .a(n_38129), .b(n_38094), .o(n_38173) );
in01s01 g743209 ( .a(FE_OCPN1624_n_37661), .o(n_37739) );
oa12s01 g743210 ( .a(n_36905), .b(n_36904), .c(n_36903), .o(n_37661) );
in01m80 g743213 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_5_), .o(n_36918) );
na02f03 g743215 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_2_), .b(delay_add_ln22_unr23_stage9_stallmux_q_2_), .o(n_36886) );
na02s06 g743217 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_4_), .b(n_35506), .o(n_37175) );
na02m20 g743218 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_3_), .b(n_35473), .o(n_37032) );
na02s20 g743219 ( .a(n_36872), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_3_), .o(n_36917) );
na02s20 g743220 ( .a(n_36873), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_4_), .o(n_36944) );
no02s01 g743221 ( .a(n_36803), .b(n_36847), .o(n_36876) );
na02s01 g743222 ( .a(n_36904), .b(n_36903), .o(n_36905) );
in01s02 g743223 ( .a(n_36846), .o(n_36889) );
na02s06 g743224 ( .a(n_36801), .b(n_36756), .o(n_36846) );
oa12m10 g743227 ( .a(n_36864), .b(n_36903), .c(n_36883), .o(n_36908) );
in01s01 g743228 ( .a(n_38128), .o(n_38129) );
ao12s01 g743229 ( .a(n_38045), .b(n_38044), .c(n_46242), .o(n_38128) );
no02m04 TIMEBOOST_cell_8586 ( .a(FE_OCP_RBN4303_n_44579), .b(n_44821), .o(TIMEBOOST_net_2780) );
in01s20 g743235 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_4_), .o(n_36873) );
in01s20 g743237 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_3_), .o(n_36872) );
no02s40 g743239 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_1_), .b(delay_add_ln22_unr23_stage9_stallmux_q_1_), .o(n_36847) );
in01s01 g743240 ( .a(n_36802), .o(n_36803) );
na02s40 g743241 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_1_), .b(delay_add_ln22_unr23_stage9_stallmux_q_1_), .o(n_36802) );
in01f04 g743242 ( .a(n_36867), .o(n_36894) );
na02f08 g743243 ( .a(n_36831), .b(n_36786), .o(n_36867) );
in01s01 g743244 ( .a(n_36832), .o(n_36833) );
in01s02 g743245 ( .a(n_36801), .o(n_36832) );
no02s06 g743246 ( .a(n_36742), .b(n_36783), .o(n_36801) );
no02s01 g743247 ( .a(n_38044), .b(n_46242), .o(n_38045) );
no02f10 TIMEBOOST_cell_1762 ( .a(TIMEBOOST_net_495), .b(FE_RN_2138_0), .o(n_25940) );
na02s01 g743250 ( .a(n_36931), .b(n_36884), .o(n_36906) );
no02s01 g743251 ( .a(n_36865), .b(n_36883), .o(n_36904) );
no02s01 g743256 ( .a(n_37992), .b(n_37189), .o(n_38044) );
na02m06 g743257 ( .a(n_35466), .b(delay_sub_ln21_unr24_stage9_stallmux_q_2_), .o(n_36884) );
in01s01 g743258 ( .a(n_36864), .o(n_36865) );
na02s20 g743259 ( .a(n_36844), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_1_), .o(n_36864) );
no02s20 g743260 ( .a(n_36844), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_1_), .o(n_36883) );
na02s06 g743261 ( .a(n_36828), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_2_), .o(n_36931) );
in01s01 g743263 ( .a(n_36831), .o(n_36842) );
no02f08 g743264 ( .a(n_36789), .b(n_36777), .o(n_36831) );
in01s01 g743265 ( .a(n_36790), .o(n_36791) );
in01s02 g743266 ( .a(n_36783), .o(n_36790) );
na02s06 g743267 ( .a(n_36761), .b(n_36692), .o(n_36783) );
ao12s01 g743268 ( .a(n_37960), .b(n_37959), .c(n_37958), .o(n_38093) );
no02f08 TIMEBOOST_cell_1758 ( .a(n_6160), .b(TIMEBOOST_net_493), .o(n_6266) );
in01s06 g743273 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_2_), .o(n_36828) );
in01s40 g743275 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_1_), .o(n_36844) );
no02s01 g743277 ( .a(n_37959), .b(n_37958), .o(n_37960) );
in01s01 g743279 ( .a(n_36789), .o(n_36798) );
na02f08 g743280 ( .a(n_36767), .b(n_36732), .o(n_36789) );
in01s02 g743281 ( .a(n_36771), .o(n_36772) );
in01m01 g743282 ( .a(n_36761), .o(n_36771) );
no02s06 g743283 ( .a(n_36725), .b(n_36743), .o(n_36761) );
oa12s02 g743284 ( .a(n_46228), .b(n_37899), .c(n_46227), .o(n_37992) );
in01s02 g743285 ( .a(n_36759), .o(n_36760) );
no02s02 g743286 ( .a(n_36711), .b(n_36743), .o(n_36759) );
in01m02 g743287 ( .a(n_36757), .o(n_36758) );
no02m02 g743288 ( .a(n_36742), .b(n_36710), .o(n_36757) );
in01s01 g743289 ( .a(n_36769), .o(n_36770) );
na02s02 g743290 ( .a(n_36724), .b(n_36756), .o(n_36769) );
no02s02 TIMEBOOST_cell_1753 ( .a(n_43179), .b(FE_OCP_RBN3375_n_43046), .o(TIMEBOOST_net_491) );
in01s01 g743292 ( .a(n_38019), .o(n_38020) );
oa12s01 g743293 ( .a(n_37923), .b(n_37922), .c(n_46247), .o(n_38019) );
in01s01 g743295 ( .a(n_37504), .o(n_36768) );
oa22s01 g743296 ( .a(n_36708), .b(delay_add_ln22_unr23_stage9_stallmux_q_0_), .c(n_35362), .d(delay_sub_ln22_unr24_stage9_stallmux_q_0_), .o(n_37504) );
na02s01 g743297 ( .a(n_37922), .b(n_46247), .o(n_37923) );
na02s40 g743298 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_0_), .b(delay_add_ln22_unr23_stage9_stallmux_q_0_), .o(n_36875) );
na02s01 g743299 ( .a(n_37899), .b(n_37898), .o(n_37959) );
in01s01 g743301 ( .a(n_36767), .o(n_36780) );
no02f08 g743302 ( .a(n_36736), .b(n_36755), .o(n_36767) );
in01s01 g743303 ( .a(n_36739), .o(n_36740) );
in01s01 g743304 ( .a(n_36725), .o(n_36739) );
na02s06 g743305 ( .a(n_36677), .b(n_36712), .o(n_36725) );
no02s06 g743306 ( .a(n_36675), .b(n_36750), .o(n_36743) );
no02s02 g743307 ( .a(n_36676), .b(FE_OCPN1947_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36711) );
no02s06 g743308 ( .a(n_36750), .b(n_36673), .o(n_36742) );
no02s02 g743309 ( .a(n_36674), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36710) );
na02s06 g743310 ( .a(n_36690), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36756) );
na02s02 g743311 ( .a(n_36750), .b(n_36691), .o(n_36724) );
na02s01 g743312 ( .a(n_37857), .b(n_37856), .o(n_37858) );
no02s02 TIMEBOOST_cell_1754 ( .a(TIMEBOOST_net_491), .b(n_43215), .o(n_43370) );
no02s02 g743315 ( .a(n_36735), .b(n_36755), .o(n_36778) );
in01m02 g743316 ( .a(n_36787), .o(n_36788) );
na02m04 TIMEBOOST_cell_8621 ( .a(TIMEBOOST_net_2797), .b(n_16379), .o(TIMEBOOST_net_1702) );
in01f02 g743318 ( .a(n_36796), .o(n_36797) );
na02f04 g743319 ( .a(n_36786), .b(n_36765), .o(n_36796) );
in01f02 g743320 ( .a(n_36737), .o(n_36738) );
na02f04 g743321 ( .a(n_36695), .b(n_36712), .o(n_36737) );
oa12s01 g743322 ( .a(n_37841), .b(n_37840), .c(n_37839), .o(n_38021) );
no02m02 TIMEBOOST_cell_1755 ( .a(n_43266), .b(n_43265), .o(TIMEBOOST_net_492) );
in01s02 g743326 ( .a(n_36722), .o(n_36723) );
in01s01 g743328 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_0_), .o(n_36708) );
na02s01 g743330 ( .a(n_37840), .b(n_37839), .o(n_37841) );
in01s01 g743331 ( .a(n_37855), .o(n_37899) );
no02s02 g743332 ( .a(n_37828), .b(n_46226), .o(n_37855) );
in01s01 g743333 ( .a(n_36753), .o(n_36754) );
in01s01 g743334 ( .a(n_36736), .o(n_36753) );
na02f08 g743335 ( .a(n_36705), .b(n_36717), .o(n_36736) );
no02f08 g743338 ( .a(n_36660), .b(n_36614), .o(n_36677) );
no02s02 g743339 ( .a(n_36704), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36735) );
no02f08 g743340 ( .a(n_36703), .b(FE_OFN5083_n_36750), .o(n_36755) );
no02m10 TIMEBOOST_cell_8693 ( .a(TIMEBOOST_net_2833), .b(n_1542), .o(TIMEBOOST_net_33) );
no02f08 g743342 ( .a(n_36715), .b(FE_OFN5084_n_36750), .o(n_36777) );
na02s06 g743343 ( .a(TIMEBOOST_net_2321), .b(n_36730), .o(n_36786) );
na02f04 g743344 ( .a(n_36731), .b(FE_OFN5084_n_36750), .o(n_36765) );
na02f04 g743345 ( .a(n_36656), .b(n_36750), .o(n_36695) );
na02s06 g743346 ( .a(n_36655), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36712) );
no02s06 TIMEBOOST_cell_1743 ( .a(n_26272), .b(n_23564), .o(TIMEBOOST_net_486) );
no02s03 TIMEBOOST_cell_1756 ( .a(TIMEBOOST_net_492), .b(FE_OCP_RBN4479_FE_OCPN913_n_43230), .o(n_43364) );
no02m02 g743350 ( .a(n_36635), .b(n_36660), .o(n_36693) );
no02f04 TIMEBOOST_cell_6757 ( .a(n_4636), .b(FE_OCP_RBN4294_n_4080), .o(TIMEBOOST_net_2136) );
ao12s01 g743353 ( .a(n_37805), .b(n_37830), .c(n_46243), .o(n_37856) );
ao12s01 g743354 ( .a(n_37803), .b(n_37830), .c(n_46232), .o(n_37857) );
no02f08 TIMEBOOST_cell_1749 ( .a(n_39142), .b(n_39216), .o(TIMEBOOST_net_489) );
in01m02 g743356 ( .a(n_36763), .o(n_36764) );
oa22m04 g743357 ( .a(n_36751), .b(TIMEBOOST_net_2319), .c(n_36701), .d(FE_OFN5084_n_36750), .o(n_36763) );
in01s01 g743358 ( .a(n_36675), .o(n_36676) );
na02s01 TIMEBOOST_cell_1224 ( .a(TIMEBOOST_net_226), .b(n_45896), .o(n_38221) );
in01s02 g743360 ( .a(n_36673), .o(n_36674) );
no02s01 TIMEBOOST_cell_1448 ( .a(n_34234), .b(TIMEBOOST_net_338), .o(n_34330) );
in01s01 g743362 ( .a(n_36690), .o(n_36691) );
no02s01 TIMEBOOST_cell_1228 ( .a(TIMEBOOST_net_228), .b(n_33409), .o(n_33525) );
in01s01 g743364 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_30_), .o(n_36636) );
no02s01 g743368 ( .a(n_37813), .b(n_37814), .o(n_37840) );
in01s01 g743369 ( .a(n_37828), .o(n_37829) );
na02s02 g743370 ( .a(n_37813), .b(n_36814), .o(n_37828) );
no02s01 g743371 ( .a(n_37830), .b(n_46243), .o(n_37805) );
no02s01 g743372 ( .a(n_37830), .b(n_46232), .o(n_37803) );
in01s01 g743373 ( .a(n_36720), .o(n_36721) );
in01s01 g743374 ( .a(n_36705), .o(n_36720) );
no02f08 g743375 ( .a(n_36689), .b(n_36579), .o(n_36705) );
no02f08 g743376 ( .a(n_36583), .b(n_36750), .o(n_36660) );
no02m02 g743377 ( .a(n_36584), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36635) );
na02s01 TIMEBOOST_cell_1223 ( .a(n_37201), .b(n_37224), .o(TIMEBOOST_net_226) );
na02s02 g743379 ( .a(n_36594), .b(n_36750), .o(n_36595) );
na02s06 g743380 ( .a(n_36612), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36692) );
no02f06 TIMEBOOST_cell_8123 ( .a(TIMEBOOST_net_2692), .b(n_21271), .o(n_21459) );
na02s02 g743382 ( .a(n_36592), .b(n_36750), .o(n_36593) );
no02s01 TIMEBOOST_cell_1447 ( .a(n_33792), .b(n_34211), .o(TIMEBOOST_net_338) );
no02m08 TIMEBOOST_cell_5653 ( .a(TIMEBOOST_net_1774), .b(n_11315), .o(n_11370) );
na02s02 TIMEBOOST_cell_5644 ( .a(n_6181), .b(n_6032), .o(TIMEBOOST_net_1770) );
in01s01 g743386 ( .a(n_36718), .o(n_36719) );
no02s02 g743387 ( .a(n_36672), .b(n_36689), .o(n_36718) );
in01s01 g743388 ( .a(n_36733), .o(n_36734) );
na02s02 g743389 ( .a(n_36717), .b(n_36688), .o(n_36733) );
in01s02 g743390 ( .a(n_36748), .o(n_36749) );
no03f40 TIMEBOOST_cell_3458 ( .a(n_27918), .b(FE_RN_1979_0), .c(FE_RN_1978_0), .o(n_27839) );
na02s02 TIMEBOOST_cell_8029 ( .a(TIMEBOOST_net_2645), .b(n_20489), .o(n_20568) );
in01s01 g743393 ( .a(n_37826), .o(n_37827) );
oa12s01 g743394 ( .a(n_37788), .b(n_37787), .c(n_46248), .o(n_37826) );
no02s04 TIMEBOOST_cell_1745 ( .a(n_26176), .b(n_23353), .o(TIMEBOOST_net_487) );
na02s01 TIMEBOOST_cell_1742 ( .a(TIMEBOOST_net_485), .b(n_39436), .o(n_39510) );
in01s01 g743397 ( .a(n_36703), .o(n_36704) );
na02m06 TIMEBOOST_cell_1534 ( .a(n_14948), .b(TIMEBOOST_net_381), .o(n_15090) );
in01m02 g743399 ( .a(n_36715), .o(n_36716) );
no02s01 TIMEBOOST_cell_1432 ( .a(TIMEBOOST_net_330), .b(n_34082), .o(n_34169) );
in01s02 g743401 ( .a(n_36730), .o(n_36731) );
no02s01 TIMEBOOST_cell_1436 ( .a(n_29721), .b(TIMEBOOST_net_332), .o(n_29758) );
in01f02 g743403 ( .a(n_36655), .o(n_36656) );
na02s04 TIMEBOOST_cell_1226 ( .a(TIMEBOOST_net_227), .b(n_33852), .o(n_33876) );
in01s02 g743405 ( .a(n_36709), .o(n_36654) );
no02m04 g743406 ( .a(n_36568), .b(n_36586), .o(n_36709) );
in01s02 g743408 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_29_), .o(n_36994) );
in01s01 g743411 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_26_), .o(n_36591) );
in01s01 g743413 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_31_), .o(n_36590) );
na02s01 g743415 ( .a(n_37787), .b(n_46248), .o(n_37788) );
ao12s02 g743416 ( .a(n_37748), .b(n_36775), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37813) );
no02s01 g743417 ( .a(n_37747), .b(n_36978), .o(n_37830) );
no02f08 g743418 ( .a(n_36626), .b(FE_OFN5083_n_36750), .o(n_36689) );
no02s02 g743419 ( .a(n_36627), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36672) );
na02f08 g743420 ( .a(n_36646), .b(FE_OCPN1940_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36717) );
na02s02 g743421 ( .a(n_36647), .b(FE_OFN5083_n_36750), .o(n_36688) );
na02s02 TIMEBOOST_cell_1533 ( .a(n_14428), .b(n_14427), .o(TIMEBOOST_net_381) );
na02s01 TIMEBOOST_cell_4886 ( .a(n_17610), .b(n_17536), .o(TIMEBOOST_net_1391) );
na02m08 g743424 ( .a(n_36667), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36732) );
no02f06 TIMEBOOST_cell_8592 ( .a(FE_OCP_RBN3008_n_15206), .b(n_14340), .o(TIMEBOOST_net_2783) );
no02s01 TIMEBOOST_cell_1431 ( .a(n_34074), .b(n_33701), .o(TIMEBOOST_net_330) );
na02s03 g743427 ( .a(n_36651), .b(FE_OFN5084_n_36750), .o(n_36652) );
no02s01 TIMEBOOST_cell_1435 ( .a(n_29078), .b(n_29306), .o(TIMEBOOST_net_332) );
no03s03 TIMEBOOST_cell_3453 ( .a(n_1521), .b(n_1422), .c(n_1543), .o(n_1557) );
in01s02 g743430 ( .a(n_36657), .o(n_36631) );
in01s01 g743431 ( .a(n_36614), .o(n_36657) );
no02f06 g743432 ( .a(n_36588), .b(n_36750), .o(n_36614) );
na02s01 TIMEBOOST_cell_5973 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_21_), .b(FE_OCP_RBN2404_n_45697), .o(TIMEBOOST_net_1838) );
no03s10 TIMEBOOST_cell_3503 ( .a(FE_RN_646_0), .b(FE_RN_648_0), .c(n_32936), .o(TIMEBOOST_net_737) );
na02s01 TIMEBOOST_cell_1225 ( .a(n_33367), .b(n_33851), .o(TIMEBOOST_net_227) );
no02s02 g743436 ( .a(TIMEBOOST_net_2325), .b(n_36567), .o(n_36568) );
no02s04 g743437 ( .a(n_36551), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36586) );
na02s01 g743438 ( .a(n_37750), .b(n_37749), .o(n_37751) );
no02m02 TIMEBOOST_cell_1738 ( .a(TIMEBOOST_net_483), .b(n_26389), .o(n_26421) );
ao12s01 g743440 ( .a(n_37681), .b(n_37680), .c(n_46244), .o(n_37789) );
in01s01 g743441 ( .a(n_37784), .o(n_37785) );
oa12s01 g743442 ( .a(n_37729), .b(n_37728), .c(n_37727), .o(n_37784) );
in01s02 g743443 ( .a(n_36594), .o(n_36566) );
in01s02 g743445 ( .a(n_36592), .o(n_36565) );
in01s02 g743447 ( .a(n_36615), .o(n_36585) );
in01m02 g743449 ( .a(n_36751), .o(n_36701) );
no02m02 TIMEBOOST_cell_8834 ( .a(TIMEBOOST_net_2278), .b(FE_OCP_RBN4384_n_5221), .o(TIMEBOOST_net_2904) );
in01s06 g743451 ( .a(n_36583), .o(n_36584) );
no02f04 TIMEBOOST_cell_1440 ( .a(n_38124), .b(TIMEBOOST_net_334), .o(n_38172) );
in01s01 g743453 ( .a(n_36612), .o(n_36613) );
no02s01 TIMEBOOST_cell_7058 ( .a(TIMEBOOST_net_2287), .b(n_20518), .o(TIMEBOOST_net_1269) );
in01s01 g743455 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_31_), .o(n_36650) );
in01s01 g743457 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_25_), .o(n_36540) );
in01s02 g743459 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_28_), .o(n_36564) );
no02s01 g743461 ( .a(n_37680), .b(n_46244), .o(n_37681) );
na02s01 g743462 ( .a(n_37728), .b(n_37727), .o(n_37729) );
in01s01 g743463 ( .a(n_37747), .o(n_37748) );
no02s02 g743464 ( .a(n_37711), .b(n_46210), .o(n_37747) );
no02s02 g743465 ( .a(n_36629), .b(FE_OFN5084_n_36750), .o(n_36630) );
na03m08 TIMEBOOST_cell_4598 ( .a(n_23002), .b(n_22938), .c(n_22971), .o(n_23137) );
no02f04 TIMEBOOST_cell_1439 ( .a(n_38034), .b(n_38011), .o(TIMEBOOST_net_334) );
na02s04 g743468 ( .a(n_36520), .b(n_36750), .o(n_36521) );
no02s10 TIMEBOOST_cell_8469 ( .a(TIMEBOOST_net_2721), .b(n_32704), .o(n_32572) );
na02s01 TIMEBOOST_cell_5573 ( .a(TIMEBOOST_net_1734), .b(n_6343), .o(n_6435) );
no02s01 g743471 ( .a(n_37712), .b(n_36941), .o(n_37787) );
oa12s01 g743472 ( .a(n_37635), .b(n_37634), .c(n_46240), .o(n_37730) );
ao12s01 g743473 ( .a(n_37676), .b(n_37713), .c(n_46238), .o(n_37750) );
ao12s01 g743474 ( .a(n_37674), .b(n_37673), .c(n_37672), .o(n_37749) );
in01s01 g743475 ( .a(n_37725), .o(n_37726) );
oa12s01 g743476 ( .a(n_37678), .b(n_37713), .c(n_46241), .o(n_37725) );
in01m02 g743477 ( .a(n_36569), .o(n_36552) );
in01s01 g743479 ( .a(n_36567), .o(n_36551) );
in01m02 g743481 ( .a(n_36632), .o(n_36611) );
in01f02 g743483 ( .a(n_36651), .o(n_36628) );
in01s01 g743487 ( .a(n_36626), .o(n_36627) );
no02s01 TIMEBOOST_cell_1426 ( .a(n_34020), .b(TIMEBOOST_net_327), .o(n_34104) );
in01s01 g743489 ( .a(n_36646), .o(n_36647) );
no02s06 TIMEBOOST_cell_4864 ( .a(n_65), .b(beta_31), .o(TIMEBOOST_net_1380) );
in01s01 g743491 ( .a(n_36667), .o(n_36668) );
no02s01 TIMEBOOST_cell_4115 ( .a(FE_OCP_RBN6074_n_44256), .b(n_35980), .o(TIMEBOOST_net_1148) );
no02s01 TIMEBOOST_cell_1204 ( .a(TIMEBOOST_net_216), .b(n_420), .o(n_466) );
in01s01 g743494 ( .a(n_37625), .o(n_36686) );
oa12s01 g743495 ( .a(n_36624), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_0_), .c(delay_add_ln22_unr23_stage9_stallmux_q_24_), .o(n_37625) );
in01s02 g743496 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_25_), .o(n_36563) );
in01s03 g743498 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_26_), .o(n_36610) );
in01s01 g743500 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_28_), .o(n_36625) );
in01s01 g743502 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_23_), .o(n_36992) );
in01s01 g743504 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_24_), .o(n_36537) );
na02s01 g743506 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_0_), .b(delay_add_ln22_unr23_stage9_stallmux_q_24_), .o(n_36624) );
no02s01 g743507 ( .a(n_37699), .b(n_37631), .o(n_37728) );
na02s01 g743508 ( .a(n_37713), .b(n_46241), .o(n_37678) );
na02s01 g743509 ( .a(n_37634), .b(n_46240), .o(n_37635) );
no02s01 g743510 ( .a(n_37713), .b(n_46238), .o(n_37676) );
no02s40 g743511 ( .a(FE_OCP_RBN6506_delay_add_ln22_unr23_stage9_stallmux_q_24_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_0_), .o(n_36903) );
in01s01 g743512 ( .a(n_37711), .o(n_37712) );
na02s02 g743513 ( .a(n_37699), .b(n_36826), .o(n_37711) );
no02s01 g743514 ( .a(n_37673), .b(n_37672), .o(n_37674) );
no02s01 TIMEBOOST_cell_1425 ( .a(n_33997), .b(n_33671), .o(TIMEBOOST_net_327) );
na02s04 g743516 ( .a(n_36549), .b(FE_OFN5083_n_36750), .o(n_36550) );
no03f04 TIMEBOOST_cell_3511 ( .a(TIMEBOOST_net_602), .b(FE_OCP_RBN5564_n_37551), .c(n_37648), .o(n_37742) );
no02s03 TIMEBOOST_cell_8746 ( .a(n_13515), .b(n_13514), .o(TIMEBOOST_net_2860) );
na02m02 TIMEBOOST_cell_4114 ( .a(TIMEBOOST_net_1147), .b(n_35948), .o(n_36038) );
na02f08 TIMEBOOST_cell_8869 ( .a(TIMEBOOST_net_2921), .b(n_26131), .o(n_26297) );
no02s01 TIMEBOOST_cell_1203 ( .a(n_448), .b(n_447), .o(TIMEBOOST_net_216) );
na02s03 g743522 ( .a(n_36489), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36510) );
na02s01 g743523 ( .a(n_37613), .b(n_37538), .o(n_37632) );
ao12s01 g743524 ( .a(n_36841), .b(n_37584), .c(n_36852), .o(n_37680) );
no02s06 g743526 ( .a(n_36462), .b(n_36000), .o(n_36508) );
in01s02 g743527 ( .a(n_36516), .o(n_36517) );
no02s01 TIMEBOOST_cell_1198 ( .a(TIMEBOOST_net_213), .b(n_37829), .o(n_37922) );
in01s03 g743529 ( .a(n_36506), .o(n_36507) );
oa12s06 g743530 ( .a(n_36008), .b(n_36474), .c(n_47265), .o(n_36506) );
in01f02 g743531 ( .a(n_36520), .o(n_36505) );
in01s02 g743533 ( .a(n_36515), .o(n_36553) );
in01s02 g743535 ( .a(n_36629), .o(n_36607) );
oa22m04 g743536 ( .a(n_36529), .b(n_36299), .c(n_36530), .d(n_36300), .o(n_36629) );
in01s01 g743541 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_21_), .o(n_36991) );
in01s01 g743543 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_22_), .o(n_36950) );
no02s01 g743545 ( .a(n_37611), .b(n_37631), .o(n_37713) );
no03m08 TIMEBOOST_cell_2231 ( .a(n_40781), .b(n_40688), .c(n_40734), .o(n_40798) );
ao12s02 g743547 ( .a(n_37612), .b(n_36727), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37699) );
na02s01 g743548 ( .a(n_37585), .b(n_46203), .o(n_37673) );
in01s01 g743550 ( .a(n_36579), .o(n_36604) );
no02s06 g743551 ( .a(n_36543), .b(FE_OFN5083_n_36750), .o(n_36579) );
in01f04 g743552 ( .a(n_36492), .o(n_36493) );
na02f08 g743553 ( .a(n_36474), .b(FE_OCPN4836_n_36034), .o(n_36492) );
no02s01 TIMEBOOST_cell_1197 ( .a(n_37814), .b(n_36854), .o(TIMEBOOST_net_213) );
no02s06 g743555 ( .a(n_36444), .b(n_36095), .o(n_36462) );
oa12s01 g743556 ( .a(n_46206), .b(n_37586), .c(n_46213), .o(n_37634) );
oa12f08 g743558 ( .a(n_36007), .b(n_36514), .c(n_36035), .o(n_36535) );
no02m08 g743560 ( .a(n_36504), .b(n_36148), .o(n_36547) );
oa12s06 g743561 ( .a(n_36199), .b(FE_OCP_RBN6151_n_36501), .c(n_36531), .o(n_36546) );
no02m08 g743562 ( .a(n_36533), .b(FE_OCP_RBN6104_n_36199), .o(n_36560) );
na02s01 TIMEBOOST_cell_1196 ( .a(TIMEBOOST_net_212), .b(n_37854), .o(n_37920) );
in01s01 g743565 ( .a(n_37613), .o(n_37614) );
ao22s01 g743566 ( .a(n_37586), .b(n_36869), .c(n_37517), .d(n_36868), .o(n_37613) );
oa22s01 g743567 ( .a(n_36398), .b(n_36238), .c(n_36399), .d(n_36239), .o(n_36449) );
in01m02 g743570 ( .a(n_36549), .o(n_36534) );
na02s06 TIMEBOOST_cell_1384 ( .a(TIMEBOOST_net_306), .b(n_18869), .o(n_19002) );
in01m02 g743572 ( .a(n_36545), .o(n_36581) );
in01s02 g743574 ( .a(n_36559), .o(n_36608) );
in01s01 g743578 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_), .o(n_36461) );
in01s01 g743583 ( .a(n_37584), .o(n_37585) );
no02s01 g743584 ( .a(n_37586), .b(n_46200), .o(n_37584) );
na02s02 TIMEBOOST_cell_1383 ( .a(n_18345), .b(n_47247), .o(TIMEBOOST_net_306) );
no03s20 TIMEBOOST_cell_4592 ( .a(n_28039), .b(FE_RN_125_0), .c(n_28282), .o(n_28319) );
no02m06 g743587 ( .a(n_36482), .b(n_36147), .o(n_36504) );
no02m08 g743588 ( .a(FE_OCP_RBN6151_n_36501), .b(n_36531), .o(n_36533) );
in01s01 g743589 ( .a(n_37611), .o(n_37612) );
na02s02 TIMEBOOST_cell_1728 ( .a(TIMEBOOST_net_478), .b(n_4098), .o(n_4173) );
in01s02 g743591 ( .a(n_36529), .o(n_36530) );
no02m06 TIMEBOOST_cell_1388 ( .a(TIMEBOOST_net_308), .b(n_7703), .o(n_7752) );
na02m06 g743595 ( .a(n_36400), .b(n_36045), .o(n_36447) );
na02s01 TIMEBOOST_cell_1195 ( .a(n_37773), .b(n_37789), .o(TIMEBOOST_net_212) );
no02f02 TIMEBOOST_cell_1730 ( .a(TIMEBOOST_net_479), .b(n_15547), .o(n_15621) );
no02s02 TIMEBOOST_cell_1731 ( .a(n_4363), .b(n_4416), .o(TIMEBOOST_net_480) );
oa22s01 g743599 ( .a(n_36412), .b(n_36257), .c(n_36413), .d(n_36256), .o(n_36460) );
oa22s01 g743600 ( .a(n_36378), .b(n_36255), .c(n_36379), .d(n_36254), .o(n_36433) );
oa22s01 g743601 ( .a(n_36382), .b(n_35860), .c(n_36383), .d(n_35859), .o(n_36432) );
oa12s06 g743604 ( .a(n_36102), .b(n_36416), .c(n_36192), .o(n_36444) );
oa22s01 g743605 ( .a(n_36437), .b(n_36364), .c(n_36438), .d(n_36363), .o(n_36487) );
in01s01 g743606 ( .a(n_36543), .o(n_36544) );
na02f04 TIMEBOOST_cell_5446 ( .a(FE_OCP_RBN6083_n_5454), .b(n_4316), .o(TIMEBOOST_net_1671) );
in01s01 g743608 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_17_), .o(n_36486) );
in01s01 g743610 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_18_), .o(n_36503) );
in01m01 g743613 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_21_), .o(n_36470) );
in01s01 g743617 ( .a(n_37517), .o(n_37586) );
oa12s01 g743618 ( .a(n_37435), .b(n_37437), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37517) );
no02m06 TIMEBOOST_cell_6016 ( .a(TIMEBOOST_net_1859), .b(n_13208), .o(n_13209) );
no02m04 TIMEBOOST_cell_6805 ( .a(FE_OCP_RBN5953_FE_OFN4772_n_44463), .b(FE_OCP_RBN3227_n_10644), .o(TIMEBOOST_net_2160) );
na02f04 g743622 ( .a(n_36381), .b(n_35899), .o(n_36400) );
no02m08 g743624 ( .a(n_36397), .b(n_36011), .o(n_36431) );
no02m04 TIMEBOOST_cell_1387 ( .a(n_7702), .b(n_7634), .o(TIMEBOOST_net_308) );
in01s02 g743626 ( .a(n_36457), .o(n_36458) );
oa12f06 g743627 ( .a(n_36105), .b(n_36410), .c(n_47266), .o(n_36457) );
in01m06 g743630 ( .a(n_36482), .o(n_36501) );
oa12m06 g743631 ( .a(n_36205), .b(n_36410), .c(n_36270), .o(n_36482) );
in01s01 g743632 ( .a(n_37538), .o(n_37539) );
ao12s01 g743633 ( .a(n_37478), .b(n_37477), .c(n_46239), .o(n_37538) );
oa22s01 g743634 ( .a(n_36347), .b(n_36259), .c(n_36348), .d(n_36258), .o(n_36415) );
oa22s01 g743635 ( .a(n_36394), .b(n_35738), .c(n_36395), .d(n_35737), .o(n_36442) );
oa22s01 g743636 ( .a(n_36349), .b(n_35779), .c(n_36350), .d(n_35778), .o(n_36414) );
in01s01 g743637 ( .a(n_36398), .o(n_36399) );
oa12s01 g743638 ( .a(n_36012), .b(n_36352), .c(n_35821), .o(n_36398) );
oa22s01 g743639 ( .a(n_36424), .b(n_36332), .c(n_36425), .d(n_36333), .o(n_36469) );
oa22s01 g743640 ( .a(n_36427), .b(n_35953), .c(n_36428), .d(n_35952), .o(n_36468) );
in01m02 g743641 ( .a(n_36514), .o(n_36481) );
na02f10 g743642 ( .a(n_36441), .b(n_36203), .o(n_36514) );
no02s01 g743644 ( .a(n_37477), .b(n_46239), .o(n_37478) );
na02f10 g743645 ( .a(n_44835), .b(n_36099), .o(n_36441) );
na02s02 g743646 ( .a(n_36410), .b(n_36103), .o(n_36483) );
no02s02 g743647 ( .a(n_44831), .b(n_36071), .o(n_36467) );
in01s01 g743648 ( .a(n_36382), .o(n_36383) );
na02s01 g743649 ( .a(n_36352), .b(n_35954), .o(n_36382) );
in01s01 g743650 ( .a(n_36412), .o(n_36413) );
na03f04 TIMEBOOST_cell_6465 ( .a(n_29864), .b(n_29894), .c(n_29890), .o(n_29989) );
in01s06 g743652 ( .a(n_36416), .o(n_36397) );
in01f08 g743653 ( .a(n_36381), .o(n_36416) );
in01s01 g743656 ( .a(n_36378), .o(n_36379) );
oa12s02 g743657 ( .a(n_35917), .b(n_36329), .c(n_35739), .o(n_36378) );
no02s06 TIMEBOOST_cell_1726 ( .a(n_25869), .b(TIMEBOOST_net_477), .o(n_26016) );
na02s01 TIMEBOOST_cell_1727 ( .a(n_4070), .b(n_3926), .o(TIMEBOOST_net_478) );
oa22s02 g743660 ( .a(n_36325), .b(n_36291), .c(n_36326), .d(n_36292), .o(n_36396) );
oa22s01 g743661 ( .a(n_36391), .b(n_36359), .c(n_36390), .d(n_36360), .o(n_36440) );
oa22s01 g743662 ( .a(n_36408), .b(n_35828), .c(n_36409), .d(n_35829), .o(n_36455) );
oa22s01 g743663 ( .a(n_36393), .b(n_35866), .c(n_36392), .d(n_35865), .o(n_36439) );
oa22s01 g743664 ( .a(n_36373), .b(n_36366), .c(n_36374), .d(n_36365), .o(n_36430) );
in01s01 g743665 ( .a(n_36437), .o(n_36438) );
oa12s01 g743666 ( .a(n_36072), .b(n_36411), .c(n_35911), .o(n_36437) );
in01s01 g743670 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_13_), .o(n_36429) );
no02s01 g743672 ( .a(n_37436), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_), .o(n_37437) );
no02s01 g743673 ( .a(n_37436), .b(n_37434), .o(n_37477) );
in01s01 g743674 ( .a(n_36427), .o(n_36428) );
na02s01 g743675 ( .a(n_36411), .b(n_36013), .o(n_36427) );
in01s01 g743676 ( .a(n_36394), .o(n_36395) );
na02s01 g743677 ( .a(n_36328), .b(n_35683), .o(n_36394) );
no03f06 TIMEBOOST_cell_7217 ( .a(TIMEBOOST_net_2251), .b(n_3955), .c(n_3877), .o(n_4212) );
in01s01 g743679 ( .a(n_36349), .o(n_36350) );
na02s01 g743680 ( .a(n_36329), .b(n_35864), .o(n_36349) );
ao12s01 g743681 ( .a(n_37434), .b(n_37363), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_), .o(n_37435) );
in01s01 g743686 ( .a(n_36347), .o(n_36348) );
oa12s02 g743687 ( .a(n_36188), .b(n_36279), .c(n_35619), .o(n_36347) );
oa12s01 g743689 ( .a(n_37383), .b(n_37382), .c(n_37381), .o(n_37541) );
oa22s01 g743690 ( .a(n_36248), .b(n_36240), .c(n_36279), .d(n_36241), .o(n_36377) );
in01s01 g743691 ( .a(n_36424), .o(n_36425) );
no03m10 TIMEBOOST_cell_3436 ( .a(n_22869), .b(FE_OCP_RBN5181_n_44061), .c(n_22803), .o(n_22965) );
in01s01 g743693 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_13_), .o(n_36466) );
na02s01 g743696 ( .a(n_37362), .b(n_46212), .o(n_37436) );
na02s01 g743697 ( .a(n_37382), .b(n_37381), .o(n_37383) );
in01s01 g743698 ( .a(n_36376), .o(n_36411) );
no02f10 g743699 ( .a(n_36346), .b(n_36331), .o(n_36376) );
in01s01 g743700 ( .a(n_36408), .o(n_36409) );
na02s01 g743701 ( .a(n_36344), .b(n_35868), .o(n_36408) );
no03m20 TIMEBOOST_cell_3435 ( .a(n_32436), .b(FE_OCP_RBN7006_n_44962), .c(n_32388), .o(n_32547) );
in01s01 g743703 ( .a(n_36327), .o(n_36328) );
no02s02 g743704 ( .a(n_36279), .b(n_35641), .o(n_36327) );
in01s01 g743705 ( .a(n_36373), .o(n_36374) );
na02s01 g743706 ( .a(n_36346), .b(n_35988), .o(n_36373) );
in01s01 g743707 ( .a(n_36392), .o(n_36393) );
ao12s01 g743708 ( .a(n_35987), .b(n_36372), .c(n_35870), .o(n_36392) );
in01s02 g743709 ( .a(n_36325), .o(n_36326) );
ao12s02 g743710 ( .a(n_35570), .b(n_36247), .c(n_35615), .o(n_36325) );
in01s01 g743711 ( .a(n_36390), .o(n_36391) );
ao12s01 g743712 ( .a(n_35744), .b(n_36372), .c(n_36303), .o(n_36390) );
ao12s01 g743713 ( .a(n_37361), .b(n_37405), .c(n_46235), .o(n_37472) );
oa12s01 g743714 ( .a(n_37359), .b(n_37405), .c(n_46233), .o(n_37540) );
oa22s01 g743715 ( .a(n_36273), .b(n_36287), .c(n_36274), .d(n_36288), .o(n_36371) );
oa22s01 g743716 ( .a(n_36277), .b(n_35638), .c(n_36247), .d(n_35639), .o(n_36345) );
in01s01 g743717 ( .a(n_36280), .o(n_36329) );
oa22s01 g743719 ( .a(n_36276), .b(n_36367), .c(n_36275), .d(n_36368), .o(n_36423) );
oa22s01 g743720 ( .a(n_36372), .b(n_36318), .c(n_36309), .d(n_36319), .o(n_36407) );
ao22s01 g743721 ( .a(n_37329), .b(n_46245), .c(n_37328), .d(n_36849), .o(n_37473) );
no02s01 g743723 ( .a(n_37342), .b(n_37434), .o(n_37382) );
in01s01 g743724 ( .a(n_37362), .o(n_37363) );
na02s01 g743725 ( .a(n_37342), .b(n_36818), .o(n_37362) );
no02s01 g743726 ( .a(n_37405), .b(n_46235), .o(n_37361) );
na02s01 g743727 ( .a(n_37405), .b(n_46233), .o(n_37359) );
in01s01 g743728 ( .a(n_36343), .o(n_36344) );
no02s01 g743729 ( .a(n_36309), .b(n_35752), .o(n_36343) );
na02f10 g743730 ( .a(n_36272), .b(n_35918), .o(n_36346) );
in01s01 g743733 ( .a(n_36248), .o(n_36279) );
in01s01 g743735 ( .a(n_36208), .o(n_36248) );
no03f06 TIMEBOOST_cell_8338 ( .a(n_19722), .b(FE_RN_2592_0), .c(FE_RN_2595_0), .o(n_19915) );
oa22s01 g743737 ( .a(n_36339), .b(n_36361), .c(n_36338), .d(n_36362), .o(n_36422) );
oa22s01 g743738 ( .a(n_36207), .b(n_35788), .c(n_36206), .d(n_35787), .o(n_36310) );
in01s01 g743739 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_11_), .o(n_36465) );
in01s01 g743742 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_11_), .o(n_36435) );
no02s01 g743744 ( .a(n_37295), .b(n_36899), .o(n_37405) );
ao12s01 g743745 ( .a(n_37294), .b(n_36557), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37342) );
in01s01 g743747 ( .a(n_36247), .o(n_36277) );
no02s02 g743748 ( .a(n_36110), .b(n_35692), .o(n_36247) );
no02s01 g743749 ( .a(n_37292), .b(n_37246), .o(n_37308) );
na02s01 g743750 ( .a(n_37305), .b(n_37304), .o(n_37307) );
no02s01 g743751 ( .a(n_37305), .b(n_37304), .o(n_37306) );
in01s01 g743752 ( .a(n_36275), .o(n_36276) );
ao12s01 g743753 ( .a(n_35754), .b(n_36109), .c(n_35873), .o(n_36275) );
in01s01 g743754 ( .a(n_37328), .o(n_37329) );
na02s01 g743755 ( .a(n_37285), .b(n_46219), .o(n_37328) );
in01s01 g743756 ( .a(n_36273), .o(n_36274) );
ao12s01 g743757 ( .a(n_36135), .b(n_36074), .c(n_36242), .o(n_36273) );
in01s01 g743760 ( .a(n_36309), .o(n_36372) );
in01s01 g743761 ( .a(n_36272), .o(n_36309) );
oa22s01 g743764 ( .a(n_36047), .b(n_36260), .c(n_36074), .d(n_36261), .o(n_36340) );
in01s01 g743765 ( .a(n_37294), .o(n_37295) );
na02s01 g743766 ( .a(n_37284), .b(n_36824), .o(n_37294) );
no02s01 g743767 ( .a(n_37284), .b(n_36793), .o(n_37285) );
no02s01 g743768 ( .a(n_36074), .b(n_36075), .o(n_36110) );
in01s01 g743769 ( .a(n_36338), .o(n_36339) );
ao12s01 g743770 ( .a(n_35669), .b(n_36324), .c(n_36304), .o(n_36338) );
in01s01 g743772 ( .a(n_36206), .o(n_36207) );
oa12s01 g743773 ( .a(n_35694), .b(n_36324), .c(n_35872), .o(n_36206) );
oa12s01 g743774 ( .a(n_37262), .b(n_37283), .c(n_46230), .o(n_37304) );
in01s01 g743775 ( .a(n_37292), .o(n_37293) );
oa12s01 g743776 ( .a(n_37260), .b(n_37283), .c(n_37259), .o(n_37292) );
oa22s01 g743777 ( .a(n_36322), .b(n_36289), .c(n_36323), .d(n_36290), .o(n_36389) );
oa22s01 g743778 ( .a(n_36369), .b(n_36316), .c(n_36370), .d(n_36317), .o(n_36421) );
oa22s01 g743779 ( .a(n_36324), .b(n_36320), .c(n_36073), .d(n_36321), .o(n_36388) );
oa12s01 g743780 ( .a(n_37264), .b(n_37283), .c(n_46234), .o(n_37305) );
na03m08 TIMEBOOST_cell_6432 ( .a(n_37697), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .c(n_37671), .o(TIMEBOOST_net_1862) );
in01s01 g743784 ( .a(n_36108), .o(n_36109) );
no02f10 g743785 ( .a(n_36046), .b(n_35693), .o(n_36108) );
no02s01 TIMEBOOST_cell_1663 ( .a(n_19649), .b(n_20135), .o(TIMEBOOST_net_446) );
na02s01 g743787 ( .a(n_37283), .b(n_46234), .o(n_37264) );
na02s01 g743788 ( .a(n_37283), .b(n_46230), .o(n_37262) );
na02s01 g743789 ( .a(n_37283), .b(n_37259), .o(n_37260) );
in01s01 g743792 ( .a(n_36047), .o(n_36074) );
in01s01 g743794 ( .a(n_36015), .o(n_36047) );
no02s01 TIMEBOOST_cell_1158 ( .a(TIMEBOOST_net_193), .b(n_41154), .o(n_41273) );
in01s01 g743796 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_9_), .o(n_36151) );
in01s01 g743798 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_), .o(n_36014) );
ao12f06 g743800 ( .a(FE_OCP_RBN6046_n_35487), .b(n_35878), .c(n_35555), .o(n_35923) );
in01s01 g743801 ( .a(n_46253), .o(n_37283) );
in01s01 g743803 ( .a(n_36369), .o(n_36370) );
na02s01 TIMEBOOST_cell_3414 ( .a(n_27509), .b(n_27561), .o(TIMEBOOST_net_998) );
in01s01 g743805 ( .a(n_36322), .o(n_36323) );
oa12s01 g743806 ( .a(n_36243), .b(n_35877), .c(n_36185), .o(n_36322) );
in01s01 g743807 ( .a(n_36324), .o(n_36073) );
in01s01 g743808 ( .a(n_36046), .o(n_36324) );
oa12f08 g743809 ( .a(n_35643), .b(n_36335), .c(n_35706), .o(n_36046) );
no02m08 TIMEBOOST_cell_1662 ( .a(TIMEBOOST_net_445), .b(n_20017), .o(n_20137) );
in01s01 g743811 ( .a(n_37246), .o(n_37247) );
oa12s01 g743812 ( .a(n_37218), .b(n_37217), .c(n_46231), .o(n_37246) );
oa22s01 g743813 ( .a(n_35876), .b(n_36262), .c(n_35877), .d(n_36263), .o(n_36337) );
oa12m01 g743814 ( .a(n_36336), .b(n_36335), .c(n_36334), .o(n_36387) );
na02s01 g743815 ( .a(n_46251), .b(n_46202), .o(n_37202) );
na02s01 g743816 ( .a(n_37217), .b(n_46231), .o(n_37218) );
no02m06 TIMEBOOST_cell_3413 ( .a(n_27568), .b(TIMEBOOST_net_997), .o(FE_RN_1283_0) );
no02m08 TIMEBOOST_cell_1626 ( .a(n_19358), .b(TIMEBOOST_net_427), .o(n_19474) );
na02s01 g743819 ( .a(n_36335), .b(n_36334), .o(n_36336) );
no02s01 TIMEBOOST_cell_1157 ( .a(n_40862), .b(n_40995), .o(TIMEBOOST_net_193) );
oa12s01 g743821 ( .a(n_35836), .b(n_35835), .c(n_35834), .o(n_35922) );
oa12s01 g743822 ( .a(n_35921), .b(n_35920), .c(n_35919), .o(n_35990) );
in01s01 g743823 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_8_), .o(n_35989) );
na02s01 g743826 ( .a(n_37168), .b(n_46202), .o(n_37217) );
no02m08 g743827 ( .a(n_36071), .b(n_47264), .o(n_36105) );
no02m06 g743828 ( .a(n_36071), .b(n_36204), .o(n_36205) );
no02s06 g743829 ( .a(n_36071), .b(n_36039), .o(n_36203) );
na02s01 g743831 ( .a(n_37190), .b(n_37021), .o(n_37191) );
na02s01 g743832 ( .a(n_35835), .b(n_35834), .o(n_35836) );
na02s01 g743833 ( .a(n_35920), .b(n_35919), .o(n_35921) );
na02f08 g743834 ( .a(n_35833), .b(n_35708), .o(n_36335) );
in01s01 g743835 ( .a(n_35876), .o(n_35877) );
in01s01 g743837 ( .a(n_35878), .o(n_35876) );
no02s01 TIMEBOOST_cell_1138 ( .a(TIMEBOOST_net_183), .b(n_37472), .o(n_37475) );
in01s01 g743840 ( .a(n_37168), .o(n_37169) );
no02s01 g743841 ( .a(n_37138), .b(n_36805), .o(n_37168) );
na02f06 g743842 ( .a(n_35832), .b(n_35707), .o(n_35833) );
no02s01 g743843 ( .a(n_36043), .b(n_35909), .o(n_36072) );
no02s01 TIMEBOOST_cell_1137 ( .a(n_37473), .b(n_37307), .o(TIMEBOOST_net_183) );
no02s01 g743845 ( .a(n_35674), .b(n_35553), .o(n_35835) );
in01s01 g743850 ( .a(n_36071), .o(n_36103) );
no02s01 g743852 ( .a(n_35832), .b(n_35621), .o(n_35920) );
oa12s01 g743853 ( .a(n_37027), .b(n_46250), .c(n_46236), .o(n_37190) );
in01s01 g743854 ( .a(n_37166), .o(n_37167) );
oa12s01 g743855 ( .a(n_37025), .b(n_46250), .c(n_46229), .o(n_37166) );
oa12s01 g743856 ( .a(n_35672), .b(n_35671), .c(n_35670), .o(n_35757) );
oa12s01 g743857 ( .a(n_35794), .b(n_35793), .c(n_35792), .o(n_35874) );
ao22s01 g743858 ( .a(n_46250), .b(n_36851), .c(n_36980), .d(n_46246), .o(n_37224) );
in01s06 g743859 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_7_), .o(n_35713) );
in01s01 g743861 ( .a(n_37898), .o(n_37189) );
no02s01 g743862 ( .a(n_37814), .b(n_36863), .o(n_37898) );
na02s01 g743863 ( .a(n_46250), .b(n_46236), .o(n_37027) );
na02s01 g743864 ( .a(n_46250), .b(n_46229), .o(n_37025) );
no02s01 g743865 ( .a(n_35987), .b(n_35827), .o(n_35988) );
no02m04 g743866 ( .a(n_36011), .b(n_35815), .o(n_36045) );
no02s04 g743867 ( .a(n_36011), .b(n_36100), .o(n_36102) );
ao12s01 g743868 ( .a(n_46250), .b(n_36434), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37138) );
in01s01 g743869 ( .a(n_35673), .o(n_35674) );
na02f08 g743870 ( .a(n_35627), .b(n_35519), .o(n_35673) );
na02s01 g743871 ( .a(n_35671), .b(n_35670), .o(n_35672) );
no02f06 g743872 ( .a(n_35712), .b(n_35622), .o(n_35832) );
in01s01 g743874 ( .a(n_36013), .o(n_36043) );
no02m08 g743875 ( .a(n_35987), .b(n_35867), .o(n_36013) );
no02s01 g743876 ( .a(n_36204), .b(n_36245), .o(n_36307) );
na02s01 g743877 ( .a(n_35793), .b(n_35792), .o(n_35794) );
no02s06 TIMEBOOST_cell_1594 ( .a(TIMEBOOST_net_411), .b(FE_OCP_RBN2930_n_34971), .o(n_35048) );
oa12s01 g743879 ( .a(n_35711), .b(n_35710), .c(n_35709), .o(n_35791) );
oa12s01 g743881 ( .a(n_36979), .b(n_36774), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37814) );
no02m10 g743882 ( .a(n_35869), .b(n_35826), .o(n_35918) );
no02s01 g743883 ( .a(n_35985), .b(n_35820), .o(n_36012) );
no02s01 g743884 ( .a(n_35872), .b(n_35751), .o(n_35873) );
no02s01 g743885 ( .a(n_35914), .b(n_35698), .o(n_35955) );
na02m10 g743889 ( .a(n_35954), .b(n_35822), .o(n_36011) );
in01s01 g743890 ( .a(n_35712), .o(n_35793) );
oa12f06 g743891 ( .a(n_35565), .b(n_35573), .c(n_35599), .o(n_35712) );
na02m06 g743893 ( .a(n_35830), .b(n_35868), .o(n_35987) );
na02m06 g743894 ( .a(n_36038), .b(n_36040), .o(n_36204) );
na02s01 g743895 ( .a(n_35710), .b(n_35709), .o(n_35711) );
no02m06 TIMEBOOST_cell_2933 ( .a(TIMEBOOST_net_757), .b(n_19335), .o(n_19434) );
in01s01 g743897 ( .a(n_46250), .o(n_36980) );
no02s02 g743899 ( .a(n_36270), .b(n_36200), .o(n_36271) );
in01s01 g743900 ( .a(n_37020), .o(n_37021) );
ao12s01 g743901 ( .a(n_36927), .b(n_36942), .c(n_46237), .o(n_37020) );
in01s01 g743902 ( .a(n_35627), .o(n_35671) );
oa12f08 g743903 ( .a(n_35484), .b(n_35538), .c(n_35502), .o(n_35627) );
oa12s01 g743904 ( .a(n_35579), .b(n_35578), .c(n_35577), .o(n_35626) );
no02s01 g743906 ( .a(n_36942), .b(n_46237), .o(n_36927) );
na02s01 g743907 ( .a(n_46249), .b(n_46211), .o(n_36941) );
na02s02 g743908 ( .a(n_36199), .b(n_36198), .o(n_36200) );
no02s01 g743909 ( .a(n_35916), .b(n_35736), .o(n_35917) );
in01s01 g743910 ( .a(n_36978), .o(n_36979) );
oa12s01 g743911 ( .a(n_46249), .b(n_36861), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_36978) );
in01s01 g743913 ( .a(n_35954), .o(n_35985) );
no02m10 g743914 ( .a(n_35916), .b(n_35783), .o(n_35954) );
no02s02 TIMEBOOST_cell_6365 ( .a(FE_OCP_RBN4396_n_16146), .b(FE_OCP_RBN6173_n_16923), .o(TIMEBOOST_net_2034) );
na02s01 g743916 ( .a(n_35578), .b(n_35577), .o(n_35579) );
in01s01 g743917 ( .a(n_35869), .o(n_35870) );
na02f06 g743919 ( .a(n_35651), .b(n_35707), .o(n_35708) );
na02s04 g743920 ( .a(n_36099), .b(n_36037), .o(n_36270) );
no02m06 g743921 ( .a(n_35649), .b(FE_OCP_RBN4904_n_44256), .o(n_35706) );
no02f08 g743922 ( .a(n_35704), .b(FE_OCP_RBN4904_n_44256), .o(n_35872) );
in01s01 g743925 ( .a(n_35868), .o(n_35914) );
na02m02 g743926 ( .a(n_35750), .b(FE_OCP_RBN4903_n_44256), .o(n_35868) );
na02s04 g743927 ( .a(n_35748), .b(FE_OCP_RBN4909_n_44222), .o(n_35830) );
na02m02 TIMEBOOST_cell_1230 ( .a(n_33388), .b(TIMEBOOST_net_229), .o(n_33434) );
in01s03 g743930 ( .a(n_36039), .o(n_36040) );
no02s06 g743931 ( .a(n_35951), .b(FE_OCP_RBN6074_n_44256), .o(n_36039) );
na03m06 TIMEBOOST_cell_7193 ( .a(n_14063), .b(n_14126), .c(TIMEBOOST_net_1524), .o(n_14326) );
no02s06 TIMEBOOST_cell_3991 ( .a(n_38770), .b(n_38778), .o(TIMEBOOST_net_1086) );
oa12s01 g743934 ( .a(n_35647), .b(n_35646), .c(n_35645), .o(n_35705) );
oa12s01 g743935 ( .a(n_35529), .b(n_35593), .c(FE_OCP_RBN3206_n_35517), .o(n_35710) );
na02s01 g743937 ( .a(n_36901), .b(n_46209), .o(n_36942) );
na02s01 g743938 ( .a(n_36915), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_0_), .o(n_36925) );
oa12s01 g743939 ( .a(n_36900), .b(n_36556), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37434) );
na02s01 g743941 ( .a(n_36901), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_36902) );
no02s06 g743945 ( .a(n_47266), .b(n_35984), .o(n_36099) );
no02s02 g743946 ( .a(n_47267), .b(n_36036), .o(n_36037) );
no02s02 g743948 ( .a(n_36098), .b(n_36148), .o(n_36199) );
na02s02 g743949 ( .a(n_36306), .b(n_36305), .o(n_36334) );
na02f04 g743950 ( .a(n_35650), .b(n_35596), .o(n_35651) );
no02s04 g743951 ( .a(n_35625), .b(n_35648), .o(n_35649) );
in01s01 g743952 ( .a(n_36320), .o(n_36321) );
na02s01 g743953 ( .a(n_36304), .b(n_35700), .o(n_36320) );
no02m08 g743954 ( .a(n_35669), .b(n_35703), .o(n_35704) );
in01s01 g743955 ( .a(n_35787), .o(n_35788) );
no02s01 g743956 ( .a(n_35751), .b(n_35754), .o(n_35787) );
in01s01 g743957 ( .a(n_36318), .o(n_36319) );
na02s01 g743958 ( .a(n_36303), .b(n_35699), .o(n_36318) );
in01s01 g743960 ( .a(n_35828), .o(n_35829) );
na02s01 g743961 ( .a(n_35831), .b(n_35747), .o(n_35828) );
na02m02 g743962 ( .a(n_35699), .b(n_35749), .o(n_35750) );
na02s02 g743963 ( .a(n_35747), .b(n_34726), .o(n_35748) );
in01s01 g743964 ( .a(n_35865), .o(n_35866) );
no02s01 g743965 ( .a(n_35827), .b(n_35826), .o(n_35865) );
in01s01 g743966 ( .a(n_35952), .o(n_35953) );
no02s01 g743967 ( .a(n_35909), .b(n_35911), .o(n_35952) );
na02s02 TIMEBOOST_cell_1229 ( .a(n_33386), .b(FE_RN_2043_0), .o(TIMEBOOST_net_229) );
in01s01 g743970 ( .a(n_36009), .o(n_36010) );
no02s02 g743971 ( .a(n_47266), .b(n_47264), .o(n_36009) );
no02s06 g743972 ( .a(n_47264), .b(n_35905), .o(n_35951) );
no02s01 g743974 ( .a(n_47267), .b(n_36035), .o(n_36069) );
in01s01 g743976 ( .a(n_36196), .o(n_36197) );
no02s01 g743977 ( .a(n_36148), .b(n_36147), .o(n_36196) );
no02s04 TIMEBOOST_cell_1205 ( .a(n_47245), .b(FE_OCPN1686_n_23097), .o(TIMEBOOST_net_217) );
no02s01 g743979 ( .a(n_35624), .b(n_35597), .o(n_35919) );
no02s02 g743980 ( .a(n_35947), .b(n_35974), .o(n_36008) );
na02m08 g743981 ( .a(n_35691), .b(n_35663), .o(n_35746) );
in01s01 g743982 ( .a(n_35916), .o(n_35864) );
oa12s08 g743983 ( .a(n_35683), .b(n_35689), .c(FE_OCP_RBN6048_n_35487), .o(n_35916) );
na02s02 g743984 ( .a(n_35976), .b(n_36034), .o(n_36100) );
no02f06 g743985 ( .a(n_35574), .b(n_35516), .o(n_35599) );
na02s01 g743986 ( .a(n_35646), .b(n_35645), .o(n_35647) );
na02s01 g743987 ( .a(n_35650), .b(n_35623), .o(n_35792) );
in01s01 g743988 ( .a(n_36367), .o(n_36368) );
no02s01 g743989 ( .a(n_36297), .b(n_35755), .o(n_36367) );
in01s01 g743990 ( .a(n_36332), .o(n_36333) );
na02s01 g743991 ( .a(n_36264), .b(n_35697), .o(n_36332) );
in01s01 g743992 ( .a(n_36365), .o(n_36366) );
no02s01 g743993 ( .a(n_36331), .b(n_36294), .o(n_36365) );
in01s01 g743994 ( .a(n_36363), .o(n_36364) );
no02s01 g743995 ( .a(n_35910), .b(n_36293), .o(n_36363) );
in01s02 g743996 ( .a(n_36032), .o(n_36033) );
no02s01 TIMEBOOST_cell_1100 ( .a(TIMEBOOST_net_164), .b(n_37410), .o(n_37525) );
in01s01 g743998 ( .a(n_36194), .o(n_36195) );
no02m20 TIMEBOOST_cell_1102 ( .a(FE_OCP_RBN5552_n_23328), .b(TIMEBOOST_net_165), .o(n_23411) );
in01s01 g744000 ( .a(n_36268), .o(n_36269) );
no02s01 TIMEBOOST_cell_7886 ( .a(n_35763), .b(FE_OCP_RBN3292_n_35539), .o(TIMEBOOST_net_2574) );
in01s01 g744002 ( .a(n_36301), .o(n_36302) );
na02s02 g744003 ( .a(n_36198), .b(n_36191), .o(n_36301) );
no02s01 g744004 ( .a(n_36192), .b(n_36097), .o(n_36193) );
ao12s01 g744005 ( .a(n_36881), .b(n_36882), .c(n_36880), .o(n_37022) );
ao12f08 g744006 ( .a(n_35535), .b(n_35537), .c(n_35536), .o(n_35538) );
oa12s01 g744007 ( .a(n_35523), .b(n_35537), .c(n_35522), .o(n_35557) );
oa12s01 g744008 ( .a(n_35536), .b(n_35537), .c(n_35535), .o(n_35578) );
in01s01 g744009 ( .a(n_36316), .o(n_36317) );
oa22s01 g744010 ( .a(FE_OCPN890_n_44223), .b(n_34593), .c(n_44222), .d(n_35648), .o(n_36316) );
in01s01 g744011 ( .a(n_36361), .o(n_36362) );
na02s01 g744012 ( .a(n_36298), .b(n_36267), .o(n_36361) );
in01s01 g744013 ( .a(n_36359), .o(n_36360) );
na02s01 g744014 ( .a(n_36295), .b(n_36265), .o(n_36359) );
in01s01 g744015 ( .a(n_36299), .o(n_36300) );
na02s01 g744016 ( .a(n_36190), .b(n_36143), .o(n_36299) );
na02s01 g744018 ( .a(n_36882), .b(n_36838), .o(n_36901) );
no02s01 g744019 ( .a(n_36882), .b(n_36880), .o(n_36881) );
in01s01 g744020 ( .a(n_36899), .o(n_36900) );
oa12s01 g744021 ( .a(n_36794), .b(n_36862), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_36899) );
oa12s01 g744022 ( .a(n_46203), .b(n_36860), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37631) );
na02s01 g744023 ( .a(n_36065), .b(n_36096), .o(n_36097) );
na02s02 g744024 ( .a(FE_OCPN890_n_44223), .b(n_35598), .o(n_36306) );
in01s01 g744025 ( .a(n_35625), .o(n_36305) );
no02s04 g744026 ( .a(n_44256), .b(n_35598), .o(n_35625) );
in01s01 g744027 ( .a(n_35707), .o(n_35624) );
na02s06 g744028 ( .a(n_44256), .b(n_34263), .o(n_35707) );
in01s01 g744029 ( .a(n_35596), .o(n_35597) );
na02s02 g744030 ( .a(n_35550), .b(n_34262), .o(n_35596) );
na02s01 g744031 ( .a(FE_OCPN890_n_44223), .b(FE_OCPUNCON1759_n_35644), .o(n_36304) );
in01s01 g744033 ( .a(n_35669), .o(n_35700) );
no02m08 g744034 ( .a(FE_OCP_RBN4904_n_44256), .b(FE_OCPUNCON1759_n_35644), .o(n_35669) );
na02s01 g744035 ( .a(FE_OCPN890_n_44223), .b(FE_RN_2661_0), .o(n_36298) );
na02s01 g744036 ( .a(n_44222), .b(n_35703), .o(n_36267) );
no02s04 g744037 ( .a(FE_OCP_RBN4902_n_44256), .b(n_34541), .o(n_35754) );
no02s06 g744038 ( .a(FE_OCP_RBN4904_n_44256), .b(n_34540), .o(n_35751) );
no02s04 g744039 ( .a(FE_OCP_RBN4902_n_44256), .b(n_35667), .o(n_35755) );
no02s01 g744040 ( .a(FE_OCPN890_n_44223), .b(n_34724), .o(n_36297) );
in01s01 g744042 ( .a(n_35699), .o(n_35744) );
na02s02 g744043 ( .a(FE_OCP_RBN4903_n_44256), .b(n_34676), .o(n_35699) );
na02s01 g744044 ( .a(FE_OCPN890_n_44223), .b(n_34712), .o(n_36303) );
na02s01 g744045 ( .a(FE_OCPN890_n_44223), .b(n_35749), .o(n_36295) );
na02s01 g744046 ( .a(n_44222), .b(n_34660), .o(n_36265) );
na02s04 g744047 ( .a(FE_OCP_RBN4904_n_44256), .b(n_34678), .o(n_35831) );
in01s01 g744048 ( .a(n_35747), .o(n_35698) );
na02s02 g744049 ( .a(FE_OCP_RBN4903_n_44256), .b(n_34677), .o(n_35747) );
in01s01 g744050 ( .a(n_35696), .o(n_35697) );
no02s04 g744051 ( .a(n_44222), .b(n_35665), .o(n_35696) );
na02s01 g744052 ( .a(n_44222), .b(n_35665), .o(n_36264) );
no02s10 g744053 ( .a(FE_OCP_RBN4909_n_44222), .b(n_34752), .o(n_35826) );
no02s02 g744054 ( .a(FE_OCP_RBN4904_n_44256), .b(n_34751), .o(n_35827) );
no02s01 g744055 ( .a(FE_OCPN890_n_44223), .b(n_34772), .o(n_36294) );
no02s03 g744056 ( .a(FE_OCP_RBN4910_n_44222), .b(n_35785), .o(n_36331) );
no02s06 g744057 ( .a(FE_OCP_RBN4910_n_44222), .b(n_35742), .o(n_35911) );
in01s01 g744058 ( .a(n_35784), .o(n_35909) );
na02s01 g744059 ( .a(FE_OCP_RBN4903_n_44256), .b(n_35742), .o(n_35784) );
no02s06 g744060 ( .a(FE_OCP_RBN4910_n_44222), .b(n_34861), .o(n_35910) );
no02s01 g744061 ( .a(FE_OCPN890_n_44223), .b(n_35824), .o(n_36293) );
no02m03 g744066 ( .a(n_35905), .b(FE_OCP_RBN4910_n_44222), .o(n_35984) );
no02s01 TIMEBOOST_cell_1099 ( .a(n_37445), .b(n_37097), .o(TIMEBOOST_net_164) );
in01s01 g744068 ( .a(n_47267), .o(n_36007) );
in01m01 g744071 ( .a(n_35948), .o(n_36035) );
na02m01 g744072 ( .a(n_35977), .b(FE_OCP_RBN4910_n_44222), .o(n_35948) );
no02s01 g744073 ( .a(FE_OCP_RBN4910_n_44222), .b(n_35006), .o(n_36036) );
no02s20 TIMEBOOST_cell_1101 ( .a(n_23378), .b(n_23022), .o(TIMEBOOST_net_165) );
no02s01 g744075 ( .a(FE_OCP_RBN6076_n_44256), .b(n_34903), .o(n_36147) );
no02s02 g744076 ( .a(FE_OCP_RBN4910_n_44222), .b(FE_OCP_RBN7038_n_34903), .o(n_36148) );
no02s01 g744077 ( .a(FE_OCP_RBN4910_n_44222), .b(FE_OCP_RBN5899_n_35005), .o(n_36098) );
no02s03 TIMEBOOST_cell_5520 ( .a(n_5947), .b(n_5963), .o(TIMEBOOST_net_1708) );
na02s01 g744079 ( .a(FE_OCP_RBN6076_n_44256), .b(FE_OCP_RBN2896_n_35003), .o(n_36198) );
na02s01 g744080 ( .a(FE_OCP_RBN4910_n_44222), .b(n_35003), .o(n_36191) );
na02s01 g744081 ( .a(FE_OCP_RBN6076_n_44256), .b(n_34996), .o(n_36143) );
na02s01 g744082 ( .a(FE_OCP_RBN4910_n_44222), .b(n_34978), .o(n_36190) );
na02s01 g744083 ( .a(n_35522), .b(n_35537), .o(n_35523) );
in01s01 g744084 ( .a(n_35622), .o(n_35623) );
no02m04 g744085 ( .a(n_35595), .b(n_35594), .o(n_35622) );
in01s01 g744086 ( .a(n_35650), .o(n_35621) );
no02f02 TIMEBOOST_cell_8765 ( .a(TIMEBOOST_net_2869), .b(n_14129), .o(n_14185) );
na02s02 g744090 ( .a(n_35901), .b(n_44040), .o(n_36192) );
na02s02 g744091 ( .a(n_44256), .b(n_34629), .o(n_35643) );
in01s01 g744092 ( .a(n_35693), .o(n_35694) );
no02s06 g744094 ( .a(n_44222), .b(n_34713), .o(n_35752) );
no02m02 g744095 ( .a(FE_OCP_RBN6076_n_44256), .b(n_35060), .o(n_36531) );
in01s01 g744096 ( .a(n_35691), .o(n_35692) );
no02f04 TIMEBOOST_cell_4999 ( .a(TIMEBOOST_net_1447), .b(n_13379), .o(n_13380) );
na02m08 g744098 ( .a(n_35612), .b(FE_OCP_RBN3168_n_44211), .o(n_35663) );
na02f04 TIMEBOOST_cell_8790 ( .a(FE_OCP_RBN3049_n_15200), .b(FE_OCP_RBN2837_n_13962), .o(TIMEBOOST_net_2882) );
na02s06 TIMEBOOST_cell_8767 ( .a(TIMEBOOST_net_2870), .b(n_38138), .o(n_38185) );
in01s01 g744101 ( .a(n_36034), .o(n_35947) );
na02s02 g744102 ( .a(n_35819), .b(FE_OCP_RBN3171_n_44211), .o(n_36034) );
no02s10 TIMEBOOST_cell_3390 ( .a(n_36011), .b(FE_RN_2485_0), .o(TIMEBOOST_net_986) );
no03m08 TIMEBOOST_cell_4670 ( .a(n_19141), .b(n_19032), .c(n_19180), .o(n_19355) );
in01s01 g744105 ( .a(n_36915), .o(n_36916) );
oa22s01 g744106 ( .a(n_36870), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_1_), .c(n_36871), .d(n_36898), .o(n_36915) );
in01s01 g744107 ( .a(n_35593), .o(n_35646) );
in01s01 g744108 ( .a(n_35574), .o(n_35593) );
ao12f06 g744109 ( .a(n_35490), .b(n_35556), .c(n_35515), .o(n_35574) );
oa12s01 g744110 ( .a(n_35552), .b(n_35551), .c(n_35556), .o(n_35592) );
na02s06 g744112 ( .a(n_35547), .b(n_35590), .o(n_35591) );
in01s01 g744113 ( .a(n_35640), .o(n_35641) );
no02s06 g744114 ( .a(n_35620), .b(n_35619), .o(n_35640) );
no02s01 g744115 ( .a(n_35729), .b(n_35690), .o(n_35782) );
no02s01 g744121 ( .a(n_47265), .b(n_35900), .o(n_35901) );
in01s01 g744122 ( .a(n_36065), .o(n_36066) );
no02s01 g744123 ( .a(n_36030), .b(n_36000), .o(n_36065) );
in01s01 g744124 ( .a(n_36262), .o(n_36263) );
na02s01 g744125 ( .a(n_36184), .b(n_36243), .o(n_36262) );
no02f02 TIMEBOOST_cell_8764 ( .a(n_14127), .b(n_13437), .o(TIMEBOOST_net_2869) );
no02s02 g744127 ( .a(n_35531), .b(n_35554), .o(n_35555) );
in01s01 g744128 ( .a(n_36260), .o(n_36261) );
na02s01 g744129 ( .a(n_36136), .b(n_36242), .o(n_36260) );
in01s01 g744130 ( .a(n_35638), .o(n_35639) );
na02s01 g744131 ( .a(n_35590), .b(n_35615), .o(n_35638) );
no03m04 TIMEBOOST_cell_6471 ( .a(n_34201), .b(n_34200), .c(FE_OCP_RBN5712_n_44102), .o(TIMEBOOST_net_1534) );
in01s01 g744133 ( .a(n_36240), .o(n_36241) );
na02s01 g744134 ( .a(n_36188), .b(n_35588), .o(n_36240) );
na02m08 g744135 ( .a(n_35615), .b(n_35611), .o(n_35612) );
in01s01 g744136 ( .a(n_35737), .o(n_35738) );
no02s01 g744137 ( .a(n_35616), .b(n_35690), .o(n_35737) );
in01s01 g744138 ( .a(n_35778), .o(n_35779) );
no02s01 g744139 ( .a(n_35739), .b(n_35736), .o(n_35778) );
no02s06 g744140 ( .a(n_35690), .b(n_35567), .o(n_35689) );
no02s06 TIMEBOOST_cell_3395 ( .a(TIMEBOOST_net_988), .b(FE_OCP_RBN6177_n_36444), .o(n_36516) );
in01s01 g744142 ( .a(n_35859), .o(n_35860) );
no02s01 g744143 ( .a(n_35821), .b(n_35820), .o(n_35859) );
na02s04 TIMEBOOST_cell_8766 ( .a(FE_OCP_RBN6571_n_44875), .b(n_37598), .o(TIMEBOOST_net_2870) );
na02s01 g744146 ( .a(n_35776), .b(n_35899), .o(n_35945) );
in01s01 g744147 ( .a(n_36004), .o(n_36005) );
no02s02 g744148 ( .a(n_47265), .b(n_35974), .o(n_36004) );
na02s01 g744149 ( .a(n_35776), .b(FE_OCP_RBN4925_n_34980), .o(n_35819) );
in01s01 g744150 ( .a(n_36139), .o(n_36140) );
no02s01 g744151 ( .a(n_36095), .b(n_36000), .o(n_36139) );
no03m02 TIMEBOOST_cell_4629 ( .a(n_18942), .b(n_18890), .c(FE_OCP_RBN7026_n_18866), .o(n_19054) );
no02s01 TIMEBOOST_cell_953 ( .a(n_99), .b(n_122), .o(TIMEBOOST_net_91) );
no02s01 g744154 ( .a(n_35575), .b(n_35533), .o(n_35834) );
oa12s01 g744155 ( .a(n_46223), .b(n_46222), .c(n_36898), .o(n_36882) );
no02s01 g744156 ( .a(n_35520), .b(n_35553), .o(n_35670) );
na02f06 g744157 ( .a(n_35517), .b(n_35545), .o(n_35573) );
na02s01 g744158 ( .a(n_35551), .b(n_35556), .o(n_35552) );
no02s01 g744159 ( .a(n_35566), .b(n_35546), .o(n_35709) );
ao12m08 g744200 ( .a(n_35265), .b(n_35532), .c(n_35285), .o(n_35550) );
ao12s01 g744201 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n_46215), .c(n_36747), .o(n_36863) );
in01s01 g744202 ( .a(n_36291), .o(n_36292) );
oa22s01 g744203 ( .a(FE_OCPN1612_n_44174), .b(n_34899), .c(FE_OCP_RBN3167_n_44211), .d(n_35611), .o(n_36291) );
in01s01 g744204 ( .a(n_36258), .o(n_36259) );
no02s01 g744205 ( .a(n_36133), .b(n_35620), .o(n_36258) );
in01s01 g744206 ( .a(n_36256), .o(n_36257) );
no02s01 g744207 ( .a(n_36132), .b(n_35617), .o(n_36256) );
in01s01 g744208 ( .a(n_36254), .o(n_36255) );
no02s01 g744209 ( .a(n_36130), .b(n_35740), .o(n_36254) );
in01s01 g744210 ( .a(n_36238), .o(n_36239) );
na02s01 g744211 ( .a(n_36090), .b(n_35780), .o(n_36238) );
in01s01 g744212 ( .a(n_35971), .o(n_35972) );
na02s01 g744213 ( .a(n_35857), .b(n_35814), .o(n_35971) );
in01s01 g744214 ( .a(n_36093), .o(n_36094) );
no02s02 g744215 ( .a(n_35900), .b(n_36001), .o(n_36093) );
in01s01 g744216 ( .a(n_36186), .o(n_36187) );
no02s01 g744217 ( .a(n_36030), .b(n_36059), .o(n_36186) );
in01s01 g744218 ( .a(n_36236), .o(n_36237) );
no02s01 TIMEBOOST_cell_5512 ( .a(FE_OCP_RBN3308_n_43022), .b(n_43005), .o(TIMEBOOST_net_1704) );
oa12f08 g744220 ( .a(n_35429), .b(n_35495), .c(n_35459), .o(n_35537) );
in01s01 g744221 ( .a(n_36289), .o(n_36290) );
na02s01 g744222 ( .a(n_36183), .b(n_36138), .o(n_36289) );
in01s01 g744223 ( .a(n_36287), .o(n_36288) );
na02s01 g744224 ( .a(n_36182), .b(n_36134), .o(n_36287) );
in01s01 g744225 ( .a(n_36234), .o(n_36235) );
na02s01 g744226 ( .a(n_36088), .b(n_36058), .o(n_36234) );
oa12s01 g744227 ( .a(n_35489), .b(n_35488), .c(n_35495), .o(n_35507) );
in01m01 g744229 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_4_), .o(n_35506) );
na02s01 g744231 ( .a(n_46203), .b(n_46214), .o(n_36841) );
no02s01 g744232 ( .a(n_36816), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_10_), .o(n_36862) );
no02s01 g744233 ( .a(n_36859), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_22_), .o(n_36861) );
no02s01 g744234 ( .a(n_36811), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_18_), .o(n_36860) );
no02s01 g744235 ( .a(n_46225), .b(n_36859), .o(n_37727) );
na02s01 g744236 ( .a(n_46209), .b(n_36838), .o(n_36880) );
in01s01 g744237 ( .a(n_36870), .o(n_36871) );
na02s01 g744238 ( .a(n_46223), .b(n_36822), .o(n_36870) );
no02s01 g744239 ( .a(n_46220), .b(n_36808), .o(n_37381) );
na02s01 g744240 ( .a(n_46219), .b(n_36820), .o(n_37259) );
na02s01 g744241 ( .a(n_46228), .b(n_36855), .o(n_37958) );
no02s01 g744242 ( .a(n_46216), .b(n_36854), .o(n_37839) );
in01s01 g744243 ( .a(n_36868), .o(n_36869) );
na02s01 g744244 ( .a(n_46206), .b(n_36810), .o(n_36868) );
na02s01 g744245 ( .a(n_46214), .b(n_36852), .o(n_37672) );
in01s01 g744246 ( .a(n_35531), .o(n_36243) );
no02s02 g744247 ( .a(n_35487), .b(n_35521), .o(n_35531) );
in01s01 g744248 ( .a(n_36184), .o(n_36185) );
na02s01 g744249 ( .a(FE_OCP_RBN6046_n_35487), .b(n_35521), .o(n_36184) );
no02s06 g744251 ( .a(n_35487), .b(n_34516), .o(n_35533) );
na02s01 g744252 ( .a(FE_OCPN1612_n_44174), .b(n_35554), .o(n_36183) );
na02s01 g744253 ( .a(FE_OCP_RBN6046_n_35487), .b(n_34893), .o(n_36138) );
na02s20 TIMEBOOST_cell_6005 ( .a(FE_OCPN6915_n_23112), .b(n_23111), .o(TIMEBOOST_net_1854) );
na02s01 g744255 ( .a(FE_OCPN1612_n_44174), .b(n_36091), .o(n_36242) );
in01s01 g744256 ( .a(n_36135), .o(n_36136) );
no02s01 g744257 ( .a(FE_OCPN1612_n_44174), .b(n_36091), .o(n_36135) );
na02s01 g744258 ( .a(FE_OCPN1612_n_44174), .b(n_34869), .o(n_36182) );
na02s01 g744259 ( .a(FE_OCP_RBN3167_n_44211), .b(n_35613), .o(n_36134) );
na02m08 g744260 ( .a(FE_OCP_RBN3170_n_44211), .b(n_34766), .o(n_35615) );
in01s01 g744261 ( .a(n_35590), .o(n_35570) );
na02s06 g744262 ( .a(FE_OCP_RBN3167_n_44211), .b(n_34765), .o(n_35590) );
na02s04 g744263 ( .a(FE_OCP_RBN3167_n_44211), .b(n_35611), .o(n_35547) );
na02s01 g744264 ( .a(FE_OCPN1612_n_44174), .b(n_35569), .o(n_36188) );
in01s01 g744265 ( .a(n_35619), .o(n_35588) );
no02s02 g744266 ( .a(FE_OCP_RBN3168_n_44211), .b(n_35569), .o(n_35619) );
no02s01 g744267 ( .a(FE_OCP_RBN6048_n_35487), .b(FE_RN_1790_0), .o(n_36133) );
no02s02 g744268 ( .a(FE_OCP_RBN3168_n_44211), .b(n_34919), .o(n_35620) );
in01s01 g744270 ( .a(n_35616), .o(n_35587) );
no02s02 g744271 ( .a(FE_OCP_RBN3171_n_44211), .b(n_34870), .o(n_35616) );
no02s01 g744272 ( .a(FE_OCP_RBN6048_n_35487), .b(n_34926), .o(n_36132) );
no02s02 g744273 ( .a(FE_OCP_RBN3171_n_44211), .b(n_35567), .o(n_35617) );
no02s06 g744274 ( .a(FE_OCP_RBN6048_n_35487), .b(n_34966), .o(n_35736) );
no02s02 g744275 ( .a(FE_OCP_RBN3171_n_44211), .b(n_34967), .o(n_35739) );
no02s01 g744276 ( .a(FE_OCP_RBN6048_n_35487), .b(n_34989), .o(n_36130) );
no02s01 g744277 ( .a(FE_OCP_RBN3171_n_44211), .b(n_35659), .o(n_35740) );
in01s01 g744278 ( .a(n_35687), .o(n_35820) );
na02s01 g744279 ( .a(FE_OCP_RBN3171_n_44211), .b(FE_OCP_DRV_N1498_n_34924), .o(n_35687) );
in01s01 g744280 ( .a(n_35732), .o(n_35821) );
na02s01 g744281 ( .a(FE_OCPN950_n_44180), .b(n_34925), .o(n_35732) );
na02s01 g744282 ( .a(FE_OCPN950_n_44180), .b(n_35684), .o(n_35780) );
na02s01 g744283 ( .a(FE_OCPN1612_n_44174), .b(n_35025), .o(n_36090) );
in01s01 g744285 ( .a(n_35776), .o(n_35815) );
na02s01 g744286 ( .a(FE_OCP_RBN3171_n_44211), .b(FE_OCP_RBN4260_n_34921), .o(n_35776) );
na02s01 g744288 ( .a(FE_OCPN950_n_44180), .b(n_35774), .o(n_35899) );
na02s01 g744290 ( .a(FE_OCPN950_n_44180), .b(FE_OCP_RBN4925_n_34980), .o(n_35857) );
na02s01 g744291 ( .a(FE_OCP_RBN3171_n_44211), .b(FE_OCP_RBN4924_n_34980), .o(n_35814) );
in01s01 g744292 ( .a(n_35856), .o(n_35974) );
na02s01 g744293 ( .a(FE_OCP_RBN3171_n_44211), .b(n_34946), .o(n_35856) );
no02s01 g744296 ( .a(FE_OCPN950_n_44180), .b(n_35897), .o(n_36001) );
no02s01 g744297 ( .a(FE_OCP_RBN3171_n_44211), .b(n_34999), .o(n_35900) );
no02s01 g744298 ( .a(FE_OCPN950_n_44180), .b(n_35090), .o(n_36095) );
no02m01 g744302 ( .a(FE_OCP_RBN3171_n_44211), .b(n_35193), .o(n_36000) );
no02s01 g744303 ( .a(FE_OCPN950_n_44180), .b(n_35132), .o(n_36059) );
no02s01 g744304 ( .a(FE_OCP_RBN3171_n_44211), .b(n_35194), .o(n_36030) );
no02f06 TIMEBOOST_cell_5511 ( .a(TIMEBOOST_net_1703), .b(FE_RN_1197_0), .o(n_21953) );
na02s01 g744306 ( .a(FE_OCPN950_n_44180), .b(FE_OCP_RBN6787_n_35130), .o(n_36096) );
na02s01 g744307 ( .a(FE_OCPN950_n_44180), .b(n_35113), .o(n_36058) );
na02s01 g744308 ( .a(FE_OCPN1612_n_44174), .b(n_35092), .o(n_36088) );
in01s01 g744311 ( .a(n_46246), .o(n_36851) );
in01s01 g744313 ( .a(n_46245), .o(n_36849) );
in01s01 g744315 ( .a(n_35519), .o(n_35520) );
na02s03 g744316 ( .a(n_35505), .b(n_35504), .o(n_35519) );
no02f04 g744317 ( .a(n_35505), .b(n_35504), .o(n_35553) );
na02s01 g744318 ( .a(n_35488), .b(n_35495), .o(n_35489) );
in01s01 g744319 ( .a(n_35565), .o(n_35566) );
na02f06 g744320 ( .a(n_35513), .b(n_34152), .o(n_35565) );
in01s01 g744321 ( .a(n_35545), .o(n_35546) );
na02m06 g744322 ( .a(n_35512), .b(FE_OCPUNCON7067_n_34151), .o(n_35545) );
no02s01 g744323 ( .a(FE_OCP_RBN3206_n_35517), .b(n_35516), .o(n_35645) );
no02s06 g744325 ( .a(FE_OCP_RBN3168_n_44211), .b(n_34895), .o(n_36075) );
in01s01 g744327 ( .a(n_35683), .o(n_35729) );
no02s01 g744329 ( .a(FE_OCPN950_n_44180), .b(n_35195), .o(n_36063) );
oa12f08 g744330 ( .a(n_35440), .b(n_35503), .c(n_35465), .o(n_35556) );
oa12s01 g744331 ( .a(n_35494), .b(n_35493), .c(n_35503), .o(n_35518) );
in01s02 g744348 ( .a(delay_sub_ln23_0_unr28_stage10_stallmux_q), .o(n_41337) );
in01s01 g744351 ( .a(n_46227), .o(n_36855) );
in01s01 g744354 ( .a(n_46225), .o(n_36826) );
in01s01 g744356 ( .a(n_46224), .o(n_36824) );
in01s01 g744359 ( .a(n_46222), .o(n_36822) );
in01s01 g744361 ( .a(n_46221), .o(n_36820) );
in01s01 g744363 ( .a(n_46220), .o(n_36818) );
in01s01 g744365 ( .a(n_46219), .o(n_36816) );
in01s01 g744368 ( .a(n_46217), .o(n_36852) );
in01s01 g744370 ( .a(n_46216), .o(n_36814) );
in01s01 g744372 ( .a(n_46215), .o(n_36854) );
in01s01 g744374 ( .a(n_46214), .o(n_36811) );
in01s01 g744376 ( .a(n_46213), .o(n_36810) );
in01s01 g744378 ( .a(n_46212), .o(n_36808) );
na02s01 g744380 ( .a(n_35854), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_36838) );
in01s01 g744381 ( .a(n_46211), .o(n_36859) );
in01s01 g744385 ( .a(n_46208), .o(n_36805) );
in01s01 g744389 ( .a(n_36793), .o(n_36794) );
ao12s01 g744390 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n_36785), .c(n_36784), .o(n_36793) );
no02s01 g744392 ( .a(n_35485), .b(n_35502), .o(n_35577) );
na02f04 g744395 ( .a(n_35501), .b(FE_OCPUNCON3484_n_35500), .o(n_35517) );
in01s01 g744397 ( .a(n_35516), .o(n_35529) );
no02m06 g744398 ( .a(n_35501), .b(FE_OCPUNCON3484_n_35500), .o(n_35516) );
na02s01 g744399 ( .a(n_35493), .b(n_35503), .o(n_35494) );
na02s01 g744400 ( .a(n_35491), .b(n_35515), .o(n_35551) );
in01m02 g744402 ( .a(n_35532), .o(n_35499) );
na02m08 g744403 ( .a(n_35471), .b(n_35468), .o(n_35532) );
ao12m10 g744445 ( .a(FE_OCP_RBN4344_n_35177), .b(n_35475), .c(n_35148), .o(n_35487) );
ao12f08 g744447 ( .a(n_35385), .b(n_35460), .c(n_35410), .o(n_35495) );
oa12s01 g744448 ( .a(n_35450), .b(n_35449), .c(n_35460), .o(n_35474) );
in01m02 g744449 ( .a(n_35512), .o(n_35513) );
na02s02 TIMEBOOST_cell_5440 ( .a(n_9964), .b(n_9624), .o(TIMEBOOST_net_1668) );
in01s02 g744452 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_3_), .o(n_35473) );
na02s01 g744456 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_), .o(n_36775) );
no02s01 g744457 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_), .o(n_36774) );
na02s01 TIMEBOOST_cell_8045 ( .a(TIMEBOOST_net_2653), .b(n_47274), .o(n_32124) );
na02f08 TIMEBOOST_cell_5439 ( .a(TIMEBOOST_net_1667), .b(n_15953), .o(n_16169) );
no02f20 TIMEBOOST_cell_968 ( .a(TIMEBOOST_net_98), .b(n_28096), .o(n_28123) );
in01s01 g744461 ( .a(n_35484), .o(n_35485) );
na02m04 g744462 ( .a(n_35470), .b(n_35469), .o(n_35484) );
no02m04 g744463 ( .a(n_35470), .b(n_35469), .o(n_35502) );
na02s01 g744464 ( .a(n_35449), .b(n_35460), .o(n_35450) );
no02s01 g744465 ( .a(n_35459), .b(n_35430), .o(n_35488) );
na02s01 g744466 ( .a(n_35536), .b(n_35446), .o(n_35522) );
in01s01 g744467 ( .a(n_35490), .o(n_35491) );
no02f04 g744468 ( .a(n_35483), .b(FE_OCPUNCON1757_n_35482), .o(n_35490) );
na02f04 g744469 ( .a(n_35483), .b(FE_OCPUNCON1757_n_35482), .o(n_35515) );
na02m08 TIMEBOOST_cell_966 ( .a(TIMEBOOST_net_97), .b(n_40936), .o(n_46947) );
na02f04 TIMEBOOST_cell_5447 ( .a(TIMEBOOST_net_1671), .b(n_5488), .o(n_5651) );
ao12f08 g744472 ( .a(n_35393), .b(n_35467), .c(n_35418), .o(n_35503) );
oa12s01 g744473 ( .a(n_35457), .b(n_35456), .c(n_35467), .o(n_35481) );
in01s01 g744474 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_), .o(n_36762) );
in01s01 g744477 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_), .o(n_36773) );
in01s01 g744481 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_2_), .o(n_35466) );
na02s06 TIMEBOOST_cell_965 ( .a(n_40878), .b(n_40934), .o(TIMEBOOST_net_97) );
no02m06 TIMEBOOST_cell_4470 ( .a(TIMEBOOST_net_1325), .b(n_39527), .o(n_39575) );
na02m04 g744485 ( .a(n_35423), .b(n_35359), .o(n_35447) );
no02f04 g744486 ( .a(n_35416), .b(n_35415), .o(n_35459) );
in01s01 g744487 ( .a(n_35429), .o(n_35430) );
na02f04 g744488 ( .a(n_35416), .b(n_35415), .o(n_35429) );
na02m06 g744489 ( .a(n_35428), .b(FE_OCP_DRV_N1484_n_35427), .o(n_35536) );
in01s01 g744490 ( .a(n_35535), .o(n_35446) );
no02f06 g744491 ( .a(n_35428), .b(FE_OCP_DRV_N1484_n_35427), .o(n_35535) );
na02s01 g744492 ( .a(n_35456), .b(n_35467), .o(n_35457) );
no02s01 g744493 ( .a(n_35441), .b(n_35465), .o(n_35493) );
no02s04 g744494 ( .a(n_35425), .b(n_35344), .o(n_35455) );
no02s06 TIMEBOOST_cell_6330 ( .a(TIMEBOOST_net_2016), .b(FE_OCP_RBN4471_n_31819), .o(n_31968) );
in01f02 g744496 ( .a(n_35475), .o(n_35443) );
na02f10 g744497 ( .a(n_35405), .b(n_35401), .o(n_35475) );
no02m20 TIMEBOOST_cell_967 ( .a(n_27999), .b(FE_RN_1890_0), .o(TIMEBOOST_net_98) );
oa22s02 g744499 ( .a(n_36684), .b(n_36176), .c(n_36683), .d(n_36177), .o(n_36729) );
no02m01 TIMEBOOST_cell_3324 ( .a(FE_OCP_RBN6203_n_31819), .b(n_30541), .o(TIMEBOOST_net_953) );
oa12f08 g744501 ( .a(n_35317), .b(n_35414), .c(n_35351), .o(n_35460) );
oa12s01 g744502 ( .a(n_35403), .b(n_35402), .c(n_35414), .o(n_35426) );
oa12m02 g744504 ( .a(n_36685), .b(n_36682), .c(n_36049), .o(n_36728) );
in01s01 g744506 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_26_), .o(n_36747) );
na02s01 g744509 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_19_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_20_), .o(n_36727) );
na02s01 g744510 ( .a(n_36745), .b(n_36744), .o(n_36746) );
in01s02 g744511 ( .a(n_35444), .o(n_35425) );
na02m08 g744512 ( .a(n_35413), .b(n_35342), .o(n_35444) );
in01s02 g744513 ( .a(n_35423), .o(n_35424) );
no02s03 g744514 ( .a(n_35413), .b(n_35283), .o(n_35423) );
na02f08 TIMEBOOST_cell_8651 ( .a(TIMEBOOST_net_2812), .b(n_26378), .o(n_26524) );
no02s10 TIMEBOOST_cell_8712 ( .a(n_17975), .b(n_17971), .o(TIMEBOOST_net_2843) );
no02m02 g744519 ( .a(n_35364), .b(n_35231), .o(n_35404) );
na02s01 g744520 ( .a(n_35402), .b(n_35414), .o(n_35403) );
na02s01 g744521 ( .a(n_35386), .b(n_35410), .o(n_35449) );
in01s01 g744522 ( .a(n_35440), .o(n_35441) );
na02f04 g744523 ( .a(n_35421), .b(FE_OCPUNCON1755_n_35420), .o(n_35440) );
no02m06 g744524 ( .a(n_35421), .b(FE_OCPUNCON1755_n_35420), .o(n_35465) );
no02f04 TIMEBOOST_cell_6851 ( .a(n_21154), .b(FE_OCP_RBN1604_n_20995), .o(TIMEBOOST_net_2183) );
oa22s01 g744526 ( .a(n_36664), .b(n_36162), .c(FE_OCP_RBN3429_n_36664), .d(n_36161), .o(n_36714) );
oa22s02 g744527 ( .a(n_36644), .b(n_36211), .c(n_36645), .d(n_36212), .o(n_36700) );
oa22m01 g744528 ( .a(n_36678), .b(n_36250), .c(n_36662), .d(n_36251), .o(n_36726) );
no02f04 TIMEBOOST_cell_7684 ( .a(n_42139), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(TIMEBOOST_net_2473) );
oa12s01 g744531 ( .a(n_35398), .b(n_35397), .c(n_35396), .o(n_35419) );
oa12s01 g744533 ( .a(n_35439), .b(n_35438), .c(n_35437), .o(n_35464) );
in01s01 g744534 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_19_), .o(n_36745) );
in01s01 g744537 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_), .o(n_36713) );
no02m08 g744540 ( .a(n_35387), .b(n_35284), .o(n_35413) );
na02m04 g744542 ( .a(n_35387), .b(n_35224), .o(n_35399) );
na02s02 TIMEBOOST_cell_5077 ( .a(TIMEBOOST_net_1486), .b(n_41701), .o(n_41771) );
na02m04 g744544 ( .a(n_35333), .b(n_35236), .o(n_35353) );
na02s02 g744546 ( .a(n_36662), .b(n_36681), .o(n_36685) );
in01s01 g744548 ( .a(n_35385), .o(n_35386) );
na02s01 g744550 ( .a(n_35397), .b(n_35396), .o(n_35398) );
na02s01 g744552 ( .a(n_35438), .b(n_35437), .o(n_35439) );
na02s01 g744553 ( .a(n_35394), .b(n_35418), .o(n_35456) );
no02m04 TIMEBOOST_cell_5256 ( .a(n_20203), .b(n_20183), .o(TIMEBOOST_net_1576) );
na02s04 TIMEBOOST_cell_6814 ( .a(TIMEBOOST_net_2164), .b(n_11025), .o(n_11137) );
na02s02 g744556 ( .a(n_35365), .b(n_35257), .o(n_35364) );
oa22s01 g744557 ( .a(n_36639), .b(n_36213), .c(n_36638), .d(n_36214), .o(n_36699) );
oa22s01 g744558 ( .a(n_36623), .b(n_36169), .c(n_36642), .d(n_36170), .o(n_36698) );
in01s02 g744559 ( .a(n_36683), .o(n_36684) );
oa12s04 g744560 ( .a(FE_OCPN1953_n_36121), .b(n_36623), .c(FE_OCPN1955_n_36050), .o(n_36683) );
ao12m02 g744561 ( .a(n_36681), .b(n_36622), .c(n_36178), .o(n_36682) );
ao12f08 g744562 ( .a(n_35363), .b(n_35328), .c(n_35330), .o(n_35414) );
oa12s01 g744564 ( .a(n_35381), .b(n_35380), .c(n_35379), .o(n_35409) );
in01s01 g744567 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_20_), .o(n_36744) );
na02m08 g744569 ( .a(n_35329), .b(n_35223), .o(n_35387) );
in01s02 g744570 ( .a(n_35365), .o(n_35352) );
in01s02 g744572 ( .a(n_35333), .o(n_35334) );
na02s04 g744573 ( .a(n_35290), .b(n_35211), .o(n_35333) );
no02s01 g744574 ( .a(n_35363), .b(n_35331), .o(n_35397) );
no02s01 g744575 ( .a(n_35318), .b(n_35351), .o(n_35402) );
na02m06 g744576 ( .a(n_35383), .b(FE_OCPUNCON1753_n_35382), .o(n_35418) );
in01s01 g744577 ( .a(n_35393), .o(n_35394) );
no02f04 g744578 ( .a(n_35383), .b(FE_OCPUNCON1753_n_35382), .o(n_35393) );
na02s01 g744579 ( .a(n_35379), .b(n_35380), .o(n_35381) );
no02s01 g744580 ( .a(n_35376), .b(n_35361), .o(n_35438) );
no02f04 g744582 ( .a(n_35296), .b(n_35152), .o(n_35332) );
oa22s02 g744583 ( .a(n_36599), .b(n_36155), .c(n_36600), .d(n_36156), .o(n_36666) );
oa22s01 g744584 ( .a(n_36598), .b(n_36052), .c(n_36619), .d(n_36053), .o(n_36680) );
oa12s02 g744586 ( .a(n_36021), .b(n_36598), .c(n_35880), .o(n_36664) );
oa22s01 g744587 ( .a(n_36601), .b(n_36219), .c(n_36577), .d(n_36220), .o(n_36663) );
in01s01 g744588 ( .a(n_36644), .o(n_36645) );
oa12s02 g744589 ( .a(n_36171), .b(n_36577), .c(n_36080), .o(n_36644) );
in01s01 g744591 ( .a(n_36662), .o(n_36678) );
no02s04 g744592 ( .a(n_36621), .b(n_36284), .o(n_36662) );
oa12s01 g744594 ( .a(n_35350), .b(n_35349), .c(FE_OCP_RBN4643_n_35121), .o(n_35378) );
in01s01 g744595 ( .a(n_35377), .o(n_35437) );
oa12f06 g744596 ( .a(n_35313), .b(n_35314), .c(n_35345), .o(n_35377) );
in01s01 g744598 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_0_), .o(n_35362) );
no02f04 g744602 ( .a(n_45327), .b(n_35294), .o(n_35296) );
in01s01 g744603 ( .a(n_35317), .o(n_35318) );
na02f06 g744604 ( .a(n_35293), .b(FE_OCP_DRV_N1424_n_35292), .o(n_35317) );
no02m08 g744605 ( .a(n_35293), .b(FE_OCP_DRV_N1424_n_35292), .o(n_35351) );
no02f06 g744606 ( .a(n_35316), .b(FE_OCP_DRV_N3510_n_35315), .o(n_35363) );
in01s01 g744607 ( .a(n_35330), .o(n_35331) );
na02f08 g744608 ( .a(n_35316), .b(FE_OCP_DRV_N3510_n_35315), .o(n_35330) );
na02s01 g744609 ( .a(n_35349), .b(FE_OCP_RBN4643_n_35121), .o(n_35350) );
in01s01 g744611 ( .a(n_36623), .o(n_36642) );
na02s03 g744612 ( .a(n_36603), .b(n_36283), .o(n_36623) );
in01s01 g744613 ( .a(n_35375), .o(n_35376) );
na02m06 g744614 ( .a(n_35325), .b(n_33905), .o(n_35375) );
in01s01 g744615 ( .a(n_35360), .o(n_35361) );
na02f08 g744618 ( .a(n_35275), .b(n_35216), .o(n_35290) );
in01f02 g744619 ( .a(n_35346), .o(n_35347) );
in01f02 g744620 ( .a(n_35329), .o(n_35346) );
oa12f06 g744621 ( .a(n_35136), .b(n_35272), .c(n_35134), .o(n_35329) );
oa22s01 g744622 ( .a(n_36571), .b(n_36164), .c(n_36572), .d(n_36165), .o(n_36641) );
oa22s01 g744623 ( .a(n_36575), .b(n_35965), .c(n_36576), .d(n_35964), .o(n_36640) );
oa22s01 g744624 ( .a(n_36574), .b(n_35992), .c(n_36596), .d(n_35993), .o(n_36661) );
in01s01 g744625 ( .a(n_36638), .o(n_36639) );
ao12s02 g744626 ( .a(n_35883), .b(n_36574), .c(n_35961), .o(n_36638) );
in01s02 g744627 ( .a(n_36621), .o(n_36622) );
no02s04 g744628 ( .a(n_36603), .b(n_36084), .o(n_36621) );
in01s01 g744629 ( .a(n_35328), .o(n_35396) );
na02f08 g744630 ( .a(n_35266), .b(n_35273), .o(n_35328) );
oa12s01 g744632 ( .a(n_35311), .b(n_35345), .c(n_35310), .o(n_35380) );
in01s01 g744634 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_), .o(n_36578) );
in01s01 g744636 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_), .o(n_36637) );
na02s02 g744639 ( .a(n_35211), .b(FE_OCP_RBN2980_n_35213), .o(n_35274) );
no02s02 g744640 ( .a(n_35256), .b(n_35213), .o(n_35257) );
in01s01 g744641 ( .a(n_35343), .o(n_35344) );
no02s02 g744642 ( .a(n_35326), .b(n_35283), .o(n_35343) );
no02s04 g744643 ( .a(n_35326), .b(n_35281), .o(n_35327) );
in01m02 g744644 ( .a(n_35358), .o(n_35359) );
in01s01 g744647 ( .a(n_36577), .o(n_36601) );
no02s02 g744648 ( .a(n_36558), .b(n_36228), .o(n_36577) );
na02m06 g744649 ( .a(n_36558), .b(n_36018), .o(n_36603) );
na02f06 g744650 ( .a(n_35251), .b(n_35121), .o(n_35273) );
no02s01 g744651 ( .a(n_35267), .b(n_35252), .o(n_35349) );
no02f06 g744652 ( .a(n_35379), .b(FE_OCP_DRV_N1428_n_35312), .o(n_35314) );
na02f06 g744653 ( .a(n_35379), .b(FE_OCPN1350_n_35312), .o(n_35313) );
na02s01 g744654 ( .a(n_35345), .b(n_35310), .o(n_35311) );
oa22s01 g744658 ( .a(n_36498), .b(n_36216), .c(n_36499), .d(n_36215), .o(n_36542) );
in01s01 g744659 ( .a(n_36599), .o(n_36600) );
oa12s02 g744660 ( .a(n_35889), .b(n_36555), .c(n_35934), .o(n_36599) );
in01s01 g744662 ( .a(n_36598), .o(n_36619) );
oa12s02 g744663 ( .a(n_36125), .b(n_36513), .c(n_35960), .o(n_36598) );
oa12s01 g744664 ( .a(n_35270), .b(n_35269), .c(n_35268), .o(n_35309) );
na02m04 TIMEBOOST_cell_4532 ( .a(TIMEBOOST_net_1356), .b(n_11189), .o(n_11307) );
na02f08 g744666 ( .a(n_35239), .b(n_35215), .o(n_35316) );
in01s01 g744667 ( .a(n_35340), .o(n_35341) );
in01m02 g744669 ( .a(n_35324), .o(n_35325) );
no02s03 TIMEBOOST_cell_6800 ( .a(TIMEBOOST_net_2157), .b(n_4680), .o(n_4954) );
na02s01 g744671 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_), .o(n_36557) );
no02s01 g744672 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_), .o(n_36556) );
no02f08 g744673 ( .a(n_35294), .b(n_35118), .o(n_35216) );
na02f04 g744675 ( .a(n_35178), .b(n_35123), .o(n_35215) );
na02f08 g744676 ( .a(n_35084), .b(n_35179), .o(n_35239) );
in01m02 g744677 ( .a(n_35288), .o(n_35289) );
in01f02 g744678 ( .a(n_35272), .o(n_35288) );
na02f08 g744679 ( .a(n_35200), .b(n_35253), .o(n_35272) );
no02f04 g744680 ( .a(n_44713), .b(n_35229), .o(n_35271) );
na03s02 TIMEBOOST_cell_4671 ( .a(n_8232), .b(TIMEBOOST_net_1064), .c(n_9111), .o(n_9419) );
no02f04 g744682 ( .a(n_35213), .b(n_35207), .o(n_35214) );
no02f06 g744684 ( .a(n_35152), .b(n_35156), .o(n_35237) );
na02s02 TIMEBOOST_cell_5499 ( .a(TIMEBOOST_net_1697), .b(n_22367), .o(n_22496) );
na02m02 TIMEBOOST_cell_4529 ( .a(n_11019), .b(n_10926), .o(TIMEBOOST_net_1355) );
na02m02 g744687 ( .a(n_35235), .b(FE_OCP_RBN2979_n_35213), .o(n_35236) );
no02s02 g744688 ( .a(n_35213), .b(n_35183), .o(n_35234) );
na02s06 g744689 ( .a(n_35287), .b(FE_OCPN6281_n_30612), .o(n_35342) );
no02m06 g744691 ( .a(n_35287), .b(FE_OCPN1376_n_30612), .o(n_35326) );
na02m02 g744692 ( .a(n_35285), .b(n_35264), .o(n_35307) );
no02m04 g744693 ( .a(n_35305), .b(n_35265), .o(n_35323) );
in01s01 g744694 ( .a(n_36575), .o(n_36576) );
na02s02 g744695 ( .a(n_36555), .b(n_35996), .o(n_36575) );
in01s01 g744697 ( .a(n_36574), .o(n_36596) );
na02s02 g744698 ( .a(n_36513), .b(n_36026), .o(n_36574) );
na02s01 g744699 ( .a(n_35269), .b(n_35268), .o(n_35270) );
in01s01 g744700 ( .a(n_35266), .o(n_35267) );
na02m06 g744701 ( .a(n_35199), .b(n_34056), .o(n_35266) );
in01s01 g744702 ( .a(n_35251), .o(n_35252) );
na02f04 g744703 ( .a(n_35198), .b(n_34055), .o(n_35251) );
no02f08 g744704 ( .a(n_35269), .b(FE_OCPN1380_n_33640), .o(n_35379) );
in01s03 g744706 ( .a(n_35211), .o(n_35256) );
oa12s06 g744707 ( .a(n_30633), .b(n_35155), .c(n_35029), .o(n_35211) );
oa22s01 g744708 ( .a(n_36477), .b(n_36217), .c(n_36478), .d(n_36218), .o(n_36528) );
oa22s01 g744709 ( .a(n_36479), .b(n_35967), .c(n_36480), .d(n_35966), .o(n_36527) );
oa22s01 g744710 ( .a(n_36495), .b(n_36172), .c(n_36494), .d(n_36173), .o(n_36573) );
in01s01 g744711 ( .a(n_36571), .o(n_36572) );
oa12s01 g744712 ( .a(n_36122), .b(n_36494), .c(n_35848), .o(n_36571) );
no02m06 g744713 ( .a(n_36513), .b(n_36054), .o(n_36558) );
oa12s01 g744714 ( .a(n_35121), .b(n_35107), .c(FE_OCP_DRV_N1478_n_35106), .o(n_35210) );
no02f06 g744717 ( .a(n_35230), .b(n_35205), .o(n_35345) );
in01s01 g744718 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_), .o(n_36541) );
no02f02 g744720 ( .a(n_35167), .b(n_35204), .o(n_35205) );
no02f04 g744721 ( .a(n_35168), .b(n_35172), .o(n_35230) );
in01s02 g744722 ( .a(n_35184), .o(n_35157) );
no02f10 g744723 ( .a(n_35122), .b(n_35123), .o(n_35184) );
in01s02 g744724 ( .a(n_35253), .o(n_35229) );
no02f08 g744725 ( .a(n_35204), .b(n_35133), .o(n_35253) );
no02m04 g744726 ( .a(n_35101), .b(n_30587), .o(n_35156) );
no02f10 g744727 ( .a(n_35155), .b(n_30546), .o(n_35294) );
in01s01 g744728 ( .a(n_35235), .o(n_35183) );
na02m08 g744729 ( .a(n_35154), .b(FE_OCPN1681_n_30614), .o(n_35235) );
no02f06 g744733 ( .a(n_35154), .b(FE_OCPN1681_n_30614), .o(n_35213) );
na02s02 g744734 ( .a(n_35177), .b(n_35148), .o(n_35201) );
no02m04 g744735 ( .a(FE_OCP_RBN4344_n_35177), .b(n_35175), .o(n_35228) );
in01s01 g744737 ( .a(n_35152), .o(n_35180) );
no02m04 g744738 ( .a(n_35102), .b(FE_OCPN1681_n_30614), .o(n_35152) );
in01m02 g744740 ( .a(n_35285), .o(n_35305) );
na02m08 g744741 ( .a(n_35220), .b(n_30633), .o(n_35285) );
in01s03 g744742 ( .a(n_35264), .o(n_35265) );
na02s03 g744744 ( .a(n_35219), .b(n_30614), .o(n_35264) );
no02m04 g744745 ( .a(n_35169), .b(n_35171), .o(n_35226) );
na02m04 g744746 ( .a(n_35224), .b(n_35223), .o(n_35225) );
na02s02 g744747 ( .a(n_36495), .b(n_35936), .o(n_36555) );
na02s04 g744750 ( .a(n_35107), .b(FE_OCP_DRV_N1478_n_35106), .o(n_35121) );
in01f04 g744751 ( .a(n_35178), .o(n_35179) );
no02m04 TIMEBOOST_cell_4979 ( .a(TIMEBOOST_net_1437), .b(FE_RN_133_0), .o(n_12641) );
no02s04 g744754 ( .a(n_35284), .b(n_35250), .o(n_35303) );
na02f04 g744756 ( .a(n_35141), .b(n_35200), .o(n_35221) );
ao12m06 g744760 ( .a(FE_OCP_DRV_N6893_FE_OCPN6281_n_30612), .b(n_35249), .c(n_35143), .o(n_35283) );
in01s01 g744761 ( .a(n_36498), .o(n_36499) );
oa12s01 g744762 ( .a(n_35970), .b(n_36464), .c(n_35938), .o(n_36498) );
na02f06 g744766 ( .a(n_36476), .b(n_36024), .o(n_36513) );
na02f06 g744767 ( .a(n_35174), .b(n_35150), .o(n_35269) );
in01m02 g744768 ( .a(n_35198), .o(n_35199) );
na02m06 TIMEBOOST_cell_5560 ( .a(n_31359), .b(n_31076), .o(TIMEBOOST_net_1728) );
in01s02 g744771 ( .a(n_35281), .o(n_35282) );
in01m04 g744772 ( .a(n_35262), .o(n_35281) );
na02s01 TIMEBOOST_cell_5982 ( .a(TIMEBOOST_net_1842), .b(n_7219), .o(n_7272) );
in01s01 g744777 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_), .o(n_36497) );
in01f04 g744781 ( .a(n_35123), .o(n_35084) );
na02f02 g744783 ( .a(n_35145), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35150) );
na02m08 g744785 ( .a(n_35100), .b(n_47233), .o(n_35177) );
no02f08 g744786 ( .a(n_35057), .b(n_30588), .o(n_35122) );
in01s02 g744788 ( .a(n_35148), .o(n_35175) );
na02m08 g744789 ( .a(n_35099), .b(n_30633), .o(n_35148) );
in01f02 g744790 ( .a(n_35146), .o(n_35147) );
na02f04 g744791 ( .a(n_35083), .b(n_35119), .o(n_35146) );
na02m06 TIMEBOOST_cell_2114 ( .a(TIMEBOOST_net_671), .b(n_35444), .o(n_35471) );
na02f04 g744793 ( .a(FE_OCP_RBN4870_n_35145), .b(n_30545), .o(n_35174) );
na02s02 TIMEBOOST_cell_5974 ( .a(TIMEBOOST_net_1838), .b(n_12431), .o(n_12666) );
no02m02 g744795 ( .a(n_35194), .b(FE_OCPN5230_n_30587), .o(n_35197) );
in01s01 g744796 ( .a(n_35204), .o(n_35172) );
no02m08 g744797 ( .a(n_35145), .b(n_30545), .o(n_35204) );
na02s06 g744798 ( .a(n_35097), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35200) );
in01s02 g744799 ( .a(n_35223), .o(n_35171) );
na02m08 g744800 ( .a(n_35143), .b(FE_OCPN5280_n_30614), .o(n_35223) );
no02s04 g744801 ( .a(n_35192), .b(FE_OCPN5230_n_30587), .o(n_35284) );
no02s04 TIMEBOOST_cell_4998 ( .a(n_13350), .b(n_13378), .o(TIMEBOOST_net_1447) );
no02m04 g744803 ( .a(FE_OCP_RBN6788_n_35130), .b(FE_OCPN1376_n_30612), .o(n_35196) );
no02s03 g744804 ( .a(n_35249), .b(FE_OCPN6281_n_30612), .o(n_35250) );
in01m04 g744805 ( .a(n_35169), .o(n_35224) );
no02s06 g744806 ( .a(n_35143), .b(FE_OCPN5280_n_30614), .o(n_35169) );
na02f02 g744807 ( .a(n_35098), .b(FE_OCPN5230_n_30587), .o(n_35141) );
in01s01 g744808 ( .a(n_36479), .o(n_36480) );
na02s01 g744809 ( .a(n_36464), .b(n_35941), .o(n_36479) );
no02s01 g744810 ( .a(n_35194), .b(n_35193), .o(n_35195) );
in01m02 g744811 ( .a(n_35139), .o(n_35140) );
no02s06 TIMEBOOST_cell_3152 ( .a(n_16011), .b(FE_OCPN1705_n_14730), .o(TIMEBOOST_net_867) );
oa22s01 g744813 ( .a(n_36450), .b(n_36175), .c(n_36451), .d(n_36174), .o(n_36496) );
in01s01 g744814 ( .a(n_36477), .o(n_36478) );
oa12s01 g744815 ( .a(n_35764), .b(n_36463), .c(n_36123), .o(n_36477) );
in01s02 g744820 ( .a(n_36494), .o(n_36495) );
in01s01 g744821 ( .a(n_36476), .o(n_36494) );
oa12m06 g744822 ( .a(n_35969), .b(n_36463), .c(n_35940), .o(n_36476) );
in01f06 g744824 ( .a(n_35102), .o(n_35155) );
in01m02 g744825 ( .a(n_35102), .o(n_35101) );
no02f06 TIMEBOOST_cell_5985 ( .a(n_28102), .b(n_28041), .o(TIMEBOOST_net_1844) );
na02m08 g744828 ( .a(n_35065), .b(n_35037), .o(n_35207) );
na02s01 TIMEBOOST_cell_5638 ( .a(n_6010), .b(n_5725), .o(TIMEBOOST_net_1767) );
in01s03 g744830 ( .a(n_35219), .o(n_35220) );
no03s08 TIMEBOOST_cell_8189 ( .a(FE_OCPN937_n_17684), .b(n_17683), .c(n_17655), .o(n_17720) );
na02f04 TIMEBOOST_cell_4482 ( .a(TIMEBOOST_net_1331), .b(n_39667), .o(n_39698) );
no02m04 TIMEBOOST_cell_4386 ( .a(TIMEBOOST_net_1283), .b(n_5011), .o(n_5121) );
na02s06 g744834 ( .a(FE_OCP_RBN2895_n_35003), .b(n_30612), .o(n_35065) );
na02s04 g744835 ( .a(n_35003), .b(n_30633), .o(n_35037) );
no02f08 g744836 ( .a(n_35029), .b(n_30546), .o(n_35118) );
no02m08 g744839 ( .a(n_34960), .b(n_30545), .o(n_35012) );
na02s08 g744840 ( .a(n_35063), .b(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35119) );
na02m02 TIMEBOOST_cell_5634 ( .a(n_40536), .b(n_40250), .o(TIMEBOOST_net_1765) );
no02f06 TIMEBOOST_cell_5387 ( .a(TIMEBOOST_net_1641), .b(n_16337), .o(n_16471) );
no02s01 TIMEBOOST_cell_5121 ( .a(TIMEBOOST_net_1508), .b(n_14455), .o(n_14492) );
no02s04 TIMEBOOST_cell_4183 ( .a(n_22304), .b(FE_OCP_RBN2118_n_22351), .o(TIMEBOOST_net_1182) );
na02m02 TIMEBOOST_cell_2112 ( .a(n_30354), .b(TIMEBOOST_net_670), .o(n_30429) );
na02m02 g744849 ( .a(n_35095), .b(n_35136), .o(n_35137) );
no02m02 g744850 ( .a(n_35134), .b(n_35096), .o(n_35135) );
no02s01 g744851 ( .a(FE_OCP_RBN5899_n_35005), .b(FE_OCP_RBN7039_n_34903), .o(n_35060) );
na02f04 g744853 ( .a(n_35009), .b(n_35059), .o(n_35078) );
in01f02 g744854 ( .a(n_35167), .o(n_35168) );
no02f02 g744855 ( .a(n_35093), .b(n_35133), .o(n_35167) );
ao12s01 g744856 ( .a(n_36419), .b(n_36420), .c(n_35797), .o(n_36464) );
oa22s01 g744857 ( .a(n_36405), .b(n_36157), .c(n_36406), .d(n_36158), .o(n_36454) );
no02f04 TIMEBOOST_cell_5177 ( .a(TIMEBOOST_net_1536), .b(n_25039), .o(n_25180) );
in01m04 g744860 ( .a(n_35099), .o(n_35100) );
na03m08 TIMEBOOST_cell_5899 ( .a(n_26880), .b(n_26963), .c(n_26962), .o(n_27041) );
in01f02 g744862 ( .a(n_35057), .o(n_35058) );
na02f06 g744863 ( .a(n_34985), .b(n_34961), .o(n_35057) );
in01m04 g744865 ( .a(n_35132), .o(n_35194) );
in01m02 g744868 ( .a(n_35097), .o(n_35098) );
na02s01 TIMEBOOST_cell_3038 ( .a(n_2895), .b(n_2894), .o(TIMEBOOST_net_810) );
no02m08 g744870 ( .a(n_35055), .b(n_35030), .o(n_35143) );
in01m04 g744871 ( .a(n_35192), .o(n_35249) );
na02s01 TIMEBOOST_cell_5981 ( .a(n_7040), .b(n_7203), .o(TIMEBOOST_net_1842) );
in01s01 g744873 ( .a(FE_OCP_RBN6787_n_35130), .o(n_36062) );
oa22s01 g744877 ( .a(n_36403), .b(n_35886), .c(n_36404), .d(n_35887), .o(n_36453) );
oa22s01 g744878 ( .a(n_46953), .b(n_36210), .c(n_36402), .d(n_36209), .o(n_36452) );
in01s01 g744879 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_8_), .o(n_36785) );
na02m04 g744881 ( .a(n_35001), .b(n_30504), .o(n_35034) );
no02s06 TIMEBOOST_cell_3226 ( .a(n_20763), .b(n_45013), .o(TIMEBOOST_net_904) );
no02s02 TIMEBOOST_cell_6304 ( .a(TIMEBOOST_net_2003), .b(n_10934), .o(n_11055) );
na02s06 g744884 ( .a(n_34955), .b(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35059) );
na02f04 g744885 ( .a(n_34933), .b(n_30588), .o(n_34985) );
na02s04 g744886 ( .a(n_34934), .b(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34961) );
na02f02 g744887 ( .a(n_34956), .b(n_30504), .o(n_35009) );
no02f04 TIMEBOOST_cell_6213 ( .a(n_35058), .b(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(TIMEBOOST_net_1958) );
in01m01 g744889 ( .a(n_35136), .o(n_35096) );
na02m04 g744890 ( .a(n_35077), .b(FE_OCPN5230_n_30587), .o(n_35136) );
in01m01 g744891 ( .a(n_35134), .o(n_35095) );
no02m04 g744892 ( .a(n_35077), .b(FE_OCPN5230_n_30587), .o(n_35134) );
no02s06 g744893 ( .a(n_35046), .b(n_30588), .o(n_35133) );
na02m04 TIMEBOOST_cell_3037 ( .a(TIMEBOOST_net_809), .b(FE_OCP_RBN6640_n_24268), .o(n_24398) );
no02m02 g744895 ( .a(n_34980), .b(n_30504), .o(n_35008) );
no02s04 g744896 ( .a(n_34999), .b(n_30546), .o(n_35030) );
no02m08 g744897 ( .a(n_35897), .b(FE_OCP_DRV_N6893_FE_OCPN6281_n_30612), .o(n_35055) );
na02s06 TIMEBOOST_cell_6924 ( .a(TIMEBOOST_net_2220), .b(n_2699), .o(n_2805) );
na02s02 TIMEBOOST_cell_6664 ( .a(TIMEBOOST_net_2089), .b(n_8077), .o(FE_RN_299_0) );
no02f02 g744900 ( .a(n_35047), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35093) );
in01s01 g744901 ( .a(n_36450), .o(n_36451) );
in01s01 g744902 ( .a(n_36463), .o(n_36450) );
no02m06 g744903 ( .a(n_36420), .b(n_36419), .o(n_36463) );
in01s01 g744905 ( .a(n_34960), .o(n_34983) );
na02m08 g744906 ( .a(n_34883), .b(n_34864), .o(n_34960) );
in01s02 g744908 ( .a(n_35029), .o(n_35053) );
na02m08 g744909 ( .a(n_34959), .b(n_34936), .o(n_35029) );
no02f08 g744910 ( .a(n_34957), .b(n_34935), .o(n_35063) );
in01s02 g744912 ( .a(n_35092), .o(n_35113) );
oa22m02 g744914 ( .a(n_34990), .b(n_34743), .c(n_34991), .d(n_34744), .o(n_35092) );
in01s01 g744915 ( .a(n_35980), .o(n_35006) );
in01s01 g744916 ( .a(n_34982), .o(n_35980) );
in01m02 g744917 ( .a(n_34982), .o(n_34981) );
oa22s06 g744927 ( .a(n_34906), .b(n_34447), .c(n_34907), .d(n_34448), .o(n_35003) );
in01s01 g744928 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_7_), .o(n_36784) );
no02m06 g744931 ( .a(n_34972), .b(n_34654), .o(n_35049) );
na02m06 g744932 ( .a(n_34835), .b(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34883) );
na02s04 g744933 ( .a(n_34836), .b(n_30588), .o(n_34864) );
na02m08 g744934 ( .a(FE_OCP_RBN7039_n_34903), .b(n_30546), .o(n_34959) );
na02s04 g744935 ( .a(n_34903), .b(FE_OFN5087_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34936) );
no02f06 g744936 ( .a(n_35977), .b(n_30504), .o(n_34957) );
no02s03 g744937 ( .a(n_34905), .b(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34935) );
no02m04 g744938 ( .a(n_36154), .b(n_36385), .o(n_36420) );
oa12m08 g744939 ( .a(n_34651), .b(FE_OCP_RBN2930_n_34971), .c(n_34993), .o(n_35026) );
no02s02 TIMEBOOST_cell_5976 ( .a(TIMEBOOST_net_1839), .b(n_23107), .o(TIMEBOOST_net_112) );
oa22s01 g744941 ( .a(n_36386), .b(n_36168), .c(n_36356), .d(n_36167), .o(n_36418) );
in01s01 g744942 ( .a(n_36405), .o(n_36406) );
oa12s01 g744943 ( .a(n_36117), .b(n_36386), .c(n_35630), .o(n_36405) );
in01s01 g744944 ( .a(n_35684), .o(n_35025) );
in01s01 g744945 ( .a(n_35001), .o(n_35684) );
in01f04 g744946 ( .a(n_35001), .o(n_35000) );
in01m02 g744948 ( .a(n_34955), .o(n_34956) );
no02m04 TIMEBOOST_cell_4389 ( .a(n_30496), .b(n_30141), .o(TIMEBOOST_net_1285) );
in01f01 g744951 ( .a(n_35046), .o(n_35047) );
na02f04 g744952 ( .a(n_34974), .b(n_34952), .o(n_35046) );
in01m04 g744959 ( .a(n_34999), .o(n_35897) );
in01s01 g744962 ( .a(n_35193), .o(n_35090) );
in01s03 g744963 ( .a(n_35075), .o(n_35193) );
no03m04 TIMEBOOST_cell_8278 ( .a(FE_OCP_RBN2780_n_8664), .b(FE_RN_1774_0), .c(n_8895), .o(FE_RN_1775_0) );
in01s02 g744966 ( .a(n_35905), .o(n_34954) );
in01s02 g744967 ( .a(n_34934), .o(n_35905) );
in01f02 g744968 ( .a(n_34934), .o(n_34933) );
in01s02 g744971 ( .a(n_34978), .o(n_34996) );
oa22m04 g744973 ( .a(n_34878), .b(n_34445), .c(FE_OCP_RBN4261_n_34878), .d(n_34446), .o(n_34978) );
in01s01 g744974 ( .a(n_36403), .o(n_36404) );
oa12s01 g744975 ( .a(n_35795), .b(n_36386), .c(n_35807), .o(n_36403) );
in01s01 g744976 ( .a(n_46953), .o(n_36402) );
na02f06 TIMEBOOST_cell_4996 ( .a(n_41313), .b(delay_sub_ln23_0_unr28_stage10_stallmux_q), .o(TIMEBOOST_net_1446) );
no02s01 TIMEBOOST_cell_5929 ( .a(FE_RN_724_0), .b(FE_RN_725_0), .o(TIMEBOOST_net_1816) );
no02s02 TIMEBOOST_cell_3043 ( .a(n_24402), .b(TIMEBOOST_net_812), .o(n_24467) );
na02f08 TIMEBOOST_cell_4388 ( .a(n_20476), .b(TIMEBOOST_net_1284), .o(FE_RN_110_0) );
no03f08 TIMEBOOST_cell_8335 ( .a(TIMEBOOST_net_874), .b(n_34769), .c(n_34362), .o(n_34905) );
na02s01 TIMEBOOST_cell_3039 ( .a(TIMEBOOST_net_810), .b(n_3633), .o(n_3736) );
na02s02 g744984 ( .a(n_34923), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34953) );
na02f02 g744985 ( .a(FE_OCP_RBN4258_n_34921), .b(n_30504), .o(n_34974) );
na02s02 g744986 ( .a(n_34921), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34952) );
no03m08 TIMEBOOST_cell_660 ( .a(n_11056), .b(n_11124), .c(n_11053), .o(n_11209) );
in01s03 g744989 ( .a(n_34906), .o(n_34907) );
no02s02 TIMEBOOST_cell_3100 ( .a(FE_RN_701_0), .b(FE_RN_702_0), .o(TIMEBOOST_net_841) );
no02m06 g744991 ( .a(n_34971), .b(n_34652), .o(n_34972) );
in01s01 g744992 ( .a(n_34990), .o(n_34991) );
in01m04 g744994 ( .a(n_34880), .o(n_34881) );
na02m06 g744995 ( .a(n_34797), .b(n_34338), .o(n_34880) );
oa22s01 g744996 ( .a(n_36314), .b(n_36159), .c(n_36313), .d(n_36160), .o(n_36384) );
in01s01 g744997 ( .a(n_35659), .o(n_34989) );
oa12s02 g744998 ( .a(n_34931), .b(n_34930), .c(n_34929), .o(n_35659) );
in01s01 g744999 ( .a(n_35824), .o(n_34861) );
in01s01 g745000 ( .a(n_34836), .o(n_35824) );
in01m02 g745001 ( .a(n_34836), .o(n_34835) );
in01m04 g745003 ( .a(n_34905), .o(n_35977) );
no02s02 TIMEBOOST_cell_6618 ( .a(TIMEBOOST_net_2066), .b(n_17971), .o(n_18054) );
no02f06 TIMEBOOST_cell_6065 ( .a(n_12902), .b(FE_OCP_RBN5580_n_12753), .o(TIMEBOOST_net_1884) );
na02f04 g745011 ( .a(n_36315), .b(n_35808), .o(n_36385) );
in01s01 g745012 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_6_), .o(n_36358) );
no02m08 TIMEBOOST_cell_5593 ( .a(TIMEBOOST_net_1744), .b(n_31953), .o(n_31971) );
na02f06 TIMEBOOST_cell_3099 ( .a(TIMEBOOST_net_840), .b(n_25528), .o(n_25640) );
na02s01 g745016 ( .a(n_34930), .b(n_34929), .o(n_34931) );
no02m10 g745018 ( .a(n_34747), .b(n_34927), .o(n_34971) );
na02m04 g745019 ( .a(n_34795), .b(FE_OCP_RBN5743_n_34278), .o(n_34797) );
na02s02 TIMEBOOST_cell_1543 ( .a(FE_OCP_RBN2078_n_14149), .b(FE_RN_1467_0), .o(TIMEBOOST_net_386) );
na02m08 TIMEBOOST_cell_4975 ( .a(TIMEBOOST_net_1435), .b(n_18019), .o(n_18106) );
na03s02 TIMEBOOST_cell_8261 ( .a(n_41345), .b(FE_OCP_RBN5676_n_41420), .c(n_41771), .o(n_41831) );
no02s06 TIMEBOOST_cell_6657 ( .a(n_7784), .b(n_8453), .o(TIMEBOOST_net_2086) );
no02m04 g745025 ( .a(n_45185), .b(n_34397), .o(n_34830) );
in01s01 TIMEBOOST_cell_5924 ( .a(TIMEBOOST_net_1812), .o(TIMEBOOST_net_1813) );
in01f02 g745028 ( .a(n_34876), .o(n_34877) );
oa12f04 g745029 ( .a(n_34506), .b(n_34786), .c(n_34535), .o(n_34876) );
oa12m04 g745030 ( .a(n_34537), .b(n_34858), .c(FE_OCP_RBN2816_n_34509), .o(n_34875) );
na02s04 TIMEBOOST_cell_3834 ( .a(TIMEBOOST_net_1007), .b(n_1551), .o(n_47027) );
oa12m08 g745033 ( .a(n_34380), .b(n_34873), .c(FE_OCPN5268_n_34852), .o(n_34874) );
no02m02 TIMEBOOST_cell_5568 ( .a(n_31014), .b(n_30938), .o(TIMEBOOST_net_1732) );
oa12f08 g745035 ( .a(n_34238), .b(n_34753), .c(n_47254), .o(n_34793) );
na02s04 TIMEBOOST_cell_8808 ( .a(n_10806), .b(n_44511), .o(TIMEBOOST_net_2891) );
in01s01 g745037 ( .a(n_35567), .o(n_34926) );
oa12s02 g745038 ( .a(n_34856), .b(n_34855), .c(n_34854), .o(n_35567) );
in01s01 g745039 ( .a(FE_OCP_DRV_N1498_n_34924), .o(n_34925) );
oa12s01 g745040 ( .a(n_34851), .b(n_34873), .c(n_34850), .o(n_34924) );
in01s02 g745044 ( .a(n_34923), .o(n_34946) );
no02m08 TIMEBOOST_cell_4988 ( .a(n_37597), .b(n_37709), .o(TIMEBOOST_net_1442) );
in01s01 g745047 ( .a(FE_OCP_RBN4260_n_34921), .o(n_35774) );
in01s01 g745051 ( .a(n_35785), .o(n_34772) );
oa12s02 g745052 ( .a(n_34718), .b(n_34717), .c(n_34716), .o(n_35785) );
in01s01 g745053 ( .a(n_35861), .o(n_35906) );
in01s01 g745054 ( .a(n_34828), .o(n_35861) );
in01s03 g745055 ( .a(n_34828), .o(n_34827) );
no03s02 TIMEBOOST_cell_7678 ( .a(n_2674), .b(n_2888), .c(FE_OCP_RBN5644_n_2674), .o(TIMEBOOST_net_2470) );
in01s01 g745058 ( .a(n_36386), .o(n_36356) );
in01s01 g745059 ( .a(n_36315), .o(n_36386) );
ao12f04 g745060 ( .a(n_35718), .b(n_36232), .c(n_35769), .o(n_36315) );
na02f40 TIMEBOOST_cell_3831 ( .a(n_27776), .b(FE_OCP_RBN7127_n_44722), .o(TIMEBOOST_net_1006) );
na02m06 TIMEBOOST_cell_4165 ( .a(n_40170), .b(n_40438), .o(TIMEBOOST_net_1173) );
na02s02 TIMEBOOST_cell_2111 ( .a(n_30176), .b(n_30143), .o(TIMEBOOST_net_670) );
na02s01 g745065 ( .a(n_34855), .b(n_34854), .o(n_34856) );
na03f08 TIMEBOOST_cell_8245 ( .a(TIMEBOOST_net_2701), .b(FE_RN_2376_0), .c(TIMEBOOST_net_223), .o(TIMEBOOST_net_2413) );
no03m08 TIMEBOOST_cell_661 ( .a(FE_RN_1121_0), .b(n_10955), .c(n_10958), .o(n_11074) );
in01s01 g745068 ( .a(n_36313), .o(n_36314) );
no02s01 g745069 ( .a(n_36233), .b(n_35654), .o(n_36313) );
na02s01 g745070 ( .a(n_34850), .b(n_34873), .o(n_34851) );
na02s01 g745071 ( .a(n_34717), .b(n_34716), .o(n_34718) );
na02m08 TIMEBOOST_cell_8487 ( .a(TIMEBOOST_net_2730), .b(n_32908), .o(n_33014) );
na02s06 g745073 ( .a(n_34711), .b(n_34281), .o(n_34730) );
na02s02 TIMEBOOST_cell_8115 ( .a(TIMEBOOST_net_2688), .b(n_11582), .o(TIMEBOOST_net_1791) );
oa12s01 g745075 ( .a(n_34817), .b(n_34897), .c(n_34846), .o(n_34930) );
oa12m04 g745077 ( .a(n_34241), .b(n_34714), .c(n_34687), .o(n_34715) );
no02m08 TIMEBOOST_cell_8727 ( .a(TIMEBOOST_net_2850), .b(n_23500), .o(n_23576) );
oa22s01 g745079 ( .a(n_36180), .b(n_35767), .c(n_36179), .d(n_35768), .o(n_36286) );
in01s01 g745080 ( .a(n_35611), .o(n_34899) );
ao12s02 g745081 ( .a(n_34825), .b(n_34824), .c(n_34823), .o(n_35611) );
in01s01 g745082 ( .a(FE_RN_1790_0), .o(n_34919) );
ao12s01 g745083 ( .a(n_34849), .b(n_34848), .c(n_34847), .o(n_34947) );
oa12s01 g745085 ( .a(n_34791), .b(n_34790), .c(n_34789), .o(n_34870) );
in01s01 g745086 ( .a(n_34966), .o(n_34967) );
ao12s01 g745087 ( .a(n_34898), .b(n_34897), .c(n_34896), .o(n_34966) );
oa12s01 g745088 ( .a(n_34686), .b(n_34714), .c(n_34685), .o(n_35742) );
in01s02 g745089 ( .a(n_34795), .o(n_34769) );
ao12f08 g745090 ( .a(n_34437), .b(n_34661), .c(n_34267), .o(n_34795) );
ao12m02 g745092 ( .a(n_34489), .b(n_34661), .c(n_34368), .o(n_34768) );
no02s01 g745093 ( .a(n_34824), .b(n_34823), .o(n_34825) );
no02s01 g745094 ( .a(n_34848), .b(n_34847), .o(n_34849) );
no02s01 g745095 ( .a(n_34897), .b(n_34896), .o(n_34898) );
na02s01 TIMEBOOST_cell_5949 ( .a(n_37357), .b(n_37049), .o(TIMEBOOST_net_1826) );
na02s01 g745097 ( .a(n_34790), .b(n_34789), .o(n_34791) );
na02s01 g745098 ( .a(n_34685), .b(n_34714), .o(n_34686) );
no02s01 g745099 ( .a(n_35613), .b(n_34706), .o(n_34895) );
no02s01 g745100 ( .a(n_35749), .b(n_34712), .o(n_34713) );
in01s01 g745101 ( .a(n_34753), .o(n_34754) );
in01f06 g745102 ( .a(n_34728), .o(n_34753) );
in01m04 g745103 ( .a(n_34728), .o(n_34727) );
in01f08 g745104 ( .a(n_34711), .o(n_34728) );
no02f10 g745105 ( .a(n_34661), .b(n_34375), .o(n_34711) );
in01s04 g745106 ( .a(n_34788), .o(n_34858) );
ao12m04 g745108 ( .a(n_34655), .b(n_34767), .c(n_34539), .o(n_34788) );
in01f08 g745109 ( .a(n_34822), .o(n_34872) );
in01f06 g745110 ( .a(n_34786), .o(n_34822) );
ao12f08 g745111 ( .a(n_34591), .b(n_34767), .c(n_34488), .o(n_34786) );
oa12s01 g745112 ( .a(n_34176), .b(n_34683), .c(n_34618), .o(n_34717) );
ao12s01 g745113 ( .a(n_34464), .b(n_34749), .c(n_34460), .o(n_34855) );
oa22s01 g745114 ( .a(n_36252), .b(n_36114), .c(n_36253), .d(n_36113), .o(n_36330) );
in01s01 g745116 ( .a(n_35665), .o(n_34726) );
oa12s01 g745117 ( .a(n_34664), .b(n_34663), .c(n_34662), .o(n_35665) );
in01s01 g745118 ( .a(n_34751), .o(n_34752) );
ao12s01 g745119 ( .a(n_34684), .b(n_34683), .c(n_34682), .o(n_34751) );
in01s01 g745120 ( .a(n_36232), .o(n_36233) );
ao12f04 g745121 ( .a(n_36126), .b(n_36127), .c(n_35724), .o(n_36232) );
in01s01 g745122 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_), .o(n_36355) );
no02s01 g745125 ( .a(n_34514), .b(n_34767), .o(n_34897) );
na02s01 g745126 ( .a(n_34663), .b(n_34662), .o(n_34664) );
no02s01 g745127 ( .a(n_34683), .b(n_34682), .o(n_34684) );
na02m06 g745128 ( .a(n_34632), .b(n_34342), .o(n_34714) );
no02s01 g745129 ( .a(n_34749), .b(n_34435), .o(n_34790) );
in01s01 g745130 ( .a(n_36179), .o(n_36180) );
no02s01 g745131 ( .a(n_36127), .b(n_36126), .o(n_36179) );
ao12s01 g745132 ( .a(n_34377), .b(n_34725), .c(n_34344), .o(n_34824) );
oa12s01 g745133 ( .a(n_34348), .b(n_34820), .c(n_34764), .o(n_34848) );
in01s01 g745138 ( .a(n_35613), .o(n_34869) );
ao12s01 g745139 ( .a(n_34785), .b(n_34784), .c(n_34783), .o(n_35613) );
in01s01 g745140 ( .a(n_34765), .o(n_34766) );
ao12s01 g745141 ( .a(n_34710), .b(n_34725), .c(n_34709), .o(n_34765) );
in01s01 g745142 ( .a(n_34894), .o(n_35569) );
ao12s01 g745143 ( .a(n_34821), .b(n_34820), .c(n_34819), .o(n_34894) );
in01s01 g745144 ( .a(FE_RN_2666_0), .o(n_34724) );
oa12s01 g745145 ( .a(n_34659), .b(n_34658), .c(n_34657), .o(n_35667) );
in01s01 g745146 ( .a(n_35749), .o(n_34660) );
ao12s01 g745147 ( .a(n_34577), .b(n_34576), .c(n_34575), .o(n_35749) );
in01s01 g745148 ( .a(n_34677), .o(n_34678) );
oa12s01 g745149 ( .a(n_34605), .b(n_34604), .c(n_34603), .o(n_34677) );
no02s01 g745150 ( .a(n_34725), .b(n_34709), .o(n_34710) );
no02s01 g745151 ( .a(n_34784), .b(n_34783), .o(n_34785) );
no02s01 g745152 ( .a(n_34576), .b(n_34575), .o(n_34577) );
na02s01 g745153 ( .a(n_34604), .b(n_34603), .o(n_34605) );
no02s01 g745154 ( .a(n_34820), .b(n_34399), .o(n_34749) );
na02s01 g745155 ( .a(n_34658), .b(n_34657), .o(n_34659) );
no02s01 g745156 ( .a(n_34574), .b(n_34287), .o(n_34683) );
no02s01 g745158 ( .a(n_34819), .b(n_34820), .o(n_34821) );
na02s01 g745159 ( .a(n_35554), .b(n_34628), .o(n_34918) );
no02m04 g745160 ( .a(n_36056), .b(n_36055), .o(n_36127) );
oa12s01 g745162 ( .a(n_36231), .b(n_36230), .c(n_36229), .o(n_36285) );
in01s01 g745163 ( .a(n_36252), .o(n_36253) );
na02s01 g745164 ( .a(n_36056), .b(n_36112), .o(n_36252) );
ao12s01 g745165 ( .a(n_34220), .b(n_34542), .c(n_34203), .o(n_34663) );
no02s01 g745166 ( .a(n_34542), .b(n_34193), .o(n_34604) );
na02s01 g745167 ( .a(n_36230), .b(n_36229), .o(n_36231) );
ao12s01 g745169 ( .a(n_34434), .b(n_34656), .c(n_34412), .o(n_34725) );
oa12s01 g745170 ( .a(n_34477), .b(n_34601), .c(n_34522), .o(n_34576) );
na02f04 TIMEBOOST_cell_6721 ( .a(n_24057), .b(n_23661), .o(TIMEBOOST_net_2118) );
oa12s01 g745173 ( .a(n_34405), .b(n_34656), .c(n_34340), .o(n_34784) );
oa12s01 g745174 ( .a(n_34187), .b(n_34494), .c(n_34128), .o(n_34658) );
in01s01 g745175 ( .a(n_35554), .o(n_34893) );
na02s01 g745176 ( .a(n_34782), .b(n_34818), .o(n_35554) );
in01s01 g745177 ( .a(n_34706), .o(n_36091) );
ao12s01 g745178 ( .a(n_34631), .b(n_34656), .c(n_34630), .o(n_34706) );
in01s01 g745179 ( .a(n_34540), .o(n_34541) );
ao12s01 g745180 ( .a(n_34467), .b(n_34494), .c(n_34466), .o(n_34540) );
in01s01 g745181 ( .a(n_34712), .o(n_34676) );
ao12s01 g745182 ( .a(n_34602), .b(n_34601), .c(n_34600), .o(n_34712) );
na02f04 g745183 ( .a(n_36230), .b(n_35604), .o(n_36056) );
in01s01 g745184 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_), .o(n_36354) );
na02s01 g745186 ( .a(n_34594), .b(n_34763), .o(n_34818) );
na02s01 g745187 ( .a(n_34595), .b(n_34762), .o(n_34782) );
no02s01 g745188 ( .a(n_34494), .b(n_34466), .o(n_34467) );
no02s01 g745189 ( .a(n_34601), .b(n_34600), .o(n_34602) );
no02s01 g745190 ( .a(n_34656), .b(n_34630), .o(n_34631) );
na02s01 g745191 ( .a(n_36283), .b(n_36221), .o(n_36284) );
in01s01 g745192 ( .a(n_34493), .o(n_34542) );
na02s06 TIMEBOOST_cell_4967 ( .a(TIMEBOOST_net_1431), .b(n_32915), .o(n_32978) );
in01s01 g745195 ( .a(FE_RN_2661_0), .o(n_35703) );
ao12s01 g745196 ( .a(n_34598), .b(n_34597), .c(n_34596), .o(n_34707) );
oa12f04 g745197 ( .a(n_35770), .b(n_35810), .c(FE_OCP_RBN3292_n_35539), .o(n_36230) );
no02s01 g745198 ( .a(n_34597), .b(n_34596), .o(n_34598) );
no02s02 g745199 ( .a(n_36228), .b(n_36023), .o(n_36283) );
na02s01 g745200 ( .a(n_35648), .b(FE_OCPUNCON3490_n_34327), .o(n_34629) );
in01s01 g745201 ( .a(n_34594), .o(n_34595) );
oa12s01 g745202 ( .a(n_34290), .b(n_34573), .c(n_34353), .o(n_34594) );
in01s01 g745203 ( .a(n_34440), .o(n_34601) );
in01s01 g745205 ( .a(n_34572), .o(n_34656) );
oa12f08 g745206 ( .a(n_34355), .b(n_34492), .c(n_34384), .o(n_34572) );
oa12s01 g745207 ( .a(n_34136), .b(n_34415), .c(n_34414), .o(n_34494) );
oa12s01 g745208 ( .a(n_36227), .b(n_36226), .c(n_36225), .o(n_36282) );
in01s01 g745209 ( .a(n_35521), .o(n_34628) );
ao22s01 g745210 ( .a(n_34573), .b(n_34378), .c(n_34518), .d(n_34379), .o(n_35521) );
in01s01 g745211 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_2_), .o(n_36353) );
no02s01 g745213 ( .a(n_34358), .b(n_34480), .o(n_34597) );
in01s01 g745214 ( .a(n_36228), .o(n_36178) );
na02f04 TIMEBOOST_cell_5629 ( .a(TIMEBOOST_net_1762), .b(n_16558), .o(n_16686) );
na02s01 g745216 ( .a(n_36226), .b(n_36225), .o(n_36227) );
no02f04 g745217 ( .a(n_36226), .b(n_35809), .o(n_35810) );
in01s01 g745218 ( .a(n_35648), .o(n_34593) );
oa12s01 g745219 ( .a(n_34521), .b(n_34520), .c(n_34519), .o(n_35648) );
ao12s01 g745220 ( .a(n_34571), .b(n_34570), .c(n_34569), .o(n_35644) );
in01s01 g745221 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_1_), .o(n_35854) );
na02s01 g745223 ( .a(n_34520), .b(n_34519), .o(n_34521) );
no02s01 g745224 ( .a(n_34570), .b(n_34569), .o(n_34571) );
in01s01 g745225 ( .a(n_34415), .o(n_34358) );
no02s02 g745227 ( .a(n_36025), .b(n_35930), .o(n_36125) );
na02s04 g745228 ( .a(n_35682), .b(n_35809), .o(n_35770) );
in01s01 g745229 ( .a(n_36250), .o(n_36251) );
na02s01 g745230 ( .a(n_36086), .b(n_36124), .o(n_36250) );
oa12s01 g745231 ( .a(n_36224), .b(n_36223), .c(n_36222), .o(n_36281) );
in01s01 g745232 ( .a(n_34573), .o(n_34518) );
in01s01 g745233 ( .a(n_34492), .o(n_34573) );
ao12f08 g745234 ( .a(n_34376), .b(n_34465), .c(n_34310), .o(n_34492) );
ao12s01 g745236 ( .a(n_34439), .b(n_34465), .c(n_34438), .o(n_34516) );
na02f04 g745237 ( .a(n_35681), .b(n_35584), .o(n_36226) );
na02m04 g745238 ( .a(n_34592), .b(n_34627), .o(n_34655) );
na02s01 g745239 ( .a(n_35853), .b(n_35795), .o(n_36419) );
no02s01 g745240 ( .a(n_35968), .b(n_35937), .o(n_35970) );
no03s01 TIMEBOOST_cell_8350 ( .a(n_31223), .b(FE_OCP_RBN4418_n_31117), .c(n_31224), .o(TIMEBOOST_net_1629) );
in01s01 g745242 ( .a(n_36025), .o(n_36026) );
na02s01 g745243 ( .a(n_35996), .b(n_35939), .o(n_36025) );
na02s01 g745244 ( .a(n_35725), .b(n_36049), .o(n_36124) );
na02s01 g745245 ( .a(n_36681), .b(FE_OCP_RBN3303_n_35539), .o(n_36086) );
na02s01 g745246 ( .a(n_36223), .b(n_36222), .o(n_36224) );
no02s01 g745247 ( .a(n_34438), .b(n_34465), .o(n_34439) );
oa12s01 g745248 ( .a(n_34119), .b(n_34275), .c(n_34149), .o(n_34520) );
ao12f08 g745249 ( .a(n_34131), .b(n_34275), .c(n_34150), .o(n_34570) );
oa12s01 g745250 ( .a(n_35657), .b(n_35656), .c(FE_OFN231_n_35655), .o(n_35726) );
in01s01 g745251 ( .a(FE_OCPUNCON3490_n_34327), .o(n_35598) );
oa12s01 g745252 ( .a(n_34265), .b(n_34275), .c(n_34264), .o(n_34327) );
in01m02 g745253 ( .a(n_35681), .o(n_35682) );
no02s02 TIMEBOOST_cell_6906 ( .a(TIMEBOOST_net_2211), .b(n_8163), .o(TIMEBOOST_net_1470) );
na02s01 g745255 ( .a(n_35656), .b(FE_OFN231_n_35655), .o(n_35657) );
na02s01 g745256 ( .a(n_36083), .b(n_36121), .o(n_36084) );
na02s01 g745257 ( .a(n_34264), .b(n_34275), .o(n_34265) );
ao12s01 g745258 ( .a(n_34747), .b(n_34675), .c(FE_OCP_RBN6668_n_34297), .o(n_34748) );
no02s02 g745259 ( .a(n_35807), .b(n_35715), .o(n_35808) );
in01m02 g745260 ( .a(n_34591), .o(n_34592) );
no02s01 TIMEBOOST_cell_8490 ( .a(n_37541), .b(n_37540), .o(TIMEBOOST_net_2732) );
no03f06 TIMEBOOST_cell_5480 ( .a(n_35146), .b(n_35184), .c(n_35147), .o(TIMEBOOST_net_1688) );
in01s01 g745263 ( .a(n_35968), .o(n_35941) );
no02s01 g745264 ( .a(n_35806), .b(FE_OCP_RBN3292_n_35539), .o(n_35968) );
na02s01 g745265 ( .a(n_35851), .b(n_35849), .o(n_35940) );
na03m06 TIMEBOOST_cell_4808 ( .a(FE_OCPN1942_n_20723), .b(n_22267), .c(FE_OCP_RBN6878_n_44267), .o(n_22381) );
no02s08 TIMEBOOST_cell_2982 ( .a(n_19105), .b(n_18708), .o(TIMEBOOST_net_782) );
no02s01 g745268 ( .a(n_35963), .b(n_35935), .o(n_36024) );
na02s01 g745269 ( .a(n_35994), .b(n_35959), .o(n_36054) );
no02s01 TIMEBOOST_cell_5930 ( .a(TIMEBOOST_net_1816), .b(n_27899), .o(FE_RN_727_0) );
ao12s01 g745271 ( .a(FE_OCP_RBN3300_n_35539), .b(n_36171), .c(n_36022), .o(n_36023) );
in01s01 g745272 ( .a(n_36176), .o(n_36177) );
oa12s01 g745273 ( .a(n_36083), .b(FE_OCP_RBN3303_n_35539), .c(n_36118), .o(n_36176) );
in01s01 g745274 ( .a(n_36681), .o(n_35725) );
no02s01 g745275 ( .a(n_35635), .b(n_35606), .o(n_36681) );
ao12s01 g745276 ( .a(n_34387), .b(n_34386), .c(n_34385), .o(n_35504) );
ao12f08 g745277 ( .a(n_34272), .b(n_34326), .c(n_34245), .o(n_34465) );
na02s01 g745278 ( .a(n_36120), .b(n_36049), .o(n_36221) );
oa12m04 g745279 ( .a(n_35561), .b(n_35605), .c(FE_OFN231_n_35655), .o(n_36222) );
na02s02 g745280 ( .a(n_35680), .b(FE_OCP_RBN3295_n_35539), .o(n_35769) );
no02s20 TIMEBOOST_cell_8698 ( .a(n_27822), .b(FE_OCP_RBN7128_n_44722), .o(TIMEBOOST_net_2836) );
in01s01 g745285 ( .a(n_36174), .o(n_36175) );
no02s01 g745286 ( .a(n_36123), .b(n_35805), .o(n_36174) );
no02s01 g745287 ( .a(n_35805), .b(n_35804), .o(n_35806) );
in01s01 g745288 ( .a(n_35966), .o(n_35967) );
no02s01 g745289 ( .a(n_35938), .b(n_35937), .o(n_35966) );
in01s01 g745290 ( .a(n_36172), .o(n_36173) );
na02s01 g745291 ( .a(n_36122), .b(n_35890), .o(n_36172) );
in01s01 g745292 ( .a(n_35935), .o(n_35936) );
na02s01 g745293 ( .a(n_35890), .b(n_35891), .o(n_35935) );
in01s01 g745294 ( .a(n_35964), .o(n_35965) );
no02s01 g745295 ( .a(n_35934), .b(n_35888), .o(n_35964) );
no02s01 g745296 ( .a(n_35888), .b(n_35839), .o(n_35889) );
na02s01 g745297 ( .a(n_35962), .b(n_35847), .o(n_35963) );
in01s01 g745298 ( .a(n_36052), .o(n_36053) );
na02s01 g745299 ( .a(n_36021), .b(n_35932), .o(n_36052) );
in01s01 g745300 ( .a(n_36219), .o(n_36220) );
na02s01 g745301 ( .a(n_36081), .b(n_36171), .o(n_36219) );
no03f08 TIMEBOOST_cell_8239 ( .a(n_13272), .b(n_13269), .c(TIMEBOOST_net_1216), .o(n_13435) );
in01s01 g745303 ( .a(n_36169), .o(n_36170) );
na02s01 g745304 ( .a(n_36119), .b(n_36121), .o(n_36169) );
na02s01 g745305 ( .a(n_36118), .b(FE_OCP_RBN3300_n_35539), .o(n_36083) );
no02s01 g745306 ( .a(n_35582), .b(n_35188), .o(n_35635) );
no02s01 g745307 ( .a(n_35581), .b(n_35187), .o(n_35606) );
na02s01 g745308 ( .a(n_36119), .b(n_36118), .o(n_36120) );
in01s01 g745309 ( .a(n_35767), .o(n_35768) );
na02s01 g745310 ( .a(n_35724), .b(n_35679), .o(n_35767) );
no02s01 g745311 ( .a(n_34386), .b(n_34385), .o(n_34387) );
no02s01 g745312 ( .a(n_35928), .b(n_35958), .o(n_35994) );
in01s01 g745313 ( .a(n_35992), .o(n_35993) );
na02s01 g745314 ( .a(n_35961), .b(n_35929), .o(n_35992) );
no02m08 TIMEBOOST_cell_2981 ( .a(TIMEBOOST_net_781), .b(n_29196), .o(n_29273) );
no02s01 g745316 ( .a(n_35562), .b(n_35605), .o(n_35656) );
in01s01 g745317 ( .a(n_36167), .o(n_36168) );
na02s01 g745318 ( .a(n_36117), .b(n_35722), .o(n_36167) );
no02f06 TIMEBOOST_cell_4547 ( .a(FE_RN_153_0), .b(n_16563), .o(TIMEBOOST_net_1364) );
no02s01 g745320 ( .a(n_35850), .b(n_35796), .o(n_35851) );
no02m10 TIMEBOOST_cell_2983 ( .a(TIMEBOOST_net_782), .b(n_19175), .o(n_19264) );
na02s01 g745322 ( .a(n_35679), .b(n_35678), .o(n_35680) );
na02s01 g745323 ( .a(n_35722), .b(n_35723), .o(n_35807) );
in01s01 g745324 ( .a(n_35886), .o(n_35887) );
na02s01 g745325 ( .a(n_35716), .b(n_35717), .o(n_35886) );
in01s01 g745327 ( .a(n_36217), .o(n_36218) );
oa22s01 g745328 ( .a(n_36049), .b(n_35804), .c(FE_OCP_RBN3301_n_35539), .d(n_35259), .o(n_36217) );
in01s01 g745329 ( .a(n_36215), .o(n_36216) );
no02s01 g745330 ( .a(n_36082), .b(n_35850), .o(n_36215) );
in01s01 g745331 ( .a(n_36164), .o(n_36165) );
oa12s01 g745332 ( .a(n_35891), .b(FE_OCP_RBN3303_n_35539), .c(n_35800), .o(n_36164) );
in01s01 g745333 ( .a(n_36213), .o(n_36214) );
oa22s01 g745334 ( .a(n_36049), .b(n_35842), .c(FE_OCP_RBN3301_n_35539), .d(n_35476), .o(n_36213) );
in01s01 g745335 ( .a(n_35959), .o(n_35960) );
na03f04 TIMEBOOST_cell_8241 ( .a(n_37717), .b(TIMEBOOST_net_197), .c(n_37761), .o(n_37791) );
na02s01 g745337 ( .a(n_35929), .b(n_35841), .o(n_35930) );
in01s01 g745338 ( .a(n_36161), .o(n_36162) );
oa12s01 g745339 ( .a(n_35927), .b(FE_OCP_RBN3303_n_35539), .c(n_35931), .o(n_36161) );
in01s01 g745340 ( .a(n_36211), .o(n_36212) );
oa22s01 g745341 ( .a(n_36049), .b(n_35525), .c(FE_OCP_RBN3303_n_35539), .d(n_36022), .o(n_36211) );
oa22s01 g745342 ( .a(n_35956), .b(n_35583), .c(FE_OCP_RBN3301_n_35539), .d(n_35559), .o(n_36223) );
oa22s01 g745343 ( .a(n_35956), .b(n_35809), .c(FE_OCP_RBN3293_n_35539), .d(n_34671), .o(n_36225) );
oa22s01 g745344 ( .a(n_35956), .b(n_36111), .c(FE_OCP_RBN3293_n_35539), .d(n_35602), .o(n_36229) );
in01s01 g745345 ( .a(n_36113), .o(n_36114) );
ao12s01 g745346 ( .a(n_36055), .b(n_35956), .c(n_35633), .o(n_36113) );
in01s01 g745347 ( .a(n_36159), .o(n_36160) );
oa12s01 g745348 ( .a(n_35719), .b(FE_OCP_RBN3293_n_35539), .c(n_35678), .o(n_36159) );
in01s01 g745349 ( .a(n_36157), .o(n_36158) );
oa12s01 g745350 ( .a(n_35723), .b(FE_OCP_RBN3293_n_35539), .c(n_35653), .o(n_36157) );
oa12f08 g745351 ( .a(n_34148), .b(n_34226), .c(n_34114), .o(n_34275) );
in01s01 g745352 ( .a(n_36155), .o(n_36156) );
oa12s01 g745353 ( .a(n_35962), .b(FE_OCP_RBN3303_n_35539), .c(n_35884), .o(n_36155) );
in01s01 g745354 ( .a(n_34262), .o(n_34263) );
oa12s01 g745355 ( .a(n_34210), .b(n_34226), .c(n_34209), .o(n_34262) );
in01s01 g745356 ( .a(n_36209), .o(n_36210) );
no02s01 g745357 ( .a(n_36079), .b(n_36154), .o(n_36209) );
in01s02 g745358 ( .a(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n_40598) );
no02m02 g745360 ( .a(n_34487), .b(n_34511), .o(n_34539) );
na02s01 g745361 ( .a(n_34463), .b(n_34351), .o(n_34464) );
in01s01 g745362 ( .a(n_35805), .o(n_35764) );
no02s01 g745363 ( .a(FE_OCP_RBN3292_n_35539), .b(n_35258), .o(n_35805) );
no02s01 g745364 ( .a(FE_OCP_RBN3292_n_35539), .b(n_35720), .o(n_35937) );
in01s01 g745365 ( .a(n_35849), .o(n_35938) );
na02s01 g745366 ( .a(FE_OCP_RBN3292_n_35539), .b(n_35720), .o(n_35849) );
no02s01 g745367 ( .a(FE_OCP_RBN3301_n_35539), .b(n_35298), .o(n_36082) );
no02s01 g745368 ( .a(FE_OCP_RBN3299_n_35539), .b(n_35763), .o(n_35850) );
na02s01 g745369 ( .a(n_36049), .b(n_35391), .o(n_36122) );
in01s01 g745370 ( .a(n_35890), .o(n_35848) );
na02s01 g745371 ( .a(FE_OCP_RBN3300_n_35539), .b(n_35371), .o(n_35890) );
na02s01 g745372 ( .a(FE_OCP_RBN3300_n_35539), .b(n_35800), .o(n_35891) );
in01s01 g745373 ( .a(n_35799), .o(n_35888) );
na02s01 g745374 ( .a(FE_OCP_RBN3299_n_35539), .b(n_35388), .o(n_35799) );
in01s01 g745375 ( .a(n_35847), .o(n_35934) );
na02s01 g745376 ( .a(FE_OCP_RBN3300_n_35539), .b(n_35389), .o(n_35847) );
na02s01 g745377 ( .a(FE_OCP_RBN3300_n_35539), .b(n_35884), .o(n_35962) );
in01s01 g745378 ( .a(n_35929), .o(n_35883) );
na02s01 g745379 ( .a(FE_OCP_RBN3299_n_35539), .b(n_35845), .o(n_35929) );
in01s01 g745380 ( .a(n_35882), .o(n_35961) );
no02s01 g745381 ( .a(FE_OCP_RBN3299_n_35539), .b(n_35845), .o(n_35882) );
no02m08 TIMEBOOST_cell_2977 ( .a(TIMEBOOST_net_779), .b(FE_OCP_RBN7037_n_18982), .o(n_19107) );
in01s01 g745383 ( .a(n_35927), .o(n_35928) );
na02s01 g745384 ( .a(FE_OCP_RBN3300_n_35539), .b(n_35931), .o(n_35927) );
na02s01 g745385 ( .a(FE_OCP_RBN3299_n_35539), .b(n_35926), .o(n_36171) );
in01s01 g745386 ( .a(n_36080), .o(n_36081) );
no02s01 g745387 ( .a(n_36049), .b(n_35926), .o(n_36080) );
na02s01 g745388 ( .a(FE_OCP_RBN3300_n_35539), .b(n_36019), .o(n_36121) );
na02s01 g745389 ( .a(n_36049), .b(n_35629), .o(n_36117) );
na02m06 g745391 ( .a(n_34433), .b(n_34409), .o(n_34462) );
na02s01 g745392 ( .a(FE_OCP_RBN3299_n_35539), .b(n_35842), .o(n_35841) );
na02s04 g745393 ( .a(n_34568), .b(n_34627), .o(n_34747) );
ao12m04 g745394 ( .a(n_34490), .b(FE_OCP_RBN6668_n_34297), .c(n_34404), .o(n_34491) );
in01s01 g745395 ( .a(n_36050), .o(n_36119) );
no02s01 g745396 ( .a(FE_OCP_RBN3300_n_35539), .b(n_36019), .o(n_36050) );
in01s01 g745397 ( .a(n_35958), .o(n_36021) );
no02s01 g745398 ( .a(FE_OCP_RBN3299_n_35539), .b(n_35840), .o(n_35958) );
na02s01 g745399 ( .a(n_34653), .b(n_34590), .o(n_34675) );
na02s01 g745400 ( .a(n_34226), .b(n_34209), .o(n_34210) );
in01s01 g745401 ( .a(n_35561), .o(n_35562) );
na02m04 g745402 ( .a(n_35543), .b(n_35542), .o(n_35561) );
in01s01 g745403 ( .a(n_35932), .o(n_35880) );
na02s01 g745404 ( .a(FE_OCP_RBN3299_n_35539), .b(n_35840), .o(n_35932) );
no02s01 g745405 ( .a(n_36049), .b(n_35240), .o(n_36123) );
no02s01 g745406 ( .a(FE_OCP_RBN3292_n_35539), .b(n_35765), .o(n_36079) );
na02s01 g745407 ( .a(n_36049), .b(n_36111), .o(n_36112) );
in01s01 g745408 ( .a(n_35634), .o(n_35724) );
no02s01 g745409 ( .a(FE_OCP_RBN3295_n_35539), .b(n_35631), .o(n_35634) );
na02s02 g745410 ( .a(FE_OCP_RBN3290_n_35539), .b(n_35583), .o(n_35584) );
no02s01 TIMEBOOST_cell_6905 ( .a(FE_OCP_RBN5609_n_7730), .b(FE_OCP_RBN4136_n_7743), .o(TIMEBOOST_net_2211) );
no02m04 g745412 ( .a(n_35543), .b(n_35542), .o(n_35605) );
na02s01 g745413 ( .a(FE_OCP_RBN3292_n_35539), .b(n_35602), .o(n_35604) );
no02s01 g745414 ( .a(FE_OCP_RBN3290_n_35539), .b(n_35633), .o(n_36055) );
in01s01 g745415 ( .a(n_35679), .o(n_35654) );
na02s01 g745416 ( .a(FE_OCP_RBN3295_n_35539), .b(n_35631), .o(n_35679) );
in01s01 g745417 ( .a(n_35718), .o(n_35719) );
no02s01 g745418 ( .a(FE_OCP_RBN3295_n_35539), .b(n_34988), .o(n_35718) );
in01s01 g745420 ( .a(n_35630), .o(n_35722) );
no02s01 g745421 ( .a(FE_OCP_RBN3295_n_35539), .b(n_35629), .o(n_35630) );
na02s01 g745422 ( .a(FE_OCP_RBN3292_n_35539), .b(n_35653), .o(n_35723) );
na02s01 g745425 ( .a(n_35675), .b(FE_OCP_RBN3295_n_35539), .o(n_35717) );
in01s01 g745426 ( .a(n_35715), .o(n_35716) );
no02s01 g745427 ( .a(FE_OCP_RBN3295_n_35539), .b(n_35675), .o(n_35715) );
no02s01 g745428 ( .a(FE_OCP_RBN3290_n_35539), .b(n_35217), .o(n_36154) );
in01s01 g745429 ( .a(n_35839), .o(n_35996) );
no02s01 g745430 ( .a(FE_OCP_RBN3300_n_35539), .b(n_35392), .o(n_35839) );
na02s01 g745431 ( .a(FE_OCP_RBN3300_n_35539), .b(n_35526), .o(n_36018) );
in01s01 g745432 ( .a(n_35581), .o(n_35582) );
ao12s01 g745433 ( .a(n_34890), .b(n_35540), .c(n_34942), .o(n_35581) );
in01s01 g745434 ( .a(n_34326), .o(n_34386) );
oa12f08 g745435 ( .a(n_34198), .b(n_34298), .c(n_34247), .o(n_34326) );
oa12s01 g745436 ( .a(n_34274), .b(n_34298), .c(n_34273), .o(n_35469) );
in01s01 g745437 ( .a(n_35796), .o(n_35797) );
no02s01 g745438 ( .a(FE_OCP_RBN3290_n_35539), .b(n_35260), .o(n_35796) );
no02s01 g745439 ( .a(n_35541), .b(n_35524), .o(n_36118) );
na02s01 g745442 ( .a(FE_OCP_RBN3295_n_35539), .b(n_35189), .o(n_35795) );
no02s01 g745443 ( .a(FE_OCP_RBN3292_n_35539), .b(n_35108), .o(n_36126) );
na02m02 g745444 ( .a(FE_OCP_RBN5773_n_34375), .b(n_34450), .o(n_34489) );
na02s01 g745445 ( .a(n_35926), .b(n_35525), .o(n_35526) );
no02s01 g745446 ( .a(n_35511), .b(n_34964), .o(n_35524) );
no02s01 g745447 ( .a(n_35540), .b(n_34965), .o(n_35541) );
na02s01 g745448 ( .a(n_34298), .b(n_34273), .o(n_34274) );
na02f08 g745449 ( .a(FE_OCP_RBN5772_n_34375), .b(n_34307), .o(n_34437) );
no02s01 g745451 ( .a(n_34704), .b(n_34649), .o(n_34705) );
na02s06 g745452 ( .a(n_34412), .b(n_34356), .o(n_34413) );
in01s06 g745454 ( .a(n_34487), .o(n_34488) );
in01s02 g745455 ( .a(n_34459), .o(n_34487) );
in01s01 g745458 ( .a(n_34463), .o(n_34435) );
na02s06 g745459 ( .a(n_34349), .b(FE_OCP_RBN4191_n_34285), .o(n_34463) );
in01s01 g745460 ( .a(n_34433), .o(n_34434) );
na02m04 g745462 ( .a(n_34297), .b(n_34345), .o(n_34409) );
no02s06 g745463 ( .a(n_34325), .b(n_34315), .o(n_34384) );
na02m06 TIMEBOOST_cell_4018 ( .a(n_25704), .b(TIMEBOOST_net_1099), .o(n_25783) );
in01s01 g745465 ( .a(n_34653), .o(n_34654) );
no02s01 TIMEBOOST_cell_2874 ( .a(n_37920), .b(n_38021), .o(TIMEBOOST_net_728) );
ao12s01 g745467 ( .a(n_35510), .b(n_35509), .c(n_35508), .o(n_36019) );
oa12f08 g745468 ( .a(n_34067), .b(n_34167), .c(n_34095), .o(n_34226) );
oa12s01 g745469 ( .a(n_34154), .b(n_34167), .c(n_34153), .o(n_35594) );
in01s01 g745479 ( .a(FE_OCP_RBN3301_n_35539), .o(n_36049) );
in01s01 g745490 ( .a(FE_OCP_RBN3300_n_35539), .o(n_35956) );
in01s04 g745506 ( .a(n_35543), .o(n_35539) );
oa12m08 g745507 ( .a(n_34943), .b(n_35496), .c(n_34941), .o(n_35543) );
ao12s01 g745508 ( .a(n_34451), .b(n_34453), .c(n_44102), .o(n_34538) );
no02s06 g745509 ( .a(n_34357), .b(n_34318), .o(n_34412) );
no02s06 g745510 ( .a(n_34377), .b(n_34316), .o(n_34356) );
no02s06 g745511 ( .a(n_34354), .b(n_34353), .o(n_34355) );
na02s06 g745513 ( .a(n_34383), .b(n_34339), .o(n_34406) );
na02m02 g745515 ( .a(n_34486), .b(n_47255), .o(n_34511) );
na02s01 g745518 ( .a(n_34651), .b(n_34650), .o(n_34652) );
na02s01 g745519 ( .a(n_34650), .b(n_34648), .o(n_34649) );
na02s06 g745521 ( .a(n_34348), .b(n_34347), .o(n_34349) );
na02m04 g745523 ( .a(n_34344), .b(n_34343), .o(n_34345) );
in01s01 g745524 ( .a(n_34378), .o(n_34379) );
no02s01 g745525 ( .a(n_34353), .b(n_34324), .o(n_34378) );
na02s01 g745526 ( .a(n_34405), .b(n_34320), .o(n_34630) );
no02s01 g745527 ( .a(n_34377), .b(n_34319), .o(n_34709) );
no02s01 g745528 ( .a(n_34764), .b(n_34321), .o(n_34819) );
no02s06 g745529 ( .a(n_34324), .b(n_34323), .o(n_34325) );
no02s01 g745530 ( .a(n_34403), .b(n_34322), .o(n_34789) );
no02s01 g745531 ( .a(n_34816), .b(n_34846), .o(n_34896) );
na02s01 g745532 ( .a(n_34380), .b(n_34374), .o(n_34850) );
na02s01 TIMEBOOST_cell_2871 ( .a(n_28650), .b(TIMEBOOST_net_726), .o(TIMEBOOST_net_234) );
na02s03 g745534 ( .a(FE_OCP_RBN4918_n_33491), .b(n_34374), .o(n_34404) );
in01s01 g745535 ( .a(n_34562), .o(n_34563) );
na02s01 g745536 ( .a(n_34509), .b(n_34537), .o(n_34562) );
na02s01 g745537 ( .a(n_34486), .b(n_34506), .o(n_34507) );
no02s01 g745538 ( .a(n_34535), .b(n_34484), .o(n_34536) );
in01s01 g745539 ( .a(n_34624), .o(n_34625) );
no02m01 g745540 ( .a(n_34993), .b(n_34704), .o(n_34624) );
na02s06 TIMEBOOST_cell_5367 ( .a(TIMEBOOST_net_1631), .b(FE_RN_1128_0), .o(n_30914) );
in01s01 g745542 ( .a(n_35511), .o(n_35540) );
na02s01 g745543 ( .a(n_35496), .b(n_34914), .o(n_35511) );
no02s01 g745544 ( .a(n_34311), .b(n_34376), .o(n_34438) );
no02s01 g745545 ( .a(n_35509), .b(n_35508), .o(n_35510) );
na02s01 g745546 ( .a(n_34167), .b(n_34153), .o(n_34154) );
in01s01 g745549 ( .a(n_34762), .o(n_34763) );
ao12s01 g745550 ( .a(n_34354), .b(FE_OCPN4855_n_34369), .c(n_34323), .o(n_34762) );
ao12s01 g745551 ( .a(n_34357), .b(FE_OCPN4855_n_34369), .c(n_34294), .o(n_34783) );
oa12s01 g745552 ( .a(n_34317), .b(FE_OCP_RBN6673_n_34297), .c(n_34343), .o(n_34823) );
in01s01 g745553 ( .a(n_34533), .o(n_34534) );
na02s02 g745554 ( .a(n_34381), .b(n_34458), .o(n_34533) );
ao12s01 g745555 ( .a(n_34402), .b(FE_OCPN4855_n_34369), .c(n_33564), .o(n_34854) );
oa12s01 g745556 ( .a(n_34383), .b(FE_OCP_RBN6665_n_34297), .c(n_34313), .o(n_34929) );
in01s01 g745557 ( .a(n_34702), .o(n_34703) );
na02s02 g745558 ( .a(n_34650), .b(n_34621), .o(n_34702) );
in01s01 g745559 ( .a(n_34558), .o(n_34559) );
na02s01 g745560 ( .a(n_47255), .b(n_34454), .o(n_34558) );
in01s01 g745561 ( .a(n_34622), .o(n_34623) );
no02m06 TIMEBOOST_cell_4205 ( .a(n_32740), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_7_), .o(TIMEBOOST_net_1193) );
in01s01 g745563 ( .a(n_34745), .o(n_34746) );
na02s01 g745564 ( .a(n_34648), .b(n_34674), .o(n_34745) );
oa12s01 g745565 ( .a(n_35480), .b(n_35479), .c(n_35478), .o(n_35926) );
ao12f08 g745566 ( .a(n_34157), .b(n_34250), .c(n_34197), .o(n_34298) );
ao12s01 g745567 ( .a(n_34249), .b(n_34248), .c(n_34250), .o(n_35427) );
oa22s01 g745568 ( .a(FE_OCPN4855_n_34369), .b(n_33545), .c(FE_OCP_RBN6672_n_34297), .d(n_34347), .o(n_34847) );
in01s01 g745569 ( .a(n_34743), .o(n_34744) );
oa22s01 g745570 ( .a(FE_OCP_RBN6667_n_34297), .b(n_34039), .c(FE_OCP_RBN6673_n_34297), .d(FE_OCP_RBN5685_FE_RN_308_0), .o(n_34743) );
in01s01 g745571 ( .a(n_34351), .o(n_34322) );
na02s03 g745572 ( .a(n_34297), .b(n_33539), .o(n_34351) );
in01s01 g745573 ( .a(n_34348), .o(n_34321) );
na02s03 g745574 ( .a(n_34297), .b(FE_OCP_DRV_N6891_n_34296), .o(n_34348) );
in01s01 g745576 ( .a(n_34320), .o(n_34340) );
na02s04 g745577 ( .a(n_34291), .b(n_34293), .o(n_34320) );
in01s01 g745578 ( .a(n_34344), .o(n_34319) );
na02s06 g745579 ( .a(n_34291), .b(n_34292), .o(n_34344) );
no02s03 g745580 ( .a(n_34297), .b(n_34294), .o(n_34357) );
in01s01 g745581 ( .a(n_34318), .o(n_34405) );
no02s04 g745582 ( .a(n_34291), .b(n_34293), .o(n_34318) );
in01s01 g745583 ( .a(n_34316), .o(n_34317) );
no02s02 g745584 ( .a(n_34297), .b(n_33426), .o(n_34316) );
no02s06 g745585 ( .a(n_34297), .b(n_34292), .o(n_34377) );
no02s02 g745586 ( .a(n_34291), .b(n_34323), .o(n_34354) );
no02s03 g745587 ( .a(n_34291), .b(n_33222), .o(n_34353) );
no02s01 g745588 ( .a(FE_OCPN4855_n_34369), .b(FE_OCP_DRV_N6891_n_34296), .o(n_34764) );
in01s01 g745589 ( .a(n_34324), .o(n_34290) );
no02s02 g745590 ( .a(n_34261), .b(FE_OCP_DRV_N1894_n_33221), .o(n_34324) );
in01s01 g745591 ( .a(n_34460), .o(n_34403) );
na02s06 g745592 ( .a(FE_OCP_RBN6666_n_34297), .b(n_33540), .o(n_34460) );
in01s01 g745593 ( .a(n_34401), .o(n_34402) );
na02s06 g745594 ( .a(FE_OCP_RBN6666_n_34297), .b(n_34350), .o(n_34401) );
in01s01 g745595 ( .a(n_34339), .o(n_34846) );
na02s06 g745596 ( .a(n_34315), .b(n_34314), .o(n_34339) );
in01s01 g745598 ( .a(n_34374), .o(n_34852) );
na02s02 g745599 ( .a(n_34297), .b(FE_OCP_RBN4916_n_33503), .o(n_34374) );
na02s06 g745600 ( .a(FE_OCP_RBN6665_n_34297), .b(n_34313), .o(n_34383) );
in01s01 g745602 ( .a(n_34380), .o(n_34372) );
na02s08 g745603 ( .a(n_34285), .b(n_33542), .o(n_34380) );
na02s01 g745604 ( .a(FE_OCP_RBN6668_n_34297), .b(FE_OCP_RBN4917_n_33491), .o(n_34458) );
na02s06 g745605 ( .a(n_34315), .b(FE_OCP_RBN4918_n_33491), .o(n_34381) );
in01s01 g745606 ( .a(n_34816), .o(n_34817) );
no02s01 g745607 ( .a(FE_OCP_RBN6665_n_34297), .b(n_34314), .o(n_34816) );
in01s01 g745608 ( .a(n_34704), .o(n_34651) );
no02s06 g745609 ( .a(FE_OCP_RBN6668_n_34297), .b(FE_OCP_RBN2553_n_33697), .o(n_34704) );
in01m01 g745610 ( .a(n_34532), .o(n_34993) );
na02s06 g745611 ( .a(FE_OCP_RBN6668_n_34297), .b(FE_OCP_RBN2553_n_33697), .o(n_34532) );
na02s02 g745613 ( .a(FE_OCP_RBN6668_n_34297), .b(FE_OCP_RBN2551_n_33664), .o(n_34509) );
in01s01 g745614 ( .a(n_34486), .o(n_34535) );
na02m01 g745615 ( .a(FE_OCP_RBN6671_n_34297), .b(n_33594), .o(n_34486) );
no02s01 g745618 ( .a(FE_OCP_RBN6668_n_34297), .b(n_33691), .o(n_34565) );
in01s01 g745619 ( .a(n_34564), .o(n_34537) );
no02s06 g745620 ( .a(FE_OCP_RBN2551_n_33664), .b(FE_OCP_RBN6668_n_34297), .o(n_34564) );
na02s01 g745621 ( .a(FE_OCP_RBN6668_n_34297), .b(n_33735), .o(n_34621) );
na02s01 g745622 ( .a(FE_OCP_RBN6672_n_34297), .b(FE_OCP_RBN2570_n_33735), .o(n_34650) );
na02s01 g745623 ( .a(FE_OCP_RBN6668_n_34297), .b(n_33581), .o(n_34506) );
no02s01 g745624 ( .a(FE_OCP_RBN6671_n_34297), .b(n_33594), .o(n_34484) );
na02s01 g745625 ( .a(FE_OCP_RBN6668_n_34297), .b(FE_OCP_RBN2544_n_33584), .o(n_34454) );
no02f08 TIMEBOOST_cell_4204 ( .a(n_6959), .b(TIMEBOOST_net_1192), .o(n_7031) );
na02s01 g745627 ( .a(FE_OCP_RBN6667_n_34297), .b(n_33964), .o(n_34674) );
na02s01 g745628 ( .a(FE_OCP_RBN6672_n_34297), .b(n_34590), .o(n_34648) );
na02s01 g745629 ( .a(n_35462), .b(n_34938), .o(n_35509) );
in01s01 g745630 ( .a(n_34310), .o(n_34311) );
na02s08 g745631 ( .a(n_34289), .b(FE_OCPN1370_n_34288), .o(n_34310) );
no02s01 g745632 ( .a(n_34248), .b(n_34250), .o(n_34249) );
no02m06 g745633 ( .a(n_34289), .b(FE_OCPN1370_n_34288), .o(n_34376) );
na02s01 g745634 ( .a(n_35479), .b(n_35478), .o(n_35480) );
no02s01 TIMEBOOST_cell_4561 ( .a(FE_OFN5083_n_36750), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_1371) );
na02f06 g745636 ( .a(n_35461), .b(n_35159), .o(n_35496) );
in01s01 g745638 ( .a(n_34398), .o(n_34399) );
na02s02 g745639 ( .a(FE_OCP_RBN6666_n_34297), .b(n_33546), .o(n_34398) );
na02s01 g745640 ( .a(FE_OCP_RBN6668_n_34297), .b(n_33662), .o(n_34627) );
no02s01 g745641 ( .a(n_35477), .b(n_35463), .o(n_35931) );
in01s01 g745642 ( .a(n_35525), .o(n_36022) );
oa22s01 g745643 ( .a(n_35451), .b(n_34962), .c(n_35452), .d(n_34963), .o(n_35525) );
ao12f08 g745644 ( .a(n_33985), .b(n_34121), .c(n_34041), .o(n_34167) );
in01s01 g745645 ( .a(FE_OCPUNCON7067_n_34151), .o(n_34152) );
oa12s01 g745646 ( .a(n_34102), .b(n_34101), .c(n_34121), .o(n_34151) );
na02s01 g745647 ( .a(n_34452), .b(n_34427), .o(n_34453) );
no02s01 g745648 ( .a(n_34272), .b(n_34246), .o(n_34385) );
no02s01 g745649 ( .a(n_35453), .b(n_34842), .o(n_35463) );
na02s01 g745650 ( .a(n_34121), .b(n_34101), .o(n_34102) );
na02s06 g745652 ( .a(n_34221), .b(n_34219), .o(n_34287) );
in01s01 g745653 ( .a(n_34450), .o(n_34451) );
no02s02 g745654 ( .a(n_34366), .b(FE_OCP_RBN5756_n_34307), .o(n_34450) );
no02s01 g745655 ( .a(n_34841), .b(n_35454), .o(n_35477) );
in01s01 g745656 ( .a(n_35461), .o(n_35462) );
no02f06 g745657 ( .a(n_35432), .b(n_34885), .o(n_35461) );
in01s04 g745687 ( .a(n_34297), .o(n_34285) );
in01m10 g745688 ( .a(n_34261), .o(n_34297) );
in01s06 g745689 ( .a(n_34291), .o(n_34315) );
in01s06 g745690 ( .a(n_34261), .o(n_34291) );
no02s01 g745693 ( .a(n_34430), .b(n_34367), .o(n_34481) );
oa12s01 g745694 ( .a(n_35436), .b(n_35435), .c(n_35434), .o(n_35840) );
na02s02 TIMEBOOST_cell_2854 ( .a(n_37561), .b(n_37057), .o(TIMEBOOST_net_718) );
oa12f06 g745696 ( .a(n_34109), .b(n_34191), .c(n_34134), .o(n_34250) );
oa12s01 g745697 ( .a(n_34190), .b(n_34189), .c(n_34191), .o(n_35415) );
oa12s01 g745698 ( .a(n_34843), .b(n_35433), .c(n_34805), .o(n_35479) );
no02f06 TIMEBOOST_cell_2853 ( .a(n_37374), .b(TIMEBOOST_net_717), .o(n_37451) );
no02m08 g745700 ( .a(n_34181), .b(n_34224), .o(n_34225) );
na02s01 g745701 ( .a(n_35435), .b(n_35434), .o(n_35436) );
in01s01 g745702 ( .a(n_35453), .o(n_35454) );
na02s01 g745703 ( .a(n_35433), .b(n_34865), .o(n_35453) );
no02s01 g745704 ( .a(n_34199), .b(n_34247), .o(n_34273) );
na02s01 g745705 ( .a(n_34189), .b(n_34191), .o(n_34190) );
in01s01 g745706 ( .a(n_34245), .o(n_34246) );
na02f06 g745707 ( .a(n_34223), .b(FE_OCPUNCON7061_n_34222), .o(n_34245) );
no02m06 g745708 ( .a(n_34223), .b(FE_OCPUNCON7061_n_34222), .o(n_34272) );
na02f04 TIMEBOOST_cell_2882 ( .a(FE_OCP_RBN5027_n_18515), .b(FE_RN_288_0), .o(TIMEBOOST_net_732) );
in01s01 g745712 ( .a(n_34367), .o(n_34368) );
na02m01 g745713 ( .a(n_34284), .b(n_34338), .o(n_34367) );
na02f04 g745714 ( .a(n_34120), .b(FE_OCP_RBN2687_n_44100), .o(n_34150) );
na02m01 TIMEBOOST_cell_4239 ( .a(n_12496), .b(n_12461), .o(TIMEBOOST_net_1210) );
no02s02 TIMEBOOST_cell_2083 ( .a(n_19565), .b(n_19641), .o(TIMEBOOST_net_656) );
na02m02 g745720 ( .a(n_34259), .b(n_44102), .o(n_34307) );
na02s03 TIMEBOOST_cell_2081 ( .a(n_34978), .b(n_30633), .o(TIMEBOOST_net_655) );
oa12f08 g745722 ( .a(n_33966), .b(n_34069), .c(n_34013), .o(n_34121) );
in01s01 g745723 ( .a(n_35842), .o(n_35476) );
na02s01 g745724 ( .a(n_35431), .b(n_35417), .o(n_35842) );
oa12s01 g745725 ( .a(n_34054), .b(n_34053), .c(n_34069), .o(n_35500) );
in01s01 g745726 ( .a(n_35451), .o(n_35452) );
in01s01 g745727 ( .a(n_35432), .o(n_35451) );
ao12f04 g745728 ( .a(n_34866), .b(n_35390), .c(n_34888), .o(n_35432) );
na02s01 g745730 ( .a(n_34429), .b(n_34428), .o(n_34430) );
in01s01 g745731 ( .a(n_34396), .o(n_34397) );
no02s01 g745732 ( .a(n_34365), .b(n_34364), .o(n_34396) );
na02m08 TIMEBOOST_cell_2881 ( .a(n_7470), .b(TIMEBOOST_net_731), .o(n_7534) );
na02f04 g745734 ( .a(n_34130), .b(n_34117), .o(n_34131) );
no02s06 g745735 ( .a(n_34162), .b(n_34522), .o(n_34186) );
na02s01 g745736 ( .a(n_34219), .b(n_34184), .o(n_34220) );
na02f10 g745737 ( .a(n_34177), .b(n_34203), .o(n_34204) );
no02s01 g745739 ( .a(n_34266), .b(n_34283), .o(n_34284) );
no02s01 g745740 ( .a(n_34149), .b(n_34100), .o(n_34264) );
na02s01 g745741 ( .a(n_34479), .b(n_34328), .o(n_34569) );
na02f02 g745742 ( .a(n_34119), .b(n_34118), .o(n_34120) );
na02s01 g745743 ( .a(n_34116), .b(n_34187), .o(n_34466) );
no02s01 g745745 ( .a(n_34478), .b(n_34522), .o(n_34600) );
no02s01 g745746 ( .a(n_34161), .b(n_34179), .o(n_34603) );
no02s01 g745747 ( .a(n_34618), .b(n_34201), .o(n_34682) );
na02f08 TIMEBOOST_cell_4238 ( .a(TIMEBOOST_net_1209), .b(n_37560), .o(n_37667) );
na02s01 TIMEBOOST_cell_8718 ( .a(n_7177), .b(n_7343), .o(TIMEBOOST_net_2846) );
na02s01 g745750 ( .a(n_34241), .b(n_34196), .o(n_34685) );
in01s01 g745751 ( .a(n_34281), .o(n_34282) );
no02s03 g745752 ( .a(n_47254), .b(n_34256), .o(n_34281) );
na02s02 g745754 ( .a(FE_OCP_RBN1813_n_33846), .b(n_34238), .o(n_34259) );
in01s01 g745755 ( .a(n_34362), .o(n_34363) );
na02s06 g745756 ( .a(n_34338), .b(FE_OCP_RBN5743_n_34278), .o(n_34362) );
na02m04 TIMEBOOST_cell_2087 ( .a(n_35075), .b(FE_OCPN6281_n_30612), .o(TIMEBOOST_net_658) );
na02s01 g745758 ( .a(n_35407), .b(n_34806), .o(n_35431) );
in01s01 g745759 ( .a(n_34198), .o(n_34199) );
na02m06 g745760 ( .a(n_34183), .b(FE_OCPUNCON4498_n_34182), .o(n_34198) );
na02s01 g745761 ( .a(n_34197), .b(n_34158), .o(n_34248) );
no02m06 g745762 ( .a(n_34183), .b(FE_OCPUNCON4498_n_34182), .o(n_34247) );
na02s01 g745763 ( .a(n_35406), .b(n_34807), .o(n_35417) );
na02s01 g745764 ( .a(n_34115), .b(n_34148), .o(n_34209) );
na02s01 g745765 ( .a(n_34069), .b(n_34053), .o(n_34054) );
in01m04 g745766 ( .a(n_34180), .o(n_34181) );
no02m08 g745767 ( .a(n_34164), .b(n_34036), .o(n_34180) );
oa12s01 g745768 ( .a(n_34130), .b(FE_OCP_RBN5713_n_44102), .c(FE_OCPN1699_n_34118), .o(n_34519) );
ao12s01 g745769 ( .a(n_34414), .b(n_44102), .c(n_33500), .o(n_34596) );
ao12s01 g745770 ( .a(n_34145), .b(n_44102), .c(n_34127), .o(n_34657) );
oa12s01 g745771 ( .a(n_34163), .b(FE_OCP_RBN5713_n_44102), .c(n_33613), .o(n_34575) );
ao12s01 g745772 ( .a(n_34178), .b(n_44102), .c(n_33632), .o(n_34662) );
in01s01 g745773 ( .a(n_34304), .o(n_34305) );
na02m01 g745774 ( .a(n_34242), .b(n_34258), .o(n_34304) );
in01s01 g745775 ( .a(n_34394), .o(n_34395) );
na02s06 TIMEBOOST_cell_2822 ( .a(n_7010), .b(n_7011), .o(TIMEBOOST_net_702) );
in01s01 g745777 ( .a(n_34447), .o(n_34448) );
oa12m01 g745778 ( .a(n_34428), .b(FE_OCP_RBN5714_n_44102), .c(n_34427), .o(n_34447) );
oa12s01 g745779 ( .a(n_35374), .b(n_35373), .c(n_35372), .o(n_35845) );
ao12s01 g745780 ( .a(n_34845), .b(n_35408), .c(n_34775), .o(n_35435) );
ao12s01 g745781 ( .a(n_34813), .b(n_35408), .c(n_34804), .o(n_35433) );
ao12s01 g745782 ( .a(n_34141), .b(n_34140), .c(n_34139), .o(n_35367) );
ao12f06 g745783 ( .a(n_34111), .b(n_34094), .c(n_34076), .o(n_34191) );
na02s02 TIMEBOOST_cell_8598 ( .a(n_26077), .b(n_23398), .o(TIMEBOOST_net_2786) );
oa22s01 g745785 ( .a(n_44102), .b(n_34200), .c(FE_OCP_RBN5712_n_44102), .d(n_33686), .o(n_34716) );
in01s01 g745786 ( .a(n_34445), .o(n_34446) );
oa22s01 g745787 ( .a(FE_OCP_RBN5715_n_44102), .b(n_34206), .c(n_44102), .d(n_34224), .o(n_34445) );
in01s01 g745788 ( .a(n_34334), .o(n_34335) );
oa22m01 g745789 ( .a(n_44102), .b(n_33895), .c(FE_OCP_RBN5714_n_44102), .d(FE_OCP_RBN1813_n_33846), .o(n_34334) );
in01s01 g745790 ( .a(n_34423), .o(n_34424) );
oa22m01 g745791 ( .a(FE_OCP_RBN5714_n_44102), .b(FE_OCP_RBN5629_n_33976), .c(n_44102), .d(n_33976), .o(n_34423) );
in01s01 g745792 ( .a(n_34303), .o(n_34365) );
na02s01 g745793 ( .a(n_44102), .b(n_33954), .o(n_34303) );
no02s01 g745794 ( .a(n_44102), .b(n_33954), .o(n_34364) );
na02m02 g745795 ( .a(n_34124), .b(n_34427), .o(n_34126) );
no02s01 TIMEBOOST_cell_8591 ( .a(TIMEBOOST_net_2782), .b(n_15491), .o(n_15635) );
in01s01 g745797 ( .a(n_34119), .o(n_34100) );
na02f01 g745798 ( .a(n_34066), .b(FE_OCPN1234_n_33341), .o(n_34119) );
in01s01 g745799 ( .a(n_34117), .o(n_34149) );
na02m01 g745801 ( .a(n_44100), .b(FE_OCPN1699_n_34118), .o(n_34130) );
in01s01 g745802 ( .a(n_34479), .o(n_34480) );
na02s01 g745803 ( .a(n_44102), .b(n_33499), .o(n_34479) );
na02s06 g745804 ( .a(FE_OCP_RBN2688_n_44100), .b(n_34122), .o(n_34328) );
in01s01 g745805 ( .a(n_34146), .o(n_34414) );
na02m02 g745806 ( .a(n_44100), .b(n_34123), .o(n_34146) );
in01s01 g745807 ( .a(n_34128), .o(n_34116) );
no02s03 g745808 ( .a(n_44100), .b(n_34098), .o(n_34128) );
na02s03 g745809 ( .a(n_44100), .b(n_34098), .o(n_34187) );
in01s01 g745810 ( .a(n_34144), .o(n_34145) );
na02m02 g745811 ( .a(n_44100), .b(n_33517), .o(n_34144) );
no02s06 g745812 ( .a(n_44102), .b(n_34143), .o(n_34522) );
in01s01 g745813 ( .a(n_34477), .o(n_34478) );
na02s01 g745814 ( .a(n_44102), .b(n_34143), .o(n_34477) );
in01s01 g745815 ( .a(n_34162), .o(n_34163) );
in01s01 g745817 ( .a(n_34203), .o(n_34179) );
in01s01 g745819 ( .a(n_34184), .o(n_34161) );
na02s02 g745820 ( .a(FE_OCP_RBN2687_n_44100), .b(n_33604), .o(n_34184) );
in01s01 g745821 ( .a(n_34177), .o(n_34178) );
na02f10 g745822 ( .a(FE_OCP_RBN5713_n_44102), .b(n_34160), .o(n_34177) );
no02s01 g745823 ( .a(n_44102), .b(n_33708), .o(n_34618) );
in01s01 g745824 ( .a(n_34201), .o(n_34176) );
no02s02 g745825 ( .a(FE_OCP_RBN2689_n_44100), .b(FE_OCP_DRV_N1414_n_33673), .o(n_34201) );
in01m01 g745827 ( .a(n_34196), .o(n_34687) );
na02f01 g745828 ( .a(n_44102), .b(n_33706), .o(n_34196) );
in01s01 g745830 ( .a(n_34241), .o(n_34239) );
na02s04 g745831 ( .a(FE_OCP_RBN5714_n_44102), .b(n_33844), .o(n_34241) );
na02s03 g745832 ( .a(FE_OCP_RBN5714_n_44102), .b(FE_OCP_RBN1812_n_33750), .o(n_34242) );
na02s01 g745833 ( .a(n_44102), .b(n_33750), .o(n_34258) );
in01m01 g745838 ( .a(n_34238), .o(n_34256) );
na02s10 g745839 ( .a(n_44102), .b(FE_OCP_RBN4912_n_33803), .o(n_34238) );
na02m02 g745840 ( .a(FE_OCP_RBN5714_n_44102), .b(n_33897), .o(n_34338) );
no02s01 g745842 ( .a(FE_OCP_RBN5714_n_44102), .b(n_33897), .o(n_34278) );
na02f08 TIMEBOOST_cell_2821 ( .a(n_37251), .b(TIMEBOOST_net_701), .o(FE_RN_636_0) );
no02s01 g745844 ( .a(n_44102), .b(n_34003), .o(n_34283) );
na02s01 g745845 ( .a(FE_OCP_RBN5714_n_44102), .b(n_34427), .o(n_34428) );
na02s01 g745846 ( .a(n_35373), .b(n_35372), .o(n_35374) );
no02s01 g745847 ( .a(n_34140), .b(n_34139), .o(n_34141) );
na02m04 g745848 ( .a(n_34138), .b(FE_OCPUNCON1747_n_34137), .o(n_34197) );
in01s01 g745849 ( .a(n_34157), .o(n_34158) );
no02m04 g745850 ( .a(n_34138), .b(FE_OCPUNCON1747_n_34137), .o(n_34157) );
na02s06 g745851 ( .a(n_34097), .b(FE_OCP_DRV_N6907_n_34096), .o(n_34148) );
in01s01 g745852 ( .a(n_34114), .o(n_34115) );
no02s01 g745854 ( .a(n_34068), .b(n_34095), .o(n_34153) );
no02s01 g745855 ( .a(n_35391), .b(n_35335), .o(n_35392) );
in01s01 g745856 ( .a(n_35406), .o(n_35407) );
in01s01 g745857 ( .a(n_35390), .o(n_35406) );
na02f04 g745858 ( .a(n_35354), .b(n_34844), .o(n_35390) );
oa12s01 g745860 ( .a(FE_OCP_RBN5714_n_44102), .b(FE_OCP_RBN5629_n_33976), .c(FE_OCP_RBN2637_n_33954), .o(n_34429) );
in01s01 g745861 ( .a(n_34135), .o(n_34136) );
ao12s02 g745862 ( .a(n_44100), .b(n_34123), .c(n_34122), .o(n_34135) );
in01s01 g745863 ( .a(n_34219), .o(n_34193) );
na02s03 g745864 ( .a(n_44102), .b(n_33614), .o(n_34219) );
in01s01 g745866 ( .a(n_34266), .o(n_34267) );
no02s01 g745867 ( .a(n_44102), .b(n_33939), .o(n_34266) );
ao12s01 g745868 ( .a(n_35357), .b(n_35356), .c(n_35355), .o(n_35884) );
ao12f08 g745870 ( .a(n_33923), .b(n_34017), .c(n_33963), .o(n_34069) );
ao12s01 g745871 ( .a(n_34016), .b(n_34015), .c(n_34017), .o(n_35482) );
in01s01 g745872 ( .a(n_35388), .o(n_35389) );
oa12s01 g745873 ( .a(n_35339), .b(n_35338), .c(n_35337), .o(n_35388) );
na02s01 g745874 ( .a(n_35338), .b(n_35337), .o(n_35339) );
no02s01 g745875 ( .a(n_35356), .b(n_35355), .o(n_35357) );
no02s01 g745876 ( .a(n_34134), .b(n_34110), .o(n_34189) );
in01s01 g745878 ( .a(n_34067), .o(n_34068) );
na02s06 g745879 ( .a(n_34052), .b(FE_OCP_DRV_N1416_n_34051), .o(n_34067) );
na02s01 g745880 ( .a(n_33986), .b(n_34041), .o(n_34101) );
no02s01 g745881 ( .a(n_34015), .b(n_34017), .o(n_34016) );
in01s01 g745882 ( .a(n_35354), .o(n_35408) );
na02f04 g745883 ( .a(n_35336), .b(n_34800), .o(n_35354) );
in01s02 g745884 ( .a(n_34124), .o(n_34113) );
oa12s01 g745886 ( .a(n_34089), .b(n_34088), .c(n_34087), .o(n_35292) );
in01s01 g745887 ( .a(n_34094), .o(n_34139) );
oa12f06 g745888 ( .a(n_34063), .b(n_34048), .c(n_34030), .o(n_34094) );
na02m04 g745889 ( .a(n_34079), .b(n_34065), .o(n_34138) );
no02m06 g745890 ( .a(n_34040), .b(n_34014), .o(n_34097) );
no02s01 g745891 ( .a(n_35336), .b(n_34759), .o(n_35373) );
in01s01 g745892 ( .a(n_35391), .o(n_35371) );
oa12s01 g745893 ( .a(n_35322), .b(n_35321), .c(n_35320), .o(n_35391) );
ao12f08 g745932 ( .a(n_33928), .b(FE_OCP_RBN6637_n_33983), .c(FE_OCP_RBN5684_FE_RN_308_0), .o(n_34066) );
na02m02 g745933 ( .a(n_34064), .b(FE_OCP_RBN2638_n_33954), .o(n_34065) );
na02m04 g745934 ( .a(n_34049), .b(n_33954), .o(n_34079) );
no02s02 g745935 ( .a(n_33983), .b(FE_OCP_RBN5685_FE_RN_308_0), .o(n_34014) );
no02m04 g745936 ( .a(FE_OCP_RBN6636_n_33983), .b(n_34039), .o(n_34040) );
no02f08 g745937 ( .a(FE_OCP_RBN5686_FE_RN_308_0), .b(n_34037), .o(n_33928) );
na02s01 g745938 ( .a(n_35321), .b(n_35320), .o(n_35322) );
no02s01 g745939 ( .a(n_34077), .b(n_34111), .o(n_34140) );
in01s01 g745940 ( .a(n_34109), .o(n_34110) );
na02s04 g745941 ( .a(n_34086), .b(n_34085), .o(n_34109) );
na02s01 g745942 ( .a(n_34088), .b(n_34087), .o(n_34089) );
no02f04 g745943 ( .a(n_34086), .b(n_34085), .o(n_34134) );
na02m06 g745944 ( .a(n_33969), .b(FE_OCPN1739_n_33968), .o(n_34041) );
in01s01 g745945 ( .a(n_33985), .o(n_33986) );
no02m06 g745946 ( .a(n_33969), .b(FE_OCPN1739_n_33968), .o(n_33985) );
no02s01 g745947 ( .a(n_35278), .b(n_34777), .o(n_35356) );
no02s01 g745948 ( .a(n_33967), .b(n_34013), .o(n_34053) );
no02f04 g745949 ( .a(n_35277), .b(n_34808), .o(n_35336) );
in01m04 g745950 ( .a(n_34083), .o(n_34084) );
in01s04 g745951 ( .a(n_34078), .o(n_34083) );
no02m08 g745952 ( .a(n_34064), .b(n_33961), .o(n_34078) );
oa12s01 g745953 ( .a(n_34699), .b(n_35299), .c(n_35070), .o(n_35338) );
ao12s01 g745954 ( .a(n_34062), .b(n_34061), .c(n_34060), .o(n_35315) );
na02f06 g745956 ( .a(n_33965), .b(n_33944), .o(n_34052) );
oa12s01 g745957 ( .a(n_33927), .b(n_33926), .c(n_33925), .o(n_35420) );
in01s01 g745958 ( .a(n_35335), .o(n_35800) );
oa12s01 g745959 ( .a(n_35280), .b(n_35299), .c(n_35279), .o(n_35335) );
na02s01 g745960 ( .a(n_35299), .b(n_35279), .o(n_35280) );
na02s01 g745961 ( .a(n_34031), .b(n_34063), .o(n_34088) );
no02s01 g745962 ( .a(n_34061), .b(n_34060), .o(n_34062) );
no02m04 g745963 ( .a(n_34059), .b(FE_OCPUNCON7059_n_34058), .o(n_34111) );
in01s01 g745964 ( .a(n_34076), .o(n_34077) );
na02m04 g745965 ( .a(n_34059), .b(FE_OCPUNCON7059_n_34058), .o(n_34076) );
no02m08 g745967 ( .a(n_33946), .b(FE_OCP_DRV_N6889_n_33945), .o(n_34013) );
in01s01 g745968 ( .a(n_33966), .o(n_33967) );
na02m04 g745970 ( .a(n_33906), .b(n_34590), .o(n_33944) );
na02s02 g745971 ( .a(n_33962), .b(n_33964), .o(n_33965) );
na02s01 g745972 ( .a(n_33963), .b(n_33924), .o(n_34015) );
na02s01 g745973 ( .a(n_33925), .b(n_33926), .o(n_33927) );
in01s01 g745974 ( .a(n_35277), .o(n_35278) );
na02f04 g745975 ( .a(n_35241), .b(n_34734), .o(n_35277) );
in01m02 g745976 ( .a(n_34064), .o(n_34049) );
na02m08 g745977 ( .a(FE_OCP_RBN5643_n_33977), .b(n_33981), .o(n_34064) );
ao12s01 g745981 ( .a(n_35247), .b(n_35246), .c(n_35245), .o(n_35720) );
in01s01 g745982 ( .a(n_35763), .o(n_35298) );
oa12s01 g745983 ( .a(n_35244), .b(n_35243), .c(n_35242), .o(n_35763) );
ao12s01 g745984 ( .a(n_34635), .b(n_35218), .c(n_34697), .o(n_35321) );
na02m08 TIMEBOOST_cell_5561 ( .a(TIMEBOOST_net_1728), .b(n_31381), .o(n_31488) );
in01s01 g745986 ( .a(n_34048), .o(n_34087) );
ao12f06 g745987 ( .a(n_34032), .b(n_33940), .c(n_33978), .o(n_34048) );
in01s02 g745988 ( .a(FE_OCP_RBN5685_FE_RN_308_0), .o(n_34039) );
no02m04 g745992 ( .a(n_33787), .b(n_33213), .o(n_33810) );
na02s06 g745994 ( .a(n_33956), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_33981) );
no02s02 g745997 ( .a(n_34427), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_34036) );
no02m02 g745998 ( .a(n_33977), .b(n_33975), .o(n_34011) );
na02s01 TIMEBOOST_cell_5530 ( .a(n_6112), .b(n_5897), .o(TIMEBOOST_net_1713) );
no02s01 g746001 ( .a(n_35246), .b(n_35245), .o(n_35247) );
na02s01 g746002 ( .a(n_35243), .b(n_35242), .o(n_35244) );
no02s01 g746003 ( .a(n_33979), .b(n_34032), .o(n_34061) );
in01s01 g746004 ( .a(n_34030), .o(n_34031) );
no02f04 g746005 ( .a(n_34010), .b(FE_OCP_DRV_N1886_n_34009), .o(n_34030) );
na02s04 g746006 ( .a(n_34010), .b(FE_OCP_DRV_N1886_n_34009), .o(n_34063) );
in01s01 g746007 ( .a(n_33923), .o(n_33924) );
no02f06 g746008 ( .a(n_33908), .b(FE_OCPN1912_n_33907), .o(n_33923) );
na02f06 g746009 ( .a(n_33908), .b(FE_OCPN1912_n_33907), .o(n_33963) );
na02s01 g746010 ( .a(n_33880), .b(n_33881), .o(n_33926) );
no02s01 g746011 ( .a(n_35259), .b(n_35258), .o(n_35260) );
in01s01 g746014 ( .a(n_34055), .o(n_34056) );
ao12s01 g746015 ( .a(n_34008), .b(n_34007), .c(n_34006), .o(n_34055) );
na02m04 TIMEBOOST_cell_5529 ( .a(TIMEBOOST_net_1712), .b(n_6023), .o(n_6105) );
oa12f06 g746017 ( .a(n_33778), .b(n_33877), .c(n_33829), .o(n_33925) );
na02f04 TIMEBOOST_cell_7769 ( .a(TIMEBOOST_net_2515), .b(n_9841), .o(n_10040) );
ao12s01 g746019 ( .a(n_33879), .b(n_33878), .c(n_33877), .o(n_35382) );
in01s01 g746020 ( .a(n_35241), .o(n_35299) );
oa12f04 g746021 ( .a(n_34742), .b(n_35191), .c(n_34695), .o(n_35241) );
na02m06 g746023 ( .a(n_33719), .b(n_33646), .o(n_33787) );
no02m06 g746024 ( .a(n_33942), .b(n_34037), .o(n_33961) );
in01s01 g746026 ( .a(n_35243), .o(n_35218) );
na02s01 g746027 ( .a(n_35191), .b(n_34669), .o(n_35243) );
na02f08 TIMEBOOST_cell_4154 ( .a(TIMEBOOST_net_1167), .b(n_17091), .o(n_17250) );
no02s01 g746029 ( .a(n_34007), .b(n_34006), .o(n_34008) );
na02s02 g746030 ( .a(n_33957), .b(n_33872), .o(n_33960) );
no02f04 g746031 ( .a(n_33959), .b(n_33958), .o(n_34032) );
in01s01 g746032 ( .a(n_33978), .o(n_33979) );
na02f04 g746033 ( .a(n_33959), .b(n_33958), .o(n_33978) );
na02m06 g746035 ( .a(n_33781), .b(n_32986), .o(n_33881) );
na02s04 g746036 ( .a(n_33833), .b(FE_OCP_RBN2552_n_33697), .o(n_33835) );
no03s02 TIMEBOOST_cell_8269 ( .a(FE_OCP_RBN5877_n_3848), .b(n_3848), .c(n_4218), .o(TIMEBOOST_net_1589) );
no02s01 g746038 ( .a(n_33877), .b(n_33878), .o(n_33879) );
na02s02 g746041 ( .a(n_33833), .b(n_33733), .o(n_33834) );
in01s01 g746042 ( .a(n_35258), .o(n_35240) );
ao12s01 g746043 ( .a(n_35164), .b(n_35163), .c(n_35162), .o(n_35258) );
in01s01 g746044 ( .a(n_35259), .o(n_35804) );
ao12s01 g746045 ( .a(n_35161), .b(n_35190), .c(n_35160), .o(n_35259) );
oa12s01 g746046 ( .a(n_34644), .b(n_35190), .c(n_35069), .o(n_35246) );
in01s02 g746047 ( .a(n_34224), .o(n_34206) );
na02m10 g746048 ( .a(n_33955), .b(n_33974), .o(n_34224) );
in01s02 g746049 ( .a(FE_OCP_RBN5627_n_33976), .o(n_34005) );
in01s02 g746058 ( .a(n_34427), .o(n_34026) );
no02m04 TIMEBOOST_cell_3894 ( .a(TIMEBOOST_net_1037), .b(n_29144), .o(TIMEBOOST_net_739) );
no02f06 g746061 ( .a(n_33784), .b(n_33809), .o(n_33908) );
in01s01 g746062 ( .a(FE_OCPUNCON7063_n_33904), .o(n_33905) );
ao12s01 g746063 ( .a(n_33832), .b(n_33831), .c(n_33830), .o(n_33904) );
in01s02 g746068 ( .a(n_33975), .o(n_34003) );
in01m02 g746069 ( .a(n_33956), .o(n_33975) );
na02m06 g746070 ( .a(n_33903), .b(n_33876), .o(n_33956) );
na02s01 TIMEBOOST_cell_8578 ( .a(n_42392), .b(n_42483), .o(TIMEBOOST_net_2776) );
no02s01 TIMEBOOST_cell_4405 ( .a(n_23353), .b(n_23398), .o(TIMEBOOST_net_1293) );
no02s03 g746074 ( .a(n_33898), .b(n_33402), .o(n_33922) );
no02f02 g746076 ( .a(n_33873), .b(n_33846), .o(n_33901) );
na02f06 g746079 ( .a(n_33735), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_33785) );
na02s04 TIMEBOOST_cell_5495 ( .a(TIMEBOOST_net_1695), .b(n_16482), .o(n_16575) );
na02s08 g746082 ( .a(n_33938), .b(n_33447), .o(n_33974) );
na02s06 g746083 ( .a(n_33937), .b(n_33448), .o(n_33955) );
no02s01 g746084 ( .a(n_35163), .b(n_35162), .o(n_35164) );
in01s04 g746088 ( .a(n_33942), .o(n_33954) );
no03s02 TIMEBOOST_cell_8736 ( .a(n_13280), .b(n_13351), .c(n_13352), .o(TIMEBOOST_net_2855) );
no02s01 g746090 ( .a(n_33831), .b(n_33830), .o(n_33832) );
no02s01 g746091 ( .a(n_33829), .b(n_33779), .o(n_33878) );
no02s01 g746092 ( .a(n_35190), .b(n_35160), .o(n_35161) );
na02f04 g746093 ( .a(n_35109), .b(n_34634), .o(n_35191) );
oa12m06 g746094 ( .a(FE_OCP_RBN4009_n_32860), .b(n_33677), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_), .o(n_33719) );
ao12s01 g746102 ( .a(n_33919), .b(n_33918), .c(FE_OCPN5228_n_33917), .o(n_34007) );
na02f04 g746103 ( .a(n_33874), .b(n_33850), .o(n_33959) );
in01s01 g746104 ( .a(n_33940), .o(n_34060) );
in01s01 g746106 ( .a(n_33964), .o(n_34590) );
na02s06 g746107 ( .a(n_33718), .b(n_33737), .o(n_33964) );
in01m02 g746108 ( .a(n_33780), .o(n_33781) );
ao12f08 g746110 ( .a(n_33731), .b(n_33777), .c(n_33830), .o(n_33877) );
in01s01 g746111 ( .a(FE_OCPN1350_n_35312), .o(n_35310) );
oa12s01 g746112 ( .a(n_33776), .b(n_33775), .c(FE_OCP_RBN4635_n_33589), .o(n_35312) );
oa12s01 g746113 ( .a(n_35112), .b(n_35111), .c(n_35110), .o(n_35675) );
in01s01 g746114 ( .a(n_35765), .o(n_35217) );
ao12s01 g746115 ( .a(n_35128), .b(n_35127), .c(n_35126), .o(n_35765) );
no02m04 TIMEBOOST_cell_1856 ( .a(TIMEBOOST_net_542), .b(FE_OCP_RBN6129_n_21804), .o(n_21927) );
no02s06 g746117 ( .a(n_33847), .b(n_33855), .o(n_33875) );
na02s03 g746118 ( .a(n_33827), .b(n_33870), .o(n_33900) );
na03s01 TIMEBOOST_cell_7329 ( .a(TIMEBOOST_net_2182), .b(n_27400), .c(FE_RN_611_0), .o(FE_RN_612_0) );
na02s02 g746121 ( .a(n_33677), .b(n_33178), .o(n_33737) );
na02s04 g746122 ( .a(n_33695), .b(n_33179), .o(n_33718) );
na02s02 TIMEBOOST_cell_7935 ( .a(TIMEBOOST_net_2598), .b(n_5351), .o(n_5493) );
oa12s04 g746125 ( .a(n_33450), .b(n_33772), .c(n_33379), .o(n_33898) );
no02s01 g746126 ( .a(n_33918), .b(FE_OCPN5228_n_33917), .o(n_33919) );
na02f02 g746127 ( .a(n_33826), .b(n_33803), .o(n_33874) );
na02f02 g746128 ( .a(FE_OCP_RBN6569_n_33803), .b(n_33849), .o(n_33850) );
in01s01 g746129 ( .a(n_33778), .o(n_33779) );
na02f04 g746130 ( .a(n_33757), .b(n_33756), .o(n_33778) );
no02m04 g746131 ( .a(n_33757), .b(FE_OCP_DRV_N1888_n_33756), .o(n_33829) );
na02s01 g746132 ( .a(n_33732), .b(n_33777), .o(n_33831) );
na02s01 g746133 ( .a(n_33775), .b(FE_OCP_RBN4635_n_33589), .o(n_33776) );
no02s01 g746134 ( .a(n_33896), .b(FE_OCP_RBN6568_n_33803), .o(n_33939) );
na02s01 g746135 ( .a(n_35653), .b(n_35125), .o(n_35189) );
na02s01 g746136 ( .a(n_35111), .b(n_35110), .o(n_35112) );
no02s01 g746137 ( .a(n_35127), .b(n_35126), .o(n_35128) );
no02f02 TIMEBOOST_cell_1859 ( .a(n_10582), .b(FE_OFN756_n_44464), .o(TIMEBOOST_net_544) );
no02f08 TIMEBOOST_cell_4122 ( .a(TIMEBOOST_net_1151), .b(n_25914), .o(n_26098) );
in01s04 g746141 ( .a(n_33937), .o(n_33938) );
no02s01 TIMEBOOST_cell_7057 ( .a(n_20124), .b(FE_OCP_RBN4337_n_20242), .o(TIMEBOOST_net_2287) );
ao12s01 g746143 ( .a(n_34670), .b(n_35089), .c(n_34638), .o(n_35163) );
in01s02 g746146 ( .a(n_33872), .o(n_33897) );
in01s01 g746152 ( .a(n_35109), .o(n_35190) );
oa12f04 g746153 ( .a(n_34701), .b(n_35045), .c(n_34639), .o(n_35109) );
na02s04 g746155 ( .a(n_33807), .b(n_33305), .o(n_33852) );
na03f08 TIMEBOOST_cell_5731 ( .a(n_18343), .b(n_18301), .c(TIMEBOOST_net_1453), .o(n_18435) );
in01m01 g746158 ( .a(n_33717), .o(n_33733) );
no02m08 g746160 ( .a(n_33697), .b(n_34037), .o(n_33717) );
in01s02 g746162 ( .a(n_33677), .o(n_33695) );
no02s01 TIMEBOOST_cell_1878 ( .a(TIMEBOOST_net_553), .b(n_36531), .o(n_36245) );
in01s01 g746167 ( .a(n_33731), .o(n_33732) );
no02s01 g746169 ( .a(n_35089), .b(n_34700), .o(n_35127) );
in01s02 g746171 ( .a(n_33827), .o(n_33847) );
na02s06 g746172 ( .a(n_33772), .b(n_33408), .o(n_33827) );
in01f01 g746173 ( .a(n_33849), .o(n_33826) );
ao12f06 g746174 ( .a(n_34037), .b(n_33752), .c(n_33728), .o(n_33849) );
no02m08 TIMEBOOST_cell_5673 ( .a(TIMEBOOST_net_1784), .b(n_26759), .o(n_26851) );
no02f04 TIMEBOOST_cell_1860 ( .a(TIMEBOOST_net_544), .b(n_10587), .o(n_10647) );
in01s01 g746181 ( .a(n_33868), .o(n_33918) );
oa12f08 g746184 ( .a(n_33590), .b(n_33591), .c(n_33711), .o(n_33830) );
ao12s01 g746185 ( .a(n_33690), .b(n_33711), .c(n_33689), .o(n_33775) );
ao12s01 g746186 ( .a(n_35088), .b(n_35087), .c(n_35086), .o(n_35653) );
ao12s01 g746187 ( .a(n_34615), .b(n_35087), .c(n_35041), .o(n_35111) );
in01s01 g746191 ( .a(n_33895), .o(n_33896) );
in01s01 g746192 ( .a(FE_OCP_RBN1813_n_33846), .o(n_33895) );
in01m02 g746194 ( .a(n_33825), .o(n_33846) );
in01m02 g746199 ( .a(n_33675), .o(n_33691) );
no02s01 TIMEBOOST_cell_1876 ( .a(TIMEBOOST_net_552), .b(n_44277), .o(n_22201) );
na02f06 g746203 ( .a(n_33157), .b(n_33622), .o(n_33648) );
in01m02 g746204 ( .a(n_33807), .o(n_33773) );
no02m08 g746205 ( .a(n_33753), .b(n_33340), .o(n_33807) );
no02m10 g746206 ( .a(n_33664), .b(n_34037), .o(n_33782) );
no02s03 g746207 ( .a(n_33664), .b(n_34037), .o(n_33663) );
in01s04 g746211 ( .a(n_33804), .o(n_33805) );
in01s04 g746212 ( .a(n_33772), .o(n_33804) );
na02s06 g746213 ( .a(n_33753), .b(n_33324), .o(n_33772) );
no02s01 g746216 ( .a(n_33711), .b(n_33689), .o(n_33690) );
in01s01 g746217 ( .a(n_35045), .o(n_35089) );
na02f04 g746218 ( .a(n_35087), .b(n_34581), .o(n_35045) );
no02s01 g746219 ( .a(n_35087), .b(n_35086), .o(n_35088) );
in01f01 g746224 ( .a(n_33771), .o(n_33803) );
oa22s01 g746226 ( .a(n_33844), .b(n_33768), .c(n_33706), .d(n_32574), .o(n_35106) );
na02s02 TIMEBOOST_cell_5500 ( .a(n_5024), .b(n_4442), .o(TIMEBOOST_net_1698) );
in01s01 g746230 ( .a(n_35629), .o(n_35125) );
oa12s01 g746231 ( .a(n_35073), .b(n_35072), .c(n_35071), .o(n_35629) );
no02m08 g746232 ( .a(n_33707), .b(n_33264), .o(n_33753) );
na02m08 g746233 ( .a(n_33549), .b(FE_OCP_DRV_N3496_n_33156), .o(n_33622) );
in01s01 g746235 ( .a(n_33752), .o(n_33769) );
na02m08 g746236 ( .a(n_33706), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_33752) );
in01s01 g746237 ( .a(n_33820), .o(n_34006) );
na02s02 g746238 ( .a(n_33706), .b(n_33768), .o(n_33820) );
in01m03 g746239 ( .a(n_33595), .o(n_33596) );
in01s01 TIMEBOOST_cell_8894 ( .a(n_1211), .o(TIMEBOOST_net_2938) );
na02s02 g746241 ( .a(n_33568), .b(n_33218), .o(n_33646) );
no02f04 g746242 ( .a(n_33642), .b(n_33594), .o(n_33621) );
na02s01 TIMEBOOST_cell_5939 ( .a(FE_RN_2557_0), .b(FE_RN_2556_0), .o(TIMEBOOST_net_1821) );
na02s01 g746244 ( .a(n_33594), .b(n_33584), .o(n_33662) );
na02s01 g746246 ( .a(n_35072), .b(n_35071), .o(n_35073) );
in01m02 g746247 ( .a(n_33729), .o(n_33730) );
na02m04 g746248 ( .a(n_33707), .b(n_33329), .o(n_33729) );
na02m04 g746249 ( .a(n_33644), .b(n_33620), .o(n_33660) );
no02m02 g746250 ( .a(n_33642), .b(n_47249), .o(n_33643) );
na03m08 TIMEBOOST_cell_8268 ( .a(n_24936), .b(n_24959), .c(n_24912), .o(n_25065) );
no02f08 g746254 ( .a(n_33618), .b(n_33592), .o(n_33711) );
ao12m04 g746255 ( .a(n_34610), .b(n_34944), .c(n_34616), .o(n_35087) );
in01m02 g746259 ( .a(n_33728), .o(n_33750) );
in01f02 g746262 ( .a(n_33687), .o(n_33688) );
no02f04 g746263 ( .a(n_33674), .b(n_33328), .o(n_33687) );
no02s01 TIMEBOOST_cell_8590 ( .a(FE_OCP_RBN6802_n_15156), .b(n_15518), .o(TIMEBOOST_net_2782) );
no02s06 g746265 ( .a(n_33529), .b(n_33080), .o(n_33550) );
na02f06 TIMEBOOST_cell_8795 ( .a(TIMEBOOST_net_2884), .b(n_24320), .o(n_24347) );
in01m02 g746267 ( .a(n_47249), .o(n_33620) );
no02s04 g746270 ( .a(n_44815), .b(FE_OCP_RBN4049_n_33491), .o(n_33592) );
no02f06 g746271 ( .a(n_44814), .b(FE_OCP_RBN4917_n_33491), .o(n_33618) );
no02s06 g746273 ( .a(n_33589), .b(n_33588), .o(n_33591) );
na02s06 g746274 ( .a(n_33589), .b(FE_OCPN1634_n_33588), .o(n_33590) );
na02s01 g746275 ( .a(n_34944), .b(n_34550), .o(n_35072) );
in01m04 g746280 ( .a(n_33549), .o(n_33568) );
ao12m08 g746281 ( .a(n_33206), .b(n_33476), .c(n_33105), .o(n_33549) );
na02f06 g746282 ( .a(n_33547), .b(n_33527), .o(n_33642) );
no02m06 g746283 ( .a(n_44815), .b(n_33528), .o(n_33644) );
in01s01 g746284 ( .a(n_33640), .o(n_35268) );
ao22s01 g746285 ( .a(FE_OCP_RBN4916_n_33503), .b(FE_OCPN1701_n_33544), .c(FE_OCP_RBN4915_n_33503), .d(n_32728), .o(n_33640) );
in01s01 g746287 ( .a(n_33706), .o(n_33844) );
na02m08 g746291 ( .a(n_33636), .b(n_33657), .o(n_33706) );
in01f04 g746296 ( .a(n_33567), .o(n_33584) );
in01s01 g746298 ( .a(n_34200), .o(n_33686) );
oa12s01 g746299 ( .a(n_33639), .b(n_33638), .c(n_33637), .o(FE_RN_2852_0) );
in01s01 g746300 ( .a(n_35678), .o(n_34988) );
ao12s01 g746301 ( .a(n_34917), .b(n_34916), .c(n_34915), .o(n_35678) );
no02f08 g746302 ( .a(n_33635), .b(n_33233), .o(n_33674) );
in01s04 g746303 ( .a(n_33529), .o(n_33530) );
in01m06 g746304 ( .a(n_33508), .o(n_33529) );
oa12m08 g746305 ( .a(n_33205), .b(n_33475), .c(n_33474), .o(n_33508) );
na02s01 g746306 ( .a(n_33638), .b(n_33637), .o(n_33639) );
no04f06 TIMEBOOST_cell_7299 ( .a(n_26058), .b(n_25994), .c(n_25972), .d(n_26057), .o(n_26249) );
in01s02 g746309 ( .a(n_33527), .o(n_33528) );
na02m06 g746310 ( .a(n_33491), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_33527) );
na02f06 g746314 ( .a(n_33503), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_33547) );
in01f02 g746315 ( .a(n_33655), .o(n_33656) );
na02s01 g746317 ( .a(n_33545), .b(n_34296), .o(n_33546) );
no02s06 g746319 ( .a(FE_OCP_RBN4915_n_33503), .b(FE_OCPN1701_n_33544), .o(n_33589) );
na02s01 g746320 ( .a(n_33613), .b(n_33534), .o(n_33614) );
no02s01 g746321 ( .a(n_34916), .b(n_34915), .o(n_34917) );
in01s01 g746322 ( .a(n_33583), .o(n_34313) );
oa12s01 g746323 ( .a(n_33526), .b(n_33525), .c(n_33524), .o(n_33583) );
in01s01 g746324 ( .a(n_34350), .o(n_33564) );
ao12s02 g746325 ( .a(n_33507), .b(n_33506), .c(n_33505), .o(n_34350) );
in01s02 g746331 ( .a(n_33594), .o(n_33581) );
no02s08 g746332 ( .a(n_33494), .b(n_33504), .o(n_33594) );
in01s01 g746333 ( .a(n_34160), .o(n_33632) );
ao12s03 g746334 ( .a(n_33562), .b(n_33561), .c(n_33560), .o(n_34160) );
in01s01 g746335 ( .a(FE_OCP_DRV_N1414_n_33673), .o(n_33708) );
ao12s01 g746336 ( .a(n_33608), .b(n_33607), .c(n_33606), .o(n_33673) );
ao12m06 g746337 ( .a(n_34867), .b(n_34868), .c(n_34545), .o(n_34944) );
oa12s01 g746338 ( .a(n_35044), .b(n_35043), .c(n_35042), .o(n_35631) );
na02s01 g746339 ( .a(n_33525), .b(n_33524), .o(n_33526) );
na02f08 g746340 ( .a(n_33558), .b(n_33198), .o(n_33635) );
no02s01 g746341 ( .a(n_33506), .b(n_33505), .o(n_33507) );
no02m08 g746342 ( .a(n_33475), .b(n_33474), .o(n_33476) );
na02m04 TIMEBOOST_cell_8851 ( .a(TIMEBOOST_net_2912), .b(n_10136), .o(n_10309) );
no02s01 g746345 ( .a(n_33561), .b(n_33560), .o(n_33562) );
no02s01 g746347 ( .a(n_33607), .b(n_33606), .o(n_33608) );
no02s01 g746348 ( .a(n_35633), .b(n_36111), .o(n_35108) );
na02s01 g746349 ( .a(n_35043), .b(n_35042), .o(n_35044) );
no02s01 g746350 ( .a(n_34868), .b(n_34867), .o(n_34916) );
na02m06 g746352 ( .a(n_33475), .b(n_33164), .o(n_33492) );
ao12s01 g746353 ( .a(n_33235), .b(n_33559), .c(n_33200), .o(n_33638) );
in01s01 g746355 ( .a(FE_OCP_RBN4916_n_33503), .o(n_33542) );
in01s01 g746359 ( .a(n_33541), .o(n_34314) );
oa12s01 g746360 ( .a(n_33490), .b(n_33489), .c(n_33488), .o(n_33541) );
in01s01 g746361 ( .a(n_33539), .o(n_33540) );
oa12s01 g746362 ( .a(n_33487), .b(n_33486), .c(n_33485), .o(n_33539) );
in01s01 g746363 ( .a(n_33545), .o(n_34347) );
oa12s01 g746364 ( .a(n_33472), .b(n_33471), .c(n_33470), .o(n_33545) );
na02m04 g746369 ( .a(n_33412), .b(n_33434), .o(n_33491) );
ao12s01 g746371 ( .a(n_33521), .b(n_33520), .c(n_33519), .o(n_33613) );
oa12s01 g746373 ( .a(n_33537), .b(n_33536), .c(n_33535), .o(n_33604) );
na02s02 TIMEBOOST_cell_6826 ( .a(TIMEBOOST_net_2170), .b(n_6338), .o(n_6465) );
na02s01 g746375 ( .a(n_33471), .b(n_33470), .o(n_33472) );
no02f06 TIMEBOOST_cell_3367 ( .a(TIMEBOOST_net_974), .b(n_44809), .o(n_36730) );
no02s01 g746379 ( .a(n_33520), .b(n_33519), .o(n_33521) );
na02s01 g746380 ( .a(n_33536), .b(n_33535), .o(n_33537) );
no02s01 g746381 ( .a(n_33559), .b(n_33219), .o(n_33607) );
na02s01 g746382 ( .a(n_33489), .b(n_33488), .o(n_33490) );
in01m02 g746383 ( .a(n_33558), .o(n_33610) );
no02f08 g746384 ( .a(n_33518), .b(n_33201), .o(n_33558) );
na02s01 g746385 ( .a(n_33486), .b(n_33485), .o(n_33487) );
no02s01 g746386 ( .a(n_34779), .b(n_34911), .o(n_35043) );
no02f06 g746387 ( .a(n_34778), .b(n_34815), .o(n_34868) );
ao12s01 g746388 ( .a(n_33220), .b(n_33501), .c(n_33152), .o(n_33561) );
ao12s01 g746390 ( .a(n_32947), .b(n_33458), .c(n_33021), .o(n_33506) );
oa12s01 g746391 ( .a(n_35021), .b(n_35020), .c(n_35019), .o(n_35633) );
no02s02 TIMEBOOST_cell_1866 ( .a(TIMEBOOST_net_547), .b(n_39977), .o(n_40081) );
no02s01 g746393 ( .a(n_33410), .b(n_33459), .o(n_33489) );
no02s01 g746394 ( .a(n_33458), .b(n_32999), .o(n_33486) );
no02m10 g746398 ( .a(n_33388), .b(n_32995), .o(n_33411) );
no02s01 g746399 ( .a(n_33501), .b(n_33203), .o(n_33536) );
in01s01 g746400 ( .a(n_33518), .o(n_33559) );
oa12s01 g746402 ( .a(n_33289), .b(n_33429), .c(n_33246), .o(n_33471) );
na02s01 TIMEBOOST_cell_3141 ( .a(TIMEBOOST_net_861), .b(n_35799), .o(n_35939) );
oa12s01 g746404 ( .a(n_33057), .b(n_33484), .c(n_33449), .o(n_33520) );
in01s01 g746405 ( .a(n_34778), .o(n_34779) );
na02f04 g746406 ( .a(n_35020), .b(n_34760), .o(n_34778) );
na02s01 g746407 ( .a(n_35020), .b(n_35019), .o(n_35021) );
in01f02 g746408 ( .a(n_33427), .o(n_33428) );
ao12f06 g746409 ( .a(n_33083), .b(n_33331), .c(n_33067), .o(n_33427) );
oa22s01 g746410 ( .a(n_33429), .b(n_33304), .c(n_33331), .d(n_33303), .o(n_34296) );
in01s01 g746411 ( .a(n_33534), .o(n_34143) );
ao12s01 g746412 ( .a(n_33483), .b(n_33484), .c(n_33482), .o(n_33534) );
in01s01 g746413 ( .a(n_33409), .o(n_33410) );
na02s01 g746414 ( .a(n_33331), .b(n_33038), .o(n_33409) );
no02s01 g746416 ( .a(n_33429), .b(n_32935), .o(n_33458) );
no02s01 g746417 ( .a(n_33484), .b(n_33482), .o(n_33483) );
oa12s02 g746419 ( .a(n_33352), .b(n_33351), .c(n_33350), .o(n_34292) );
in01s01 g746420 ( .a(n_34123), .o(n_33500) );
ao12s01 g746421 ( .a(n_33457), .b(n_33456), .c(n_33455), .o(n_34123) );
ao12s01 g746422 ( .a(n_33425), .b(n_33424), .c(n_33423), .o(n_34098) );
in01s01 g746423 ( .a(n_34127), .o(n_33517) );
oa12s01 g746424 ( .a(n_33469), .b(n_33468), .c(n_33467), .o(n_34127) );
oa12f04 g746425 ( .a(n_34617), .b(n_34646), .c(n_34473), .o(n_35020) );
oa22s01 g746427 ( .a(n_33308), .b(n_33262), .c(n_33307), .d(n_33263), .o(FE_RN_2733_0) );
in01s01 g746428 ( .a(n_33426), .o(n_34343) );
oa22s01 g746429 ( .a(n_33346), .b(n_33302), .c(n_33347), .d(n_33301), .o(n_33426) );
na02s01 g746430 ( .a(n_33351), .b(n_33350), .o(n_33352) );
no02s01 g746431 ( .a(n_33456), .b(n_33455), .o(n_33457) );
na02s01 g746432 ( .a(n_33468), .b(n_33467), .o(n_33469) );
no02s01 g746433 ( .a(n_33424), .b(n_33423), .o(n_33425) );
no02s02 g746434 ( .a(n_34892), .b(n_34913), .o(n_34943) );
in01s01 g746437 ( .a(n_33331), .o(n_33429) );
in01s01 g746442 ( .a(n_36111), .o(n_35602) );
oa12s01 g746443 ( .a(n_35018), .b(n_35017), .c(n_35016), .o(n_36111) );
no02s06 TIMEBOOST_cell_1807 ( .a(FE_RN_1310_0), .b(FE_RN_1311_0), .o(TIMEBOOST_net_518) );
no02s01 g746445 ( .a(n_33382), .b(n_33380), .o(n_33424) );
in01s01 g746448 ( .a(n_33307), .o(n_33308) );
ao12s01 g746449 ( .a(n_33252), .b(n_33291), .c(n_33210), .o(n_33307) );
in01s01 g746450 ( .a(n_33346), .o(n_33347) );
no02s04 TIMEBOOST_cell_1721 ( .a(n_20372), .b(n_19245), .o(TIMEBOOST_net_475) );
ao12s01 g746452 ( .a(n_33401), .b(FE_OCP_RBN7021_n_33330), .c(n_33036), .o(n_33456) );
no02s01 g746453 ( .a(n_33381), .b(n_33190), .o(n_33468) );
no02f04 g746454 ( .a(n_35017), .b(n_34645), .o(n_34646) );
na02s01 g746455 ( .a(n_35017), .b(n_35016), .o(n_35018) );
oa22s01 g746456 ( .a(n_33291), .b(n_33265), .c(n_33255), .d(n_33266), .o(n_34293) );
ao12s01 g746457 ( .a(n_33345), .b(n_33344), .c(n_33343), .o(n_34118) );
in01s01 g746458 ( .a(n_34122), .o(n_33499) );
ao12s02 g746459 ( .a(n_33454), .b(FE_OCP_RBN7021_n_33330), .c(n_33452), .o(n_34122) );
ao12s01 g746460 ( .a(n_34666), .b(n_34942), .c(n_34891), .o(n_34892) );
no02s01 TIMEBOOST_cell_1831 ( .a(n_31770), .b(n_31871), .o(TIMEBOOST_net_530) );
no02s01 g746462 ( .a(n_33344), .b(n_33343), .o(n_33345) );
no02f08 g746463 ( .a(n_33330), .b(n_33143), .o(n_33382) );
na02s01 g746464 ( .a(n_34844), .b(n_34776), .o(n_34845) );
in01s01 g746465 ( .a(n_34964), .o(n_34965) );
na02s01 g746466 ( .a(n_34942), .b(n_44262), .o(n_34964) );
no02s01 g746467 ( .a(FE_OCP_RBN7021_n_33330), .b(n_33452), .o(n_33454) );
no02m04 TIMEBOOST_cell_1695 ( .a(n_20076), .b(FE_OCPN1316_n_20265), .o(TIMEBOOST_net_462) );
na02f04 g746469 ( .a(n_34553), .b(n_34498), .o(n_35017) );
na02s04 g746470 ( .a(n_34554), .b(n_34645), .o(n_34617) );
na02s02 g746471 ( .a(n_34940), .b(n_44262), .o(n_34941) );
no02m06 TIMEBOOST_cell_1715 ( .a(n_38953), .b(n_44925), .o(TIMEBOOST_net_472) );
in01s01 g746473 ( .a(n_35187), .o(n_35188) );
oa12s01 g746474 ( .a(n_34940), .b(n_34891), .c(n_34666), .o(n_35187) );
in01s01 g746475 ( .a(n_35809), .o(n_34671) );
na02s02 g746476 ( .a(n_34552), .b(n_34587), .o(n_35809) );
oa22s02 g746477 ( .a(n_33223), .b(n_33261), .c(n_33224), .d(n_33260), .o(n_34323) );
na02s01 g746478 ( .a(n_34721), .b(n_34740), .o(n_34759) );
no02s01 g746479 ( .a(n_34812), .b(n_34809), .o(n_34843) );
na02s01 g746480 ( .a(n_34642), .b(n_34640), .o(n_34670) );
na02s01 g746481 ( .a(n_34814), .b(n_34810), .o(n_34942) );
na02s01 g746482 ( .a(n_34865), .b(n_34811), .o(n_34866) );
in01s01 g746483 ( .a(n_34844), .o(n_34813) );
no02s01 g746484 ( .a(n_34741), .b(n_34777), .o(n_34844) );
no02s01 g746485 ( .a(n_34668), .b(n_34698), .o(n_34742) );
in01m02 g746486 ( .a(n_34553), .o(n_34554) );
na02f04 g746487 ( .a(n_34529), .b(n_34499), .o(n_34553) );
no02s02 g746488 ( .a(n_34700), .b(n_34641), .o(n_34701) );
na02s01 g746489 ( .a(n_34891), .b(n_34666), .o(n_34940) );
no02s01 g746491 ( .a(n_34814), .b(n_34810), .o(n_34890) );
na02s01 g746492 ( .a(n_34529), .b(n_34525), .o(n_34552) );
na02s01 g746493 ( .a(n_34500), .b(n_34526), .o(n_34587) );
in01s01 g746494 ( .a(n_33291), .o(n_33255) );
in01s01 g746495 ( .a(n_33273), .o(n_33291) );
ao12f08 g746496 ( .a(FE_OCPN3552_n_33225), .b(n_33207), .c(n_32923), .o(n_33273) );
oa12s01 g746497 ( .a(n_33079), .b(n_33306), .c(n_33032), .o(n_33344) );
ao12f08 g746499 ( .a(n_33082), .b(n_33306), .c(n_33106), .o(n_33330) );
oa22s01 g746501 ( .a(n_33306), .b(n_33101), .c(n_33272), .d(n_33100), .o(n_33341) );
in01s01 g746502 ( .a(n_35559), .o(n_35583) );
ao12s01 g746503 ( .a(n_34528), .b(n_34527), .c(n_35542), .o(n_35559) );
in01s01 g746504 ( .a(n_33223), .o(n_33224) );
na02s01 g746505 ( .a(n_33207), .b(n_32918), .o(n_33223) );
no02s01 g746506 ( .a(n_34527), .b(n_35542), .o(n_34528) );
in01s01 g746507 ( .a(FE_OCP_DRV_N1894_n_33221), .o(n_33222) );
ao12s01 g746508 ( .a(n_33167), .b(n_33168), .c(n_33166), .o(n_33221) );
oa12s01 g746509 ( .a(n_35159), .b(n_34666), .c(n_34889), .o(n_35508) );
in01s01 g746510 ( .a(n_34913), .o(n_34914) );
ao12s01 g746511 ( .a(n_34666), .b(n_34938), .c(n_34889), .o(n_34913) );
oa12s01 g746512 ( .a(n_34421), .b(n_34420), .c(n_34419), .o(n_34814) );
ao12s01 g746513 ( .a(n_34443), .b(n_34442), .c(n_34441), .o(n_34891) );
in01s01 g746514 ( .a(n_34812), .o(n_34865) );
ao12s01 g746515 ( .a(n_34666), .b(n_34776), .c(n_34738), .o(n_34812) );
oa12s01 g746516 ( .a(n_34810), .b(n_34809), .c(n_34299), .o(n_34811) );
no02s01 g746517 ( .a(n_34803), .b(n_34840), .o(n_34888) );
in01s01 g746518 ( .a(n_34777), .o(n_34721) );
ao12s01 g746519 ( .a(n_34666), .b(n_34699), .c(n_34733), .o(n_34777) );
ao12s01 g746520 ( .a(n_34666), .b(n_34740), .c(n_34739), .o(n_34741) );
ao12s01 g746521 ( .a(n_34473), .b(n_34697), .c(n_34696), .o(n_34698) );
in01s01 g746522 ( .a(n_34668), .o(n_34669) );
ao12s01 g746523 ( .a(n_34473), .b(n_34644), .c(n_34643), .o(n_34668) );
in01s01 g746524 ( .a(n_34529), .o(n_34500) );
oa12m04 g746525 ( .a(n_34417), .b(n_34475), .c(n_35542), .o(n_34529) );
na02s02 g746526 ( .a(n_34551), .b(FE_OCP_RBN6728_n_34388), .o(n_34616) );
in01s01 g746527 ( .a(n_34642), .o(n_34700) );
oa12s01 g746528 ( .a(FE_OCP_RBN6728_n_34388), .b(n_34615), .c(n_34614), .o(n_34642) );
ao12s01 g746529 ( .a(n_34473), .b(n_34640), .c(n_34582), .o(n_34641) );
na02s06 g746531 ( .a(n_33450), .b(n_33377), .o(n_33451) );
no02s01 g746532 ( .a(n_33168), .b(n_33166), .o(n_33167) );
no02s01 g746533 ( .a(n_35070), .b(n_34637), .o(n_35279) );
no02s01 g746534 ( .a(n_34808), .b(n_34692), .o(n_35355) );
in01s01 g746535 ( .a(n_34806), .o(n_34807) );
na02s01 g746536 ( .a(n_34775), .b(n_34776), .o(n_34806) );
no02s01 g746537 ( .a(n_35069), .b(n_34586), .o(n_35160) );
no02s01 g746538 ( .a(n_34475), .b(n_34418), .o(n_34527) );
no02s01 g746539 ( .a(n_34546), .b(n_34496), .o(n_34915) );
in01s01 g746540 ( .a(n_34841), .o(n_34842) );
no02s01 g746541 ( .a(n_34805), .b(n_34809), .o(n_34841) );
in01s01 g746542 ( .a(n_34525), .o(n_34526) );
na02s01 g746543 ( .a(n_34499), .b(n_34498), .o(n_34525) );
no02s01 g746544 ( .a(n_34608), .b(n_34544), .o(n_35126) );
in01s01 g746545 ( .a(n_34962), .o(n_34963) );
na02s01 g746546 ( .a(n_34886), .b(n_34938), .o(n_34962) );
na02s01 g746547 ( .a(n_34693), .b(n_34697), .o(n_35242) );
na02s01 g746548 ( .a(n_34420), .b(n_34419), .o(n_34421) );
no02s01 g746549 ( .a(n_34442), .b(n_34441), .o(n_34443) );
na02s01 g746550 ( .a(n_34889), .b(n_34666), .o(n_35159) );
in01s01 g746551 ( .a(n_34803), .o(n_34804) );
na02s01 g746552 ( .a(n_34757), .b(n_34775), .o(n_34803) );
na02s01 g746553 ( .a(n_34839), .b(n_34756), .o(n_34840) );
na02s01 g746554 ( .a(n_34694), .b(n_34693), .o(n_34695) );
na02s01 g746555 ( .a(n_34550), .b(n_34585), .o(n_34551) );
na02s01 g746556 ( .a(n_34606), .b(n_34638), .o(n_34639) );
na02s01 g746557 ( .a(n_35041), .b(n_34549), .o(n_35086) );
na02s01 g746558 ( .a(n_34912), .b(n_34760), .o(n_35019) );
in01s01 g746559 ( .a(n_33306), .o(n_33272) );
oa12f08 g746560 ( .a(n_33052), .b(n_33254), .c(n_33012), .o(n_33306) );
ao12s01 g746561 ( .a(n_34607), .b(n_34810), .c(n_33865), .o(n_35162) );
oa22s01 g746562 ( .a(n_34810), .b(n_34080), .c(n_34666), .d(n_34733), .o(n_35337) );
ao12s01 g746563 ( .a(n_34801), .b(n_34810), .c(n_34155), .o(n_35372) );
ao12s01 g746564 ( .a(n_34758), .b(n_34810), .c(n_34229), .o(n_35434) );
oa12s01 g746565 ( .a(n_34839), .b(n_34666), .c(n_34774), .o(n_35478) );
ao12s01 g746566 ( .a(n_33237), .b(n_33254), .c(n_33236), .o(n_34096) );
ao12s01 g746567 ( .a(n_34815), .b(n_34810), .c(n_34497), .o(n_35042) );
ao22s01 g746568 ( .a(n_34666), .b(n_34579), .c(n_34810), .d(n_34614), .o(n_35110) );
oa12s01 g746569 ( .a(n_34694), .b(n_34666), .c(n_34696), .o(n_35320) );
oa22s01 g746570 ( .a(n_34810), .b(n_33993), .c(n_34666), .d(n_34643), .o(n_35245) );
oa12s01 g746571 ( .a(n_34609), .b(n_34666), .c(n_34585), .o(n_35071) );
oa22s01 g746572 ( .a(n_34810), .b(n_34645), .c(n_34666), .d(n_33685), .o(n_35016) );
no02s02 g746575 ( .a(FE_OCP_RBN6566_n_33368), .b(n_33300), .o(n_33408) );
no02s01 g746576 ( .a(n_33236), .b(n_33254), .o(n_33237) );
no02s01 g746577 ( .a(n_34810), .b(n_34547), .o(n_35069) );
no02s06 g746578 ( .a(FE_OCP_RBN5585_n_33368), .b(n_33327), .o(n_33450) );
na02s01 g746579 ( .a(n_34666), .b(n_34580), .o(n_35041) );
no02s01 g746580 ( .a(n_34810), .b(n_34613), .o(n_35070) );
in01s01 g746581 ( .a(n_34615), .o(n_34549) );
no02s01 g746582 ( .a(n_34473), .b(n_34580), .o(n_34615) );
na02s01 g746583 ( .a(n_34810), .b(n_34802), .o(n_34938) );
in01s01 g746584 ( .a(n_34885), .o(n_34886) );
no02s01 g746585 ( .a(n_34810), .b(n_34802), .o(n_34885) );
na02s01 g746586 ( .a(n_34612), .b(n_34227), .o(n_34776) );
no02s01 g746587 ( .a(n_34666), .b(n_34735), .o(n_34809) );
in01s01 g746588 ( .a(n_34757), .o(n_34758) );
na02s01 g746589 ( .a(n_34666), .b(n_34738), .o(n_34757) );
na02s01 g746590 ( .a(n_34666), .b(n_34228), .o(n_34775) );
na02s01 g746591 ( .a(n_34666), .b(n_34774), .o(n_34839) );
in01s01 g746592 ( .a(n_34756), .o(n_34805) );
na02s01 g746593 ( .a(n_34666), .b(n_34735), .o(n_34756) );
in01s01 g746594 ( .a(n_34699), .o(n_34637) );
na02s01 g746595 ( .a(n_34612), .b(n_34613), .o(n_34699) );
in01s01 g746596 ( .a(n_34740), .o(n_34692) );
na02s01 g746597 ( .a(n_34612), .b(n_34667), .o(n_34740) );
in01s01 g746598 ( .a(n_34800), .o(n_34801) );
na02s01 g746599 ( .a(n_34666), .b(n_34739), .o(n_34800) );
na02s01 g746600 ( .a(FE_OCP_RBN6725_n_34388), .b(n_34611), .o(n_34697) );
in01s01 g746601 ( .a(n_34644), .o(n_34586) );
na02s01 g746602 ( .a(FE_OCP_RBN6726_n_34388), .b(n_34547), .o(n_34644) );
na02s01 g746603 ( .a(n_34473), .b(n_34696), .o(n_34694) );
in01s01 g746604 ( .a(n_34635), .o(n_34693) );
no02s01 g746605 ( .a(n_34612), .b(n_34611), .o(n_34635) );
in01s01 g746606 ( .a(n_34609), .o(n_34610) );
na02s01 g746607 ( .a(n_34473), .b(n_34585), .o(n_34609) );
no02s02 g746608 ( .a(FE_OCP_RBN6728_n_34388), .b(n_34497), .o(n_34815) );
na02s02 g746609 ( .a(n_34388), .b(n_33910), .o(n_34499) );
no02m04 g746610 ( .a(n_34390), .b(n_34389), .o(n_34475) );
in01s01 g746611 ( .a(n_34417), .o(n_34418) );
na02m04 g746612 ( .a(n_34390), .b(n_34389), .o(n_34417) );
na02s02 g746613 ( .a(FE_OCP_RBN6726_n_34388), .b(n_33911), .o(n_34498) );
na02s02 g746614 ( .a(n_34473), .b(n_34474), .o(n_34760) );
in01s01 g746615 ( .a(n_34545), .o(n_34546) );
na02s02 g746616 ( .a(n_34473), .b(n_34472), .o(n_34545) );
in01s02 g746617 ( .a(n_34496), .o(n_34550) );
no02s01 g746618 ( .a(n_34473), .b(n_34472), .o(n_34496) );
in01s01 g746619 ( .a(n_34638), .o(n_34608) );
na02s01 g746620 ( .a(n_34473), .b(n_34523), .o(n_34638) );
in01s01 g746621 ( .a(n_34606), .o(n_34607) );
na02s01 g746622 ( .a(n_34473), .b(n_34582), .o(n_34606) );
in01s01 g746623 ( .a(n_34544), .o(n_34640) );
no02s01 g746624 ( .a(n_34473), .b(n_34523), .o(n_34544) );
no02s01 g746625 ( .a(n_34612), .b(n_34667), .o(n_34808) );
in01s01 g746626 ( .a(n_34911), .o(n_34912) );
no02s01 g746627 ( .a(n_34666), .b(n_34474), .o(n_34911) );
oa22s01 g746629 ( .a(n_33068), .b(n_32893), .c(n_33113), .d(n_32894), .o(n_34288) );
ao12s01 g746630 ( .a(n_34333), .b(n_34359), .c(n_34332), .o(n_34889) );
ao12s01 g746631 ( .a(n_33990), .b(n_34359), .c(n_33971), .o(n_34420) );
oa12s01 g746632 ( .a(n_33760), .b(n_34300), .c(n_33703), .o(n_34442) );
oa12s01 g746633 ( .a(n_34473), .b(n_34580), .c(n_34579), .o(n_34581) );
no02s02 g746634 ( .a(n_34473), .b(n_33972), .o(n_34867) );
oa12s01 g746635 ( .a(n_34473), .b(n_34643), .c(n_33992), .o(n_34634) );
oa12s01 g746636 ( .a(n_34666), .b(n_34733), .c(n_34073), .o(n_34734) );
na02s06 g746637 ( .a(n_33205), .b(n_33065), .o(n_33206) );
no02s06 g746639 ( .a(n_33340), .b(n_33269), .o(n_33368) );
no02s01 g746640 ( .a(n_34359), .b(n_34332), .o(n_34333) );
oa12f08 g746641 ( .a(n_32988), .b(n_33204), .c(n_32954), .o(n_33254) );
oa22s01 g746642 ( .a(n_33204), .b(n_33011), .c(n_33162), .d(n_33010), .o(n_34051) );
in01s02 g746663 ( .a(n_34666), .o(n_34810) );
in01s03 g746675 ( .a(n_34612), .o(n_34666) );
in01s01 g746679 ( .a(n_34473), .o(n_34612) );
in01s04 g746686 ( .a(FE_OCP_RBN6726_n_34388), .o(n_34473) );
in01s04 g746688 ( .a(n_34390), .o(n_34388) );
na02s04 TIMEBOOST_cell_8884 ( .a(n_22288), .b(FE_OCP_RBN3721_n_20621), .o(TIMEBOOST_net_2929) );
oa12s01 g746690 ( .a(n_34331), .b(n_34330), .c(n_34329), .o(n_34802) );
no02s04 g746691 ( .a(n_33328), .b(n_33253), .o(n_33329) );
no02s06 g746692 ( .a(FE_OCP_RBN2484_FE_RN_657_0), .b(n_32997), .o(n_33205) );
no02s02 g746693 ( .a(FE_OCP_RBN2483_FE_RN_657_0), .b(n_32996), .o(n_33164) );
na02s06 g746694 ( .a(n_33290), .b(n_33217), .o(n_33340) );
in01s01 g746695 ( .a(n_34359), .o(n_34300) );
no02s01 g746696 ( .a(n_34276), .b(n_33815), .o(n_34359) );
na02s01 g746697 ( .a(n_34330), .b(n_34329), .o(n_34331) );
in01s01 g746698 ( .a(n_33113), .o(n_33068) );
ao12s01 g746700 ( .a(n_33026), .b(n_33039), .c(n_33025), .o(n_34222) );
na02s01 TIMEBOOST_cell_6816 ( .a(TIMEBOOST_net_2165), .b(FE_OCPN1612_n_44174), .o(n_36236) );
in01s01 g746702 ( .a(n_34774), .o(n_34299) );
ao12s01 g746703 ( .a(n_34253), .b(n_34252), .c(n_34251), .o(n_34774) );
no02m02 g746705 ( .a(n_33083), .b(n_32963), .o(n_33386) );
no02s01 g746706 ( .a(n_33039), .b(n_33025), .o(n_33026) );
in01s02 g746710 ( .a(n_33290), .o(n_33328) );
no02s06 g746711 ( .a(n_33270), .b(n_33202), .o(n_33290) );
no02f06 g746712 ( .a(n_34233), .b(n_33991), .o(n_34276) );
no02s01 g746713 ( .a(n_34252), .b(n_34251), .o(n_34253) );
in01s01 g746714 ( .a(n_33204), .o(n_33162) );
oa12f08 g746715 ( .a(n_33007), .b(n_33145), .c(n_32968), .o(n_33204) );
no02s01 TIMEBOOST_cell_1881 ( .a(n_35785), .b(FE_OCP_RBN4904_n_44256), .o(TIMEBOOST_net_555) );
ao12s01 g746717 ( .a(n_33111), .b(n_33145), .c(n_33110), .o(n_33968) );
ao12s01 g746718 ( .a(n_34232), .b(n_34231), .c(n_34230), .o(n_34735) );
na02m08 g746719 ( .a(n_33022), .b(n_32978), .o(n_33083) );
no02s01 g746721 ( .a(n_33110), .b(n_33145), .o(n_33111) );
na02s01 g746722 ( .a(n_33234), .b(n_33097), .o(n_33235) );
in01s04 g746723 ( .a(n_33270), .o(n_33609) );
na02m08 g746724 ( .a(n_33189), .b(n_33234), .o(n_33270) );
in01s01 g746725 ( .a(n_34233), .o(n_34234) );
na02f06 g746726 ( .a(n_34212), .b(n_33740), .o(n_34233) );
no02s01 g746727 ( .a(n_34212), .b(n_34211), .o(n_34252) );
no02s01 g746728 ( .a(n_34231), .b(n_34230), .o(n_34232) );
oa12f08 g746729 ( .a(n_32821), .b(n_32980), .c(n_32788), .o(n_33039) );
oa22s01 g746730 ( .a(n_32951), .b(n_32831), .c(n_32980), .d(n_32832), .o(n_34182) );
in01s01 g746731 ( .a(n_34738), .o(n_34229) );
ao12s01 g746732 ( .a(n_34173), .b(n_34172), .c(n_34171), .o(n_34738) );
na02s01 g746733 ( .a(n_33144), .b(n_33099), .o(n_33190) );
na02s01 g746734 ( .a(n_33188), .b(n_33107), .o(n_33220) );
in01s01 g746735 ( .a(n_33022), .o(n_33459) );
no02m06 TIMEBOOST_cell_8054 ( .a(n_6321), .b(n_6244), .o(TIMEBOOST_net_2658) );
in01s01 g746737 ( .a(n_33234), .o(n_33219) );
no02m08 g746738 ( .a(n_33203), .b(n_33109), .o(n_33234) );
no02s04 g746739 ( .a(n_33037), .b(n_33023), .o(n_33067) );
no02f06 g746740 ( .a(n_34174), .b(n_33739), .o(n_34212) );
no02s01 g746741 ( .a(n_34172), .b(n_34171), .o(n_34173) );
oa12f08 g746742 ( .a(n_32925), .b(n_33066), .c(n_32967), .o(n_33145) );
oa22s01 g746743 ( .a(n_33016), .b(n_32984), .c(n_33066), .d(n_32983), .o(n_33945) );
in01s01 g746744 ( .a(n_34227), .o(n_34228) );
oa12s01 g746745 ( .a(n_34170), .b(n_34169), .c(n_34168), .o(n_34227) );
no02s02 TIMEBOOST_cell_1874 ( .a(TIMEBOOST_net_551), .b(n_10770), .o(n_10808) );
no02s01 g746747 ( .a(n_33185), .b(n_33155), .o(n_33218) );
na02s02 g746748 ( .a(n_33378), .b(n_33376), .o(n_33406) );
in01s01 g746750 ( .a(n_32980), .o(n_32951) );
ao12f08 g746751 ( .a(n_32743), .b(n_32924), .c(n_32775), .o(n_32980) );
in01s01 g746752 ( .a(n_33037), .o(n_33038) );
na02s04 g746753 ( .a(n_32977), .b(n_33021), .o(n_33037) );
na02f06 g746755 ( .a(n_34132), .b(n_33681), .o(n_34174) );
no02s01 g746756 ( .a(n_34132), .b(n_33705), .o(n_34172) );
na02s01 g746757 ( .a(n_34169), .b(n_34168), .o(n_34170) );
oa12s02 g746758 ( .a(FE_OCP_RBN4017_n_33034), .b(n_33253), .c(delay_add_ln22_unr20_stage8_stallmux_q_25_), .o(n_33217) );
oa12m06 g746759 ( .a(FE_OCP_RBN4019_n_33034), .b(FE_OCP_RBN5562_n_33097), .c(delay_add_ln22_unr20_stage8_stallmux_q_21_), .o(n_33189) );
ao12m06 g746760 ( .a(FE_OCP_RBN4013_n_33034), .b(n_33107), .c(n_32222), .o(n_33109) );
in01s01 g746761 ( .a(n_33203), .o(n_33188) );
no02m06 g746762 ( .a(n_33103), .b(FE_OCP_RBN4013_n_33034), .o(n_33203) );
ao12s02 g746763 ( .a(FE_OCP_RBN4015_n_33034), .b(n_33199), .c(n_32336), .o(n_33202) );
ao12s02 g746764 ( .a(FE_OCP_RBN4021_n_33034), .b(n_33305), .c(n_32355), .o(n_33269) );
in01s01 g746765 ( .a(n_33143), .o(n_33144) );
no02s04 TIMEBOOST_cell_8777 ( .a(TIMEBOOST_net_2875), .b(n_3016), .o(TIMEBOOST_net_1552) );
no02s02 TIMEBOOST_cell_8564 ( .a(TIMEBOOST_net_1262), .b(n_3718), .o(TIMEBOOST_net_2769) );
ao12s01 g746772 ( .a(n_32899), .b(n_32924), .c(n_32898), .o(n_34137) );
ao12s01 g746774 ( .a(FE_OCP_RBN4007_n_32860), .b(n_32959), .c(n_32991), .o(n_32997) );
oa12s01 g746775 ( .a(FE_OCP_RBN2451_n_32860), .b(n_33063), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_27_), .o(n_33065) );
in01s01 g746776 ( .a(n_34739), .o(n_34155) );
ao12s01 g746777 ( .a(n_34108), .b(n_34107), .c(n_34106), .o(n_34739) );
no02s06 g746779 ( .a(n_32948), .b(n_33252), .o(n_33274) );
in01s02 g746780 ( .a(n_32976), .o(n_32977) );
na02s04 g746781 ( .a(n_32934), .b(n_32942), .o(n_32976) );
na02s02 g746782 ( .a(n_32941), .b(n_32939), .o(n_33023) );
in01s01 g746783 ( .a(n_33378), .o(n_33379) );
no02s01 g746784 ( .a(n_33855), .b(n_33338), .o(n_33378) );
na02s02 g746785 ( .a(n_33326), .b(n_33325), .o(n_33327) );
no02s01 g746786 ( .a(n_33259), .b(n_33323), .o(n_33324) );
no02f08 g746787 ( .a(n_33033), .b(n_33056), .o(n_33106) );
na02f08 g746788 ( .a(n_33077), .b(n_33078), .o(n_33082) );
na02m08 g746790 ( .a(n_33200), .b(n_33150), .o(n_33201) );
na02s01 g746791 ( .a(n_32911), .b(n_32916), .o(n_32947) );
in01s01 g746792 ( .a(n_33184), .o(n_33185) );
no02s01 g746793 ( .a(n_33158), .b(n_33075), .o(n_33184) );
no02s02 g746794 ( .a(n_33104), .b(n_33098), .o(n_33105) );
in01s02 g746795 ( .a(n_32974), .o(n_32975) );
no02s01 g746796 ( .a(n_32963), .b(n_32962), .o(n_32974) );
no03s04 TIMEBOOST_cell_8347 ( .a(FE_OCP_RBN3347_n_47269), .b(n_46424), .c(n_11247), .o(n_11296) );
no02s02 TIMEBOOST_cell_5270 ( .a(n_9089), .b(FE_OCP_RBN5812_n_9014), .o(TIMEBOOST_net_1583) );
no02s01 g746800 ( .a(n_32973), .b(n_32972), .o(n_33488) );
no02m04 g746801 ( .a(n_33102), .b(delay_add_ln22_unr20_stage8_stallmux_q_17_), .o(n_33103) );
no02f08 TIMEBOOST_cell_8170 ( .a(FE_RN_1183_0), .b(n_21529), .o(TIMEBOOST_net_2716) );
in01s01 g746803 ( .a(n_33404), .o(n_33405) );
na02s02 g746804 ( .a(n_33325), .b(n_33339), .o(n_33404) );
in01s01 g746805 ( .a(n_33215), .o(n_33216) );
na02s06 g746806 ( .a(n_33199), .b(n_33198), .o(n_33215) );
in01s01 g746807 ( .a(n_33267), .o(n_33268) );
no02s01 g746808 ( .a(n_33253), .b(n_33231), .o(n_33267) );
in01s01 g746809 ( .a(n_33321), .o(n_33322) );
na02s01 g746810 ( .a(n_33305), .b(n_33851), .o(n_33321) );
na02s01 g746812 ( .a(n_33377), .b(n_33376), .o(n_33402) );
no02s01 g746813 ( .a(n_32961), .b(n_32897), .o(n_33485) );
in01s01 g746814 ( .a(n_33303), .o(n_33304) );
na02s01 g746815 ( .a(n_33247), .b(n_33289), .o(n_33303) );
in01s01 g746816 ( .a(n_33265), .o(n_33266) );
no02s01 g746817 ( .a(n_33211), .b(n_33252), .o(n_33265) );
no02s01 g746818 ( .a(n_32914), .b(n_32920), .o(n_33350) );
na02s01 g746819 ( .a(n_32919), .b(n_32918), .o(n_33166) );
no02s01 g746822 ( .a(n_33158), .b(n_33137), .o(n_33196) );
in01s01 g746823 ( .a(n_33080), .o(n_33081) );
no02s01 g746824 ( .a(n_33104), .b(n_33063), .o(n_33080) );
in01s01 g746825 ( .a(n_33019), .o(n_33020) );
no02s06 g746826 ( .a(n_32957), .b(n_32996), .o(n_33019) );
in01s01 g746827 ( .a(n_33182), .o(n_33183) );
na02s02 g746828 ( .a(n_33157), .b(n_33156), .o(n_33182) );
in01s01 g746829 ( .a(n_33100), .o(n_33101) );
na02s01 g746830 ( .a(n_33079), .b(n_33078), .o(n_33100) );
na02s01 g746831 ( .a(n_33077), .b(n_33055), .o(n_33343) );
no02s01 g746832 ( .a(n_33401), .b(n_33061), .o(n_33452) );
na02s01 g746833 ( .a(n_33053), .b(n_33099), .o(n_33423) );
no02s01 g746834 ( .a(n_33449), .b(n_33102), .o(n_33482) );
no02s01 g746835 ( .a(n_33181), .b(n_33058), .o(n_33535) );
no02s01 g746836 ( .a(n_33151), .b(FE_OCP_RBN5561_n_33097), .o(n_33606) );
ao12s01 g746837 ( .a(n_32940), .b(FE_OCPN865_n_32892), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_21_), .o(n_33524) );
in01s01 g746838 ( .a(n_33250), .o(n_33251) );
ao12s02 g746839 ( .a(n_33233), .b(FE_OCP_RBN4017_n_33034), .c(delay_add_ln22_unr20_stage8_stallmux_q_23_), .o(n_33250) );
in01s01 g746840 ( .a(n_33287), .o(n_33288) );
ao12s02 g746841 ( .a(n_33264), .b(FE_OCP_RBN4017_n_33034), .c(delay_add_ln22_unr20_stage8_stallmux_q_25_), .o(n_33287) );
in01s01 g746842 ( .a(n_33366), .o(n_33367) );
ao12s01 g746843 ( .a(n_33323), .b(FE_OCP_RBN4017_n_33034), .c(delay_add_ln22_unr20_stage8_stallmux_q_27_), .o(n_33366) );
ao12s01 g746844 ( .a(n_32943), .b(FE_OCPN865_n_32892), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_19_), .o(n_33505) );
in01s01 g746845 ( .a(n_33262), .o(n_33263) );
ao12s01 g746846 ( .a(n_32948), .b(FE_OCPN865_n_32892), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_13_), .o(n_33262) );
in01s01 g746847 ( .a(n_33301), .o(n_33302) );
ao12s01 g746848 ( .a(n_32949), .b(FE_OCPN865_n_32892), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_15_), .o(n_33301) );
in01s01 g746849 ( .a(n_33260), .o(n_33261) );
ao12s01 g746850 ( .a(n_33225), .b(FE_OCPN865_n_32892), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_11_), .o(n_33260) );
no02s01 g746851 ( .a(n_32898), .b(n_32924), .o(n_32899) );
ao12s02 g746853 ( .a(n_32995), .b(FE_OCP_RBN2451_n_32860), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_23_), .o(n_33017) );
in01s01 g746854 ( .a(n_33059), .o(n_33060) );
na02s02 TIMEBOOST_cell_8703 ( .a(TIMEBOOST_net_2838), .b(n_1560), .o(n_1638) );
in01s01 g746856 ( .a(n_33140), .o(n_33141) );
ao12s01 g746857 ( .a(n_33098), .b(FE_OCP_RBN2451_n_32860), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_27_), .o(n_33140) );
ao12s01 g746858 ( .a(n_33159), .b(FE_OCP_RBN2477_n_33034), .c(delay_add_ln22_unr20_stage8_stallmux_q_15_), .o(n_33467) );
ao12s01 g746859 ( .a(n_33186), .b(FE_OCP_RBN2477_n_33034), .c(delay_add_ln22_unr20_stage8_stallmux_q_19_), .o(n_33560) );
ao12s01 g746860 ( .a(n_33149), .b(FE_OCP_RBN4019_n_33034), .c(delay_add_ln22_unr20_stage8_stallmux_q_21_), .o(n_33637) );
no02f06 g746861 ( .a(n_34081), .b(n_33951), .o(n_34132) );
no02s01 g746862 ( .a(n_34107), .b(n_34106), .o(n_34108) );
in01s01 g746863 ( .a(n_33066), .o(n_33016) );
oa12f08 g746864 ( .a(n_32905), .b(n_32994), .c(n_32868), .o(n_33066) );
in01s01 g746865 ( .a(n_33447), .o(n_33448) );
ao22m01 g746866 ( .a(FE_OCP_RBN4016_n_33034), .b(n_32335), .c(FE_OCP_RBN2477_n_33034), .d(delay_add_ln22_unr20_stage8_stallmux_q_31_), .o(n_33447) );
oa22s01 g746867 ( .a(FE_OCPN865_n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_17_), .c(FE_OCP_RBN4008_n_32860), .d(n_32362), .o(n_33470) );
oa12s01 g746868 ( .a(n_32877), .b(n_32876), .c(n_32875), .o(n_34085) );
in01s01 g746869 ( .a(n_33178), .o(n_33179) );
oa22s01 g746870 ( .a(FE_OCP_RBN4009_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_), .c(FE_OCP_RBN4008_n_32860), .d(n_33155), .o(n_33178) );
oa22s01 g746872 ( .a(FE_OCP_RBN4009_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_31_), .c(FE_OCP_RBN4008_n_32860), .d(n_32542), .o(n_33213) );
ao12s01 g746873 ( .a(n_32971), .b(n_32994), .c(n_32970), .o(n_33907) );
no02s01 TIMEBOOST_cell_1873 ( .a(n_10768), .b(n_10290), .o(TIMEBOOST_net_551) );
oa22s01 g746875 ( .a(FE_OCP_RBN2477_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_13_), .c(FE_OCP_RBN4016_n_33034), .d(n_32083), .o(n_33455) );
oa22s01 g746876 ( .a(FE_OCP_RBN2477_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_17_), .c(FE_OCP_RBN4016_n_33034), .d(n_32171), .o(n_33519) );
oa12s01 g746877 ( .a(n_34105), .b(n_34104), .c(n_34103), .o(n_34667) );
na02s01 g746878 ( .a(FE_OCP_RBN4022_n_33034), .b(n_32354), .o(n_33376) );
in01s01 g746879 ( .a(n_33855), .o(n_33870) );
no02s02 g746880 ( .a(FE_OCP_RBN4018_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_28_), .o(n_33855) );
in01s01 g746881 ( .a(n_33338), .o(n_33339) );
no02s01 g746882 ( .a(FE_OCP_RBN4018_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_29_), .o(n_33338) );
na02s01 g746883 ( .a(FE_OCP_RBN4018_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_30_), .o(n_33377) );
na02s01 g746884 ( .a(FE_OCP_RBN4018_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_29_), .o(n_33325) );
in01s01 g746885 ( .a(n_33326), .o(n_33300) );
na02s02 g746886 ( .a(FE_OCP_RBN4018_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_28_), .o(n_33326) );
no02s02 g746887 ( .a(FE_OCP_RBN4015_n_33034), .b(n_32283), .o(n_33253) );
na02s06 g746889 ( .a(FE_OCP_RBN2469_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_20_), .o(n_33097) );
in01s01 g746890 ( .a(n_33107), .o(n_33058) );
na02m06 g746891 ( .a(FE_OCP_RBN2468_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_18_), .o(n_33107) );
in01s02 g746892 ( .a(n_33057), .o(n_33102) );
na02s04 g746893 ( .a(FE_OCP_RBN4003_n_33015), .b(delay_add_ln22_unr20_stage8_stallmux_q_16_), .o(n_33057) );
na02s04 g746895 ( .a(FE_OCP_RBN2469_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_22_), .o(n_33199) );
na02s02 g746896 ( .a(FE_OCP_RBN4017_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_26_), .o(n_33305) );
in01s01 g746897 ( .a(n_33259), .o(n_33851) );
no02s01 g746898 ( .a(FE_OCP_RBN4017_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_26_), .o(n_33259) );
no02s01 g746899 ( .a(FE_OCP_RBN4017_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_27_), .o(n_33323) );
no02s02 g746900 ( .a(FE_OCP_RBN4017_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_25_), .o(n_33264) );
no02s06 g746901 ( .a(FE_OCP_RBN4017_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_23_), .o(n_33233) );
in01s01 g746902 ( .a(n_33061), .o(n_33036) );
no02s02 g746903 ( .a(n_33015), .b(n_32082), .o(n_33061) );
in01m04 g746904 ( .a(n_33055), .o(n_33056) );
na02m06 g746905 ( .a(FE_OCP_RBN4002_n_33015), .b(delay_add_ln22_unr20_stage8_stallmux_q_11_), .o(n_33055) );
na02s03 g746906 ( .a(n_33015), .b(n_31855), .o(n_33077) );
na02s02 g746908 ( .a(FE_OCP_RBN4002_n_33015), .b(delay_add_ln22_unr20_stage8_stallmux_q_14_), .o(n_33099) );
in01s01 g746909 ( .a(n_33160), .o(n_33053) );
no02s03 g746910 ( .a(FE_OCP_RBN4003_n_33015), .b(delay_add_ln22_unr20_stage8_stallmux_q_14_), .o(n_33160) );
no02s02 g746911 ( .a(FE_OCP_RBN4003_n_33015), .b(delay_add_ln22_unr20_stage8_stallmux_q_15_), .o(n_33159) );
no02m06 g746912 ( .a(FE_OCP_RBN2469_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_19_), .o(n_33186) );
in01s01 g746913 ( .a(n_33181), .o(n_33152) );
no02s06 g746914 ( .a(FE_OCP_RBN2468_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_18_), .o(n_33181) );
in01s06 g746915 ( .a(n_33151), .o(n_33200) );
no02s08 g746916 ( .a(FE_OCP_RBN4019_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_20_), .o(n_33151) );
in01s04 g746917 ( .a(n_33149), .o(n_33150) );
no02s08 g746918 ( .a(FE_OCP_RBN4019_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_21_), .o(n_33149) );
na02s06 g746919 ( .a(FE_OCP_RBN4015_n_33034), .b(n_32303), .o(n_33198) );
no02s02 g746921 ( .a(FE_OCP_RBN4017_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_24_), .o(n_33231) );
no02s01 g746922 ( .a(FE_OCP_RBN2477_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_12_), .o(n_33401) );
no02s01 g746923 ( .a(FE_OCP_RBN2477_n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_16_), .o(n_33449) );
no02s03 g746924 ( .a(n_32860), .b(n_32464), .o(n_32963) );
no02s03 g746925 ( .a(FE_OCP_RBN5548_FE_OCPN4833_n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_22_), .o(n_32962) );
in01s01 g746927 ( .a(n_32897), .o(n_32916) );
in01s01 g746929 ( .a(n_32915), .o(n_32972) );
na02s06 g746930 ( .a(FE_OCP_RBN5548_FE_OCPN4833_n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_20_), .o(n_32915) );
no02s03 g746931 ( .a(n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_15_), .o(n_32949) );
in01s01 g746933 ( .a(n_32914), .o(n_32944) );
no02s06 g746934 ( .a(n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_14_), .o(n_32914) );
no02s06 g746935 ( .a(n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_12_), .o(n_33252) );
no02s06 g746936 ( .a(n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_13_), .o(n_32948) );
ao12f08 g746937 ( .a(n_32719), .b(n_32834), .c(n_32722), .o(n_32924) );
na02s06 g746938 ( .a(n_32862), .b(n_32861), .o(n_32919) );
in01s01 g746939 ( .a(n_32879), .o(n_32918) );
no02m04 g746940 ( .a(n_32862), .b(n_32861), .o(n_32879) );
no02s01 g746941 ( .a(n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_11_), .o(n_33225) );
in01s01 g746942 ( .a(n_32920), .o(n_32895) );
no02m03 g746943 ( .a(n_32857), .b(n_32275), .o(n_32920) );
in01s01 g746944 ( .a(n_32961), .o(n_33021) );
no02s06 g746945 ( .a(FE_OCP_RBN2452_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_18_), .o(n_32961) );
in01s01 g746946 ( .a(n_32942), .o(n_32943) );
na02s02 g746947 ( .a(n_32857), .b(n_32348), .o(n_32942) );
in01s01 g746948 ( .a(n_32941), .o(n_32973) );
na02s02 g746949 ( .a(n_32857), .b(n_32381), .o(n_32941) );
in01s01 g746950 ( .a(n_32939), .o(n_32940) );
na02s02 g746951 ( .a(n_32857), .b(n_32912), .o(n_32939) );
in01m04 g746952 ( .a(n_33079), .o(n_33033) );
na02m06 g746953 ( .a(n_33014), .b(delay_add_ln22_unr20_stage8_stallmux_q_10_), .o(n_33079) );
in01m04 g746954 ( .a(n_33032), .o(n_33078) );
no02m06 g746955 ( .a(n_33014), .b(delay_add_ln22_unr20_stage8_stallmux_q_10_), .o(n_33032) );
na02s01 g746956 ( .a(FE_OCPN865_n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_), .o(n_33289) );
in01s01 g746957 ( .a(n_33246), .o(n_33247) );
no02s01 g746958 ( .a(FE_OCPN865_n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_), .o(n_33246) );
in01s01 g746959 ( .a(n_33210), .o(n_33211) );
na02s01 g746960 ( .a(FE_OCPN865_n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_12_), .o(n_33210) );
in01s01 g746961 ( .a(n_32893), .o(n_32894) );
na02s01 g746962 ( .a(FE_RN_1716_0), .b(n_32878), .o(n_32893) );
na02s01 g746963 ( .a(n_32876), .b(n_32875), .o(n_32877) );
no02s06 g746964 ( .a(FE_OCP_RBN2451_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_23_), .o(n_32995) );
in01s01 g746965 ( .a(n_33136), .o(n_33137) );
na02s01 g746966 ( .a(FE_OCP_RBN4009_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_29_), .o(n_33136) );
no02s01 g746967 ( .a(FE_OCP_RBN4009_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_29_), .o(n_33158) );
in01s01 g746968 ( .a(n_33075), .o(n_33157) );
no02s01 g746969 ( .a(FE_OCP_RBN4009_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_28_), .o(n_33075) );
na02s01 g746970 ( .a(FE_OCP_RBN4009_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_28_), .o(n_33156) );
in01s01 g746971 ( .a(n_32959), .o(n_32996) );
na02s06 g746972 ( .a(FE_OCP_RBN2451_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_24_), .o(n_32959) );
no02s02 g746973 ( .a(FE_OCP_RBN4007_n_32860), .b(n_32540), .o(n_33063) );
no02f02 g746974 ( .a(FE_OCP_RBN2451_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_25_), .o(n_33474) );
no02s06 g746976 ( .a(FE_OCP_RBN2451_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_24_), .o(n_32957) );
no02s01 g746977 ( .a(FE_OCP_RBN2451_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_26_), .o(n_33104) );
no02s01 g746978 ( .a(FE_OCP_RBN2451_n_32860), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_27_), .o(n_33098) );
no03f04 TIMEBOOST_cell_2515 ( .a(TIMEBOOST_net_290), .b(n_13433), .c(n_13483), .o(n_13552) );
na02s01 g746980 ( .a(n_33013), .b(n_33052), .o(n_33236) );
no02s01 g746981 ( .a(n_32970), .b(n_32994), .o(n_32971) );
in01s06 g746982 ( .a(n_32911), .o(n_32999) );
na02s06 g746983 ( .a(FE_OCP_RBN2452_n_32860), .b(n_32363), .o(n_32911) );
in01s01 g746984 ( .a(n_32936), .o(n_33276) );
no02s03 g746985 ( .a(n_32857), .b(n_32319), .o(n_32936) );
in01s01 g746986 ( .a(n_32934), .o(n_32935) );
na02s02 g746987 ( .a(n_32857), .b(n_32347), .o(n_32934) );
in01s01 g746990 ( .a(n_34081), .o(n_34082) );
na02f06 g746991 ( .a(n_34075), .b(n_33667), .o(n_34081) );
no02s01 g746992 ( .a(n_34075), .b(n_34074), .o(n_34107) );
na02s01 g746993 ( .a(n_34104), .b(n_34103), .o(n_34105) );
in01s01 g746994 ( .a(n_34613), .o(n_34073) );
oa12s01 g746995 ( .a(n_34023), .b(n_34022), .c(n_34021), .o(n_34613) );
in01s01 g746996 ( .a(n_34733), .o(n_34080) );
ao12s01 g746997 ( .a(n_34044), .b(n_34043), .c(n_34042), .o(n_34733) );
na02m06 g746998 ( .a(n_32822), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_9_), .o(n_32878) );
no02m04 g747000 ( .a(n_32822), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_9_), .o(n_32835) );
na02s06 g747001 ( .a(n_32990), .b(n_32989), .o(n_33052) );
in01s01 g747002 ( .a(n_33012), .o(n_33013) );
no02s06 g747003 ( .a(n_32990), .b(n_32989), .o(n_33012) );
na02s01 g747004 ( .a(n_32834), .b(n_32736), .o(n_32876) );
na02s01 g747005 ( .a(n_32833), .b(n_32801), .o(n_33025) );
in01s01 g747006 ( .a(n_33010), .o(n_33011) );
na02s01 g747007 ( .a(n_32988), .b(n_32955), .o(n_33010) );
in01m10 g747037 ( .a(n_32863), .o(n_32860) );
in01s10 g747045 ( .a(n_32863), .o(n_32857) );
no02m06 g747047 ( .a(n_34019), .b(n_33950), .o(n_34075) );
na02s01 g747048 ( .a(n_34022), .b(n_34021), .o(n_34023) );
no02s01 g747049 ( .a(n_34043), .b(n_34042), .o(n_34044) );
oa12f08 g747050 ( .a(n_32884), .b(n_32931), .c(n_32846), .o(n_32994) );
in01s01 TIMEBOOST_cell_8897 ( .a(TIMEBOOST_net_2940), .o(TIMEBOOST_net_2941) );
na02m06 g747083 ( .a(n_32792), .b(n_32762), .o(n_32862) );
no02m08 TIMEBOOST_cell_8113 ( .a(TIMEBOOST_net_2687), .b(n_27168), .o(n_27357) );
ao12s01 g747085 ( .a(n_32798), .b(n_32799), .c(n_32797), .o(n_34058) );
in01s01 g747086 ( .a(n_32985), .o(n_32986) );
ao22s01 g747087 ( .a(n_32904), .b(n_32931), .c(n_32903), .d(n_32888), .o(n_32985) );
no03m08 TIMEBOOST_cell_5778 ( .a(TIMEBOOST_net_1537), .b(FE_OCP_RBN2635_n_29371), .c(n_29673), .o(n_29751) );
ao12s01 g747089 ( .a(n_33996), .b(n_33995), .c(n_33994), .o(n_34696) );
oa12s01 g747090 ( .a(n_34001), .b(n_34000), .c(n_33999), .o(n_34611) );
na02f04 TIMEBOOST_cell_8791 ( .a(TIMEBOOST_net_2882), .b(n_15240), .o(n_15429) );
na02s04 g747093 ( .a(n_32889), .b(n_32683), .o(n_32908) );
no02s06 TIMEBOOST_cell_8785 ( .a(TIMEBOOST_net_2879), .b(TIMEBOOST_net_1081), .o(n_4472) );
in01s01 g747095 ( .a(n_32800), .o(n_32801) );
no02s06 g747096 ( .a(n_32794), .b(n_32793), .o(n_32800) );
na02f08 g747097 ( .a(n_32799), .b(n_32735), .o(n_32834) );
na02s06 g747098 ( .a(n_32794), .b(n_32793), .o(n_32833) );
oa12m04 g747099 ( .a(FE_RN_223_0), .b(n_32714), .c(FE_OCPN1904_n_32554), .o(n_32762) );
in01s01 g747101 ( .a(n_32954), .o(n_32955) );
no02m08 g747102 ( .a(n_32927), .b(delay_add_ln22_unr20_stage8_stallmux_q_8_), .o(n_32954) );
na02m08 g747103 ( .a(n_32927), .b(delay_add_ln22_unr20_stage8_stallmux_q_8_), .o(n_32988) );
in01s01 g747104 ( .a(n_32831), .o(n_32832) );
na02s01 g747105 ( .a(n_32789), .b(n_32821), .o(n_32831) );
no02s01 g747106 ( .a(n_32797), .b(n_32799), .o(n_32798) );
na02s01 g747107 ( .a(n_32969), .b(n_33007), .o(n_33110) );
na02s01 g747108 ( .a(n_34000), .b(n_33999), .o(n_34001) );
in01s01 g747109 ( .a(n_34019), .o(n_34020) );
na02f04 g747110 ( .a(n_33998), .b(n_33624), .o(n_34019) );
no02s01 g747111 ( .a(n_33998), .b(n_33997), .o(n_34043) );
no02s01 g747112 ( .a(n_33995), .b(n_33994), .o(n_33996) );
na03f04 TIMEBOOST_cell_2390 ( .a(FE_OCP_RBN5621_n_18986), .b(n_17732), .c(n_19075), .o(n_19114) );
no02s02 TIMEBOOST_cell_1739 ( .a(FE_OCPN3574_n_30345), .b(n_30882), .o(TIMEBOOST_net_484) );
oa12s01 g747115 ( .a(n_33445), .b(n_33953), .c(n_33572), .o(n_34022) );
ao12s06 g747116 ( .a(FE_RN_256_0), .b(n_32721), .c(FE_OCP_RBN3984_n_32791), .o(n_32761) );
na03f08 TIMEBOOST_cell_6508 ( .a(TIMEBOOST_net_884), .b(n_15409), .c(FE_OCP_RBN6005_n_15704), .o(n_15911) );
no02s02 TIMEBOOST_cell_2137 ( .a(FE_OCP_RBN6159_n_39816), .b(n_39599), .o(TIMEBOOST_net_683) );
in01s01 g747120 ( .a(n_32788), .o(n_32789) );
no03s03 TIMEBOOST_cell_5703 ( .a(n_12402), .b(n_12416), .c(n_12401), .o(TIMEBOOST_net_1421) );
in01m08 g747124 ( .a(n_32889), .o(n_32928) );
na02s06 g747126 ( .a(n_32953), .b(n_32952), .o(n_33007) );
in01s01 g747127 ( .a(n_32968), .o(n_32969) );
no02s06 g747128 ( .a(n_32953), .b(n_32952), .o(n_32968) );
na02s01 g747129 ( .a(n_32708), .b(n_32775), .o(n_32898) );
in01s01 g747130 ( .a(n_32983), .o(n_32984) );
no02s01 g747131 ( .a(n_32926), .b(n_32967), .o(n_32983) );
na02s01 g747132 ( .a(n_33953), .b(n_33464), .o(n_33995) );
oa12f08 g747133 ( .a(n_32733), .b(n_32774), .c(n_32695), .o(n_32799) );
in01s01 g747134 ( .a(n_32931), .o(n_32888) );
ao12f08 g747135 ( .a(n_32814), .b(n_32845), .c(n_32885), .o(n_32931) );
oa12m08 g747136 ( .a(n_32854), .b(n_32856), .c(n_32853), .o(n_32927) );
oa22s01 g747137 ( .a(n_32755), .b(n_32734), .c(n_32756), .d(n_32774), .o(n_34009) );
oa12s01 g747138 ( .a(n_32887), .b(n_32886), .c(n_32885), .o(n_33756) );
no02m04 g747139 ( .a(n_33953), .b(n_33602), .o(n_33998) );
oa12s01 g747140 ( .a(n_33391), .b(n_33952), .c(n_33884), .o(n_34000) );
in01s01 g747141 ( .a(n_34643), .o(n_33993) );
ao12s01 g747142 ( .a(n_33934), .b(n_33952), .c(n_33933), .o(n_34643) );
no02s08 TIMEBOOST_cell_8475 ( .a(TIMEBOOST_net_2724), .b(FE_RN_1830_0), .o(n_12129) );
in01s04 g747149 ( .a(n_32708), .o(n_32743) );
in01s06 g747151 ( .a(n_32870), .o(n_32871) );
na02s10 g747152 ( .a(FE_OCP_RBN3991_FE_RN_1579_0), .b(n_32856), .o(n_32870) );
na02m08 g747153 ( .a(n_32856), .b(n_32853), .o(n_32854) );
in01s01 g747154 ( .a(n_32925), .o(n_32926) );
na02m08 g747155 ( .a(n_32906), .b(delay_add_ln22_unr20_stage8_stallmux_q_6_), .o(n_32925) );
no02m08 g747156 ( .a(n_32906), .b(delay_add_ln22_unr20_stage8_stallmux_q_6_), .o(n_32967) );
na02s01 g747157 ( .a(n_32720), .b(n_32701), .o(n_32875) );
na02s01 g747158 ( .a(n_32867), .b(n_32905), .o(n_32970) );
na02s01 g747159 ( .a(n_32886), .b(n_32885), .o(n_32887) );
na02m04 g747160 ( .a(n_33553), .b(n_33888), .o(n_33953) );
no02s01 g747161 ( .a(n_33952), .b(n_33933), .o(n_33934) );
na02s03 TIMEBOOST_cell_8034 ( .a(FE_OCP_RBN6791_n_20242), .b(n_20608), .o(TIMEBOOST_net_2648) );
na02s01 TIMEBOOST_cell_3975 ( .a(FE_OFN5092_delay_sub_ln23_0_unr25_stage9_stallmux_q), .b(n_38778), .o(TIMEBOOST_net_1078) );
ao12s01 g747164 ( .a(n_32759), .b(FE_OCP_DRV_N1882_n_32758), .c(n_32757), .o(n_33958) );
ao12s01 g747165 ( .a(n_32850), .b(n_32849), .c(n_32848), .o(n_33714) );
in01s01 g747166 ( .a(n_34547), .o(n_33992) );
oa12s01 g747167 ( .a(n_33932), .b(n_33931), .c(n_33930), .o(n_34547) );
ao12s01 g747168 ( .a(n_33894), .b(n_33893), .c(n_33892), .o(n_34580) );
ao12s01 g747169 ( .a(n_33891), .b(n_33890), .c(n_33889), .o(n_34523) );
ao12m08 g747170 ( .a(n_32573), .b(n_46413), .c(FE_OCPN1902_n_32712), .o(n_32741) );
no02m08 TIMEBOOST_cell_3974 ( .a(TIMEBOOST_net_1077), .b(n_14721), .o(n_14891) );
na02f06 TIMEBOOST_cell_6715 ( .a(FE_OCP_RBN5824_n_14552), .b(FE_OCP_RBN2744_n_14114), .o(TIMEBOOST_net_2115) );
in01s01 g747179 ( .a(n_32719), .o(n_32720) );
no02s06 g747180 ( .a(n_32702), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_5_), .o(n_32719) );
na02s01 g747181 ( .a(n_32702), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_5_), .o(n_32701) );
in01m06 g747183 ( .a(n_32867), .o(n_32868) );
na02m06 g747184 ( .a(n_32827), .b(delay_add_ln22_unr20_stage8_stallmux_q_5_), .o(n_32867) );
na02s01 g747186 ( .a(n_32736), .b(n_32735), .o(n_32797) );
in01s01 g747187 ( .a(n_32903), .o(n_32904) );
na02s01 g747188 ( .a(n_32884), .b(n_32847), .o(n_32903) );
na02s01 g747189 ( .a(n_33931), .b(n_33930), .o(n_33932) );
in01s01 g747190 ( .a(n_32774), .o(n_32734) );
ao12f08 g747191 ( .a(n_32718), .b(n_32668), .c(n_32653), .o(n_32774) );
oa12f08 g747192 ( .a(n_32786), .b(n_32817), .c(n_32848), .o(n_32885) );
no02s01 g747193 ( .a(n_32758), .b(n_32757), .o(n_32759) );
no02s01 g747194 ( .a(n_32849), .b(n_32848), .o(n_32850) );
no02s01 g747195 ( .a(n_33893), .b(n_33892), .o(n_33894) );
no02s01 g747196 ( .a(n_33890), .b(n_33889), .o(n_33891) );
in01s01 g747197 ( .a(n_33888), .o(n_33952) );
na03m04 TIMEBOOST_cell_8418 ( .a(n_11303), .b(n_11304), .c(n_11349), .o(TIMEBOOST_net_1776) );
in01s01 g747199 ( .a(n_34614), .o(n_34579) );
oa12s01 g747200 ( .a(n_33799), .b(n_33798), .c(n_33797), .o(n_34614) );
ao12s01 g747201 ( .a(n_33796), .b(n_33795), .c(n_33794), .o(n_34585) );
ao12s01 g747202 ( .a(n_33914), .b(n_33913), .c(n_33912), .o(n_34472) );
in01s01 g747203 ( .a(n_34582), .o(n_33865) );
ao12s01 g747204 ( .a(n_33802), .b(n_33801), .c(n_33800), .o(n_34582) );
na02s06 g747207 ( .a(n_46413), .b(FE_OCP_RBN6521_n_32706), .o(n_32672) );
oa12s08 g747209 ( .a(n_32597), .b(n_32643), .c(FE_OCPN3542_n_32436), .o(n_32698) );
na02s06 g747210 ( .a(n_32671), .b(n_32670), .o(n_32735) );
in01s01 g747211 ( .a(n_32697), .o(n_32736) );
no02f06 g747212 ( .a(n_32671), .b(n_32670), .o(n_32697) );
in01s10 g747213 ( .a(n_32851), .o(n_32830) );
in01s01 g747215 ( .a(n_32846), .o(n_32847) );
no02m08 g747216 ( .a(n_32829), .b(delay_add_ln22_unr20_stage8_stallmux_q_4_), .o(n_32846) );
na02m08 g747217 ( .a(n_32829), .b(delay_add_ln22_unr20_stage8_stallmux_q_4_), .o(n_32884) );
no02s01 g747218 ( .a(n_32669), .b(n_32718), .o(n_32758) );
in01s01 g747219 ( .a(n_32755), .o(n_32756) );
na02s01 g747220 ( .a(n_32696), .b(n_32733), .o(n_32755) );
na02s01 g747221 ( .a(n_32845), .b(n_32813), .o(n_32886) );
no02s01 g747222 ( .a(n_32787), .b(n_32817), .o(n_32849) );
no02s01 g747223 ( .a(n_33801), .b(n_33800), .o(n_33802) );
no02s01 TIMEBOOST_cell_8132 ( .a(n_32444), .b(n_32411), .o(TIMEBOOST_net_2697) );
na02s01 g747225 ( .a(n_33798), .b(n_33797), .o(n_33799) );
no02s01 g747226 ( .a(n_33795), .b(n_33794), .o(n_33796) );
no02s01 g747227 ( .a(n_33913), .b(n_33912), .o(n_33914) );
no02s01 g747228 ( .a(n_34497), .b(n_33929), .o(n_33972) );
no02m08 TIMEBOOST_cell_3337 ( .a(TIMEBOOST_net_959), .b(n_26987), .o(n_27017) );
no02m08 g747230 ( .a(n_32627), .b(n_32626), .o(n_32702) );
oa12s01 g747233 ( .a(n_32694), .b(n_32693), .c(n_32692), .o(n_33917) );
in01s01 g747234 ( .a(FE_OCPN1634_n_33588), .o(n_33689) );
oa12s01 g747235 ( .a(n_32812), .b(n_32811), .c(n_32810), .o(n_33588) );
oa12s01 g747236 ( .a(n_33395), .b(n_33723), .c(n_33421), .o(n_33893) );
oa12s01 g747237 ( .a(n_33465), .b(n_33725), .c(n_33462), .o(n_33890) );
no02m08 g747238 ( .a(n_32617), .b(n_32548), .o(n_32627) );
no02m08 g747242 ( .a(n_32655), .b(n_32654), .o(n_32718) );
in01s01 g747243 ( .a(n_32668), .o(n_32669) );
na02m08 g747244 ( .a(n_32655), .b(n_32654), .o(n_32668) );
in01s01 g747245 ( .a(n_32695), .o(n_32696) );
no02m08 g747246 ( .a(n_32667), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_3_), .o(n_32695) );
na02m08 g747247 ( .a(n_32667), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_3_), .o(n_32733) );
in01s06 g747248 ( .a(n_32815), .o(n_32816) );
no02s10 g747249 ( .a(FE_OCP_RBN3988_n_32772), .b(FE_OCPN4520_n_32820), .o(n_32815) );
in01m06 g747250 ( .a(n_32813), .o(n_32814) );
na02m08 g747251 ( .a(n_32784), .b(delay_add_ln22_unr20_stage8_stallmux_q_3_), .o(n_32813) );
in01s01 g747253 ( .a(n_32786), .o(n_32787) );
na02f08 g747254 ( .a(n_32773), .b(delay_add_ln22_unr20_stage8_stallmux_q_2_), .o(n_32786) );
no02f08 g747255 ( .a(n_32773), .b(delay_add_ln22_unr20_stage8_stallmux_q_2_), .o(n_32817) );
na02s01 g747256 ( .a(n_32693), .b(n_32692), .o(n_32694) );
na02s01 g747257 ( .a(n_32811), .b(n_32810), .o(n_32812) );
in01m02 g747258 ( .a(n_33764), .o(n_33765) );
na02m04 g747259 ( .a(n_33748), .b(n_33495), .o(n_33764) );
no02s01 g747260 ( .a(n_33724), .b(n_33481), .o(n_33798) );
no02s01 g747261 ( .a(n_33722), .b(n_33394), .o(n_33795) );
no02s01 g747262 ( .a(n_33748), .b(n_33556), .o(n_33801) );
oa12s01 g747263 ( .a(n_33296), .b(n_45753), .c(n_33840), .o(n_33913) );
oa12s01 g747264 ( .a(n_33887), .b(n_45753), .c(n_33885), .o(n_34497) );
in01s10 g747270 ( .a(n_32617), .o(n_32643) );
in01s01 g747275 ( .a(n_33724), .o(n_33725) );
no02s01 g747276 ( .a(n_45753), .b(n_33444), .o(n_33724) );
in01s01 g747277 ( .a(n_33722), .o(n_33723) );
no02s01 g747278 ( .a(n_45753), .b(n_33335), .o(n_33722) );
na02s01 g747279 ( .a(n_45753), .b(n_33885), .o(n_33887) );
na02s04 TIMEBOOST_cell_8527 ( .a(TIMEBOOST_net_2750), .b(n_14068), .o(n_14176) );
no02m04 g747281 ( .a(n_45753), .b(n_33497), .o(n_33748) );
in01s01 g747282 ( .a(n_32653), .o(n_32757) );
ao22s01 g747288 ( .a(n_32616), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_), .c(n_32638), .d(n_31260), .o(n_32693) );
ao12s01 g747289 ( .a(n_32751), .b(n_32770), .c(delay_add_ln22_unr20_stage8_stallmux_q_1_), .o(n_32811) );
in01s01 g747290 ( .a(n_34645), .o(n_33685) );
oa12s02 g747291 ( .a(n_33631), .b(n_33630), .c(n_33629), .o(n_34645) );
no02s04 TIMEBOOST_cell_8678 ( .a(TIMEBOOST_net_1187), .b(n_36615), .o(TIMEBOOST_net_2826) );
no02s06 TIMEBOOST_cell_1568 ( .a(TIMEBOOST_net_398), .b(n_8176), .o(n_8266) );
no02s20 g747297 ( .a(n_32754), .b(n_32731), .o(n_32752) );
no02s01 g747298 ( .a(n_32770), .b(delay_add_ln22_unr20_stage8_stallmux_q_1_), .o(n_32751) );
na02s10 g747299 ( .a(n_32855), .b(n_32690), .o(n_32853) );
na02s01 g747300 ( .a(n_33630), .b(n_33629), .o(n_33631) );
oa12s08 g747301 ( .a(n_32791), .b(FE_OCP_RBN6527_n_44962), .c(n_32529), .o(n_32711) );
in01s08 g747302 ( .a(n_32597), .o(n_32598) );
no02s02 TIMEBOOST_cell_3867 ( .a(FE_OCP_RBN6562_n_33208), .b(n_33256), .o(TIMEBOOST_net_1024) );
ao12s10 g747305 ( .a(n_32554), .b(FE_OCP_RBN4633_n_44962), .c(delay_xor_ln21_unr21_stage8_stallmux_q_9_), .o(n_32579) );
no02s02 TIMEBOOST_cell_7080 ( .a(TIMEBOOST_net_2298), .b(n_31835), .o(TIMEBOOST_net_2016) );
in01s06 g747307 ( .a(n_32716), .o(n_32717) );
oa12s10 g747308 ( .a(n_32689), .b(n_32688), .c(FE_OCP_RBN6526_n_44962), .o(n_32716) );
in01s08 g747309 ( .a(n_32729), .o(n_32730) );
no02m20 g747310 ( .a(n_32666), .b(n_32818), .o(n_32729) );
no02m06 g747311 ( .a(n_33627), .b(n_33628), .o(n_45753) );
in01s01 g747312 ( .a(n_34474), .o(n_33929) );
ao12s01 g747313 ( .a(n_33864), .b(n_33863), .c(n_33862), .o(n_34474) );
in01s01 g747314 ( .a(n_33910), .o(n_33911) );
ao12s01 g747315 ( .a(n_33843), .b(n_33842), .c(n_33841), .o(n_33910) );
no02s40 g747317 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_9_), .b(FE_OCP_RBN4633_n_44962), .o(n_32554) );
in01m08 g747318 ( .a(FE_OCP_RBN3984_n_32791), .o(n_32553) );
na02m40 g747319 ( .a(n_32529), .b(FE_OCP_RBN6527_n_44962), .o(n_32791) );
no02m80 g747321 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_6_), .b(FE_OCP_RBN7015_n_44962), .o(n_32706) );
no02m06 TIMEBOOST_cell_2123 ( .a(n_43468), .b(n_43637), .o(TIMEBOOST_net_676) );
na03f08 TIMEBOOST_cell_8140 ( .a(n_23443), .b(n_23503), .c(n_23517), .o(TIMEBOOST_net_2701) );
na02m40 g747327 ( .a(FE_OCP_RBN6526_n_44962), .b(n_32624), .o(n_32855) );
in01s10 g747328 ( .a(n_32754), .o(n_32715) );
no02s80 g747330 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_6_), .b(FE_OCP_RBN4633_n_44962), .o(n_32818) );
na02s40 g747331 ( .a(n_32688), .b(FE_OCP_RBN6526_n_44962), .o(n_32689) );
na02s20 g747332 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_8_), .b(FE_OCP_RBN4633_n_44962), .o(n_32690) );
no02s20 g747333 ( .a(n_32637), .b(FE_OCP_RBN6526_n_44962), .o(n_32666) );
no02s01 g747336 ( .a(n_33863), .b(n_33862), .o(n_33864) );
no02s01 g747337 ( .a(n_33842), .b(n_33841), .o(n_33843) );
in01m08 g747338 ( .a(n_32551), .o(n_32552) );
na03f06 TIMEBOOST_cell_2278 ( .a(n_23393), .b(n_23373), .c(n_23374), .o(FE_RN_2366_0) );
in01s01 g747342 ( .a(n_32682), .o(n_32683) );
oa12s03 g747343 ( .a(n_32665), .b(FE_OCP_RBN4633_n_44962), .c(delay_xor_ln22_unr21_stage8_stallmux_q_10_), .o(n_32682) );
in01m10 g747346 ( .a(n_32663), .o(n_32664) );
no02m06 TIMEBOOST_cell_1890 ( .a(TIMEBOOST_net_559), .b(n_11148), .o(n_11223) );
na02m08 TIMEBOOST_cell_5154 ( .a(FE_RN_294_0), .b(n_25041), .o(TIMEBOOST_net_1525) );
oa12s01 g747350 ( .a(n_33579), .b(n_33578), .c(n_33359), .o(n_33630) );
in01s01 g747351 ( .a(n_32638), .o(n_32616) );
in01s01 g747353 ( .a(FE_OCPN1701_n_33544), .o(n_32728) );
ao12s01 g747354 ( .a(n_32662), .b(n_32661), .c(delay_add_ln22_unr20_stage8_stallmux_q_0_), .o(n_33544) );
in01s01 g747356 ( .a(n_33768), .o(n_32574) );
oa22s01 g747357 ( .a(FE_OCPN6909_n_32525), .b(n_30905), .c(n_32432), .d(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .o(n_33768) );
oa22s08 g747359 ( .a(FE_OCP_RBN4633_n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_10_), .c(n_32402), .d(FE_OCP_RBN6527_n_44962), .o(n_32549) );
in01m40 g747361 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_8_), .o(n_32529) );
in01s20 g747363 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_6_), .o(n_32440) );
in01m40 g747365 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_8_), .o(n_32624) );
in01s20 g747367 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_6_), .o(n_32637) );
in01s80 g747369 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_9_), .o(n_32688) );
in01s20 g747371 ( .a(n_32577), .o(n_32599) );
in01s03 g747373 ( .a(n_32600), .o(n_32439) );
no02m80 g747374 ( .a(FE_OCP_RBN7008_n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_4_), .o(n_32600) );
na02m06 TIMEBOOST_cell_8829 ( .a(TIMEBOOST_net_2901), .b(n_4204), .o(n_4538) );
no02s01 g747377 ( .a(FE_OCPN6909_n_32525), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .o(n_32692) );
no02s01 g747378 ( .a(n_32661), .b(delay_add_ln22_unr20_stage8_stallmux_q_0_), .o(n_32662) );
na02s40 g747379 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_10_), .b(FE_OCP_RBN4633_n_44962), .o(n_32665) );
no02s40 g747381 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_4_), .b(FE_OCP_RBN4633_n_44962), .o(n_32635) );
na02s10 g747382 ( .a(n_32630), .b(delay_add_ln22_unr20_stage8_stallmux_q_0_), .o(n_32810) );
no02m06 TIMEBOOST_cell_8867 ( .a(TIMEBOOST_net_2920), .b(TIMEBOOST_net_2676), .o(n_25889) );
na02s01 g747384 ( .a(n_33578), .b(n_33702), .o(n_33842) );
in01s06 g747385 ( .a(n_32547), .o(n_32548) );
no02s02 TIMEBOOST_cell_3869 ( .a(n_37416), .b(n_37152), .o(TIMEBOOST_net_1025) );
in01s04 g747387 ( .a(n_32572), .o(n_32573) );
no02m04 TIMEBOOST_cell_1658 ( .a(TIMEBOOST_net_443), .b(n_8895), .o(FE_RN_1778_0) );
in01s03 g747389 ( .a(n_32651), .o(n_32652) );
ao12m06 g747390 ( .a(n_32634), .b(FE_OCP_RBN4633_n_44962), .c(delay_xor_ln22_unr21_stage8_stallmux_q_7_), .o(n_32651) );
in01m08 g747391 ( .a(n_32678), .o(n_32679) );
no02s01 TIMEBOOST_cell_4861 ( .a(TIMEBOOST_net_1378), .b(n_37094), .o(n_37142) );
na03m08 TIMEBOOST_cell_8316 ( .a(TIMEBOOST_net_658), .b(n_35193), .c(n_30546), .o(n_35192) );
no02f04 TIMEBOOST_cell_1787 ( .a(FE_RN_2649_0), .b(n_15644), .o(TIMEBOOST_net_508) );
oa12s01 g747395 ( .a(n_33747), .b(n_33746), .c(n_33745), .o(n_34389) );
in01s10 g747396 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_10_), .o(n_32402) );
in01s20 g747400 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_4_), .o(n_32389) );
in01m03 g747402 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_10_), .o(n_32623) );
in01m80 g747404 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_2_), .o(n_32615) );
in01s20 g747407 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_4_), .o(n_32622) );
no02m20 g747409 ( .a(n_32595), .b(n_32522), .o(n_32523) );
na02m20 g747410 ( .a(n_32578), .b(n_32582), .o(n_32601) );
na02s20 g747412 ( .a(n_32687), .b(n_32632), .o(n_32649) );
in01s06 g747413 ( .a(n_32704), .o(n_32709) );
no02s40 g747414 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_7_), .b(FE_OCP_RBN4633_n_44962), .o(n_32704) );
no02m80 g747419 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_5_), .b(FE_OCP_RBN7015_n_44962), .o(n_32436) );
no02s04 TIMEBOOST_cell_3868 ( .a(TIMEBOOST_net_1024), .b(n_33361), .o(n_33397) );
na02m08 TIMEBOOST_cell_2895 ( .a(TIMEBOOST_net_738), .b(n_2222), .o(n_2303) );
in01m01 g747422 ( .a(n_32634), .o(n_32621) );
no02f06 g747423 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_7_), .b(FE_OCP_RBN4633_n_44962), .o(n_32634) );
no02m80 g747424 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_5_), .b(FE_OCP_RBN7015_n_44962), .o(n_32820) );
na02s06 TIMEBOOST_cell_3910 ( .a(TIMEBOOST_net_1045), .b(n_44875), .o(n_38050) );
na02s01 g747426 ( .a(n_33746), .b(n_33516), .o(n_33578) );
na02s01 g747427 ( .a(n_33746), .b(n_33745), .o(n_33747) );
in01f08 g747428 ( .a(n_32520), .o(n_32521) );
in01m10 g747430 ( .a(n_32472), .o(n_32473) );
in01s10 g747432 ( .a(n_32659), .o(n_32660) );
no02s02 g747436 ( .a(n_33815), .b(n_33763), .o(n_33816) );
na02m04 g747438 ( .a(n_33746), .b(n_33360), .o(n_33533) );
in01s01 g747445 ( .a(FE_OCPN6909_n_32525), .o(n_32432) );
oa22s10 g747446 ( .a(n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_0_), .c(FE_OCP_RBN7005_n_44962), .d(n_32387), .o(n_32525) );
in01s01 g747447 ( .a(n_32630), .o(n_32661) );
na02s03 TIMEBOOST_cell_5140 ( .a(FE_OCP_RBN2868_n_9188), .b(FE_OFN4771_n_8309), .o(TIMEBOOST_net_1518) );
in01s01 g747449 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_27_), .o(n_32355) );
in01s01 g747452 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_30_), .o(n_32354) );
in01s20 g747454 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_7_), .o(n_32399) );
in01s20 g747456 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_5_), .o(n_32388) );
in01s20 g747459 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_5_), .o(n_32613) );
in01s01 g747461 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_), .o(n_33155) );
no02s04 TIMEBOOST_cell_1592 ( .a(TIMEBOOST_net_410), .b(n_34858), .o(n_34901) );
no02s20 g747466 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_0_), .b(n_44962), .o(n_32568) );
in01m20 g747467 ( .a(n_32578), .o(n_32595) );
na02f80 g747468 ( .a(n_32367), .b(n_44962), .o(n_32578) );
no02s40 g747472 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_0_), .b(FE_OCP_RBN7005_n_44962), .o(n_32522) );
na02s40 g747473 ( .a(n_32387), .b(n_44962), .o(n_32582) );
in01m20 g747474 ( .a(n_32433), .o(n_32602) );
na02s80 g747479 ( .a(n_32543), .b(n_44962), .o(n_32687) );
no02s80 g747481 ( .a(FE_OCP_RBN7008_n_44962), .b(delay_xor_ln22_unr21_stage8_stallmux_q_3_), .o(n_32731) );
oa12s02 g747484 ( .a(n_33721), .b(n_33682), .c(n_33571), .o(n_33815) );
na02m06 g747485 ( .a(n_33446), .b(n_33363), .o(n_33746) );
in01s01 g747492 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_23_), .o(n_32336) );
in01s01 g747495 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_31_), .o(n_32335) );
in01f80 g747497 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_1_), .o(n_32367) );
in01s40 g747499 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_0_), .o(n_32387) );
in01s80 g747504 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_0_), .o(n_32543) );
in01s80 g747506 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_1_), .o(n_32564) );
in01s01 g747511 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_25_), .o(n_32991) );
in01s01 g747513 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_31_), .o(n_32542) );
in01s01 g747515 ( .a(n_33721), .o(n_34211) );
no02s02 g747516 ( .a(n_33705), .b(n_33654), .o(n_33721) );
no02f02 TIMEBOOST_cell_4011 ( .a(n_20290), .b(n_20189), .o(TIMEBOOST_net_1096) );
in01m02 g747526 ( .a(n_32546), .o(n_32513) );
in01s01 g747530 ( .a(n_32519), .o(n_32469) );
no02s02 g747534 ( .a(n_33814), .b(n_33793), .o(n_35542) );
in01s01 g747538 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_26_), .o(n_32540) );
no02f04 TIMEBOOST_cell_4010 ( .a(n_35271), .b(TIMEBOOST_net_1095), .o(n_35324) );
no02s01 g747542 ( .a(n_33397), .b(n_33759), .o(n_33814) );
no02s01 g747543 ( .a(n_33375), .b(n_33758), .o(n_33793) );
no02s02 g747544 ( .a(n_33556), .b(n_33515), .o(n_33557) );
in01s02 g747545 ( .a(n_33672), .o(n_33705) );
no02s02 g747546 ( .a(n_34074), .b(n_33603), .o(n_33672) );
in01f02 g747553 ( .a(n_32311), .o(n_32286) );
in01s02 g747557 ( .a(n_32310), .o(n_32285) );
in01m02 g747561 ( .a(n_32517), .o(n_32466) );
in01s01 g747566 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_22_), .o(n_32303) );
in01s01 g747568 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_24_), .o(n_32283) );
in01s01 g747570 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_22_), .o(n_32464) );
in01s01 g747572 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_21_), .o(n_32912) );
in01s01 g747575 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_1_), .o(n_36898) );
na02s02 g747577 ( .a(n_33361), .b(n_33362), .o(n_33363) );
no02s01 g747578 ( .a(n_33481), .b(n_33440), .o(n_33465) );
in01s02 g747579 ( .a(n_33498), .o(n_33556) );
no02s02 g747580 ( .a(n_33481), .b(n_33442), .o(n_33498) );
oa12s02 g747581 ( .a(n_33480), .b(n_33479), .c(FE_OCP_RBN2532_n_33372), .o(n_34074) );
in01s01 g747582 ( .a(n_33397), .o(n_33375) );
no02s02 TIMEBOOST_cell_4003 ( .a(n_3214), .b(n_2913), .o(TIMEBOOST_net_1092) );
ao12s06 g747585 ( .a(n_31947), .b(n_32324), .c(n_31898), .o(n_32382) );
oa12s02 g747586 ( .a(n_32068), .b(n_45755), .c(n_47272), .o(n_32349) );
no02s02 g747587 ( .a(n_32333), .b(n_47271), .o(n_32366) );
in01s01 g747588 ( .a(n_32364), .o(n_32365) );
no02s01 TIMEBOOST_cell_1422 ( .a(n_24792), .b(TIMEBOOST_net_325), .o(n_24904) );
oa12s06 g747590 ( .a(n_31727), .b(n_45517), .c(n_31594), .o(n_32226) );
no02m08 g747591 ( .a(n_32200), .b(FE_OCPN3586_n_31704), .o(n_32244) );
oa12s04 g747592 ( .a(n_31681), .b(n_32223), .c(n_32197), .o(n_32225) );
no02s04 g747593 ( .a(n_32198), .b(n_31703), .o(n_32243) );
ao12s04 g747594 ( .a(n_31706), .b(n_32190), .c(n_31702), .o(n_32242) );
no02s01 TIMEBOOST_cell_1512 ( .a(n_3213), .b(TIMEBOOST_net_370), .o(n_3454) );
in01s02 g747602 ( .a(n_32395), .o(n_32468) );
ao12s01 g747604 ( .a(n_33571), .b(n_33704), .c(n_33762), .o(n_33763) );
ao12s01 g747605 ( .a(n_34072), .b(n_34071), .c(n_34070), .o(n_35655) );
in01s01 g747606 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_19_), .o(n_32222) );
in01s01 g747609 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_19_), .o(n_32348) );
in01s01 g747611 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_20_), .o(n_32381) );
na02s06 g747613 ( .a(n_32362), .b(n_32276), .o(n_32363) );
na02s01 g747614 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_17_), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_), .o(n_32347) );
no02s01 g747615 ( .a(n_34071), .b(n_34070), .o(n_34072) );
no02s01 TIMEBOOST_cell_1421 ( .a(n_24132), .b(n_24151), .o(TIMEBOOST_net_325) );
no02s02 g747617 ( .a(n_45755), .b(n_47272), .o(n_32333) );
no02s08 g747618 ( .a(n_45517), .b(n_31594), .o(n_32200) );
no02s04 g747619 ( .a(n_32223), .b(n_32197), .o(n_32198) );
na02s03 g747620 ( .a(n_32191), .b(n_31841), .o(n_32241) );
no02s01 TIMEBOOST_cell_1511 ( .a(n_3229), .b(n_2654), .o(TIMEBOOST_net_370) );
no02s01 g747622 ( .a(n_33394), .b(n_33393), .o(n_33395) );
no02s01 g747623 ( .a(n_33812), .b(n_33761), .o(n_33813) );
oa12s02 g747624 ( .a(n_33374), .b(n_33356), .c(FE_OCP_RBN2532_n_33372), .o(n_33481) );
in01s01 g747625 ( .a(n_33997), .o(n_33480) );
na02s02 g747626 ( .a(n_33419), .b(n_33464), .o(n_33997) );
no02s01 g747627 ( .a(n_33420), .b(n_33418), .o(n_33445) );
na02s01 TIMEBOOST_cell_8806 ( .a(n_42339), .b(n_42413), .o(TIMEBOOST_net_2890) );
oa12f04 g747631 ( .a(n_32070), .b(n_32300), .c(n_31869), .o(n_32330) );
no02f06 g747632 ( .a(n_32301), .b(n_32055), .o(n_32346) );
in01s02 g747633 ( .a(n_32219), .o(n_32220) );
no02s01 TIMEBOOST_cell_1508 ( .a(TIMEBOOST_net_368), .b(n_3533), .o(n_3582) );
oa12f06 g747637 ( .a(n_31788), .b(n_32169), .c(n_32168), .o(n_32196) );
no02f06 g747638 ( .a(n_32170), .b(n_31763), .o(n_32218) );
no02m06 g747640 ( .a(n_32151), .b(n_31787), .o(n_32195) );
in01f02 g747641 ( .a(n_32255), .o(n_32240) );
in01m02 g747647 ( .a(n_32384), .o(n_32358) );
oa22f04 g747648 ( .a(n_32277), .b(n_32133), .c(n_32278), .d(n_32132), .o(n_32384) );
in01m02 g747649 ( .a(n_32380), .o(n_32428) );
in01f02 g747651 ( .a(n_32394), .o(n_32463) );
ao22f04 g747652 ( .a(FE_OCP_RBN5218_n_32279), .b(n_32099), .c(n_32279), .d(n_32100), .o(n_32394) );
oa12s01 g747653 ( .a(n_33299), .b(n_33298), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n_33337) );
na02s02 g747654 ( .a(n_33443), .b(n_33463), .o(n_33497) );
in01s01 g747655 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_17_), .o(n_32171) );
in01s01 g747658 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_17_), .o(n_32362) );
na02s01 g747662 ( .a(n_33298), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n_33299) );
no02f06 g747663 ( .a(n_32300), .b(n_31869), .o(n_32301) );
no02f06 g747665 ( .a(n_32169), .b(n_32168), .o(n_32170) );
no02m06 g747666 ( .a(n_32150), .b(n_32149), .o(n_32151) );
in01s01 g747667 ( .a(n_33760), .o(n_33761) );
no02s01 g747668 ( .a(n_33700), .b(n_33990), .o(n_33760) );
in01s01 g747669 ( .a(n_33297), .o(n_34070) );
no02s01 TIMEBOOST_cell_1507 ( .a(n_3532), .b(n_2731), .o(TIMEBOOST_net_368) );
oa22s01 g747676 ( .a(n_32061), .b(n_31894), .c(FE_OCP_RBN6224_n_32061), .d(n_31893), .o(n_32147) );
oa22s01 g747677 ( .a(n_32111), .b(n_31769), .c(n_32112), .d(n_31768), .o(n_32192) );
in01s02 g747679 ( .a(n_32190), .o(n_32191) );
in01s06 g747680 ( .a(n_32223), .o(n_32190) );
na02s10 g747681 ( .a(n_32089), .b(n_31879), .o(n_32223) );
oa22s01 g747682 ( .a(n_32236), .b(n_32209), .c(n_32237), .d(n_32208), .o(n_32281) );
oa22s01 g747683 ( .a(n_32260), .b(n_31989), .c(n_32261), .d(n_31988), .o(n_32325) );
in01s02 g747685 ( .a(n_32324), .o(n_32343) );
no02s06 TIMEBOOST_cell_4078 ( .a(TIMEBOOST_net_1129), .b(FE_OCP_RBN6019_n_46959), .o(n_30829) );
ao12m08 g747690 ( .a(n_32108), .b(n_32238), .c(n_32021), .o(n_32280) );
no02s01 g747691 ( .a(n_33812), .b(n_33989), .o(n_34441) );
oa12s01 g747692 ( .a(n_33699), .b(n_33571), .c(n_33684), .o(n_34419) );
in01s01 g747693 ( .a(n_33443), .o(n_33444) );
no02s02 g747694 ( .a(n_33358), .b(n_33421), .o(n_33443) );
no02m08 TIMEBOOST_cell_1718 ( .a(TIMEBOOST_net_473), .b(n_38956), .o(n_39163) );
ao12s01 g747696 ( .a(FE_OCP_RBN2532_n_33372), .b(n_33513), .c(n_33512), .o(n_33515) );
in01s01 g747697 ( .a(n_33394), .o(n_33374) );
no02s06 TIMEBOOST_cell_1804 ( .a(TIMEBOOST_net_516), .b(n_11205), .o(n_11275) );
ao12s01 g747699 ( .a(FE_OCP_RBN2532_n_33372), .b(n_33390), .c(n_33441), .o(n_33442) );
ao12s02 g747700 ( .a(FE_OCP_RBN2531_n_33372), .b(n_33532), .c(n_33227), .o(n_33603) );
in01s01 g747701 ( .a(n_33420), .o(n_33464) );
ao12s01 g747702 ( .a(FE_OCP_RBN2532_n_33372), .b(n_33391), .c(n_33552), .o(n_33420) );
oa12s01 g747703 ( .a(n_33372), .b(n_33418), .c(n_33169), .o(n_33419) );
ao12s01 g747704 ( .a(n_33571), .b(n_33653), .c(n_33720), .o(n_33654) );
in01s01 g747705 ( .a(n_33703), .o(n_33704) );
ao12s01 g747706 ( .a(n_33571), .b(n_33684), .c(n_33683), .o(n_33703) );
ao12s01 g747707 ( .a(n_33991), .b(FE_OCP_RBN2534_n_33372), .c(n_33743), .o(n_34329) );
ao12s01 g747708 ( .a(n_33951), .b(n_33372), .c(n_33670), .o(n_34168) );
na02s06 TIMEBOOST_cell_1355 ( .a(n_19534), .b(n_18032), .o(TIMEBOOST_net_292) );
na02f20 g747715 ( .a(FE_OCP_RBN6387_n_32238), .b(n_32107), .o(n_32279) );
na02m10 g747716 ( .a(n_32088), .b(n_31683), .o(n_32090) );
na02s10 g747717 ( .a(n_32088), .b(n_31808), .o(n_32089) );
in01m04 g747719 ( .a(n_32150), .o(n_32145) );
no02s02 g747720 ( .a(n_32088), .b(n_32086), .o(n_32087) );
no02m10 g747721 ( .a(n_32088), .b(n_32086), .o(n_32150) );
no02s01 g747722 ( .a(n_33741), .b(n_33792), .o(n_34251) );
no02s01 g747723 ( .a(n_33680), .b(n_33599), .o(n_34171) );
no02s01 g747724 ( .a(n_33625), .b(n_33671), .o(n_34042) );
no02s01 g747725 ( .a(n_33671), .b(n_33626), .o(n_33479) );
na02s01 g747726 ( .a(n_33702), .b(n_33516), .o(n_33745) );
na02s01 g747727 ( .a(n_33373), .b(n_33601), .o(n_33994) );
no02s01 g747728 ( .a(n_33668), .b(n_33701), .o(n_34106) );
no02s01 g747729 ( .a(n_33421), .b(n_33393), .o(n_33794) );
no02s01 g747730 ( .a(n_33840), .b(n_33317), .o(n_33885) );
na02s01 g747731 ( .a(n_33417), .b(n_33312), .o(n_33629) );
no02s01 g747732 ( .a(n_33884), .b(n_33353), .o(n_33933) );
no02s01 g747733 ( .a(n_33258), .b(n_33242), .o(n_33298) );
no02s01 g747734 ( .a(n_33239), .b(FE_OCP_RBN2534_n_33372), .o(n_33812) );
in01s01 g747735 ( .a(n_33699), .o(n_33700) );
na02s01 g747736 ( .a(n_33684), .b(n_33571), .o(n_33699) );
na02s01 g747737 ( .a(n_33357), .b(n_33334), .o(n_33358) );
no02s02 g747738 ( .a(n_33414), .b(n_33462), .o(n_33463) );
na02s01 g747739 ( .a(n_33417), .b(n_33415), .o(n_33416) );
no02s01 g747740 ( .a(n_33393), .b(n_32902), .o(n_33356) );
no02m04 TIMEBOOST_cell_8656 ( .a(n_36716), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_2815) );
na02s01 g747742 ( .a(n_33601), .b(n_33600), .o(n_33602) );
no02s01 g747743 ( .a(n_33670), .b(n_33372), .o(n_33951) );
no02s01 g747744 ( .a(FE_OCP_RBN2534_n_33372), .b(n_33743), .o(n_33991) );
no02s01 g747745 ( .a(n_33792), .b(n_33743), .o(n_33682) );
no02s01 g747746 ( .a(n_33990), .b(n_33970), .o(n_34332) );
no02s01 g747747 ( .a(n_33762), .b(n_33571), .o(n_33989) );
no02s01 g747748 ( .a(n_33440), .b(n_33462), .o(n_33797) );
no02s01 g747749 ( .a(n_33496), .b(n_33461), .o(n_33800) );
in01m03 g747751 ( .a(n_32300), .o(n_32296) );
oa12f10 g747752 ( .a(n_32027), .b(n_32188), .c(n_31949), .o(n_32300) );
oa12f10 g747755 ( .a(n_31810), .b(n_32000), .c(n_31686), .o(n_32169) );
oa22s01 g747756 ( .a(n_32002), .b(n_31912), .c(n_32001), .d(n_31913), .o(n_32085) );
oa22s01 g747757 ( .a(n_32032), .b(n_31737), .c(n_32033), .d(n_31736), .o(n_32113) );
oa12f06 g747759 ( .a(n_31747), .b(n_32000), .c(n_31554), .o(n_32143) );
oa22s01 g747760 ( .a(n_32214), .b(n_32180), .c(n_32215), .d(FE_OCP_RBN3428_n_32180), .o(n_32263) );
oa22s01 g747761 ( .a(n_32216), .b(n_32137), .c(FE_OCP_RBN6227_n_32216), .d(n_32136), .o(n_32262) );
in01m03 g747762 ( .a(n_32277), .o(n_32278) );
oa12f06 g747763 ( .a(n_32028), .b(n_32188), .c(n_31902), .o(n_32277) );
ao12s01 g747764 ( .a(n_33950), .b(n_33372), .c(n_33626), .o(n_34103) );
in01s01 g747765 ( .a(n_33758), .o(n_33759) );
oa22s01 g747766 ( .a(n_33571), .b(n_33362), .c(n_33372), .d(n_33396), .o(n_33758) );
oa12s01 g747767 ( .a(n_33413), .b(n_33571), .c(n_33441), .o(n_33889) );
oa12s01 g747768 ( .a(n_33738), .b(n_33571), .c(n_33720), .o(n_34230) );
oa12s01 g747769 ( .a(n_33600), .b(n_33571), .c(n_33554), .o(n_34021) );
oa22s01 g747770 ( .a(n_33372), .b(n_33114), .c(n_33571), .d(n_33552), .o(n_33999) );
oa12s01 g747771 ( .a(n_33817), .b(n_33571), .c(n_33512), .o(n_33930) );
oa12s01 g747772 ( .a(n_33357), .b(n_33571), .c(n_33314), .o(n_33892) );
oa22s01 g747773 ( .a(n_33372), .b(n_33576), .c(n_33571), .d(n_33415), .o(n_33862) );
oa12s01 g747774 ( .a(n_33293), .b(n_33571), .c(n_33279), .o(n_33841) );
oa22s01 g747775 ( .a(n_33372), .b(n_33316), .c(n_33571), .d(n_33310), .o(n_33912) );
oa22s01 g747776 ( .a(n_33571), .b(n_33240), .c(n_33372), .d(n_33256), .o(n_34071) );
in01s01 g747779 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_), .o(n_32276) );
in01s40 g747781 ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38778) );
no02s01 g747783 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_12_), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_13_), .o(n_32319) );
in01s01 g747784 ( .a(n_32260), .o(n_32261) );
na02s01 g747785 ( .a(n_31971), .b(n_32188), .o(n_32260) );
in01s01 g747786 ( .a(n_32111), .o(n_32112) );
na02s01 g747787 ( .a(n_32000), .b(n_31688), .o(n_32111) );
in01s01 g747788 ( .a(n_33970), .o(n_33971) );
no02s01 g747789 ( .a(n_33571), .b(n_33683), .o(n_33970) );
no02s01 g747790 ( .a(FE_OCP_RBN2532_n_33372), .b(n_33438), .o(n_33671) );
no02s01 g747791 ( .a(n_33372), .b(n_33336), .o(n_33884) );
in01s01 g747792 ( .a(n_33418), .o(n_33373) );
no02s01 g747793 ( .a(FE_OCP_RBN2505_n_33226), .b(n_33354), .o(n_33418) );
in01s01 g747794 ( .a(n_33653), .o(n_33599) );
na02s01 g747795 ( .a(FE_OCP_RBN2534_n_33372), .b(n_33573), .o(n_33653) );
in01s01 g747796 ( .a(n_33317), .o(n_33296) );
no02s02 g747797 ( .a(FE_OCP_RBN6561_n_33208), .b(n_33281), .o(n_33317) );
no02s02 g747798 ( .a(FE_OCP_RBN2505_n_33226), .b(n_32900), .o(n_33393) );
na02s01 g747799 ( .a(n_33372), .b(n_33370), .o(n_33702) );
no02s01 g747800 ( .a(n_33372), .b(n_32802), .o(n_33840) );
no02s01 g747801 ( .a(n_33372), .b(n_32901), .o(n_33421) );
no02s02 g747802 ( .a(n_33208), .b(n_32585), .o(n_33258) );
no02s02 g747803 ( .a(n_33191), .b(n_32584), .o(n_33242) );
no02s01 g747804 ( .a(n_33170), .b(FE_OCP_RBN2534_n_33372), .o(n_33990) );
in01s01 g747805 ( .a(n_33740), .o(n_33741) );
na02s01 g747806 ( .a(n_33571), .b(n_33651), .o(n_33740) );
no02s01 g747807 ( .a(n_33372), .b(n_33626), .o(n_33950) );
in01s01 g747808 ( .a(n_33624), .o(n_33625) );
na02s01 g747809 ( .a(n_33571), .b(n_33438), .o(n_33624) );
na02s01 g747810 ( .a(n_33512), .b(FE_OCP_RBN2532_n_33372), .o(n_33817) );
na02s01 g747811 ( .a(FE_OCP_RBN2505_n_33226), .b(n_33314), .o(n_33357) );
in01s01 g747812 ( .a(n_33413), .o(n_33414) );
na02s01 g747813 ( .a(FE_OCP_RBN2532_n_33372), .b(n_33441), .o(n_33413) );
no02s01 g747814 ( .a(n_33372), .b(n_33371), .o(n_33462) );
na02s06 TIMEBOOST_cell_1799 ( .a(n_30197), .b(n_30223), .o(TIMEBOOST_net_514) );
no02f06 TIMEBOOST_cell_4002 ( .a(n_4697), .b(TIMEBOOST_net_1091), .o(n_4851) );
in01s01 g747817 ( .a(n_33313), .o(n_33516) );
no02s01 g747818 ( .a(FE_OCP_RBN2503_n_33226), .b(n_33370), .o(n_33313) );
in01s01 g747819 ( .a(n_33311), .o(n_33312) );
no02s01 g747820 ( .a(FE_OCP_RBN2502_n_33226), .b(n_33294), .o(n_33311) );
in01s01 g747821 ( .a(n_33293), .o(n_33359) );
na02s01 g747822 ( .a(FE_OCP_RBN6561_n_33208), .b(n_33279), .o(n_33293) );
na02s01 g747823 ( .a(FE_OCP_RBN2502_n_33226), .b(n_33294), .o(n_33417) );
in01s01 g747824 ( .a(n_33495), .o(n_33496) );
na02s01 g747825 ( .a(FE_OCP_RBN2532_n_33372), .b(n_33437), .o(n_33495) );
in01s01 g747826 ( .a(n_33461), .o(n_33513) );
no02s02 g747827 ( .a(n_33437), .b(FE_OCP_RBN2532_n_33372), .o(n_33461) );
in01s01 g747828 ( .a(n_33390), .o(n_33440) );
na02s02 g747829 ( .a(n_33372), .b(n_33371), .o(n_33390) );
in01s01 g747830 ( .a(n_33601), .o(n_33572) );
na02s01 g747831 ( .a(FE_OCP_RBN2532_n_33372), .b(n_33354), .o(n_33601) );
na02s01 g747832 ( .a(FE_OCP_RBN2532_n_33372), .b(n_33554), .o(n_33600) );
in01s01 g747833 ( .a(n_33667), .o(n_33668) );
na02s01 g747834 ( .a(n_33571), .b(n_33511), .o(n_33667) );
in01s01 g747835 ( .a(n_33680), .o(n_33681) );
no02s01 g747836 ( .a(FE_OCP_RBN2534_n_33372), .b(n_33573), .o(n_33680) );
in01s01 g747837 ( .a(n_33738), .o(n_33739) );
na02s01 g747838 ( .a(n_33571), .b(n_33720), .o(n_33738) );
in01s01 g747839 ( .a(n_33701), .o(n_33532) );
no02s01 g747840 ( .a(FE_OCP_RBN2532_n_33372), .b(n_33511), .o(n_33701) );
in01s01 g747841 ( .a(n_33391), .o(n_33353) );
na02s01 g747842 ( .a(FE_OCP_RBN2506_n_33226), .b(n_33336), .o(n_33391) );
no02s01 g747843 ( .a(n_33571), .b(n_33651), .o(n_33792) );
no02m20 g747845 ( .a(n_32188), .b(n_31970), .o(n_32238) );
oa12s01 g747848 ( .a(n_31611), .b(n_32003), .c(n_31605), .o(n_32061) );
oa22s01 g747849 ( .a(n_32187), .b(n_32211), .c(n_32186), .d(n_32210), .o(n_32259) );
in01s01 g747850 ( .a(n_32236), .o(n_32237) );
oa12s01 g747851 ( .a(n_32104), .b(n_32189), .c(n_31903), .o(n_32236) );
in01s01 g747852 ( .a(n_33762), .o(n_33239) );
ao12s01 g747853 ( .a(n_33194), .b(n_33193), .c(n_33192), .o(n_33762) );
ao12s01 g747854 ( .a(n_33132), .b(n_33131), .c(n_33130), .o(n_33684) );
oa12s01 g747855 ( .a(FE_OCP_RBN2532_n_33372), .b(n_33552), .c(n_33027), .o(n_33553) );
in01s01 g747856 ( .a(n_33334), .o(n_33335) );
oa12s01 g747857 ( .a(FE_OCP_RBN2505_n_33226), .b(n_33310), .c(n_33281), .o(n_33334) );
oa12s02 g747858 ( .a(n_33372), .b(n_32777), .c(n_33370), .o(n_33579) );
in01s01 g747859 ( .a(n_33227), .o(n_33670) );
ao12s01 g747860 ( .a(n_33173), .b(n_33172), .c(n_33171), .o(n_33227) );
oa12s01 g747861 ( .a(n_33129), .b(n_33128), .c(n_33127), .o(n_33743) );
in01s01 g747862 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_13_), .o(n_32083) );
in01s01 g747865 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_14_), .o(n_32275) );
no02s01 g747868 ( .a(n_33193), .b(n_33192), .o(n_33194) );
no02s01 g747869 ( .a(n_33131), .b(n_33130), .o(n_33132) );
no02s01 g747870 ( .a(n_33172), .b(n_33171), .o(n_33173) );
na02s01 g747871 ( .a(n_33128), .b(n_33127), .o(n_33129) );
na02s01 g747873 ( .a(n_32189), .b(n_31861), .o(n_32216) );
in01s01 g747874 ( .a(n_32032), .o(n_32033) );
na02s01 g747875 ( .a(n_32003), .b(n_31548), .o(n_32032) );
in01s01 g747876 ( .a(n_32214), .o(n_32215) );
oa12s02 g747877 ( .a(n_32138), .b(n_32110), .c(FE_OCP_RBN3409_n_32072), .o(n_32214) );
na02f20 g747881 ( .a(n_32142), .b(n_31932), .o(n_32188) );
in01s01 g747882 ( .a(n_32001), .o(n_32002) );
ao12s01 g747883 ( .a(n_31794), .b(n_31938), .c(n_31862), .o(n_32001) );
oa22s01 g747888 ( .a(n_31884), .b(FE_OCP_RBN6187_n_31916), .c(n_31883), .d(n_31916), .o(n_31999) );
oa22s01 g747889 ( .a(n_31938), .b(n_31895), .c(n_31956), .d(n_31896), .o(n_32029) );
oa22s01 g747890 ( .a(n_32109), .b(n_32161), .c(n_32110), .d(n_32162), .o(n_32235) );
oa12s01 g747891 ( .a(n_33126), .b(n_33125), .c(n_33124), .o(n_33626) );
ao12s01 g747892 ( .a(n_33120), .b(n_33119), .c(n_33118), .o(n_33651) );
in01s03 g747923 ( .a(FE_OCP_RBN2534_n_33372), .o(n_33571) );
in01s06 g747935 ( .a(FE_OCP_RBN2505_n_33226), .o(n_33372) );
in01s04 g747943 ( .a(n_33191), .o(n_33208) );
in01s01 g747945 ( .a(n_33683), .o(n_33170) );
ao12s01 g747946 ( .a(n_33093), .b(n_33092), .c(n_33091), .o(n_33683) );
in01s01 g747947 ( .a(n_33169), .o(n_33554) );
oa12s01 g747948 ( .a(n_33090), .b(n_33089), .c(n_33088), .o(n_33169) );
ao12s01 g747949 ( .a(n_33117), .b(n_33116), .c(n_33115), .o(n_33511) );
ao12s01 g747950 ( .a(n_33123), .b(n_33122), .c(n_33121), .o(n_33720) );
no02s01 g747951 ( .a(n_33092), .b(n_33091), .o(n_33093) );
na02s01 g747952 ( .a(n_33125), .b(n_33124), .o(n_33126) );
na02s01 g747953 ( .a(n_33089), .b(n_33088), .o(n_33090) );
no02s01 g747954 ( .a(n_33122), .b(n_33121), .o(n_33123) );
no02f08 TIMEBOOST_cell_3992 ( .a(TIMEBOOST_net_1086), .b(n_38785), .o(n_38806) );
no02s01 g747956 ( .a(n_33119), .b(n_33118), .o(n_33120) );
no02s01 g747957 ( .a(n_33116), .b(n_33115), .o(n_33117) );
in01s01 g747958 ( .a(n_32142), .o(n_32189) );
in01s01 g747960 ( .a(n_31959), .o(n_32003) );
no02f20 g747961 ( .a(n_31593), .b(n_31908), .o(n_31959) );
no02f08 TIMEBOOST_cell_1686 ( .a(n_26007), .b(TIMEBOOST_net_457), .o(n_26163) );
ao12s01 g747963 ( .a(n_32646), .b(n_33041), .c(n_32555), .o(n_33172) );
ao12s01 g747964 ( .a(n_32724), .b(n_33029), .c(n_32490), .o(n_33128) );
ao12s01 g747965 ( .a(n_32776), .b(n_33048), .c(n_32452), .o(n_33131) );
in01s01 g747966 ( .a(n_32186), .o(n_32187) );
ao12s02 g747967 ( .a(n_31848), .b(n_32139), .c(n_32060), .o(n_32186) );
oa22s01 g747968 ( .a(n_31914), .b(n_31937), .c(n_31936), .d(n_31915), .o(n_31998) );
oa22s01 g747969 ( .a(n_31881), .b(n_31608), .c(n_31882), .d(n_31609), .o(n_31958) );
oa22s01 g747970 ( .a(n_32184), .b(n_32182), .c(n_32185), .d(n_32183), .o(n_32252) );
oa22s01 g747971 ( .a(n_32079), .b(n_32163), .c(n_32060), .d(n_32164), .o(n_32234) );
ao12s01 g747972 ( .a(n_33086), .b(n_33085), .c(n_33084), .o(n_33354) );
ao12s01 g747973 ( .a(n_33044), .b(n_33043), .c(n_33042), .o(n_33438) );
in01s01 g747974 ( .a(n_33552), .o(n_33114) );
ao12s01 g747975 ( .a(n_33047), .b(n_33046), .c(n_33045), .o(n_33552) );
oa12s01 g747976 ( .a(n_33071), .b(n_33070), .c(n_33069), .o(n_33573) );
in01s01 g747977 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_12_), .o(n_32082) );
no02s01 g747980 ( .a(n_33048), .b(n_33146), .o(n_33092) );
no02s01 g747981 ( .a(n_33046), .b(n_33045), .o(n_33047) );
na02s01 g747982 ( .a(n_33030), .b(n_32723), .o(n_33119) );
na02s01 g747983 ( .a(n_33040), .b(n_32645), .o(n_33116) );
no02s01 g747984 ( .a(n_33085), .b(n_33084), .o(n_33086) );
in01s01 g747985 ( .a(n_31883), .o(n_31884) );
ao12s01 g747986 ( .a(n_31560), .b(n_31813), .c(n_31613), .o(n_31883) );
in01s01 g747987 ( .a(n_33072), .o(n_33073) );
na02s06 g747988 ( .a(n_33048), .b(n_32563), .o(n_33072) );
no02s01 g747989 ( .a(n_33043), .b(n_33042), .o(n_33044) );
na02s01 g747990 ( .a(n_33070), .b(n_33069), .o(n_33071) );
ao12s01 g747991 ( .a(n_32456), .b(n_33000), .c(n_32487), .o(n_33089) );
in01s01 g747994 ( .a(n_32109), .o(n_32110) );
in01s01 g747995 ( .a(n_32081), .o(n_32109) );
na02s10 TIMEBOOST_cell_1336 ( .a(n_24072), .b(TIMEBOOST_net_282), .o(n_24147) );
in01s01 g747998 ( .a(n_31938), .o(n_31956) );
in01s01 g747999 ( .a(n_31908), .o(n_31938) );
na03f40 TIMEBOOST_cell_7432 ( .a(FE_OCP_RBN5507_n_44061), .b(FE_OCP_RBN2271_delay_xor_ln22_unr15_stage6_stallmux_q_5_), .c(FE_OCP_RBN6530_n_22822), .o(TIMEBOOST_net_2347) );
no02s02 TIMEBOOST_cell_1673 ( .a(n_34768), .b(n_34396), .o(TIMEBOOST_net_451) );
no03s08 TIMEBOOST_cell_2150 ( .a(n_17054), .b(n_16503), .c(n_17158), .o(n_17713) );
na02s01 TIMEBOOST_cell_7847 ( .a(TIMEBOOST_net_2554), .b(FE_OCP_RBN4359_n_10100), .o(n_10521) );
no02s01 g748004 ( .a(n_33004), .b(n_32489), .o(n_33005) );
in01s01 g748005 ( .a(n_33029), .o(n_33030) );
no02s01 g748006 ( .a(n_33004), .b(n_32506), .o(n_33029) );
na02s01 g748007 ( .a(n_33003), .b(n_32605), .o(n_33043) );
in01s01 g748008 ( .a(n_33040), .o(n_33041) );
na02s01 g748009 ( .a(n_32982), .b(n_32556), .o(n_33040) );
no02s01 g748010 ( .a(n_32981), .b(n_33028), .o(n_33070) );
na02s01 g748011 ( .a(n_33001), .b(n_32455), .o(n_33085) );
in01s01 g748013 ( .a(n_32060), .o(n_32079) );
no02s02 g748014 ( .a(n_31975), .b(n_31837), .o(n_32060) );
no02s06 g748015 ( .a(n_33004), .b(n_32560), .o(n_33048) );
oa12s01 g748016 ( .a(n_32485), .b(n_44347), .c(n_32414), .o(n_33046) );
na02s08 TIMEBOOST_cell_1335 ( .a(n_23665), .b(n_23707), .o(TIMEBOOST_net_282) );
in01s01 g748018 ( .a(n_32184), .o(n_32185) );
oa12s01 g748019 ( .a(n_32075), .b(n_31954), .c(n_32077), .o(n_32184) );
in01s01 g748020 ( .a(n_31936), .o(n_31937) );
ao12s01 g748021 ( .a(n_31823), .b(n_31777), .c(n_31897), .o(n_31936) );
in01s01 g748022 ( .a(n_31881), .o(n_31882) );
oa12s01 g748023 ( .a(n_31751), .b(n_31777), .c(n_31612), .o(n_31881) );
no02m08 TIMEBOOST_cell_5197 ( .a(TIMEBOOST_net_1546), .b(n_14608), .o(n_14770) );
oa22s01 g748025 ( .a(n_31777), .b(n_31919), .c(n_31748), .d(n_31920), .o(n_31996) );
oa22s01 g748026 ( .a(n_32178), .b(n_31972), .c(n_31954), .d(FE_OCP_RBN6226_n_32178), .o(n_32251) );
in01s01 g748027 ( .a(n_33336), .o(n_33027) );
oa22s01 g748028 ( .a(n_44346), .b(n_32530), .c(n_44347), .d(n_32531), .o(n_33336) );
in01s01 g748029 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_11_), .o(n_31855) );
in01s01 g748032 ( .a(n_33003), .o(n_32982) );
na02s01 g748033 ( .a(n_32535), .b(n_44346), .o(n_33003) );
in01s01 g748034 ( .a(n_33000), .o(n_33001) );
no02s01 g748035 ( .a(n_44347), .b(n_32502), .o(n_33000) );
na02m08 g748036 ( .a(n_32107), .b(n_32024), .o(n_32108) );
na02f10 g748037 ( .a(n_31708), .b(n_31751), .o(n_31813) );
in01s01 g748038 ( .a(n_31974), .o(n_31975) );
na02f10 g748039 ( .a(n_31935), .b(n_31766), .o(n_31974) );
na02s06 g748040 ( .a(n_32107), .b(n_31969), .o(n_32106) );
in01s01 g748041 ( .a(n_33004), .o(n_32981) );
na02s06 g748042 ( .a(n_32966), .b(n_32607), .o(n_33004) );
no02s01 TIMEBOOST_cell_3963 ( .a(FE_OCP_RBN5714_n_44102), .b(n_33975), .o(TIMEBOOST_net_1072) );
no02s10 g748045 ( .a(n_32086), .b(n_31653), .o(n_31880) );
no02s08 g748046 ( .a(n_32086), .b(n_31744), .o(n_31879) );
no02s01 TIMEBOOST_cell_1174 ( .a(n_28592), .b(TIMEBOOST_net_201), .o(n_28693) );
oa22s01 g748048 ( .a(n_31668), .b(n_31556), .c(n_31669), .d(n_31557), .o(n_31750) );
in01s01 g748052 ( .a(n_31748), .o(n_31777) );
in01s01 g748053 ( .a(n_31708), .o(n_31748) );
ao12f08 g748054 ( .a(n_31499), .b(n_31614), .c(n_31521), .o(n_31708) );
oa22s01 g748055 ( .a(n_31876), .b(n_31838), .c(n_31877), .d(n_31839), .o(n_31955) );
in01s01 g748057 ( .a(n_31954), .o(n_31972) );
in01s01 g748058 ( .a(n_31935), .o(n_31954) );
ao12f08 g748059 ( .a(n_31754), .b(n_31853), .c(n_31799), .o(n_31935) );
ao12s01 g748060 ( .a(n_32883), .b(n_32882), .c(n_32881), .o(n_33512) );
in01s01 g748062 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_10_), .o(n_32861) );
no02s01 g748064 ( .a(n_32882), .b(n_32881), .o(n_32883) );
no02m06 g748065 ( .a(n_31994), .b(n_31966), .o(n_32028) );
na02s20 g748066 ( .a(n_31666), .b(n_31810), .o(n_32086) );
in01m08 g748067 ( .a(n_32026), .o(n_32027) );
no02s01 TIMEBOOST_cell_8576 ( .a(n_21778), .b(n_21779), .o(TIMEBOOST_net_2775) );
in01s01 g748071 ( .a(n_33314), .o(n_32902) );
ao12s01 g748072 ( .a(n_32842), .b(n_32841), .c(n_32840), .o(n_33314) );
ao12s01 g748073 ( .a(n_32866), .b(n_32865), .c(n_32864), .o(n_33441) );
na02f04 TIMEBOOST_cell_1706 ( .a(TIMEBOOST_net_467), .b(n_15392), .o(n_45501) );
na02s01 g748075 ( .a(n_32843), .b(n_32781), .o(n_32882) );
no02s01 g748076 ( .a(n_32841), .b(n_32840), .o(n_32842) );
no02s01 g748077 ( .a(n_32865), .b(n_32864), .o(n_32866) );
no02s03 g748078 ( .a(n_31746), .b(n_31735), .o(n_31747) );
no02s20 g748079 ( .a(n_31746), .b(n_31687), .o(n_31810) );
na02s02 g748080 ( .a(n_31745), .b(n_31776), .o(n_31854) );
na02f06 g748081 ( .a(n_31875), .b(n_31836), .o(n_31934) );
in01s02 g748083 ( .a(n_31971), .o(n_31994) );
na02s01 TIMEBOOST_cell_8779 ( .a(TIMEBOOST_net_2876), .b(n_11211), .o(n_11261) );
no02s06 g748086 ( .a(n_31968), .b(n_31951), .o(n_32024) );
ao12s04 g748087 ( .a(n_32628), .b(n_32809), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_15_), .o(n_32826) );
oa22s01 g748089 ( .a(n_31550), .b(n_31525), .c(n_31551), .d(n_31524), .o(n_31670) );
in01s01 g748090 ( .a(n_31668), .o(n_31669) );
in01s01 g748091 ( .a(n_31614), .o(n_31668) );
ao12f08 g748092 ( .a(n_31468), .b(n_31506), .c(n_31519), .o(n_31614) );
oa22s01 g748093 ( .a(n_31785), .b(n_31774), .c(n_31784), .d(n_31775), .o(n_31878) );
in01s01 g748094 ( .a(n_31876), .o(n_31877) );
in01s01 g748095 ( .a(n_31853), .o(n_31876) );
ao12f08 g748096 ( .a(n_31698), .b(n_31742), .c(n_31756), .o(n_31853) );
in01s01 g748097 ( .a(n_32900), .o(n_32901) );
ao12s01 g748098 ( .a(n_32839), .b(n_32838), .c(n_32837), .o(n_32900) );
in01s01 g748099 ( .a(n_33310), .o(n_33316) );
ao12s01 g748100 ( .a(n_32808), .b(n_32807), .c(n_32806), .o(n_33310) );
oa12s01 g748101 ( .a(n_32825), .b(n_32824), .c(n_32823), .o(n_33371) );
ao12s01 g748102 ( .a(n_32805), .b(n_32804), .c(n_32803), .o(n_33437) );
in01s01 g748103 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_9_), .o(n_32989) );
no02s06 g748106 ( .a(n_32809), .b(n_32421), .o(n_32843) );
no02s01 g748107 ( .a(n_32807), .b(n_32806), .o(n_32808) );
no02s01 g748108 ( .a(n_32804), .b(n_32803), .o(n_32805) );
no02s01 g748109 ( .a(n_32838), .b(n_32837), .o(n_32839) );
na02f08 g748111 ( .a(n_31563), .b(n_31549), .o(n_31667) );
in01s01 g748112 ( .a(n_31746), .o(n_31688) );
in01s01 g748114 ( .a(n_31744), .o(n_31745) );
oa12s04 g748115 ( .a(n_31652), .b(FE_OCPN943_n_31466), .c(n_31606), .o(n_31744) );
na02s01 g748116 ( .a(n_32824), .b(n_32823), .o(n_32825) );
ao12s01 g748117 ( .a(n_32458), .b(n_32778), .c(n_32484), .o(n_32841) );
na02m10 g748120 ( .a(n_31930), .b(n_31948), .o(n_31970) );
na02f04 g748121 ( .a(n_31807), .b(n_31783), .o(n_31875) );
na02s10 TIMEBOOST_cell_6589 ( .a(FE_OCP_RBN3965_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(FE_RN_198_0), .o(TIMEBOOST_net_2052) );
no02s01 TIMEBOOST_cell_1173 ( .a(n_28176), .b(n_28055), .o(TIMEBOOST_net_201) );
in01s02 g748125 ( .a(n_31968), .o(n_31969) );
na02s02 TIMEBOOST_cell_5648 ( .a(n_6215), .b(n_6332), .o(TIMEBOOST_net_1772) );
no02m04 TIMEBOOST_cell_4049 ( .a(n_24895), .b(n_24751), .o(TIMEBOOST_net_1115) );
na02s02 g748129 ( .a(n_31743), .b(n_31808), .o(n_31809) );
no02s01 TIMEBOOST_cell_1613 ( .a(n_2760), .b(n_2875), .o(TIMEBOOST_net_421) );
no02s06 g748131 ( .a(n_32782), .b(n_32418), .o(n_32809) );
no02s01 g748132 ( .a(n_32768), .b(n_32603), .o(n_32783) );
na02s01 g748133 ( .a(n_32782), .b(n_32781), .o(n_32804) );
no02s01 g748134 ( .a(n_32769), .b(n_32796), .o(n_32824) );
na02s01 g748135 ( .a(n_32779), .b(n_32586), .o(n_32838) );
na02m06 g748136 ( .a(n_31805), .b(n_31851), .o(n_31852) );
no02s01 g748137 ( .a(n_31953), .b(n_32103), .o(n_32104) );
no02s20 g748138 ( .a(n_31903), .b(n_31872), .o(n_31932) );
in01f08 g748139 ( .a(n_31948), .o(n_31949) );
no02m10 g748140 ( .a(n_31902), .b(n_31931), .o(n_31948) );
no02m06 g748141 ( .a(n_31929), .b(n_31868), .o(n_31930) );
in01s01 g748142 ( .a(n_31990), .o(n_31991) );
no02s06 g748143 ( .a(n_47271), .b(n_31967), .o(n_31990) );
in01s01 g748144 ( .a(n_32163), .o(n_32164) );
na02s01 g748145 ( .a(n_31805), .b(n_32139), .o(n_32163) );
no02f02 TIMEBOOST_cell_5312 ( .a(n_20271), .b(n_20236), .o(TIMEBOOST_net_1604) );
in01s01 g748147 ( .a(n_32161), .o(n_32162) );
na02s01 g748148 ( .a(n_32138), .b(n_32072), .o(n_32161) );
in01s01 g748149 ( .a(n_32136), .o(n_32137) );
no02s01 g748150 ( .a(n_31903), .b(n_32103), .o(n_32136) );
in01s01 g748151 ( .a(n_31988), .o(n_31989) );
no02s01 g748152 ( .a(n_31902), .b(n_31966), .o(n_31988) );
no02m02 TIMEBOOST_cell_8552 ( .a(n_8127), .b(n_46991), .o(TIMEBOOST_net_2763) );
in01s02 g748155 ( .a(n_32101), .o(n_32102) );
no02s02 g748156 ( .a(n_31869), .b(n_32055), .o(n_32101) );
na02s03 TIMEBOOST_cell_4560 ( .a(n_32279), .b(TIMEBOOST_net_1370), .o(FE_RN_2698_0) );
in01s02 g748158 ( .a(n_32099), .o(n_32100) );
no02s03 g748159 ( .a(n_32326), .b(n_32020), .o(n_32099) );
na02s01 TIMEBOOST_cell_1162 ( .a(TIMEBOOST_net_195), .b(n_37730), .o(n_37731) );
in01s01 g748161 ( .a(n_32057), .o(n_32058) );
no02s01 g748162 ( .a(n_31947), .b(n_31863), .o(n_32057) );
in01s01 g748163 ( .a(n_32134), .o(n_32135) );
no02s02 g748164 ( .a(n_47271), .b(n_47272), .o(n_32134) );
no02f06 TIMEBOOST_cell_8846 ( .a(n_30200), .b(n_30508), .o(TIMEBOOST_net_2910) );
no02s06 TIMEBOOST_cell_1484 ( .a(TIMEBOOST_net_356), .b(n_2855), .o(n_3626) );
oa12s01 g748168 ( .a(n_32403), .b(n_32780), .c(n_32483), .o(n_32807) );
in01s01 g748169 ( .a(n_32210), .o(n_32211) );
na02s01 g748170 ( .a(n_32119), .b(n_31851), .o(n_32210) );
in01s01 g748171 ( .a(n_32208), .o(n_32209) );
no02s01 g748172 ( .a(n_32098), .b(n_32118), .o(n_32208) );
in01s02 g748173 ( .a(n_32132), .o(n_32133) );
no02s01 TIMEBOOST_cell_4007 ( .a(n_30614), .b(n_30633), .o(TIMEBOOST_net_1094) );
na03f04 TIMEBOOST_cell_7247 ( .a(n_19636), .b(FE_OCP_RBN5665_n_19101), .c(n_19672), .o(n_19808) );
in01s01 g748177 ( .a(n_32128), .o(n_32129) );
no02s01 TIMEBOOST_cell_3394 ( .a(n_36066), .b(n_36063), .o(TIMEBOOST_net_988) );
in01s01 g748179 ( .a(n_32126), .o(n_32127) );
no02s01 g748180 ( .a(n_31967), .b(n_32046), .o(n_32126) );
in01s01 g748181 ( .a(n_32124), .o(n_32125) );
na02s02 TIMEBOOST_cell_4565 ( .a(n_40532), .b(n_40221), .o(TIMEBOOST_net_1373) );
no02s06 g748183 ( .a(n_31684), .b(n_31704), .o(n_31808) );
na03m06 TIMEBOOST_cell_8318 ( .a(FE_RN_1912_0), .b(FE_RN_1913_0), .c(n_4095), .o(n_47009) );
no02s06 g748187 ( .a(n_31607), .b(FE_OCPN943_n_31466), .o(n_31687) );
na02s10 g748188 ( .a(n_31520), .b(n_31558), .o(n_31666) );
na02s01 g748189 ( .a(n_31730), .b(n_31705), .o(n_31776) );
in01s01 g748190 ( .a(n_31524), .o(n_31525) );
in01s01 g748191 ( .a(n_31506), .o(n_31524) );
oa12f08 g748192 ( .a(n_31467), .b(n_31447), .c(n_31424), .o(n_31506) );
oa22s01 g748193 ( .a(n_31497), .b(n_31471), .c(n_31498), .d(n_31472), .o(n_31561) );
in01s01 g748194 ( .a(n_31774), .o(n_31775) );
in01s01 g748195 ( .a(n_31742), .o(n_31774) );
ao12f08 g748196 ( .a(n_31648), .b(n_31678), .c(n_31697), .o(n_31742) );
in01s01 g748197 ( .a(n_32182), .o(n_32183) );
oa22s01 g748198 ( .a(FE_OCP_RBN6880_n_31819), .b(n_30299), .c(FE_OCP_RBN6881_n_31819), .d(n_30327), .o(n_32182) );
oa22s01 g748200 ( .a(FE_OCP_RBN6879_n_31819), .b(n_30573), .c(FE_OCP_RBN3414_FE_OCPN891_n_31944), .d(n_30593), .o(n_32180) );
in01s01 g748201 ( .a(n_32122), .o(n_32123) );
in01s01 TIMEBOOST_cell_4567 ( .a(TIMEBOOST_net_1374), .o(state_cordic_1_) );
oa22s01 g748203 ( .a(n_31713), .b(n_31700), .c(n_31714), .d(n_31701), .o(n_31806) );
in01s01 g748204 ( .a(n_33281), .o(n_32802) );
ao12s01 g748205 ( .a(n_32764), .b(n_32780), .c(n_32763), .o(n_33281) );
oa12s01 g748206 ( .a(n_32767), .b(n_32766), .c(n_32765), .o(n_33294) );
oa22s01 g748208 ( .a(FE_OCP_RBN6880_n_31819), .b(n_32076), .c(FE_OCP_RBN6881_n_31819), .d(n_30326), .o(n_32178) );
no02s01 TIMEBOOST_cell_7033 ( .a(FE_OCP_RBN2921_n_3878), .b(n_4316), .o(TIMEBOOST_net_2275) );
in01s01 g748212 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_8_), .o(n_32793) );
in01s01 g748214 ( .a(n_32768), .o(n_32769) );
na02s01 g748215 ( .a(n_32750), .b(n_32533), .o(n_32768) );
in01s01 g748216 ( .a(n_32778), .o(n_32779) );
no02s01 g748217 ( .a(n_32780), .b(n_32501), .o(n_32778) );
na02s01 g748218 ( .a(n_32766), .b(n_32765), .o(n_32767) );
no02s01 g748219 ( .a(n_32780), .b(n_32763), .o(n_32764) );
no02s01 g748220 ( .a(FE_OCP_RBN6880_n_31819), .b(n_32076), .o(n_32077) );
na02s01 g748221 ( .a(FE_OCP_RBN6880_n_31819), .b(n_32076), .o(n_32075) );
na03m02 TIMEBOOST_cell_2501 ( .a(n_3169), .b(n_3167), .c(TIMEBOOST_net_408), .o(n_3272) );
na02s01 g748223 ( .a(FE_OCP_RBN6880_n_31819), .b(n_31740), .o(n_32139) );
in01s01 g748225 ( .a(n_31805), .o(n_31848) );
na02s01 g748227 ( .a(FE_OCP_RBN6879_n_31819), .b(n_30522), .o(n_32119) );
na02s04 g748228 ( .a(n_31765), .b(FE_OCPN1276_n_31773), .o(n_31851) );
na02s01 g748229 ( .a(FE_OCP_RBN6879_n_31819), .b(FE_RN_1883_0), .o(n_32138) );
na02s01 g748231 ( .a(FE_OCP_RBN6203_n_31819), .b(n_30592), .o(n_32072) );
na02f04 TIMEBOOST_cell_7773 ( .a(TIMEBOOST_net_2517), .b(n_10325), .o(n_10483) );
no02s01 g748233 ( .a(FE_OCP_RBN6203_n_31819), .b(n_31770), .o(n_32103) );
no02s10 g748237 ( .a(FE_OCP_RBN3388_n_31819), .b(n_30426), .o(n_31903) );
no02s01 g748238 ( .a(FE_OCP_RBN3413_FE_OCPN891_n_31944), .b(n_30554), .o(n_32098) );
no02s10 g748239 ( .a(FE_OCP_RBN3388_n_31819), .b(FE_OCPN5254_n_31871), .o(n_31872) );
no02s01 g748240 ( .a(FE_OCP_RBN6879_n_31819), .b(FE_OCPN5254_n_31871), .o(n_32118) );
in01s01 g748241 ( .a(n_31847), .o(n_31966) );
na02s03 g748242 ( .a(n_31783), .b(FE_OCPN5107_n_31804), .o(n_31847) );
no02s06 g748246 ( .a(FE_OCP_RBN3388_n_31819), .b(FE_OCPN5107_n_31804), .o(n_31902) );
na02f08 TIMEBOOST_cell_4006 ( .a(TIMEBOOST_net_1093), .b(n_35034), .o(n_35145) );
no02s06 g748248 ( .a(FE_OCP_RBN3388_n_31819), .b(n_44437), .o(n_31931) );
no02s06 g748252 ( .a(FE_OCP_RBN2105_n_30465), .b(n_31835), .o(n_31869) );
in01s01 g748254 ( .a(n_32055), .o(n_32070) );
no02m01 g748255 ( .a(n_31783), .b(n_30465), .o(n_31868) );
no02s02 g748256 ( .a(FE_OCP_RBN3388_n_31819), .b(n_30465), .o(n_32055) );
na02m04 TIMEBOOST_cell_1165 ( .a(FE_OCP_RBN4034_n_37690), .b(n_37622), .o(TIMEBOOST_net_197) );
no02s06 g748258 ( .a(FE_OCP_RBN3388_n_31819), .b(n_31864), .o(n_31929) );
in01s01 g748260 ( .a(n_32020), .o(n_32052) );
na02s01 TIMEBOOST_cell_1161 ( .a(n_37614), .b(n_37539), .o(TIMEBOOST_net_195) );
no02s06 g748262 ( .a(FE_OCP_RBN6203_n_31819), .b(FE_OCP_RBN6001_n_30534), .o(n_32020) );
no02m03 g748263 ( .a(FE_OCP_RBN6879_n_31819), .b(n_30557), .o(n_32326) );
no02m04 TIMEBOOST_cell_6384 ( .a(TIMEBOOST_net_2043), .b(n_26020), .o(TIMEBOOST_net_1745) );
na02s02 g748265 ( .a(FE_OCPN6901_FE_OCP_RBN4472_n_31819), .b(FE_OCP_RBN6812_n_30608), .o(n_32051) );
in01s01 g748267 ( .a(n_31863), .o(n_31898) );
no02s02 g748268 ( .a(n_31835), .b(FE_OCP_RBN6022_n_46959), .o(n_31863) );
no02s06 g748272 ( .a(FE_OCP_RBN3391_n_31819), .b(FE_OCP_RBN6021_n_46959), .o(n_31947) );
na02s01 TIMEBOOST_cell_3393 ( .a(n_36445), .b(TIMEBOOST_net_987), .o(n_36490) );
no02s06 g748274 ( .a(FE_OCP_RBN3391_n_31819), .b(FE_OCP_RBN6024_n_30711), .o(n_31992) );
in01s01 g748278 ( .a(n_47271), .o(n_32068) );
no02s01 g748281 ( .a(FE_OCP_RBN4472_n_31819), .b(n_46957), .o(n_32046) );
no02m01 g748282 ( .a(FE_OCP_RBN3391_n_31819), .b(FE_OCP_RBN6055_n_46957), .o(n_31967) );
na02f06 TIMEBOOST_cell_4564 ( .a(TIMEBOOST_net_1372), .b(n_36521), .o(n_36583) );
na02m06 TIMEBOOST_cell_4566 ( .a(TIMEBOOST_net_1373), .b(n_40555), .o(n_40579) );
na02s01 g748287 ( .a(FE_OCP_RBN4472_n_31819), .b(FE_OCP_RBN6084_n_31010), .o(n_32044) );
no02s01 g748288 ( .a(n_31612), .b(n_31559), .o(n_31613) );
na02s06 g748289 ( .a(n_31522), .b(n_31501), .o(n_31523) );
no02s01 g748290 ( .a(n_31591), .b(n_31610), .o(n_31611) );
in01m06 g748292 ( .a(n_31685), .o(n_31686) );
na02f06 TIMEBOOST_cell_1462 ( .a(n_24754), .b(TIMEBOOST_net_345), .o(n_24829) );
na02f04 TIMEBOOST_cell_5643 ( .a(TIMEBOOST_net_1769), .b(n_6156), .o(n_6267) );
in01s02 g748297 ( .a(n_31706), .o(n_31738) );
na02s06 g748298 ( .a(n_31681), .b(n_31682), .o(n_31706) );
in01s01 g748299 ( .a(n_31919), .o(n_31920) );
na02s01 g748300 ( .a(n_31824), .b(n_31897), .o(n_31919) );
in01s01 g748301 ( .a(n_31608), .o(n_31609) );
no02s01 g748302 ( .a(n_31560), .b(n_31559), .o(n_31608) );
na02s04 TIMEBOOST_cell_5645 ( .a(TIMEBOOST_net_1770), .b(n_6208), .o(n_6313) );
in01s01 g748304 ( .a(n_31895), .o(n_31896) );
na02s01 g748305 ( .a(n_31793), .b(n_31862), .o(n_31895) );
in01s01 g748306 ( .a(n_31736), .o(n_31737) );
no02s01 g748307 ( .a(n_31605), .b(n_31610), .o(n_31736) );
in01s01 g748309 ( .a(n_31768), .o(n_31769) );
no02s01 g748310 ( .a(n_31554), .b(n_31735), .o(n_31768) );
in01s01 g748311 ( .a(n_31802), .o(n_31803) );
no02s06 g748312 ( .a(n_31763), .b(n_32168), .o(n_31802) );
na02f06 TIMEBOOST_cell_1456 ( .a(TIMEBOOST_net_342), .b(n_29481), .o(n_29532) );
in01m02 g748314 ( .a(n_31842), .o(n_31843) );
no02m02 g748315 ( .a(n_31787), .b(n_32149), .o(n_31842) );
na02s06 g748316 ( .a(n_31553), .b(n_30757), .o(n_31558) );
in01s02 g748317 ( .a(n_31800), .o(n_31801) );
no02m02 g748318 ( .a(FE_OCPN3586_n_31704), .b(n_31594), .o(n_31800) );
no02s02 g748319 ( .a(n_31594), .b(FE_OCP_RBN3141_n_30849), .o(n_31606) );
in01s01 g748320 ( .a(n_31840), .o(n_31841) );
no02s02 g748321 ( .a(n_32197), .b(n_31703), .o(n_31840) );
na02s01 g748322 ( .a(n_31702), .b(FE_OCPN908_n_46956), .o(n_31705) );
in01s01 g748323 ( .a(n_31556), .o(n_31557) );
na02s01 g748324 ( .a(n_31521), .b(n_31500), .o(n_31556) );
in01s01 g748325 ( .a(n_31838), .o(n_31839) );
na02s01 g748326 ( .a(n_31755), .b(n_31799), .o(n_31838) );
na02s06 g748327 ( .a(n_32750), .b(n_32604), .o(n_32782) );
na02s04 g748328 ( .a(n_31765), .b(n_30300), .o(n_31766) );
in01s01 g748329 ( .a(n_31836), .o(n_31837) );
in01s01 g748331 ( .a(n_31953), .o(n_31861) );
oa12s01 g748338 ( .a(n_31522), .b(FE_OCP_RBN6874_n_31520), .c(FE_OCP_DRV_N3516_n_31504), .o(n_31916) );
in01s01 g748339 ( .a(n_31893), .o(n_31894) );
no02s01 g748340 ( .a(n_31664), .b(n_31791), .o(n_31893) );
in01s02 g748341 ( .a(n_31833), .o(n_31834) );
na02s01 TIMEBOOST_cell_6110 ( .a(TIMEBOOST_net_1906), .b(n_42522), .o(n_42563) );
in01s02 g748343 ( .a(n_31831), .o(n_31832) );
no02s02 TIMEBOOST_cell_1482 ( .a(n_42105), .b(TIMEBOOST_net_355), .o(n_42145) );
in01s01 g748345 ( .a(n_31829), .o(n_31830) );
na02s02 g748346 ( .a(n_31759), .b(n_31725), .o(n_31829) );
in01s01 g748347 ( .a(n_31796), .o(n_31797) );
na02s03 TIMEBOOST_cell_8743 ( .a(TIMEBOOST_net_2858), .b(n_41792), .o(n_41816) );
in01s01 g748349 ( .a(n_31858), .o(n_31859) );
na02s02 TIMEBOOST_cell_1486 ( .a(TIMEBOOST_net_357), .b(n_24653), .o(n_46963) );
in01s01 g748351 ( .a(n_31914), .o(n_31915) );
oa22s01 g748352 ( .a(FE_OCP_RBN6874_n_31520), .b(n_30350), .c(FE_OCP_RBN6872_n_31520), .d(n_30324), .o(n_31914) );
in01s01 g748353 ( .a(n_31912), .o(n_31913) );
oa22s01 g748354 ( .a(FE_OCP_RBN6875_n_31520), .b(n_30527), .c(FE_OCP_RBN6872_n_31520), .d(n_30506), .o(n_31912) );
in01s01 g748355 ( .a(n_31827), .o(n_31828) );
na03f08 TIMEBOOST_cell_6480 ( .a(n_24181), .b(FE_RN_85_0), .c(FE_OFN743_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_RN_86_0) );
in01s01 g748357 ( .a(n_33279), .o(n_32777) );
ao12s01 g748358 ( .a(n_32727), .b(n_32726), .c(n_32725), .o(n_33279) );
in01s01 g748359 ( .a(n_33415), .o(n_33576) );
ao12s01 g748360 ( .a(n_32749), .b(n_32748), .c(n_32747), .o(n_33415) );
in01s02 g748361 ( .a(n_31825), .o(n_31826) );
na02s02 g748362 ( .a(n_31729), .b(n_31760), .o(n_31825) );
in01s01 g748363 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_7_), .o(n_32952) );
no02s01 g748367 ( .a(n_32748), .b(n_32747), .o(n_32749) );
no02s01 g748368 ( .a(n_32726), .b(n_32725), .o(n_32727) );
in01s01 g748369 ( .a(n_32750), .o(n_32780) );
ao12s06 g748370 ( .a(n_32442), .b(n_32674), .c(n_32588), .o(n_32750) );
na02s01 g748371 ( .a(FE_OCP_RBN6874_n_31520), .b(n_31795), .o(n_31897) );
in01s01 g748372 ( .a(n_31823), .o(n_31824) );
no02s01 g748373 ( .a(FE_OCP_RBN6874_n_31520), .b(n_31795), .o(n_31823) );
in01s01 g748374 ( .a(n_31501), .o(n_31560) );
in01s01 g748376 ( .a(n_31477), .o(n_31559) );
na02s06 g748378 ( .a(n_31476), .b(FE_OCP_DRV_N3516_n_31504), .o(n_31522) );
in01s01 g748379 ( .a(n_31793), .o(n_31794) );
na02s01 g748380 ( .a(FE_OCP_RBN6872_n_31520), .b(n_30505), .o(n_31793) );
na02s01 g748381 ( .a(FE_OCP_RBN6875_n_31520), .b(n_30526), .o(n_31862) );
in01s01 g748382 ( .a(n_31475), .o(n_31610) );
na02s02 g748383 ( .a(n_31449), .b(n_31448), .o(n_31475) );
no02s06 g748387 ( .a(n_31518), .b(n_31448), .o(n_31605) );
no02s01 g748388 ( .a(FE_OCP_RBN6875_n_31520), .b(n_31502), .o(n_31791) );
no02s03 g748389 ( .a(n_31518), .b(n_30553), .o(n_31664) );
na02f04 TIMEBOOST_cell_1455 ( .a(n_29428), .b(n_25738), .o(TIMEBOOST_net_342) );
no02s01 g748391 ( .a(FE_OCPN943_n_31466), .b(FE_OCP_RBN1845_n_30492), .o(n_31735) );
no02m03 g748395 ( .a(n_31520), .b(n_30492), .o(n_31554) );
no02s01 g748396 ( .a(FE_OCP_RBN3370_n_31520), .b(n_30637), .o(n_31764) );
na02m02 TIMEBOOST_cell_1461 ( .a(n_24618), .b(n_22207), .o(TIMEBOOST_net_345) );
no02s06 TIMEBOOST_cell_2793 ( .a(TIMEBOOST_net_687), .b(n_6715), .o(n_6710) );
in01s02 g748400 ( .a(n_31763), .o(n_31788) );
no02s06 g748402 ( .a(n_31730), .b(FE_OCP_RBN2106_n_30619), .o(n_31763) );
in01s02 g748403 ( .a(n_31553), .o(n_32168) );
na02s06 g748404 ( .a(n_31520), .b(FE_OCP_RBN2106_n_30619), .o(n_31553) );
na02f02 TIMEBOOST_cell_8773 ( .a(TIMEBOOST_net_2873), .b(n_14379), .o(n_14475) );
no02s01 TIMEBOOST_cell_1481 ( .a(n_41617), .b(n_41599), .o(TIMEBOOST_net_355) );
in01s02 g748409 ( .a(n_31787), .o(n_31821) );
no02f01 g748410 ( .a(FE_OCP_RBN3368_n_31520), .b(n_30643), .o(n_31787) );
no02s02 g748411 ( .a(n_31520), .b(FE_OCP_RBN3080_n_30643), .o(n_32149) );
na02s01 g748412 ( .a(n_31730), .b(FE_OCP_RBN1859_n_30731), .o(n_31729) );
na02s01 g748413 ( .a(FE_OCP_RBN6139_n_31520), .b(n_30731), .o(n_31760) );
no02s03 g748417 ( .a(n_30814), .b(n_31466), .o(n_31594) );
in01s01 g748420 ( .a(FE_OCPN3586_n_31704), .o(n_31727) );
no02s01 g748421 ( .a(n_31518), .b(n_46958), .o(n_31704) );
na02s01 g748422 ( .a(n_31730), .b(FE_OCP_RBN3141_n_30849), .o(n_31725) );
na02s02 TIMEBOOST_cell_5639 ( .a(TIMEBOOST_net_1767), .b(n_6048), .o(n_6154) );
na02s01 g748424 ( .a(FE_OCP_RBN6139_n_31520), .b(n_30906), .o(n_31759) );
no02s06 g748425 ( .a(FE_OCP_RBN6875_n_31520), .b(n_31655), .o(n_32197) );
in01s01 g748428 ( .a(n_31681), .o(n_31703) );
na02s02 g748429 ( .a(n_31476), .b(n_31655), .o(n_31681) );
na03s02 TIMEBOOST_cell_8742 ( .a(n_41695), .b(n_41696), .c(FE_OCP_RBN5673_n_41420), .o(TIMEBOOST_net_2858) );
na02m01 g748431 ( .a(n_30954), .b(FE_OCPN943_n_31466), .o(n_31682) );
no02s02 TIMEBOOST_cell_1483 ( .a(n_2805), .b(n_2227), .o(TIMEBOOST_net_356) );
na02s02 TIMEBOOST_cell_1485 ( .a(n_24422), .b(n_24574), .o(TIMEBOOST_net_357) );
na03m04 TIMEBOOST_cell_4622 ( .a(n_13145), .b(n_13148), .c(n_13230), .o(n_13367) );
no03s02 TIMEBOOST_cell_8223 ( .a(n_24560), .b(FE_OCPN1669_n_23941), .c(FE_OCPN1668_n_23941), .o(TIMEBOOST_net_1871) );
na02s01 g748436 ( .a(n_31730), .b(n_31107), .o(n_31721) );
in01s01 g748437 ( .a(n_31550), .o(n_31551) );
na02s01 g748438 ( .a(n_31519), .b(n_31469), .o(n_31550) );
na02f04 g748439 ( .a(n_31474), .b(FE_OCP_DRV_N1496_n_31473), .o(n_31521) );
in01s01 g748440 ( .a(n_31499), .o(n_31500) );
no02s04 g748441 ( .a(n_31474), .b(FE_OCP_DRV_N1496_n_31473), .o(n_31499) );
in01s01 g748442 ( .a(n_31784), .o(n_31785) );
na02s01 g748443 ( .a(n_31699), .b(n_31756), .o(n_31784) );
in01s01 g748444 ( .a(n_31754), .o(n_31755) );
no02m06 g748445 ( .a(n_31720), .b(FE_OCPN1938_n_31719), .o(n_31754) );
na02m06 g748446 ( .a(n_31720), .b(FE_OCPN1938_n_31719), .o(n_31799) );
ao12s01 g748447 ( .a(n_32587), .b(n_32677), .c(n_32482), .o(n_32766) );
in01s08 g748451 ( .a(n_31783), .o(n_31835) );
in01m10 g748452 ( .a(n_31765), .o(n_31783) );
in01f08 g748453 ( .a(n_31718), .o(n_31765) );
in01m10 g748492 ( .a(n_31783), .o(n_31819) );
oa12f06 g748495 ( .a(n_31494), .b(n_31589), .c(FE_OCP_RBN3273_n_31239), .o(n_31718) );
in01s01 g748497 ( .a(n_31549), .o(n_31612) );
no02s06 g748499 ( .a(n_31518), .b(n_30528), .o(n_31593) );
in01s01 g748501 ( .a(n_31548), .o(n_31591) );
na02s06 g748502 ( .a(n_31520), .b(n_30525), .o(n_31548) );
in01s01 g748503 ( .a(n_31652), .o(n_31653) );
oa12s02 g748504 ( .a(n_31520), .b(FE_OCP_RBN1859_n_30731), .c(FE_OCP_RBN3079_n_30643), .o(n_31652) );
na02m02 g748505 ( .a(n_31476), .b(n_30803), .o(n_31683) );
in01s01 g748507 ( .a(n_31702), .o(n_31716) );
na02s02 g748508 ( .a(n_31518), .b(n_30989), .o(n_31702) );
in01s01 g748509 ( .a(n_31471), .o(n_31472) );
in01s01 g748510 ( .a(n_31447), .o(n_31471) );
ao12f08 g748511 ( .a(n_31332), .b(n_31426), .c(n_31382), .o(n_31447) );
oa22s01 g748512 ( .a(n_31402), .b(n_31385), .c(n_31401), .d(n_31426), .o(n_31470) );
in01s01 g748513 ( .a(n_31700), .o(n_31701) );
in01s01 g748514 ( .a(n_31678), .o(n_31700) );
ao12f08 g748515 ( .a(n_31491), .b(n_31546), .c(n_31489), .o(n_31678) );
oa22s01 g748516 ( .a(n_31585), .b(n_31647), .c(n_31586), .d(n_31646), .o(n_31715) );
no02s01 g748517 ( .a(n_32675), .b(n_32606), .o(n_32748) );
na02s01 g748518 ( .a(n_32676), .b(n_32497), .o(n_32726) );
in01s01 g748519 ( .a(n_31468), .o(n_31469) );
no02m04 g748520 ( .a(n_31446), .b(FE_OCP_DRV_N1492_n_31445), .o(n_31468) );
na02m06 g748521 ( .a(n_31446), .b(FE_OCP_DRV_N1492_n_31445), .o(n_31519) );
in01s01 g748522 ( .a(n_31497), .o(n_31498) );
na02s01 g748523 ( .a(n_31467), .b(n_31425), .o(n_31497) );
in01s01 g748524 ( .a(n_31698), .o(n_31699) );
no02s06 g748525 ( .a(n_31677), .b(FE_OCPN1936_n_31676), .o(n_31698) );
na02s08 g748526 ( .a(n_31677), .b(FE_OCPN1936_n_31676), .o(n_31756) );
in01s01 g748527 ( .a(n_31713), .o(n_31714) );
na02s01 g748528 ( .a(n_31697), .b(n_31649), .o(n_31713) );
in01s02 g748529 ( .a(FE_OCPN943_n_31466), .o(n_31730) );
in01m10 g748551 ( .a(n_31466), .o(n_31520) );
in01m08 g748552 ( .a(n_31449), .o(n_31466) );
in01m10 g748559 ( .a(n_31476), .o(n_31518) );
in01m10 g748560 ( .a(n_31449), .o(n_31476) );
no02f20 g748561 ( .a(n_31202), .b(n_31386), .o(n_31449) );
no03m04 TIMEBOOST_cell_8516 ( .a(n_38057), .b(n_38007), .c(n_37974), .o(TIMEBOOST_net_2745) );
oa22s01 g748563 ( .a(n_31335), .b(n_31331), .c(n_31334), .d(n_31330), .o(n_31405) );
no02f06 g748564 ( .a(n_31588), .b(n_31547), .o(n_31720) );
oa22s01 g748565 ( .a(n_31545), .b(n_31487), .c(n_31544), .d(n_31486), .o(n_31673) );
oa12s01 g748566 ( .a(n_32657), .b(n_32658), .c(n_32656), .o(n_33370) );
na02s01 g748570 ( .a(n_32746), .b(n_32558), .o(n_32776) );
in01s01 g748571 ( .a(n_32676), .o(n_32677) );
na02s01 g748572 ( .a(n_32658), .b(n_32447), .o(n_32676) );
na02s01 g748573 ( .a(n_32658), .b(n_32656), .o(n_32657) );
no02f04 g748574 ( .a(n_31587), .b(FE_OCPN5262_n_27536), .o(n_31589) );
no02f02 g748575 ( .a(n_31515), .b(n_31361), .o(n_31547) );
no02s02 g748576 ( .a(n_31587), .b(n_31360), .o(n_31588) );
no02f10 g748577 ( .a(n_31383), .b(n_31201), .o(n_31386) );
in01s01 g748578 ( .a(n_31426), .o(n_31385) );
ao12f08 g748579 ( .a(n_31300), .b(n_31270), .c(n_31272), .o(n_31426) );
in01s01 g748580 ( .a(n_31424), .o(n_31425) );
no02f06 g748581 ( .a(n_31404), .b(FE_OCPN1320_n_31403), .o(n_31424) );
na02f06 g748582 ( .a(n_31404), .b(FE_OCPN1272_n_31403), .o(n_31467) );
na02m02 g748583 ( .a(n_31336), .b(n_31245), .o(n_31365) );
na02m04 TIMEBOOST_cell_7715 ( .a(TIMEBOOST_net_2488), .b(n_29616), .o(TIMEBOOST_net_360) );
in01s01 g748585 ( .a(n_31648), .o(n_31649) );
no02m04 g748586 ( .a(n_31584), .b(FE_OCPUNCON7073_n_31583), .o(n_31648) );
in01s01 g748587 ( .a(n_31585), .o(n_31586) );
in01s01 g748588 ( .a(n_31546), .o(n_31585) );
ao12f08 g748589 ( .a(n_31462), .b(n_31440), .c(n_31442), .o(n_31546) );
na02s06 g748590 ( .a(n_31584), .b(FE_OCPUNCON7073_n_31583), .o(n_31697) );
in01s01 g748591 ( .a(n_32674), .o(n_32675) );
na02s06 g748592 ( .a(n_32658), .b(n_32500), .o(n_32674) );
na02s01 g748595 ( .a(n_32723), .b(n_32491), .o(n_32724) );
in01s01 g748596 ( .a(n_33146), .o(n_32746) );
na02s02 g748597 ( .a(n_32538), .b(n_32723), .o(n_33146) );
na02s03 g748600 ( .a(n_31492), .b(FE_OCPN5262_n_27536), .o(n_31494) );
in01s01 g748603 ( .a(n_31401), .o(n_31402) );
na02s01 g748604 ( .a(n_31382), .b(n_31333), .o(n_31401) );
na02s06 g748605 ( .a(n_32611), .b(n_32562), .o(n_32658) );
in01m04 g748606 ( .a(n_31515), .o(n_31587) );
no02f08 g748607 ( .a(n_31492), .b(n_31237), .o(n_31515) );
in01m06 g748609 ( .a(n_31336), .o(n_31383) );
oa12f06 g748610 ( .a(n_31109), .b(n_31273), .c(n_31136), .o(n_31336) );
oa12s01 g748611 ( .a(n_31302), .b(n_31301), .c(n_31308), .o(n_31363) );
in01s01 g748612 ( .a(n_31334), .o(n_31335) );
oa12s01 g748613 ( .a(n_31271), .b(n_31308), .c(n_31268), .o(n_31334) );
oa22s01 g748615 ( .a(n_31438), .b(n_31419), .c(n_31437), .d(n_31420), .o(n_31514) );
in01s01 g748616 ( .a(n_31544), .o(n_31545) );
oa12s01 g748617 ( .a(n_31441), .b(n_31438), .c(n_31356), .o(n_31544) );
in01s01 g748618 ( .a(n_31646), .o(n_31647) );
oa22s01 g748619 ( .a(n_31485), .b(n_31490), .c(n_31484), .d(n_29966), .o(n_31646) );
ao12s02 g748623 ( .a(n_33028), .b(n_32453), .c(n_46107), .o(n_32723) );
na02s04 g748627 ( .a(n_31443), .b(n_31236), .o(n_31463) );
na02m06 g748632 ( .a(n_31273), .b(n_31083), .o(n_31305) );
in01s01 g748633 ( .a(n_31332), .o(n_31333) );
no02m04 g748634 ( .a(n_31304), .b(n_31303), .o(n_31332) );
na02f04 g748635 ( .a(n_31304), .b(n_31303), .o(n_31382) );
na02f08 g748636 ( .a(n_31308), .b(n_31271), .o(n_31272) );
na02s01 g748637 ( .a(n_31308), .b(n_31301), .o(n_31302) );
no02m06 g748638 ( .a(n_31488), .b(n_31490), .o(n_31491) );
na02m06 g748639 ( .a(n_31488), .b(n_31490), .o(n_31489) );
na02f08 g748640 ( .a(n_31421), .b(n_31441), .o(n_31442) );
oa12s04 g748641 ( .a(FE_OCP_RBN2311_delay_sub_ln23_unr25_stage8_stallmux_q_1_), .b(n_32610), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_), .o(n_32611) );
no02s01 TIMEBOOST_cell_4874 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_12_), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_11_), .o(TIMEBOOST_net_1385) );
in01s01 g748643 ( .a(n_33362), .o(n_33396) );
oa12s01 g748644 ( .a(n_32590), .b(n_32610), .c(n_32589), .o(n_33362) );
na02s01 g748645 ( .a(n_32645), .b(n_32448), .o(n_32646) );
no02m04 TIMEBOOST_cell_6951 ( .a(n_8128), .b(FE_OCP_RBN2670_n_46991), .o(TIMEBOOST_net_2234) );
oa12s02 g748647 ( .a(n_32645), .b(n_32424), .c(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_33028) );
na02s01 g748648 ( .a(n_32610), .b(n_32589), .o(n_32590) );
na02f08 g748649 ( .a(n_31400), .b(n_31130), .o(n_31443) );
no02m06 g748653 ( .a(n_31209), .b(n_30995), .o(n_31246) );
na02m08 g748654 ( .a(n_31209), .b(n_31030), .o(n_31273) );
no02f08 g748655 ( .a(n_31269), .b(n_31268), .o(n_31270) );
in01s01 g748656 ( .a(n_31330), .o(n_31331) );
no02s01 g748657 ( .a(n_31269), .b(n_31300), .o(n_31330) );
no02f06 g748658 ( .a(n_31439), .b(n_31356), .o(n_31440) );
in01s01 g748659 ( .a(n_31486), .o(n_31487) );
no02s01 g748660 ( .a(n_31439), .b(n_31462), .o(n_31486) );
oa12s01 g748663 ( .a(n_31205), .b(n_31204), .c(n_31203), .o(n_31267) );
in01s01 g748664 ( .a(n_31484), .o(n_31485) );
in01s01 g748665 ( .a(n_31488), .o(n_31484) );
na02s02 TIMEBOOST_cell_4531 ( .a(n_11129), .b(n_11015), .o(TIMEBOOST_net_1356) );
in01s01 g748667 ( .a(n_31437), .o(n_31438) );
in01s01 g748669 ( .a(n_31421), .o(n_31437) );
ao12f08 g748670 ( .a(n_31297), .b(n_31399), .c(n_31352), .o(n_31421) );
oa22s01 g748671 ( .a(n_31357), .b(n_31375), .c(n_31399), .d(n_31376), .o(n_31435) );
in01s01 g748673 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_4_), .o(n_32670) );
no02s01 g748675 ( .a(n_32537), .b(n_32559), .o(n_32563) );
na02s02 g748676 ( .a(n_32509), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_), .o(n_32562) );
in01s01 g748677 ( .a(n_32781), .o(n_32628) );
no02s02 g748678 ( .a(n_32796), .b(n_32494), .o(n_32781) );
ao12s02 g748679 ( .a(n_44042), .b(n_32451), .c(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_32645) );
oa12s08 g748680 ( .a(n_32446), .b(n_32539), .c(n_32508), .o(n_32610) );
no02f08 g748681 ( .a(n_31329), .b(n_31075), .o(n_31400) );
na02s04 g748682 ( .a(n_31358), .b(n_31077), .o(n_31381) );
na02m04 TIMEBOOST_cell_4530 ( .a(TIMEBOOST_net_1355), .b(n_11071), .o(n_11212) );
no02m08 g748684 ( .a(n_31142), .b(n_30996), .o(n_31209) );
in01f04 g748685 ( .a(n_31208), .o(n_31300) );
na02f03 g748686 ( .a(n_31207), .b(FE_OCP_DRV_N5155_n_31206), .o(n_31208) );
no02f06 g748687 ( .a(n_31207), .b(FE_OCP_DRV_N5155_n_31206), .o(n_31269) );
na02s01 g748689 ( .a(n_31204), .b(n_31203), .o(n_31205) );
na02s01 g748690 ( .a(n_31271), .b(n_31183), .o(n_31301) );
no02m06 g748691 ( .a(n_31380), .b(n_29843), .o(n_31462) );
no02f04 g748692 ( .a(n_31379), .b(n_29842), .o(n_31439) );
ao12s01 g748693 ( .a(n_32561), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_30_), .o(n_33192) );
na02s01 g748694 ( .a(n_32505), .b(n_32510), .o(n_32560) );
ao12s01 g748695 ( .a(n_32559), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_29_), .o(n_33130) );
no02s02 g748696 ( .a(n_32557), .b(n_32536), .o(n_32607) );
oa22s02 g748697 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_6_), .c(n_32587), .d(n_32496), .o(n_32588) );
oa12s01 g748698 ( .a(n_32495), .b(n_32532), .c(n_32499), .o(n_32606) );
ao12s01 g748699 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n_32558), .c(n_32462), .o(n_32608) );
in01m01 g748700 ( .a(n_31360), .o(n_31361) );
in01s01 g748702 ( .a(n_33240), .o(n_33256) );
oa22s01 g748703 ( .a(n_32460), .b(n_32479), .c(n_32539), .d(n_32480), .o(n_33240) );
no02s01 g748705 ( .a(n_32408), .b(n_32507), .o(n_32510) );
no02s01 g748706 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_29_), .o(n_32559) );
no02s01 g748707 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_30_), .o(n_32561) );
oa12s01 g748708 ( .a(n_32586), .b(n_32493), .c(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_32796) );
in01s01 g748709 ( .a(n_44042), .o(n_32605) );
no02s02 g748711 ( .a(n_32539), .b(n_32508), .o(n_32509) );
in01m02 g748712 ( .a(n_31244), .o(n_31245) );
no02m08 g748713 ( .a(n_31201), .b(n_31202), .o(n_31244) );
in01s01 g748714 ( .a(n_31268), .o(n_31183) );
no02f04 g748715 ( .a(n_31165), .b(FE_OCP_DRV_N5153_n_31164), .o(n_31268) );
na02f04 g748716 ( .a(n_31165), .b(FE_OCP_DRV_N5153_n_31164), .o(n_31271) );
no02s01 g748717 ( .a(n_31162), .b(n_31163), .o(n_31204) );
in01s01 g748718 ( .a(n_31419), .o(n_31420) );
na02s01 g748719 ( .a(n_31441), .b(n_31377), .o(n_31419) );
ao12s01 g748720 ( .a(n_32507), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_27_), .o(n_33127) );
no02s10 TIMEBOOST_cell_8713 ( .a(TIMEBOOST_net_2843), .b(FE_RN_5_0), .o(n_18096) );
na02f08 TIMEBOOST_cell_8531 ( .a(TIMEBOOST_net_2752), .b(FE_RN_18_0), .o(TIMEBOOST_net_2226) );
in01f02 g748723 ( .a(n_31160), .o(n_31161) );
in01f02 g748724 ( .a(n_31142), .o(n_31160) );
no02f08 g748725 ( .a(n_31062), .b(n_31063), .o(n_31142) );
in01m02 g748726 ( .a(n_31358), .o(n_31359) );
in01m02 g748727 ( .a(n_31329), .o(n_31358) );
no02f06 g748728 ( .a(n_31242), .b(n_31243), .o(n_31329) );
oa12s01 g748729 ( .a(n_46107), .b(n_32405), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_27_), .o(n_32538) );
in01s01 g748731 ( .a(n_31141), .o(n_31203) );
oa12f04 g748732 ( .a(n_31035), .b(n_31086), .c(n_31138), .o(n_31141) );
oa12s01 g748733 ( .a(n_31140), .b(n_31139), .c(n_31138), .o(n_31182) );
in01m02 g748734 ( .a(n_31379), .o(n_31380) );
no02m04 TIMEBOOST_cell_3412 ( .a(n_27229), .b(FE_RN_1282_0), .o(TIMEBOOST_net_997) );
in01s01 g748736 ( .a(n_31399), .o(n_31357) );
ao12f08 g748737 ( .a(n_31230), .b(n_31353), .c(n_31296), .o(n_31399) );
oa12s01 g748738 ( .a(n_31355), .b(n_31354), .c(n_31353), .o(n_31397) );
in01s01 g748739 ( .a(n_32584), .o(n_32585) );
oa12s01 g748740 ( .a(n_32504), .b(n_32503), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n_32584) );
in01s01 g748743 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_29_), .o(n_32462) );
in01s01 g748746 ( .a(n_32505), .o(n_32506) );
no02s01 g748747 ( .a(n_32489), .b(n_32461), .o(n_32505) );
no02s01 g748748 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_27_), .o(n_32507) );
no02s01 g748749 ( .a(n_32537), .b(n_32449), .o(n_33091) );
na02s01 g748750 ( .a(n_32503), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n_32504) );
na02f06 TIMEBOOST_cell_3411 ( .a(TIMEBOOST_net_996), .b(n_36611), .o(n_36703) );
na02s20 TIMEBOOST_cell_8465 ( .a(n_36910), .b(TIMEBOOST_net_2719), .o(n_36921) );
ao12f04 g748755 ( .a(FE_OCPN5286_n_30708), .b(n_31241), .c(n_31027), .o(n_31243) );
ao12f08 g748756 ( .a(n_27246), .b(n_31061), .c(n_30889), .o(n_31063) );
no02m10 g748757 ( .a(n_31112), .b(n_27366), .o(n_31202) );
no02s06 g748758 ( .a(n_31111), .b(n_27536), .o(n_31201) );
no02f04 g748759 ( .a(n_31056), .b(FE_OFN4733_n_29677), .o(n_31163) );
no02m06 g748760 ( .a(n_31057), .b(n_29678), .o(n_31162) );
na02s01 g748761 ( .a(n_31139), .b(n_31138), .o(n_31140) );
in01s01 g748763 ( .a(n_31356), .o(n_31377) );
no02m06 g748764 ( .a(n_31328), .b(n_31327), .o(n_31356) );
na02m06 g748765 ( .a(n_31328), .b(n_31327), .o(n_31441) );
na02s01 g748766 ( .a(n_31354), .b(n_31353), .o(n_31355) );
in01s01 g748767 ( .a(n_31375), .o(n_31376) );
na02s01 g748768 ( .a(n_31352), .b(n_31298), .o(n_31375) );
ao12s01 g748769 ( .a(n_32425), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_23_), .o(n_33171) );
in01s01 g748770 ( .a(n_32535), .o(n_32536) );
no02m04 TIMEBOOST_cell_8657 ( .a(TIMEBOOST_net_2815), .b(n_36777), .o(n_36787) );
in01s01 g748772 ( .a(n_32533), .o(n_32534) );
na02s01 TIMEBOOST_cell_2918 ( .a(n_38093), .b(n_38020), .o(TIMEBOOST_net_750) );
no02s06 TIMEBOOST_cell_1556 ( .a(TIMEBOOST_net_392), .b(n_3419), .o(n_4528) );
in01s01 g748775 ( .a(n_32587), .o(n_32532) );
ao12s02 g748776 ( .a(n_32498), .b(n_32481), .c(n_32497), .o(n_32587) );
ao12s01 g748777 ( .a(n_32461), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_25_), .o(n_33121) );
in01s01 g748778 ( .a(n_32539), .o(n_32460) );
ao12s10 g748779 ( .a(n_32376), .b(n_32423), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n_32539) );
oa12f08 g748780 ( .a(n_30857), .b(n_31061), .c(n_30943), .o(n_31062) );
oa12f04 g748781 ( .a(n_30962), .b(n_31241), .c(n_31081), .o(n_31242) );
ao12s01 g748782 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n_32495), .c(n_31887), .o(n_32496) );
ao12s01 g748783 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n_32416), .c(n_32157), .o(n_32494) );
no03s40 TIMEBOOST_cell_3464 ( .a(n_17547), .b(FE_RN_271_0), .c(FE_RN_270_0), .o(n_17617) );
na02f08 TIMEBOOST_cell_7849 ( .a(TIMEBOOST_net_2555), .b(n_16056), .o(n_16231) );
oa12s01 g748788 ( .a(n_31263), .b(n_31262), .c(n_31261), .o(n_31326) );
in01s01 g748789 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_2_), .o(n_32654) );
no02s01 g748792 ( .a(n_32445), .b(n_32459), .o(n_32556) );
na02s01 g748793 ( .a(n_32586), .b(n_32457), .o(n_32458) );
na02s01 g748794 ( .a(n_32455), .b(n_32454), .o(n_32456) );
no02s01 g748795 ( .a(n_32409), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_11_), .o(n_32493) );
na02s01 g748796 ( .a(n_32407), .b(n_32357), .o(n_32453) );
in01s01 g748797 ( .a(n_32425), .o(n_32426) );
no02s01 g748798 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_23_), .o(n_32425) );
no02s01 g748799 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_25_), .o(n_32461) );
in01s01 g748800 ( .a(n_32537), .o(n_32452) );
no02s01 g748801 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_28_), .o(n_32537) );
no02s01 g748802 ( .a(n_32390), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_23_), .o(n_32424) );
no02s02 g748803 ( .a(n_32417), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_19_), .o(n_32492) );
na02s01 g748804 ( .a(n_32318), .b(n_32450), .o(n_32451) );
in01s01 g748805 ( .a(n_32558), .o(n_32449) );
na02s01 g748806 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_28_), .o(n_32558) );
na02s01 g748807 ( .a(n_32491), .b(n_32490), .o(n_33118) );
no02s01 g748808 ( .a(n_32489), .b(n_32488), .o(n_33069) );
na02s01 g748809 ( .a(n_32454), .b(n_32487), .o(n_33084) );
na02s01 g748810 ( .a(n_32450), .b(n_32412), .o(n_33042) );
no02s01 g748811 ( .a(n_32603), .b(n_32486), .o(n_32823) );
na02s01 g748812 ( .a(n_32420), .b(n_32419), .o(n_32803) );
no02s01 g748813 ( .a(n_32410), .b(n_32499), .o(n_32765) );
na02s01 g748814 ( .a(n_32448), .b(n_32555), .o(n_33115) );
in01s01 g748815 ( .a(n_32530), .o(n_32531) );
na02s01 g748816 ( .a(n_32485), .b(n_32415), .o(n_32530) );
na02s01 g748817 ( .a(n_32457), .b(n_32484), .o(n_32837) );
no02s01 g748818 ( .a(n_32483), .b(n_32404), .o(n_32763) );
na02s01 g748819 ( .a(n_32482), .b(n_32481), .o(n_32725) );
na02s01 g748820 ( .a(n_32497), .b(n_32447), .o(n_32656) );
na02s01 g748821 ( .a(n_32377), .b(n_32423), .o(n_32503) );
in01s01 g748822 ( .a(n_32479), .o(n_32480) );
na02s01 g748823 ( .a(n_32392), .b(n_32446), .o(n_32479) );
no02m08 TIMEBOOST_cell_7861 ( .a(TIMEBOOST_net_2561), .b(TIMEBOOST_net_867), .o(n_16241) );
no02m04 g748825 ( .a(n_31015), .b(n_30937), .o(n_31060) );
na02s04 g748826 ( .a(n_31200), .b(n_31236), .o(n_31237) );
na02s06 g748828 ( .a(FE_OCP_RBN6840_FE_RN_2660_0), .b(n_31200), .o(n_31234) );
no03s08 TIMEBOOST_cell_843 ( .a(n_17239), .b(n_16973), .c(n_17244), .o(TIMEBOOST_net_36) );
no02m04 g748830 ( .a(FE_OCP_RBN3230_n_31107), .b(FE_OCPN5262_n_27536), .o(n_31158) );
no02s01 g748831 ( .a(n_31036), .b(n_31086), .o(n_31139) );
na02m06 g748832 ( .a(n_31265), .b(FE_OCP_DRV_N5151_n_31264), .o(n_31352) );
in01s01 g748833 ( .a(n_31297), .o(n_31298) );
no02f04 g748834 ( .a(n_31265), .b(FE_OCP_DRV_N5151_n_31264), .o(n_31297) );
na02s01 g748835 ( .a(n_31262), .b(n_31261), .o(n_31263) );
na02s01 g748836 ( .a(n_31296), .b(n_31231), .o(n_31354) );
ao12s01 g748837 ( .a(n_32445), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_21_), .o(n_33124) );
ao12s01 g748838 ( .a(n_32444), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_11_), .o(n_32840) );
ao12s01 g748839 ( .a(n_32443), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_13_), .o(n_32864) );
ao12s01 g748840 ( .a(n_32442), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_7_), .o(n_32747) );
ao12s01 g748841 ( .a(n_32441), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_19_), .o(n_33088) );
in01s02 g748844 ( .a(n_31232), .o(n_31233) );
na02f02 g748845 ( .a(n_31241), .b(n_31032), .o(n_31232) );
ao12f04 g748846 ( .a(n_30947), .b(n_31053), .c(n_31011), .o(n_31138) );
in01m02 g748847 ( .a(n_31056), .o(n_31057) );
in01m04 g748849 ( .a(n_31111), .o(n_31112) );
oa12s01 g748851 ( .a(n_31055), .b(n_31054), .c(n_31053), .o(n_31110) );
na02m06 g748852 ( .a(n_31199), .b(n_31180), .o(n_31328) );
oa12f08 g748853 ( .a(n_31196), .b(n_31177), .c(n_31151), .o(n_31353) );
oa22s01 g748854 ( .a(n_32316), .b(n_31579), .c(FE_OCP_RBN3463_n_32316), .d(n_31578), .o(n_32379) );
oa22s01 g748855 ( .a(n_32314), .b(n_31635), .c(n_32315), .d(n_31636), .o(n_32378) );
oa22s01 g748856 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .c(n_32271), .d(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_33045) );
oa22s01 g748857 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_15_), .c(n_32422), .d(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_32881) );
oa22s01 g748858 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_), .c(n_32034), .d(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_32806) );
oa22s01 g748859 ( .a(n_31778), .b(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .c(FE_OCP_RBN2311_delay_sub_ln23_unr25_stage8_stallmux_q_1_), .d(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_), .o(n_32589) );
in01s01 g748860 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_1_), .o(n_32684) );
in01s01 g748863 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_), .o(n_31260) );
in01s06 g748865 ( .a(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37709) );
in01s01 g748868 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_25_), .o(n_32357) );
no02s01 g748871 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_24_), .o(n_32489) );
na02s01 g748872 ( .a(n_32375), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_32555) );
in01s01 g748873 ( .a(n_32420), .o(n_32421) );
na02s01 g748874 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_14_), .o(n_32420) );
in01s01 g748875 ( .a(n_32418), .o(n_32419) );
no02s01 g748876 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_14_), .o(n_32418) );
na02s02 g748877 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_5_), .o(n_32481) );
no02s01 g748878 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_19_), .o(n_32441) );
in01s01 g748879 ( .a(n_32376), .o(n_32377) );
no02s10 g748880 ( .a(n_32356), .b(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .o(n_32376) );
in01s01 g748881 ( .a(n_32454), .o(n_32417) );
na02s01 g748882 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_18_), .o(n_32454) );
in01s01 g748883 ( .a(n_32416), .o(n_32486) );
na02s01 g748884 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_12_), .o(n_32416) );
in01s01 g748885 ( .a(n_32414), .o(n_32415) );
no02s01 g748886 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .o(n_32414) );
no02s01 g748887 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_), .o(n_32483) );
in01s01 g748888 ( .a(n_32413), .o(n_32487) );
no02s01 g748889 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_18_), .o(n_32413) );
in01s01 g748890 ( .a(n_32459), .o(n_32412) );
no02s01 g748891 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_20_), .o(n_32459) );
no02s01 g748892 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_21_), .o(n_32445) );
no02s01 g748893 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_11_), .o(n_32444) );
in01s01 g748894 ( .a(n_32411), .o(n_32484) );
no02s01 g748895 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_10_), .o(n_32411) );
no02s01 g748896 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_13_), .o(n_32443) );
no02s01 g748897 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_12_), .o(n_32603) );
no02s02 g748898 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_7_), .o(n_32442) );
in01s01 g748899 ( .a(n_32508), .o(n_32392) );
no02s06 g748900 ( .a(FE_OCP_RBN2311_delay_sub_ln23_unr25_stage8_stallmux_q_1_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_2_), .o(n_32508) );
na02s10 g748901 ( .a(n_32356), .b(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .o(n_32423) );
na02s03 g748902 ( .a(FE_OCP_RBN2311_delay_sub_ln23_unr25_stage8_stallmux_q_1_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_2_), .o(n_32446) );
no02s01 g748903 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_6_), .o(n_32499) );
in01s01 g748904 ( .a(n_32498), .o(n_32482) );
no02s02 g748905 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_5_), .o(n_32498) );
in01s01 g748906 ( .a(n_32391), .o(n_32447) );
no02s01 g748907 ( .a(FE_OCP_RBN2311_delay_sub_ln23_unr25_stage8_stallmux_q_1_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_4_), .o(n_32391) );
na02s02 g748908 ( .a(FE_OCP_RBN2311_delay_sub_ln23_unr25_stage8_stallmux_q_1_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_4_), .o(n_32497) );
in01s01 g748909 ( .a(n_32495), .o(n_32410) );
na02s02 g748910 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_6_), .o(n_32495) );
in01s01 g748911 ( .a(n_32457), .o(n_32409) );
na02s02 g748912 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_10_), .o(n_32457) );
in01s01 g748913 ( .a(n_32408), .o(n_32490) );
no02s01 g748914 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_26_), .o(n_32408) );
in01s01 g748915 ( .a(n_32407), .o(n_32488) );
na02s01 g748916 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_24_), .b(n_46107), .o(n_32407) );
in01s01 g748917 ( .a(n_32390), .o(n_32448) );
no02s01 g748918 ( .a(n_32375), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_32390) );
in01s01 g748919 ( .a(n_32450), .o(n_32406) );
na02s01 g748920 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_20_), .o(n_32450) );
in01s01 g748921 ( .a(n_32491), .o(n_32405) );
na02s01 g748922 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_26_), .b(n_46107), .o(n_32491) );
na02s01 g748923 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .o(n_32485) );
in01s01 g748924 ( .a(n_32403), .o(n_32404) );
na02s01 g748925 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_), .o(n_32403) );
na02f10 g748926 ( .a(n_30967), .b(n_30913), .o(n_31061) );
in01m02 g748927 ( .a(n_31014), .o(n_31015) );
no02m02 g748928 ( .a(n_30967), .b(n_30890), .o(n_31014) );
na02f08 g748929 ( .a(n_31132), .b(n_31050), .o(n_31241) );
na02s04 g748930 ( .a(FE_OCP_RBN6091_n_31153), .b(n_31070), .o(n_31199) );
na02m02 g748931 ( .a(n_31153), .b(n_31071), .o(n_31180) );
no02s06 g748932 ( .a(n_31082), .b(n_31108), .o(n_31109) );
no02s04 g748934 ( .a(n_31136), .b(n_31108), .o(n_31156) );
na02s04 g748937 ( .a(n_31101), .b(n_27366), .o(n_31200) );
in01s01 g748938 ( .a(n_31035), .o(n_31036) );
na02s01 g748941 ( .a(n_31054), .b(n_31053), .o(n_31055) );
in01s01 g748942 ( .a(n_31230), .o(n_31231) );
no02m06 g748943 ( .a(n_31198), .b(FE_OCPN5124_n_31197), .o(n_31230) );
na02m06 g748944 ( .a(n_31198), .b(FE_OCPN5124_n_31197), .o(n_31296) );
na02s01 g748945 ( .a(n_31196), .b(n_31152), .o(n_31262) );
oa12s01 g748946 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_), .o(n_32586) );
ao12s01 g748947 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .o(n_32502) );
ao12s01 g748948 ( .a(FE_OCP_RBN2328_delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_), .o(n_32501) );
na02s01 g748949 ( .a(n_32313), .b(n_46107), .o(n_32455) );
na02s02 TIMEBOOST_cell_4507 ( .a(n_6138), .b(n_5899), .o(TIMEBOOST_net_1344) );
na02s06 TIMEBOOST_cell_850 ( .a(n_6802), .b(TIMEBOOST_net_39), .o(n_6883) );
no02f08 TIMEBOOST_cell_3330 ( .a(n_31852), .b(n_31934), .o(TIMEBOOST_net_956) );
oa12s01 g748958 ( .a(n_31150), .b(n_31149), .c(n_31148), .o(n_31193) );
oa22s01 g748959 ( .a(n_32273), .b(n_31577), .c(n_32272), .d(n_31576), .o(n_32342) );
in01s01 g748962 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_21_), .o(n_32318) );
no02f10 g748967 ( .a(n_30919), .b(n_30858), .o(n_30967) );
in01f02 g748968 ( .a(n_30949), .o(n_30950) );
na02f04 g748969 ( .a(n_30919), .b(n_30744), .o(n_30949) );
no02m06 TIMEBOOST_cell_5521 ( .a(TIMEBOOST_net_1708), .b(n_6037), .o(n_6132) );
in01s01 g748973 ( .a(n_31132), .o(n_31153) );
no02m08 g748974 ( .a(n_31079), .b(n_30963), .o(n_31132) );
no02s06 g748975 ( .a(FE_OCP_RBN6841_n_31023), .b(n_27518), .o(n_31136) );
no02s03 g748976 ( .a(n_31023), .b(FE_OCPN1679_n_27315), .o(n_31108) );
na02s02 TIMEBOOST_cell_5528 ( .a(n_5957), .b(n_5688), .o(TIMEBOOST_net_1712) );
na02s04 g748978 ( .a(FE_OCP_RBN6832_n_31073), .b(FE_OCPN5262_n_27536), .o(n_31130) );
na02s02 g748979 ( .a(n_31073), .b(n_27518), .o(n_31105) );
na02s01 g748980 ( .a(n_30948), .b(n_31011), .o(n_31054) );
na03s04 TIMEBOOST_cell_849 ( .a(n_6801), .b(n_6645), .c(n_6831), .o(TIMEBOOST_net_39) );
in01s01 g748982 ( .a(n_31151), .o(n_31152) );
no02f06 g748983 ( .a(n_31126), .b(FE_OCP_DRV_N5149_n_31125), .o(n_31151) );
na02f06 g748984 ( .a(n_31126), .b(FE_OCP_DRV_N5149_n_31125), .o(n_31196) );
na02s01 g748985 ( .a(n_31149), .b(n_31148), .o(n_31150) );
ao12s01 g748987 ( .a(n_31454), .b(n_32295), .c(n_31511), .o(n_32316) );
in01s01 g748988 ( .a(n_32314), .o(n_32315) );
oa12s01 g748989 ( .a(n_31458), .b(n_32295), .c(n_31483), .o(n_32314) );
na02f04 TIMEBOOST_cell_5470 ( .a(n_39593), .b(FE_RN_1873_0), .o(TIMEBOOST_net_1683) );
in01s02 g748992 ( .a(n_31082), .o(n_31083) );
ao12s06 g748993 ( .a(FE_OCPN1340_n_27246), .b(n_31029), .c(n_30939), .o(n_31082) );
oa12f04 g748995 ( .a(n_30877), .b(n_30942), .c(n_31003), .o(n_31053) );
in01s01 g748996 ( .a(FE_OCP_RBN6084_n_31010), .o(n_31034) );
oa12s01 g749000 ( .a(n_30946), .b(n_30945), .c(n_30944), .o(n_31008) );
oa12s01 g749001 ( .a(n_31005), .b(n_31004), .c(n_31003), .o(n_31051) );
in01s02 g749004 ( .a(n_31099), .o(n_31100) );
in01s01 g749007 ( .a(n_31177), .o(n_31261) );
no02f08 g749008 ( .a(n_31095), .b(n_31094), .o(n_31177) );
oa12s01 g749009 ( .a(n_31124), .b(n_31123), .c(n_31122), .o(n_31176) );
oa22s01 g749010 ( .a(FE_OCP_RBN3438_n_32232), .b(n_31633), .c(n_32232), .d(n_31634), .o(n_32274) );
oa22s01 g749011 ( .a(n_32249), .b(n_31574), .c(n_32250), .d(n_31573), .o(n_32294) );
oa22s01 g749012 ( .a(n_32269), .b(n_31537), .c(n_32295), .d(n_31538), .o(n_32341) );
in01s01 g749014 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_22_), .o(n_32375) );
in01s01 g749017 ( .a(n_32312), .o(n_32313) );
no02s01 g749018 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .o(n_32312) );
na02f10 g749019 ( .a(n_30834), .b(n_30743), .o(n_30919) );
no02s02 g749025 ( .a(n_30961), .b(n_31025), .o(n_31032) );
na02m06 TIMEBOOST_cell_8486 ( .a(n_32928), .b(n_32682), .o(TIMEBOOST_net_2730) );
na02s06 g749027 ( .a(n_31029), .b(FE_OCPN1340_n_27246), .o(n_31030) );
na02s02 g749028 ( .a(n_30960), .b(n_27131), .o(n_31007) );
no02m04 g749029 ( .a(n_31026), .b(n_31025), .o(n_31027) );
na02s02 g749030 ( .a(n_31022), .b(n_30992), .o(n_31077) );
no02s02 g749031 ( .a(n_31075), .b(n_31074), .o(n_31076) );
in01s01 g749032 ( .a(n_30947), .o(n_30948) );
no02f02 g749033 ( .a(n_30918), .b(n_30917), .o(n_30947) );
na02s04 g749034 ( .a(n_30918), .b(FE_OCP_DRV_N1480_n_30917), .o(n_31011) );
na02s01 g749035 ( .a(n_30945), .b(n_30944), .o(n_30946) );
na02s01 g749036 ( .a(n_31004), .b(n_31003), .o(n_31005) );
no02f06 g749037 ( .a(n_31093), .b(n_31148), .o(n_31095) );
na02s01 g749038 ( .a(n_31123), .b(n_31122), .o(n_31124) );
no02s01 g749039 ( .a(n_31093), .b(n_31094), .o(n_31149) );
in01m01 g749040 ( .a(n_32292), .o(n_32293) );
oa12m02 g749041 ( .a(n_31543), .b(n_32231), .c(n_31541), .o(n_32292) );
oa12m04 g749043 ( .a(n_30855), .b(n_30883), .c(n_29896), .o(n_31001) );
na02s06 TIMEBOOST_cell_3849 ( .a(n_7107), .b(n_7106), .o(TIMEBOOST_net_1015) );
oa22s01 g749052 ( .a(n_32207), .b(n_31615), .c(n_32206), .d(n_31616), .o(n_32258) );
oa22s01 g749053 ( .a(n_32227), .b(n_31430), .c(n_32245), .d(n_31429), .o(n_32291) );
in01s01 g749054 ( .a(n_32272), .o(n_32273) );
oa12s01 g749055 ( .a(n_31387), .b(n_32227), .c(n_31411), .o(n_32272) );
in01s01 g749056 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .o(n_32271) );
in01s01 g749061 ( .a(n_32295), .o(n_32269) );
no02s02 g749062 ( .a(n_32230), .b(n_31542), .o(n_32295) );
na02s04 g749064 ( .a(n_30940), .b(n_30915), .o(n_30998) );
no02s04 g749065 ( .a(n_30996), .b(n_30995), .o(n_30997) );
no02m04 g749066 ( .a(n_30888), .b(n_30887), .o(n_30889) );
in01s01 g749067 ( .a(n_31075), .o(n_31022) );
no02s04 g749068 ( .a(n_30991), .b(n_27366), .o(n_31075) );
na02m08 TIMEBOOST_cell_8581 ( .a(TIMEBOOST_net_2777), .b(TIMEBOOST_net_655), .o(n_35099) );
no03s10 TIMEBOOST_cell_6516 ( .a(n_10826), .b(n_10778), .c(FE_OCPN4845_FE_OFN4779_n_44490), .o(n_10919) );
no02s02 g749071 ( .a(n_31021), .b(FE_OCP_DRV_N6897_FE_OCPN1679_n_27315), .o(n_31074) );
na02s01 g749072 ( .a(n_30991), .b(n_27366), .o(n_30992) );
in01m02 g749073 ( .a(n_31070), .o(n_31071) );
no02s01 g749077 ( .a(n_30878), .b(n_30942), .o(n_31004) );
na02s01 g749078 ( .a(n_30954), .b(n_31655), .o(n_30989) );
no02f04 g749079 ( .a(n_30978), .b(n_29555), .o(n_31093) );
no02m06 g749080 ( .a(n_30979), .b(n_29556), .o(n_31094) );
in01s01 g749081 ( .a(n_32249), .o(n_32250) );
oa12s01 g749082 ( .a(n_31569), .b(n_32205), .c(n_31409), .o(n_32249) );
in01f04 g749083 ( .a(n_30863), .o(n_30864) );
in01f04 g749084 ( .a(n_30834), .o(n_30863) );
oa12f08 g749085 ( .a(n_30751), .b(n_30750), .c(FE_OCPN5130_FE_OFN1198_n_27014), .o(n_30834) );
in01m02 g749087 ( .a(n_31018), .o(n_31048) );
in01s01 g749089 ( .a(n_30987), .o(n_30988) );
na02s06 TIMEBOOST_cell_4550 ( .a(TIMEBOOST_net_1365), .b(n_32241), .o(n_32305) );
in01s01 g749091 ( .a(n_30961), .o(n_30962) );
ao12s02 g749092 ( .a(FE_OCPN1404_n_30823), .b(n_30910), .c(n_30824), .o(n_30961) );
ao12m06 g749094 ( .a(n_30741), .b(n_30773), .c(FE_OCPN1298_n_30134), .o(n_30885) );
in01s06 g749097 ( .a(n_30960), .o(n_31029) );
na02f06 TIMEBOOST_cell_1112 ( .a(FE_RN_1656_0), .b(TIMEBOOST_net_170), .o(n_23348) );
ao12s01 g749100 ( .a(n_30833), .b(n_30862), .c(n_30832), .o(n_30945) );
in01s03 g749104 ( .a(n_46956), .o(n_31017) );
in01f04 g749107 ( .a(n_31026), .o(n_31081) );
na02f08 g749108 ( .a(n_30879), .b(n_30912), .o(n_31026) );
oa12s01 g749110 ( .a(n_31016), .b(n_31046), .c(n_31045), .o(n_31123) );
oa22s01 g749111 ( .a(n_32201), .b(n_31617), .c(n_32202), .d(n_31618), .o(n_32257) );
oa22s01 g749112 ( .a(n_32158), .b(n_31315), .c(n_32176), .d(n_31316), .o(n_32248) );
oa12s01 g749114 ( .a(n_31394), .b(n_32158), .c(n_31220), .o(n_32232) );
oa22s01 g749115 ( .a(n_32203), .b(n_31625), .c(n_32204), .d(n_31626), .o(n_32256) );
na02s02 TIMEBOOST_cell_7934 ( .a(n_5280), .b(n_4867), .o(TIMEBOOST_net_2598) );
no02m04 g749119 ( .a(n_30882), .b(FE_OCPN4853_n_29502), .o(n_30883) );
in01s02 g749120 ( .a(n_30996), .o(n_30940) );
no02s06 g749121 ( .a(n_30914), .b(n_27366), .o(n_30996) );
no02s06 g749122 ( .a(n_30939), .b(FE_OCPN1340_n_27246), .o(n_30995) );
na02s02 g749123 ( .a(n_30914), .b(n_27518), .o(n_30915) );
in01s02 g749124 ( .a(n_30937), .o(n_30938) );
na02s04 g749125 ( .a(n_30913), .b(n_30852), .o(n_30937) );
na02f06 TIMEBOOST_cell_1111 ( .a(n_23249), .b(FE_RN_1657_0), .o(TIMEBOOST_net_170) );
na02s04 TIMEBOOST_cell_4492 ( .a(TIMEBOOST_net_1336), .b(n_5866), .o(n_5972) );
na02s04 g749128 ( .a(n_30849), .b(n_27014), .o(n_30879) );
na02f06 g749129 ( .a(FE_OCP_RBN3140_n_30849), .b(FE_OCPN5300_n_27130), .o(n_30912) );
no02s06 g749130 ( .a(n_30847), .b(FE_OCPN5300_n_27130), .o(n_30963) );
na02m08 g749131 ( .a(n_30958), .b(FE_OCPN1340_n_27246), .o(n_31050) );
no02m06 g749133 ( .a(n_30958), .b(FE_OCP_DRV_N6897_FE_OCPN1679_n_27315), .o(n_31025) );
na02m04 TIMEBOOST_cell_7748 ( .a(n_25316), .b(n_24582), .o(TIMEBOOST_net_2505) );
na02m02 g749136 ( .a(n_30936), .b(FE_OCP_RBN5335_FE_RN_1144_0), .o(n_30956) );
no02f03 g749137 ( .a(n_30860), .b(FE_OCPN5242_n_30859), .o(n_30942) );
in01s01 g749138 ( .a(n_30877), .o(n_30878) );
na02f02 g749139 ( .a(n_30860), .b(FE_OCPN5252_n_30859), .o(n_30877) );
no02s01 g749140 ( .a(n_30862), .b(n_30832), .o(n_30833) );
na02s01 g749141 ( .a(n_31046), .b(n_31045), .o(n_31016) );
in01s01 g749143 ( .a(n_32206), .o(n_32207) );
ao12s01 g749144 ( .a(n_31529), .b(n_32116), .c(n_31570), .o(n_32206) );
in01m02 g749145 ( .a(n_32230), .o(n_32231) );
no02m04 g749146 ( .a(n_32205), .b(n_31453), .o(n_32230) );
in01s02 g749147 ( .a(n_30875), .o(n_30876) );
no02f08 TIMEBOOST_cell_7043 ( .a(n_39600), .b(n_45840), .o(TIMEBOOST_net_2280) );
in01s02 g749149 ( .a(n_30890), .o(n_30857) );
no02m04 g749150 ( .a(n_30772), .b(FE_OCPN5288_n_27315), .o(n_30890) );
oa12f06 g749151 ( .a(n_30747), .b(n_30714), .c(FE_OCPN5294_n_30584), .o(n_30751) );
in01m04 g749152 ( .a(n_30888), .o(n_30943) );
na02m08 g749153 ( .a(n_30774), .b(n_30749), .o(n_30888) );
in01s01 g749156 ( .a(FE_OCP_RBN6063_n_30908), .o(n_30955) );
na02s06 g749159 ( .a(n_30828), .b(n_30808), .o(n_30908) );
in01s06 g749162 ( .a(n_30933), .o(n_30954) );
na02s08 g749164 ( .a(n_30830), .b(n_30856), .o(n_30933) );
in01s02 g749165 ( .a(n_30991), .o(n_31021) );
no02m10 TIMEBOOST_cell_4298 ( .a(n_34164), .b(TIMEBOOST_net_1239), .o(n_34261) );
in01m02 g749167 ( .a(n_30978), .o(n_30979) );
oa22s01 g749169 ( .a(FE_OCP_RBN4490_n_32152), .b(n_31623), .c(n_32152), .d(n_31624), .o(n_32229) );
oa22s02 g749170 ( .a(n_32174), .b(n_31389), .c(n_32175), .d(n_31388), .o(n_32247) );
oa22s01 g749171 ( .a(n_32116), .b(n_31627), .c(n_32154), .d(n_31628), .o(n_32228) );
in01s01 g749173 ( .a(n_32227), .o(n_32245) );
oa12s02 g749174 ( .a(n_31513), .b(n_32115), .c(n_31432), .o(n_32227) );
in01s01 g749175 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_15_), .o(n_32422) );
in01s01 g749178 ( .a(n_32203), .o(n_32204) );
in01s01 g749179 ( .a(n_32205), .o(n_32203) );
no02m06 g749180 ( .a(n_32114), .b(n_31512), .o(n_32205) );
na02s06 g749181 ( .a(n_30347), .b(n_30807), .o(n_30856) );
na02s03 g749182 ( .a(n_30806), .b(n_30348), .o(n_30830) );
na02s03 g749183 ( .a(n_30801), .b(FE_OCPN4853_n_29502), .o(n_30855) );
in01f02 g749185 ( .a(n_30750), .o(n_30776) );
no02f08 g749186 ( .a(n_30714), .b(FE_OCP_RBN7045_FE_RN_1462_0), .o(n_30750) );
na02m08 g749188 ( .a(n_30800), .b(n_30319), .o(n_30882) );
no02s06 g749189 ( .a(n_30771), .b(FE_OCP_DRV_N7081_n_27130), .o(n_30858) );
na02s08 g749190 ( .a(n_30829), .b(FE_OCPN5288_n_27315), .o(n_30913) );
na02m06 g749191 ( .a(FE_OCP_RBN6023_n_30711), .b(n_27131), .o(n_30774) );
na02s04 g749192 ( .a(n_30711), .b(n_27014), .o(n_30749) );
in01s02 g749193 ( .a(n_30887), .o(n_30852) );
no02m04 g749194 ( .a(n_30829), .b(FE_OCPN5288_n_27315), .o(n_30887) );
na02s01 TIMEBOOST_cell_4486 ( .a(TIMEBOOST_net_1333), .b(n_5798), .o(n_5895) );
na02s06 g749197 ( .a(n_30818), .b(FE_OCPN1402_FE_OFN1196_n_27014), .o(n_30936) );
na02s02 g749198 ( .a(n_30820), .b(FE_OCPN1340_n_27246), .o(n_30851) );
no02m06 TIMEBOOST_cell_3107 ( .a(n_10422), .b(TIMEBOOST_net_844), .o(n_10551) );
na02s03 g749200 ( .a(n_30763), .b(FE_OCPN1928_n_30385), .o(n_30808) );
na02s02 g749201 ( .a(n_30739), .b(FE_OCPN1927_n_30385), .o(n_30828) );
na02m08 g749202 ( .a(n_30739), .b(n_45489), .o(n_30773) );
no02s02 g749203 ( .a(n_30771), .b(FE_OCP_RBN6016_n_30625), .o(n_30772) );
no02m06 TIMEBOOST_cell_6298 ( .a(TIMEBOOST_net_2000), .b(n_10970), .o(n_11128) );
in01s04 g749206 ( .a(n_30914), .o(n_30939) );
na02f04 g749210 ( .a(n_30713), .b(n_30683), .o(n_30862) );
in01s01 g749219 ( .a(FE_OCP_RBN3141_n_30849), .o(n_30906) );
no02m06 TIMEBOOST_cell_3144 ( .a(FE_RN_670_0), .b(FE_RN_669_0), .o(TIMEBOOST_net_863) );
in01s01 g749225 ( .a(n_32201), .o(n_32202) );
oa12s01 g749226 ( .a(n_31283), .b(n_32156), .c(n_31368), .o(n_32201) );
in01s01 g749228 ( .a(n_32158), .o(n_32176) );
oa12s01 g749229 ( .a(n_31418), .b(n_32094), .c(n_31313), .o(n_32158) );
in01f02 g749230 ( .a(n_30847), .o(n_30910) );
in01s01 g749233 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .o(n_30905) );
in01s01 g749235 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_13_), .o(n_32157) );
in01s02 g749238 ( .a(n_32174), .o(n_32175) );
na02s04 g749239 ( .a(n_32156), .b(n_31374), .o(n_32174) );
in01s01 g749241 ( .a(n_32116), .o(n_32154) );
na02s01 g749242 ( .a(n_32094), .b(n_31457), .o(n_32116) );
in01s01 g749243 ( .a(n_32114), .o(n_32115) );
no02s06 g749244 ( .a(n_32094), .b(n_31456), .o(n_32114) );
in01s04 g749245 ( .a(n_30806), .o(n_30807) );
no02s06 g749246 ( .a(n_30765), .b(FE_OCP_DRV_N3512_n_30318), .o(n_30806) );
na02f01 g749247 ( .a(n_30652), .b(n_30537), .o(n_30683) );
na02f02 g749248 ( .a(n_30653), .b(n_30559), .o(n_30713) );
no02f08 g749249 ( .a(n_30630), .b(n_30659), .o(n_30714) );
in01m02 g749251 ( .a(n_30904), .o(n_30926) );
no02m08 g749252 ( .a(n_30843), .b(n_30841), .o(n_30904) );
in01s02 g749255 ( .a(n_30766), .o(n_30767) );
na02m04 g749256 ( .a(n_30744), .b(n_30743), .o(n_30766) );
na02m02 g749257 ( .a(n_30824), .b(FE_OCPN1404_n_30823), .o(n_30825) );
no02m04 TIMEBOOST_cell_6287 ( .a(n_10054), .b(n_10134), .o(TIMEBOOST_net_1995) );
no02s06 TIMEBOOST_cell_5395 ( .a(TIMEBOOST_net_1645), .b(TIMEBOOST_net_484), .o(n_46956) );
na02s02 TIMEBOOST_cell_4394 ( .a(TIMEBOOST_net_1287), .b(n_4604), .o(n_4782) );
na02s02 TIMEBOOST_cell_1095 ( .a(n_23437), .b(n_23059), .o(TIMEBOOST_net_162) );
no02m06 g749264 ( .a(n_30677), .b(n_45489), .o(n_30741) );
na02s01 g749265 ( .a(FE_OCP_RBN1859_n_30731), .b(FE_OCP_RBN3079_n_30643), .o(n_30803) );
ao12s02 g749267 ( .a(n_31527), .b(n_32063), .c(n_31571), .o(n_32152) );
in01s02 g749268 ( .a(n_30800), .o(n_30801) );
na02m08 g749269 ( .a(n_30272), .b(n_30765), .o(n_30800) );
in01f02 g749270 ( .a(n_30869), .o(n_30870) );
no02f04 g749271 ( .a(n_30843), .b(n_30760), .o(n_30869) );
in01s02 g749273 ( .a(n_30739), .o(n_30763) );
na02s02 TIMEBOOST_cell_3278 ( .a(FE_RN_574_0), .b(n_20973), .o(TIMEBOOST_net_930) );
in01s01 g749281 ( .a(n_30842), .o(n_31655) );
in01s02 g749282 ( .a(n_30820), .o(n_30842) );
ao22s02 g749283 ( .a(n_30670), .b(n_30320), .c(n_30698), .d(n_30321), .o(n_30820) );
oa22s01 g749286 ( .a(n_32006), .b(n_31619), .c(n_32007), .d(n_31620), .o(n_32093) );
oa22s01 g749287 ( .a(n_32063), .b(n_31629), .c(n_32035), .d(n_31630), .o(n_32173) );
in01s01 g749288 ( .a(n_30771), .o(n_30737) );
na02m08 g749289 ( .a(n_30656), .b(n_30629), .o(n_30771) );
na02s06 g749290 ( .a(n_32063), .b(n_31318), .o(n_32156) );
no02m08 g749291 ( .a(n_30294), .b(n_30670), .o(n_30765) );
in01f02 g749292 ( .a(n_30657), .o(n_30658) );
in01f01 g749293 ( .a(n_30630), .o(n_30657) );
na02f06 g749294 ( .a(n_30611), .b(n_30537), .o(n_30630) );
in01m02 g749296 ( .a(n_30841), .o(n_30867) );
na02m08 g749297 ( .a(n_30621), .b(n_30817), .o(n_30841) );
na02m06 g749298 ( .a(FE_OCP_RBN6813_n_30608), .b(n_27014), .o(n_30656) );
na02s04 g749299 ( .a(n_30608), .b(n_27062), .o(n_30629) );
na02s06 g749300 ( .a(n_30625), .b(FE_OFN1198_n_27014), .o(n_30743) );
na02m02 TIMEBOOST_cell_4495 ( .a(n_11081), .b(n_10987), .o(TIMEBOOST_net_1338) );
no02f06 TIMEBOOST_cell_4480 ( .a(TIMEBOOST_net_1330), .b(n_25915), .o(TIMEBOOST_net_1151) );
na02m02 g749303 ( .a(FE_OCP_RBN6016_n_30625), .b(n_27131), .o(n_30744) );
no02f02 g749305 ( .a(FE_OCP_RBN7044_FE_RN_1462_0), .b(n_30659), .o(n_30706) );
no02m02 g749307 ( .a(n_30727), .b(FE_OCPN1402_FE_OFN1196_n_27014), .o(n_30760) );
na02s02 g749309 ( .a(n_30655), .b(FE_OCPN5105_n_30371), .o(n_30678) );
in01s02 g749310 ( .a(n_30676), .o(n_30677) );
no02m08 g749311 ( .a(n_30655), .b(n_30343), .o(n_30676) );
na02f04 g749314 ( .a(n_30758), .b(n_29441), .o(n_30799) );
in01m03 g749316 ( .a(n_30735), .o(n_30736) );
no02m06 g749317 ( .a(n_30650), .b(n_30261), .o(n_30735) );
na02s06 g749318 ( .a(n_32008), .b(n_31390), .o(n_32094) );
in01f01 g749319 ( .a(n_30652), .o(n_30653) );
na02f01 g749320 ( .a(n_30585), .b(n_30611), .o(n_30652) );
na02f04 g749322 ( .a(n_30791), .b(n_30817), .o(n_30865) );
oa12s01 g749323 ( .a(n_30673), .b(n_30672), .c(n_30671), .o(n_30734) );
na02f08 g749332 ( .a(n_30586), .b(n_30566), .o(n_30747) );
in01s06 g749339 ( .a(n_46958), .o(n_30814) );
oa12s01 g749342 ( .a(n_31122), .b(n_30693), .c(n_29229), .o(n_30813) );
oa22s01 g749343 ( .a(n_31977), .b(n_31568), .c(n_31978), .d(n_31567), .o(n_32065) );
oa22s01 g749344 ( .a(n_31979), .b(n_31369), .c(n_31980), .d(n_31370), .o(n_32064) );
no02m08 g749346 ( .a(n_30674), .b(n_30701), .o(n_30824) );
no02m04 g749349 ( .a(n_30624), .b(n_30262), .o(n_30650) );
na02s06 g749351 ( .a(n_30644), .b(FE_OCPN1332_n_30281), .o(n_30675) );
no02s06 g749352 ( .a(n_30580), .b(FE_OCPN5294_n_30584), .o(n_30659) );
na02f04 g749353 ( .a(n_30542), .b(FE_OCPN5130_FE_OFN1198_n_27014), .o(n_30611) );
na02f08 g749354 ( .a(n_30540), .b(n_30790), .o(n_30586) );
na02m04 g749355 ( .a(n_30541), .b(FE_OCPN5130_FE_OFN1198_n_27014), .o(n_30566) );
na02f02 g749357 ( .a(n_30543), .b(n_30584), .o(n_30585) );
no02s04 g749358 ( .a(n_30643), .b(FE_OFN1196_n_27014), .o(n_30674) );
no02m08 g749359 ( .a(FE_OCP_RBN3079_n_30643), .b(FE_OCPN1677_n_27062), .o(n_30701) );
na02m08 g749360 ( .a(n_30723), .b(FE_OCPN1402_FE_OFN1196_n_27014), .o(n_30817) );
na02f04 g749361 ( .a(n_30724), .b(FE_RN_1313_0), .o(n_30791) );
na02m08 g749364 ( .a(n_30349), .b(n_30582), .o(n_30655) );
na02s01 g749365 ( .a(n_30672), .b(n_30671), .o(n_30673) );
na02f04 g749366 ( .a(n_30622), .b(n_30671), .o(n_30944) );
in01s04 g749367 ( .a(n_30758), .o(n_31122) );
no02f04 g749368 ( .a(n_30692), .b(n_29228), .o(n_30758) );
in01s04 g749371 ( .a(n_32035), .o(n_32063) );
in01s02 g749373 ( .a(n_32008), .o(n_32035) );
oa12f06 g749374 ( .a(n_31348), .b(n_31981), .c(n_31341), .o(n_32008) );
in01s01 g749376 ( .a(n_30670), .o(n_30698) );
na03m80 TIMEBOOST_cell_5690 ( .a(n_32615), .b(n_44962), .c(n_32632), .o(TIMEBOOST_net_686) );
in01m04 g749378 ( .a(n_30609), .o(n_30610) );
no02m06 g749379 ( .a(n_30544), .b(n_30278), .o(n_30609) );
in01s01 g749394 ( .a(n_30729), .o(n_30757) );
in01s01 g749395 ( .a(n_30697), .o(n_30729) );
in01s01 g749400 ( .a(n_32006), .o(n_32007) );
oa12s01 g749401 ( .a(n_31343), .b(n_31981), .c(n_31279), .o(n_32006) );
in01s01 g749403 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_), .o(n_32034) );
in01s01 g749405 ( .a(n_31979), .o(n_31980) );
na02s01 g749406 ( .a(n_31981), .b(n_31276), .o(n_31979) );
in01m04 g749408 ( .a(n_30624), .o(n_30644) );
na02m08 g749409 ( .a(n_30603), .b(n_30295), .o(n_30624) );
no02m06 g749410 ( .a(n_30514), .b(n_30277), .o(n_30544) );
na02s06 g749412 ( .a(n_30535), .b(n_30292), .o(n_30564) );
in01s01 g749413 ( .a(n_31977), .o(n_31978) );
oa12s01 g749414 ( .a(n_31572), .b(n_31911), .c(n_31321), .o(n_31977) );
oa12f04 g749415 ( .a(n_30217), .b(n_30578), .c(FE_OCPN1270_n_30577), .o(n_30605) );
no02m02 TIMEBOOST_cell_6084 ( .a(TIMEBOOST_net_1893), .b(n_38615), .o(TIMEBOOST_net_1515) );
no02s04 TIMEBOOST_cell_7686 ( .a(n_8512), .b(n_8575), .o(TIMEBOOST_net_2474) );
in01s02 g749419 ( .a(n_30582), .o(n_30601) );
na02f04 TIMEBOOST_cell_7992 ( .a(FE_OCP_RBN6069_n_26140), .b(n_26124), .o(TIMEBOOST_net_2627) );
in01s01 g749421 ( .a(n_30622), .o(n_30672) );
na02s10 TIMEBOOST_cell_948 ( .a(TIMEBOOST_net_88), .b(n_17827), .o(n_17971) );
na02f06 g749424 ( .a(n_30515), .b(n_30502), .o(n_30580) );
in01f01 g749425 ( .a(n_30542), .o(n_30543) );
in01s01 g749428 ( .a(n_30541), .o(n_31864) );
in01f04 g749429 ( .a(n_30541), .o(n_30540) );
no02m06 TIMEBOOST_cell_6118 ( .a(TIMEBOOST_net_1910), .b(n_19642), .o(n_19752) );
in01s01 g749438 ( .a(n_30692), .o(n_30693) );
in01m02 g749440 ( .a(n_30723), .o(n_30724) );
na02m04 TIMEBOOST_cell_4534 ( .a(TIMEBOOST_net_1357), .b(n_11161), .o(n_11278) );
oa22s01 g749442 ( .a(n_31939), .b(n_31621), .c(n_31940), .d(n_31622), .o(n_32005) );
oa22s01 g749443 ( .a(n_31941), .b(n_31631), .c(n_31911), .d(n_31632), .o(n_32004) );
no02s02 TIMEBOOST_cell_6015 ( .a(n_13111), .b(n_13197), .o(TIMEBOOST_net_1859) );
no02m04 g749445 ( .a(n_30578), .b(n_30263), .o(n_30576) );
no03f08 TIMEBOOST_cell_8444 ( .a(n_26328), .b(n_44443), .c(TIMEBOOST_net_2044), .o(n_26531) );
no02f08 TIMEBOOST_cell_3155 ( .a(TIMEBOOST_net_868), .b(n_42843), .o(n_42896) );
na03s10 TIMEBOOST_cell_947 ( .a(n_17802), .b(n_17894), .c(n_17930), .o(TIMEBOOST_net_88) );
na02f04 g749449 ( .a(FE_OCP_RBN2104_n_30465), .b(FE_OFN1199_n_27014), .o(n_30515) );
na02s04 g749450 ( .a(n_30465), .b(n_30466), .o(n_30502) );
in01s01 g749452 ( .a(n_30537), .o(n_30559) );
na02f06 g749453 ( .a(n_30500), .b(FE_OCPN5130_FE_OFN1198_n_27014), .o(n_30537) );
in01s01 g749455 ( .a(n_30621), .o(n_30640) );
na02m06 g749456 ( .a(n_30575), .b(FE_OCPN1402_FE_OFN1196_n_27014), .o(n_30621) );
na02m02 TIMEBOOST_cell_4533 ( .a(n_11096), .b(n_10921), .o(TIMEBOOST_net_1357) );
na02m04 TIMEBOOST_cell_4496 ( .a(TIMEBOOST_net_1338), .b(n_11130), .o(n_11252) );
in01s04 g749460 ( .a(n_30514), .o(n_30535) );
na02s08 g749461 ( .a(n_30467), .b(n_30210), .o(n_30514) );
na02f08 g749462 ( .a(n_31888), .b(n_31323), .o(n_31981) );
na02s04 TIMEBOOST_cell_3098 ( .a(n_25168), .b(n_25143), .o(TIMEBOOST_net_840) );
na02m08 TIMEBOOST_cell_4919 ( .a(TIMEBOOST_net_1407), .b(n_7060), .o(n_7127) );
oa12s02 g749467 ( .a(FE_OCP_RBN6747_n_30170), .b(n_30471), .c(FE_OCPN1238_n_30470), .o(n_30501) );
na02m06 TIMEBOOST_cell_1080 ( .a(TIMEBOOST_net_154), .b(n_12516), .o(FE_RN_1390_0) );
in01s01 g749469 ( .a(FE_OCP_RBN6001_n_30534), .o(n_30557) );
na02m06 g749472 ( .a(n_30455), .b(n_30469), .o(n_30534) );
na02m20 TIMEBOOST_cell_802 ( .a(TIMEBOOST_net_15), .b(n_22769), .o(n_22822) );
oa22s01 g749476 ( .a(n_31909), .b(n_31319), .c(n_31910), .d(n_31320), .o(n_31976) );
oa22s01 g749477 ( .a(n_31886), .b(n_31564), .c(n_31885), .d(n_31565), .o(n_31960) );
no02s01 TIMEBOOST_cell_8696 ( .a(n_37118), .b(n_37119), .o(TIMEBOOST_net_2835) );
na02f04 TIMEBOOST_cell_5633 ( .a(TIMEBOOST_net_1764), .b(n_16670), .o(n_16810) );
no02s03 TIMEBOOST_cell_4273 ( .a(FE_RN_778_0), .b(n_1976), .o(TIMEBOOST_net_1227) );
na02s06 TIMEBOOST_cell_1079 ( .a(FE_RN_1387_0), .b(FE_RN_1388_0), .o(TIMEBOOST_net_154) );
na02m02 g749483 ( .a(n_30452), .b(n_30240), .o(n_30455) );
na02m04 g749484 ( .a(n_30471), .b(n_30239), .o(n_30469) );
in01s01 g749486 ( .a(n_31911), .o(n_31941) );
in01s01 g749487 ( .a(n_31888), .o(n_31911) );
oa12f06 g749488 ( .a(n_31350), .b(n_31782), .c(n_31286), .o(n_31888) );
in01m04 g749489 ( .a(n_30558), .o(n_30578) );
oa12f08 g749490 ( .a(n_30203), .b(n_30498), .c(n_30202), .o(n_30558) );
in01m04 g749491 ( .a(n_30453), .o(n_30454) );
no02f08 g749492 ( .a(n_30411), .b(n_30050), .o(n_30453) );
in01s02 g749493 ( .a(n_30467), .o(n_30468) );
in01m02 g749495 ( .a(n_30510), .o(n_30511) );
in01f01 g749496 ( .a(n_30500), .o(n_30510) );
na02f06 g749501 ( .a(n_30410), .b(n_30429), .o(n_30465) );
in01s01 g749507 ( .a(n_31599), .o(n_30637) );
in01s01 g749508 ( .a(n_30598), .o(n_31599) );
in01s02 g749509 ( .a(n_30598), .o(n_30597) );
na02s20 TIMEBOOST_cell_804 ( .a(TIMEBOOST_net_16), .b(n_11786), .o(n_11927) );
in01s01 g749514 ( .a(n_31939), .o(n_31940) );
no02s04 TIMEBOOST_cell_5496 ( .a(n_10563), .b(n_10525), .o(TIMEBOOST_net_1696) );
in01s01 g749516 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_7_), .o(n_31887) );
in01s01 g749518 ( .a(n_31909), .o(n_31910) );
na02s01 g749519 ( .a(n_31816), .b(n_31292), .o(n_31909) );
no02m04 TIMEBOOST_cell_3125 ( .a(TIMEBOOST_net_853), .b(n_34858), .o(n_34923) );
no02f06 TIMEBOOST_cell_3101 ( .a(n_25868), .b(TIMEBOOST_net_841), .o(n_25904) );
na04s01 TIMEBOOST_cell_8411 ( .a(n_27031), .b(n_26886), .c(n_26887), .d(n_27032), .o(n_27094) );
in01f03 g749523 ( .a(n_30530), .o(n_30508) );
na02f08 g749524 ( .a(n_30498), .b(n_30071), .o(n_30530) );
no02f04 g749525 ( .a(n_30409), .b(n_30116), .o(n_30411) );
na02f04 g749526 ( .a(n_30409), .b(n_30144), .o(n_30410) );
in01s01 g749530 ( .a(n_31885), .o(n_31886) );
no02s01 g749531 ( .a(n_31781), .b(n_31509), .o(n_31885) );
in01m04 g749532 ( .a(n_30452), .o(n_30471) );
na02s01 TIMEBOOST_cell_8844 ( .a(n_42826), .b(n_42825), .o(TIMEBOOST_net_2909) );
in01s01 g749534 ( .a(FE_OCPN5254_n_31871), .o(n_30554) );
oa12s01 g749535 ( .a(n_30495), .b(n_30494), .c(n_30493), .o(n_31871) );
oa22s01 g749536 ( .a(n_31752), .b(n_31535), .c(n_31780), .d(n_31534), .o(n_31856) );
in01s01 g749537 ( .a(n_31815), .o(n_31816) );
in01s01 g749538 ( .a(n_31782), .o(n_31815) );
na02f06 g749539 ( .a(n_31709), .b(n_31212), .o(n_31782) );
no02s01 g749540 ( .a(n_31780), .b(n_31510), .o(n_31781) );
in01s02 g749541 ( .a(n_30496), .o(n_30497) );
na02m06 g749542 ( .a(n_30437), .b(n_30120), .o(n_30496) );
na02f08 g749543 ( .a(n_30436), .b(n_30114), .o(n_30498) );
na02s01 g749544 ( .a(n_30494), .b(n_30493), .o(n_30495) );
no02s01 g749547 ( .a(n_30527), .b(n_30526), .o(n_30528) );
na02s01 g749548 ( .a(n_30527), .b(n_30526), .o(n_30525) );
oa12f02 g749549 ( .a(n_30051), .b(n_45631), .c(n_30356), .o(n_30379) );
na02m04 TIMEBOOST_cell_6796 ( .a(TIMEBOOST_net_2155), .b(n_5076), .o(n_5255) );
na02m08 TIMEBOOST_cell_6603 ( .a(FE_OCP_RBN984_n_22822), .b(n_22931), .o(TIMEBOOST_net_2059) );
in01s01 g749552 ( .a(n_30428), .o(n_31804) );
in01s01 g749555 ( .a(n_31502), .o(n_30553) );
ao12s01 g749556 ( .a(n_30490), .b(n_30489), .c(n_30488), .o(n_31502) );
in01s01 g749562 ( .a(n_30573), .o(n_30593) );
oa12s01 g749563 ( .a(n_30487), .b(n_30486), .c(n_30485), .o(n_30573) );
in01s01 g749564 ( .a(n_31770), .o(n_30426) );
ao12s01 g749565 ( .a(n_30378), .b(n_30377), .c(n_30376), .o(n_31770) );
oa22s01 g749566 ( .a(n_31692), .b(n_31532), .c(n_31693), .d(n_31533), .o(n_31779) );
in01m02 g749568 ( .a(n_30436), .o(n_30437) );
no02f08 g749569 ( .a(n_30405), .b(n_30010), .o(n_30436) );
no02s01 g749570 ( .a(n_30489), .b(n_30488), .o(n_30490) );
na02s02 TIMEBOOST_cell_6825 ( .a(n_6290), .b(n_5852), .o(TIMEBOOST_net_2170) );
in01m04 g749572 ( .a(n_30354), .o(n_30355) );
na02f08 g749573 ( .a(n_30302), .b(n_30046), .o(n_30354) );
na02s01 g749574 ( .a(n_30486), .b(n_30485), .o(n_30487) );
no02s01 g749575 ( .a(n_30377), .b(n_30376), .o(n_30378) );
in01s01 g749576 ( .a(n_31780), .o(n_31752) );
in01s01 g749577 ( .a(n_31709), .o(n_31780) );
ao12f06 g749578 ( .a(n_31186), .b(n_31672), .c(n_31257), .o(n_31709) );
ao12s01 g749579 ( .a(n_30017), .b(n_30285), .c(n_30021), .o(n_30494) );
in01s01 g749580 ( .a(n_30527), .o(n_30506) );
ao12s01 g749581 ( .a(n_30449), .b(n_30448), .c(n_30447), .o(n_30527) );
oa12s01 g749582 ( .a(n_30408), .b(n_30407), .c(n_30406), .o(n_31448) );
in01s01 g749584 ( .a(n_31692), .o(n_31693) );
na02s01 g749585 ( .a(n_31672), .b(n_31221), .o(n_31692) );
na02s01 g749586 ( .a(n_30407), .b(n_30406), .o(n_30408) );
no02s01 g749587 ( .a(n_30448), .b(n_30447), .o(n_30449) );
na02s01 g749588 ( .a(n_30286), .b(n_30016), .o(n_30377) );
in01m02 g749589 ( .a(n_30424), .o(n_30425) );
in01m02 g749590 ( .a(n_30405), .o(n_30424) );
ao12f08 g749591 ( .a(n_30054), .b(n_30375), .c(n_29987), .o(n_30405) );
na02s01 g749592 ( .a(n_30374), .b(n_30020), .o(n_30489) );
oa12f08 g749597 ( .a(n_30055), .b(n_30483), .c(n_30022), .o(n_30302) );
oa12s01 g749598 ( .a(n_30421), .b(n_30483), .c(n_30443), .o(n_30486) );
in01s01 g749599 ( .a(FE_OCPN1276_n_31773), .o(n_30522) );
ao12s01 g749600 ( .a(n_30462), .b(n_30461), .c(n_30460), .o(n_31773) );
in01s01 g749601 ( .a(FE_RN_1883_0), .o(n_30592) );
oa12s01 g749602 ( .a(n_30484), .b(n_30483), .c(n_30482), .o(n_30572) );
oa12s01 g749603 ( .a(n_31581), .b(n_31582), .c(n_31580), .o(n_31671) );
na02f06 g749604 ( .a(n_31582), .b(n_31222), .o(n_31672) );
na02s01 g749605 ( .a(n_31582), .b(n_31580), .o(n_31581) );
no02s01 g749606 ( .a(n_30375), .b(n_30019), .o(n_30407) );
na02s01 g749607 ( .a(n_29982), .b(n_30375), .o(n_30374) );
no02s01 g749608 ( .a(n_30461), .b(n_30460), .o(n_30462) );
in01s01 g749609 ( .a(n_30285), .o(n_30286) );
no02s01 g749610 ( .a(n_30483), .b(n_29953), .o(n_30285) );
na02s01 g749611 ( .a(n_30483), .b(n_30482), .o(n_30484) );
na02s01 g749612 ( .a(n_30299), .b(n_32076), .o(n_30300) );
ao12s01 g749614 ( .a(n_30383), .b(n_30445), .c(n_30423), .o(n_30448) );
ao12s01 g749615 ( .a(n_30459), .b(n_30458), .c(n_30457), .o(n_31504) );
in01s01 g749616 ( .a(n_30526), .o(n_30505) );
ao12s01 g749617 ( .a(n_30446), .b(n_30445), .c(n_30444), .o(n_30526) );
oa12s01 g749618 ( .a(n_31645), .b(n_31644), .c(n_31643), .o(n_31691) );
na02s01 g749620 ( .a(n_31644), .b(n_31643), .o(n_31645) );
no02s01 g749621 ( .a(n_30458), .b(n_30457), .o(n_30459) );
no02s01 g749622 ( .a(n_30445), .b(n_30444), .o(n_30446) );
no02f08 g749623 ( .a(n_30298), .b(n_29915), .o(n_30375) );
na02f06 g749624 ( .a(n_31461), .b(n_31169), .o(n_31582) );
ao12s01 g749625 ( .a(n_29986), .b(n_30250), .c(n_29920), .o(n_30461) );
oa12f08 g749626 ( .a(n_29963), .b(n_30180), .c(n_29988), .o(n_30483) );
in01s01 g749627 ( .a(n_30299), .o(n_30327) );
oa12s01 g749628 ( .a(n_30227), .b(n_30226), .c(n_30225), .o(n_30299) );
oa22s01 g749630 ( .a(n_30204), .b(n_30015), .c(n_30250), .d(n_30014), .o(n_31740) );
na02f04 g749631 ( .a(n_31433), .b(n_31460), .o(n_31461) );
na02s01 g749632 ( .a(n_31434), .b(n_31536), .o(n_31644) );
na02s01 g749635 ( .a(n_30226), .b(n_30225), .o(n_30227) );
oa12s01 g749636 ( .a(n_29965), .b(n_30283), .c(n_29899), .o(n_30458) );
in01s01 g749637 ( .a(n_30298), .o(n_30445) );
oa12f08 g749638 ( .a(n_29929), .b(n_30283), .c(n_29967), .o(n_30298) );
oa12s01 g749640 ( .a(n_30266), .b(n_30283), .c(n_30265), .o(n_30322) );
oa12s01 g749641 ( .a(n_31642), .b(n_31641), .c(n_31640), .o(n_31690) );
in01s01 g749642 ( .a(n_31433), .o(n_31434) );
no02f04 g749643 ( .a(n_31396), .b(n_31143), .o(n_31433) );
na02s01 g749644 ( .a(n_31641), .b(n_31640), .o(n_31642) );
in01s01 g749645 ( .a(n_30250), .o(n_30204) );
in01s01 g749646 ( .a(n_30180), .o(n_30250) );
oa12f08 g749647 ( .a(n_29989), .b(n_30080), .c(n_29962), .o(n_30180) );
na02s01 g749648 ( .a(n_30283), .b(n_30265), .o(n_30266) );
in01s01 g749649 ( .a(n_30324), .o(n_30350) );
oa12s01 g749650 ( .a(n_30249), .b(n_30248), .c(n_30247), .o(n_30324) );
in01s01 g749651 ( .a(n_32076), .o(n_30326) );
na02s01 g749652 ( .a(n_30179), .b(n_30155), .o(n_32076) );
oa12s01 g749653 ( .a(n_29984), .b(n_30154), .c(n_29916), .o(n_30226) );
in01s01 g749654 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_), .o(n_31778) );
na02s01 g749656 ( .a(n_30248), .b(n_30247), .o(n_30249) );
na02s01 g749657 ( .a(n_30154), .b(n_30012), .o(n_30155) );
na02s01 g749658 ( .a(n_30121), .b(n_30013), .o(n_30179) );
ao12s01 g749659 ( .a(n_31542), .b(n_31459), .c(n_31311), .o(n_31543) );
in01s01 g749660 ( .a(n_31396), .o(n_31641) );
ao12f04 g749661 ( .a(n_31258), .b(n_31295), .c(FE_OCP_RBN4419_n_31117), .o(n_31396) );
na02f08 g749662 ( .a(n_30178), .b(n_29969), .o(n_30283) );
na02f08 g749663 ( .a(n_30149), .b(n_29968), .o(n_30178) );
na02s01 g749664 ( .a(n_30150), .b(n_29925), .o(n_30248) );
no02s01 g749665 ( .a(n_31512), .b(n_31392), .o(n_31513) );
in01s01 g749666 ( .a(n_30154), .o(n_30121) );
in01s01 g749667 ( .a(n_30080), .o(n_30154) );
ao12f08 g749668 ( .a(n_29888), .b(n_30057), .c(n_29955), .o(n_30080) );
in01s01 g749669 ( .a(n_30224), .o(n_31795) );
oa12s01 g749670 ( .a(n_30153), .b(n_30152), .c(n_30151), .o(n_30224) );
oa12s01 g749671 ( .a(n_30026), .b(n_30057), .c(n_30025), .o(n_31719) );
oa12s01 g749672 ( .a(n_31639), .b(n_31638), .c(n_31637), .o(n_31689) );
na02f04 g749674 ( .a(n_31259), .b(n_31294), .o(n_31295) );
na02s01 g749675 ( .a(n_31638), .b(n_31637), .o(n_31639) );
na02s01 g749676 ( .a(n_30152), .b(n_30151), .o(n_30153) );
in01s01 g749677 ( .a(n_30149), .o(n_30150) );
no02f08 g749678 ( .a(n_30079), .b(n_29862), .o(n_30149) );
na02s01 g749679 ( .a(n_30057), .b(n_30025), .o(n_30026) );
na02s01 g749680 ( .a(n_31458), .b(n_31481), .o(n_31459) );
na02s01 g749681 ( .a(n_31482), .b(n_31540), .o(n_31541) );
oa12s02 g749682 ( .a(n_31347), .b(n_31457), .c(n_31456), .o(n_31512) );
in01s06 g749683 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_1_), .o(n_32356) );
in01s01 g749685 ( .a(n_31259), .o(n_31638) );
no02m06 g749686 ( .a(n_31191), .b(n_31114), .o(n_31259) );
no02m04 g749687 ( .a(n_31192), .b(n_31294), .o(n_31258) );
no02s01 g749688 ( .a(n_31395), .b(n_31346), .o(n_31418) );
na02s01 g749689 ( .a(n_31412), .b(n_31391), .o(n_31542) );
in01s01 g749690 ( .a(n_31482), .o(n_31483) );
no02s01 g749691 ( .a(n_31455), .b(n_31454), .o(n_31482) );
oa12f08 g749692 ( .a(FE_OCP_RBN6706_n_29787), .b(n_29970), .c(n_29859), .o(n_30057) );
oa12s01 g749693 ( .a(n_30024), .b(n_30056), .c(n_30023), .o(n_31473) );
in01s01 g749694 ( .a(n_30079), .o(n_30152) );
oa12f08 g749695 ( .a(n_29872), .b(n_30056), .c(n_29832), .o(n_30079) );
ao12s01 g749696 ( .a(n_29931), .b(n_29970), .c(n_29930), .o(n_31676) );
in01s01 g749697 ( .a(n_31578), .o(n_31579) );
ao12s01 g749698 ( .a(n_31455), .b(n_31417), .c(n_31311), .o(n_31578) );
na02s01 g749699 ( .a(n_31415), .b(n_31431), .o(n_31453) );
oa12s01 g749700 ( .a(n_31229), .b(n_31228), .c(n_31227), .o(n_31293) );
oa12s01 g749701 ( .a(n_31311), .b(n_31417), .c(n_31416), .o(n_31458) );
in01s01 g749702 ( .a(n_31635), .o(n_31636) );
oa12s01 g749703 ( .a(n_31540), .b(n_31481), .c(FE_OCP_RBN4417_n_31117), .o(n_31635) );
in01s02 g749704 ( .a(n_31191), .o(n_31192) );
no02m06 g749705 ( .a(n_31147), .b(n_31088), .o(n_31191) );
na02s01 g749706 ( .a(n_31228), .b(n_31227), .o(n_31229) );
na02s01 g749707 ( .a(n_30056), .b(n_30023), .o(n_30024) );
no02s01 g749708 ( .a(n_29930), .b(n_29970), .o(n_29931) );
no02s01 g749709 ( .a(n_31414), .b(n_31407), .o(n_31415) );
no02s01 g749710 ( .a(n_31349), .b(n_31224), .o(n_31351) );
no02m06 TIMEBOOST_cell_6194 ( .a(TIMEBOOST_net_1948), .b(n_35197), .o(n_35287) );
no02s02 g749712 ( .a(n_31290), .b(n_31342), .o(n_31348) );
in01s01 g749713 ( .a(n_31395), .o(n_31457) );
na02s02 g749714 ( .a(n_31325), .b(n_31374), .o(n_31395) );
ao12s02 g749715 ( .a(n_31346), .b(n_31255), .c(n_31311), .o(n_31347) );
no02s01 g749716 ( .a(n_31417), .b(n_31311), .o(n_31455) );
na02s01 g749717 ( .a(n_31481), .b(FE_OCP_RBN4417_n_31117), .o(n_31540) );
in01s01 g749718 ( .a(n_31576), .o(n_31577) );
ao12s01 g749719 ( .a(n_31414), .b(n_31311), .c(n_31410), .o(n_31576) );
oa12s01 g749720 ( .a(n_31175), .b(n_31174), .c(n_186), .o(n_31226) );
na02s01 TIMEBOOST_cell_8044 ( .a(n_30955), .b(FE_OCP_RBN6204_n_31819), .o(TIMEBOOST_net_2653) );
oa12s01 g749722 ( .a(n_31311), .b(n_31411), .c(n_31410), .o(n_31412) );
na02s01 g749723 ( .a(n_31174), .b(n_186), .o(n_31175) );
in01s01 g749724 ( .a(n_31431), .o(n_31432) );
no02s01 g749725 ( .a(n_31408), .b(n_31409), .o(n_31431) );
no02s01 g749726 ( .a(n_31410), .b(n_31311), .o(n_31414) );
in01s01 g749727 ( .a(n_31537), .o(n_31538) );
na02s01 g749728 ( .a(n_31428), .b(n_31511), .o(n_31537) );
in01s01 g749729 ( .a(n_31147), .o(n_31228) );
ao12f04 g749730 ( .a(n_31118), .b(n_31066), .c(n_179), .o(n_31147) );
oa12f08 g749731 ( .a(n_29828), .b(n_29875), .c(n_29784), .o(n_29970) );
ao12s01 g749732 ( .a(n_29906), .b(n_29905), .c(n_29904), .o(n_31445) );
na02f08 g749733 ( .a(n_29903), .b(n_29815), .o(n_30056) );
oa12s01 g749734 ( .a(n_29874), .b(n_29875), .c(n_29873), .o(n_31583) );
in01s01 g749735 ( .a(n_31391), .o(n_31392) );
oa12s01 g749736 ( .a(n_31311), .b(n_31372), .c(n_31371), .o(n_31391) );
na02s02 g749737 ( .a(n_31190), .b(FE_OCP_RBN4424_n_31117), .o(n_31257) );
in01s01 g749738 ( .a(n_31292), .o(n_31349) );
oa12s01 g749739 ( .a(FE_OCP_RBN4423_n_31117), .b(n_31509), .c(n_31256), .o(n_31292) );
na02s01 TIMEBOOST_cell_772 ( .a(TIMEBOOST_net_0), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_), .o(n_36434) );
ao12s01 g749741 ( .a(FE_OCP_RBN4417_n_31117), .b(n_31289), .c(n_31288), .o(n_31290) );
no02s01 g749742 ( .a(n_31317), .b(n_31345), .o(n_31390) );
oa12s01 g749743 ( .a(FE_OCP_RBN4425_n_31117), .b(n_31324), .c(n_30920), .o(n_31325) );
in01s01 g749744 ( .a(n_31633), .o(n_31634) );
oa12s01 g749745 ( .a(n_31393), .b(FE_OCP_RBN4416_n_31117), .c(n_31281), .o(n_31633) );
in01s01 g749746 ( .a(n_31573), .o(n_31574) );
ao12s01 g749747 ( .a(n_31408), .b(n_31311), .c(n_31372), .o(n_31573) );
oa12s01 g749748 ( .a(n_31121), .b(n_31120), .c(n_31119), .o(n_31417) );
ao12s01 g749749 ( .a(n_31092), .b(n_31091), .c(n_31090), .o(n_31481) );
no02s01 g749750 ( .a(n_31091), .b(n_31090), .o(n_31092) );
na02s01 g749751 ( .a(n_31120), .b(n_31119), .o(n_31121) );
ao12m06 g749752 ( .a(n_29951), .b(n_29961), .c(n_29857), .o(n_30055) );
ao12s02 g749753 ( .a(n_30211), .b(n_30242), .c(n_30134), .o(n_30297) );
no02s03 g749754 ( .a(n_30177), .b(n_30175), .o(n_30223) );
no02s01 g749755 ( .a(n_29905), .b(n_29904), .o(n_29906) );
na02f08 g749756 ( .a(n_29905), .b(n_29814), .o(n_29903) );
oa12m04 g749757 ( .a(n_29954), .b(n_29964), .c(n_29896), .o(n_30054) );
ao12f01 g749758 ( .a(FE_OCP_RBN5785_n_30071), .b(n_30119), .c(n_29869), .o(n_30203) );
oa12s01 g749759 ( .a(n_30295), .b(n_30243), .c(n_29846), .o(n_30296) );
na02s01 g749760 ( .a(n_29875), .b(n_29873), .o(n_29874) );
na02s01 TIMEBOOST_cell_771 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_5_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_), .o(TIMEBOOST_net_0) );
no02s01 g749762 ( .a(n_31118), .b(n_31067), .o(n_31174) );
na02s01 g749763 ( .a(n_31115), .b(n_31089), .o(n_31227) );
no02s01 g749764 ( .a(n_31321), .b(n_31322), .o(n_31323) );
na02s01 g749765 ( .a(n_31312), .b(n_31344), .o(n_31345) );
in01s01 g749766 ( .a(n_31319), .o(n_31320) );
na02s01 g749767 ( .a(n_31287), .b(n_31187), .o(n_31319) );
na02s01 g749768 ( .a(n_31221), .b(n_31189), .o(n_31190) );
in01s01 g749769 ( .a(n_31631), .o(n_31632) );
na02s01 g749770 ( .a(n_31572), .b(n_31280), .o(n_31631) );
na02s01 g749771 ( .a(n_31287), .b(n_31285), .o(n_31286) );
in01s01 g749772 ( .a(n_31369), .o(n_31370) );
na02s01 g749773 ( .a(n_31339), .b(n_31289), .o(n_31369) );
no02s01 g749774 ( .a(n_31342), .b(n_31219), .o(n_31343) );
na02s01 g749775 ( .a(n_31339), .b(n_31340), .o(n_31341) );
in01s01 g749776 ( .a(n_31629), .o(n_31630) );
na02s01 g749777 ( .a(n_31571), .b(n_31526), .o(n_31629) );
in01s01 g749778 ( .a(n_31317), .o(n_31318) );
na02s01 g749779 ( .a(n_31571), .b(n_31284), .o(n_31317) );
in01s01 g749780 ( .a(n_31388), .o(n_31389) );
no02s01 g749781 ( .a(n_31368), .b(n_31324), .o(n_31388) );
in01s01 g749782 ( .a(n_31429), .o(n_31430) );
no02s01 g749783 ( .a(n_31407), .b(n_31411), .o(n_31429) );
no02s01 g749784 ( .a(n_31249), .b(n_31324), .o(n_31283) );
in01s01 g749785 ( .a(n_31627), .o(n_31628) );
na02s01 g749786 ( .a(n_31570), .b(n_31528), .o(n_31627) );
in01s01 g749787 ( .a(n_31315), .o(n_31316) );
na02s01 g749788 ( .a(n_31394), .b(n_31254), .o(n_31315) );
in01s01 g749789 ( .a(n_31313), .o(n_31314) );
na02s01 g749790 ( .a(n_31570), .b(n_31282), .o(n_31313) );
na02s01 g749791 ( .a(n_31281), .b(FE_OCP_RBN4416_n_31117), .o(n_31393) );
na02s01 g749792 ( .a(n_31254), .b(n_31281), .o(n_31255) );
in01s01 g749793 ( .a(n_31625), .o(n_31626) );
na02s01 g749794 ( .a(n_31338), .b(n_31569), .o(n_31625) );
no02s01 g749795 ( .a(n_31372), .b(n_31311), .o(n_31408) );
na02s01 g749796 ( .a(n_31311), .b(n_31416), .o(n_31511) );
in01s01 g749797 ( .a(n_31454), .o(n_31428) );
no02s01 g749798 ( .a(n_31311), .b(n_31416), .o(n_31454) );
na02s01 g749799 ( .a(n_31536), .b(n_31144), .o(n_31640) );
na02s01 g749800 ( .a(n_31222), .b(n_31221), .o(n_31580) );
in01s01 g749801 ( .a(n_31534), .o(n_31535) );
no02s01 g749802 ( .a(n_31510), .b(n_31509), .o(n_31534) );
oa22s01 g749803 ( .a(n_29835), .b(n_29848), .c(n_29811), .d(n_29796), .o(n_31403) );
oa12s01 g749804 ( .a(n_31460), .b(n_31311), .c(n_31145), .o(n_31643) );
in01s01 g749805 ( .a(n_31532), .o(n_31533) );
oa12s01 g749806 ( .a(n_31185), .b(n_31530), .c(n_31189), .o(n_31532) );
in01s01 g749807 ( .a(n_31623), .o(n_31624) );
oa12s01 g749808 ( .a(n_31284), .b(FE_OCP_RBN4417_n_31117), .c(n_31216), .o(n_31623) );
in01s01 g749809 ( .a(n_31621), .o(n_31622) );
na02s01 g749810 ( .a(n_31285), .b(n_31508), .o(n_31621) );
in01s01 g749811 ( .a(n_31567), .o(n_31568) );
ao12s01 g749812 ( .a(n_31322), .b(n_31311), .c(n_31251), .o(n_31567) );
in01s01 g749813 ( .a(n_31619), .o(n_31620) );
oa12s01 g749814 ( .a(n_31340), .b(FE_OCP_RBN4417_n_31117), .c(n_31288), .o(n_31619) );
in01s01 g749815 ( .a(n_31617), .o(n_31618) );
oa12s01 g749816 ( .a(n_31344), .b(FE_OCP_RBN4417_n_31117), .c(n_31277), .o(n_31617) );
in01s01 g749817 ( .a(n_31615), .o(n_31616) );
oa12s01 g749818 ( .a(n_31282), .b(FE_OCP_RBN4416_n_31117), .c(n_31275), .o(n_31615) );
oa12s01 g749819 ( .a(n_30977), .b(n_30976), .c(n_30975), .o(n_31410) );
oa22s01 g749820 ( .a(n_31311), .b(n_31294), .c(n_31530), .d(n_30392), .o(n_31637) );
in01s01 g749821 ( .a(n_31564), .o(n_31565) );
oa22s01 g749822 ( .a(n_31311), .b(n_31256), .c(n_31530), .d(n_31211), .o(n_31564) );
in01s04 g749823 ( .a(FE_OCPN1947_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36750) );
na02s01 g749825 ( .a(n_30976), .b(n_30975), .o(n_30977) );
no02f08 g749826 ( .a(n_29834), .b(n_29848), .o(n_29905) );
no02s02 g749827 ( .a(FE_OCP_RBN4419_n_31117), .b(n_31172), .o(n_31509) );
na02s01 g749828 ( .a(FE_OCP_RBN4422_n_31117), .b(n_31253), .o(n_31572) );
in01s01 g749829 ( .a(n_31528), .o(n_31529) );
na02s01 g749830 ( .a(n_31311), .b(n_30968), .o(n_31528) );
no02m04 g749831 ( .a(n_31044), .b(n_31043), .o(n_31118) );
in01s01 g749832 ( .a(n_31254), .o(n_31220) );
na02s01 g749833 ( .a(FE_OCP_RBN4425_n_31117), .b(n_31038), .o(n_31254) );
no02s01 g749834 ( .a(n_31311), .b(n_30474), .o(n_31510) );
na02s01 g749835 ( .a(FE_OCP_RBN4419_n_31117), .b(n_31116), .o(n_31536) );
in01s01 g749836 ( .a(n_31224), .o(n_31187) );
no02s01 g749837 ( .a(FE_OCP_RBN4418_n_31117), .b(n_31171), .o(n_31224) );
na02s01 g749838 ( .a(FE_OCP_RBN4418_n_31117), .b(n_31171), .o(n_31287) );
in01s01 g749839 ( .a(n_31185), .o(n_31186) );
na02s01 g749840 ( .a(FE_OCP_RBN4419_n_31117), .b(n_31189), .o(n_31185) );
na02s01 g749841 ( .a(FE_OCP_RBN4415_n_31117), .b(n_30416), .o(n_31221) );
na02s01 g749842 ( .a(FE_OCP_RBN4415_n_31117), .b(n_31145), .o(n_31460) );
in01s01 g749843 ( .a(n_31143), .o(n_31144) );
no02s02 g749844 ( .a(FE_OCP_RBN4419_n_31117), .b(n_31116), .o(n_31143) );
in01s01 g749845 ( .a(n_31066), .o(n_31067) );
na02m04 g749846 ( .a(n_31044), .b(n_31043), .o(n_31066) );
in01s01 g749847 ( .a(n_31088), .o(n_31089) );
no02s06 g749848 ( .a(n_31040), .b(n_30102), .o(n_31088) );
in01s01 g749849 ( .a(n_31114), .o(n_31115) );
no02s02 g749850 ( .a(n_31064), .b(n_30103), .o(n_31114) );
na02s01 g749851 ( .a(FE_OCP_RBN4419_n_31117), .b(n_30417), .o(n_31222) );
na02s01 g749852 ( .a(n_31311), .b(n_31223), .o(n_31508) );
na02s01 g749853 ( .a(FE_OCP_RBN4418_n_31117), .b(n_30615), .o(n_31285) );
in01s01 g749854 ( .a(n_31321), .o(n_31280) );
no02s01 g749855 ( .a(FE_OCP_RBN4422_n_31117), .b(n_31253), .o(n_31321) );
no02s01 g749856 ( .a(FE_OCP_RBN4425_n_31117), .b(n_31251), .o(n_31322) );
in01s01 g749857 ( .a(n_31289), .o(n_31219) );
na02s01 g749858 ( .a(FE_OCP_RBN4425_n_31117), .b(n_31184), .o(n_31289) );
in01s01 g749859 ( .a(n_31279), .o(n_31339) );
no02s01 g749860 ( .a(FE_OCP_RBN4425_n_31117), .b(n_31184), .o(n_31279) );
na02s01 g749861 ( .a(FE_OCP_RBN4417_n_31117), .b(n_31288), .o(n_31340) );
in01s01 g749862 ( .a(n_31526), .o(n_31527) );
na02s01 g749863 ( .a(n_31311), .b(n_30718), .o(n_31526) );
na02s01 g749864 ( .a(FE_OCP_RBN4417_n_31117), .b(n_31210), .o(n_31571) );
na02s01 g749865 ( .a(FE_OCP_RBN4417_n_31117), .b(n_31216), .o(n_31284) );
no02s01 g749866 ( .a(FE_OCP_RBN4416_n_31117), .b(n_31214), .o(n_31324) );
in01s01 g749867 ( .a(n_31312), .o(n_31368) );
na02s01 g749868 ( .a(FE_OCP_RBN4416_n_31117), .b(n_31214), .o(n_31312) );
na02s01 g749869 ( .a(FE_OCP_RBN4417_n_31117), .b(n_31277), .o(n_31344) );
na02s01 g749870 ( .a(FE_OCP_RBN4416_n_31117), .b(n_31213), .o(n_31570) );
in01s01 g749871 ( .a(n_31407), .o(n_31387) );
no02s01 g749872 ( .a(n_31311), .b(n_30971), .o(n_31407) );
na02s01 g749873 ( .a(FE_OCP_RBN4416_n_31117), .b(n_31275), .o(n_31282) );
na02s01 g749874 ( .a(FE_OCP_RBN4416_n_31117), .b(n_31039), .o(n_31394) );
na02s01 g749875 ( .a(n_31311), .b(n_31371), .o(n_31569) );
in01s01 g749876 ( .a(n_31409), .o(n_31338) );
no02s01 g749877 ( .a(n_31311), .b(n_31371), .o(n_31409) );
no02s01 g749878 ( .a(FE_OCP_RBN4416_n_31117), .b(n_30970), .o(n_31411) );
na02f04 g749879 ( .a(n_29968), .b(n_29902), .o(n_29969) );
na03f08 TIMEBOOST_cell_8205 ( .a(n_28003), .b(n_28042), .c(n_28072), .o(n_28188) );
no02s02 TIMEBOOST_cell_8874 ( .a(n_31194), .b(n_31074), .o(TIMEBOOST_net_2924) );
ao12s01 g749883 ( .a(n_30438), .b(n_31065), .c(n_30061), .o(n_31120) );
no02m06 g749884 ( .a(n_29841), .b(n_29926), .o(n_29988) );
in01s02 g749885 ( .a(n_30176), .o(n_30177) );
na02s03 g749886 ( .a(n_29857), .b(n_30078), .o(n_30176) );
no02s06 TIMEBOOST_cell_6696 ( .a(TIMEBOOST_net_2105), .b(TIMEBOOST_net_1261), .o(n_8100) );
oa12f08 g749888 ( .a(n_29807), .b(n_29816), .c(n_29775), .o(n_29875) );
in01s01 g749889 ( .a(n_31490), .o(n_29966) );
no02s02 g749890 ( .a(n_29871), .b(n_29847), .o(n_31490) );
oa12s01 g749891 ( .a(n_31042), .b(n_31065), .c(n_31041), .o(n_31416) );
na02s01 g749892 ( .a(FE_OCP_RBN4419_n_31117), .b(n_30432), .o(n_31169) );
oa12s01 g749893 ( .a(FE_OCP_RBN4419_n_31117), .b(n_31211), .c(n_31172), .o(n_31212) );
in01s01 g749894 ( .a(n_31276), .o(n_31342) );
oa12s01 g749895 ( .a(FE_OCP_RBN4425_n_31117), .b(n_31251), .c(n_31253), .o(n_31276) );
in01s01 g749896 ( .a(n_31249), .o(n_31374) );
ao12s01 g749897 ( .a(FE_OCP_RBN4417_n_31117), .b(n_31216), .c(n_31210), .o(n_31249) );
ao12s01 g749898 ( .a(FE_OCP_RBN4416_n_31117), .b(n_31275), .c(n_31213), .o(n_31346) );
ao22s01 g749899 ( .a(n_30922), .b(n_30412), .c(n_30921), .d(n_30413), .o(n_31281) );
oa12s01 g749900 ( .a(n_30974), .b(n_30973), .c(n_30972), .o(n_31372) );
ao12s01 g749901 ( .a(n_30184), .b(n_30969), .c(n_30186), .o(n_31091) );
no02s04 g749902 ( .a(n_29897), .b(n_29928), .o(n_29929) );
no02s01 g749903 ( .a(n_30019), .b(n_30018), .o(n_30020) );
no02m04 g749904 ( .a(n_29960), .b(n_29958), .o(n_29987) );
na02s02 g749905 ( .a(n_30196), .b(n_30138), .o(n_30202) );
na02s01 g749907 ( .a(n_30216), .b(n_30245), .o(n_30246) );
na02s01 g749908 ( .a(n_29968), .b(n_29901), .o(n_30247) );
na02f02 g749909 ( .a(n_29901), .b(n_29925), .o(n_29902) );
na02s01 g749910 ( .a(n_29965), .b(n_29870), .o(n_30265) );
no03s08 TIMEBOOST_cell_8187 ( .a(FE_OCP_RBN2444_n_1675), .b(FE_RN_239_0), .c(n_1517), .o(n_1725) );
na02s01 g749912 ( .a(n_30384), .b(n_30423), .o(n_30444) );
no02s01 g749913 ( .a(n_29960), .b(n_30018), .o(n_30406) );
no02s04 g749914 ( .a(n_30018), .b(FE_OCP_RBN5603_n_29056), .o(n_29964) );
in01s02 g749915 ( .a(n_30147), .o(n_30148) );
na02s03 g749916 ( .a(n_30120), .b(n_30011), .o(n_30147) );
in01s01 g749917 ( .a(n_30200), .o(n_30201) );
no02s01 g749918 ( .a(n_30172), .b(n_30171), .o(n_30200) );
no02s01 g749920 ( .a(n_30577), .b(n_30244), .o(n_30263) );
na02m01 g749921 ( .a(n_30077), .b(n_29327), .o(n_30119) );
no02s01 g749923 ( .a(n_30262), .b(n_30261), .o(n_30281) );
in01s01 g749924 ( .a(n_30320), .o(n_30321) );
no02s01 g749925 ( .a(n_30318), .b(n_30294), .o(n_30320) );
no02s01 g749926 ( .a(n_30262), .b(n_30214), .o(n_30243) );
no02s06 g749927 ( .a(n_29918), .b(n_29986), .o(n_29963) );
no02s02 g749929 ( .a(n_30195), .b(n_30050), .o(n_30197) );
no02s01 g749930 ( .a(n_30278), .b(n_30279), .o(n_30280) );
na02s01 g749932 ( .a(n_30016), .b(n_29985), .o(n_30017) );
na02s01 g749933 ( .a(n_31065), .b(n_31041), .o(n_31042) );
na02s01 g749934 ( .a(n_30973), .b(n_30972), .o(n_30974) );
na02m08 g749935 ( .a(n_29868), .b(n_29984), .o(n_29962) );
no02s02 TIMEBOOST_cell_3981 ( .a(n_4238), .b(n_3082), .o(TIMEBOOST_net_1081) );
no02s04 g749937 ( .a(n_29893), .b(n_29892), .o(n_29926) );
na02s06 g749938 ( .a(n_29985), .b(FE_OCP_RBN5023_n_29080), .o(n_29961) );
no02s01 g749940 ( .a(n_30356), .b(n_30076), .o(n_30145) );
na02s01 g749941 ( .a(n_30213), .b(FE_OCP_RBN4156_n_29378), .o(n_30242) );
na02s03 g749942 ( .a(n_30051), .b(FE_OCP_RBN3710_n_29055), .o(n_30078) );
na02m04 TIMEBOOST_cell_2073 ( .a(n_14326), .b(FE_OCP_RBN4189_n_13765), .o(TIMEBOOST_net_651) );
na02s01 g749945 ( .a(n_30349), .b(n_30371), .o(n_30369) );
in01s01 g749946 ( .a(n_30239), .o(n_30240) );
no02s02 g749947 ( .a(n_30470), .b(FE_OCP_RBN6746_n_30170), .o(n_30239) );
in01s01 g749948 ( .a(n_30143), .o(n_30144) );
no02s01 g749949 ( .a(n_30050), .b(n_30116), .o(n_30143) );
no02s02 g749951 ( .a(n_30277), .b(n_30278), .o(n_30292) );
na02s01 g749953 ( .a(n_30372), .b(n_30344), .o(n_30403) );
no02s01 g749954 ( .a(n_29895), .b(n_29865), .o(n_30225) );
in01s01 g749955 ( .a(n_30014), .o(n_30015) );
no02s01 g749956 ( .a(n_29986), .b(n_29893), .o(n_30014) );
no02s01 g749957 ( .a(n_30443), .b(n_30422), .o(n_30482) );
na02s01 g749958 ( .a(n_30021), .b(n_29985), .o(n_30376) );
in01s01 g749959 ( .a(n_29834), .o(n_29835) );
no02f08 g749960 ( .a(n_29795), .b(n_29810), .o(n_29834) );
na02s01 g749961 ( .a(n_29833), .b(n_29872), .o(n_30023) );
na02s01 g749962 ( .a(n_29925), .b(n_29863), .o(n_30151) );
no02s01 g749963 ( .a(n_29816), .b(n_29827), .o(n_29871) );
no02s01 g749964 ( .a(n_29780), .b(n_29826), .o(n_29847) );
in01s01 g749965 ( .a(n_30012), .o(n_30013) );
na02s01 g749966 ( .a(n_29984), .b(n_29890), .o(n_30012) );
ao12s01 g749967 ( .a(n_29928), .b(n_29869), .c(n_29898), .o(n_30457) );
oa12s01 g749968 ( .a(n_29959), .b(n_29896), .c(FE_OCP_RBN2049_n_29056), .o(n_30488) );
in01s02 g749969 ( .a(n_30141), .o(n_30142) );
na02s02 g749970 ( .a(n_30114), .b(n_30053), .o(n_30141) );
in01s02 g749971 ( .a(n_30220), .o(n_30221) );
na02s01 g749972 ( .a(n_30196), .b(n_30113), .o(n_30220) );
in01s01 g749973 ( .a(n_30259), .o(n_30260) );
no02s02 g749974 ( .a(n_30173), .b(n_30194), .o(n_30259) );
in01s01 g749975 ( .a(n_30275), .o(n_30276) );
na02s01 g749976 ( .a(n_30245), .b(n_30215), .o(n_30275) );
ao12s01 g749977 ( .a(n_30318), .b(n_29869), .c(n_29530), .o(n_30319) );
ao12s01 g749978 ( .a(n_30161), .b(n_30925), .c(n_30062), .o(n_30976) );
in01s01 g749983 ( .a(n_31311), .o(n_31530) );
in01s03 g749999 ( .a(FE_OCP_RBN4418_n_31117), .o(n_31311) );
in01s06 g750012 ( .a(n_31064), .o(n_31117) );
in01s04 g750013 ( .a(n_31040), .o(n_31064) );
in01m04 g750014 ( .a(n_31044), .o(n_31040) );
na02s02 TIMEBOOST_cell_5572 ( .a(n_6204), .b(n_6281), .o(TIMEBOOST_net_1734) );
no02s01 g750017 ( .a(n_30198), .b(n_30212), .o(n_30273) );
in01s01 g750018 ( .a(n_30218), .o(n_30219) );
no02m01 g750019 ( .a(n_30195), .b(n_30108), .o(n_30218) );
in01s01 g750020 ( .a(n_30316), .o(n_30317) );
no02s02 g750021 ( .a(n_30279), .b(n_30258), .o(n_30316) );
oa12s01 g750022 ( .a(n_29919), .b(n_29922), .c(n_28995), .o(n_30460) );
ao12s01 g750023 ( .a(n_29957), .b(FE_OCPN1298_n_30134), .c(FE_OCP_RBN5024_n_29080), .o(n_30493) );
oa22s01 g750025 ( .a(FE_OCPN1298_n_30134), .b(n_29553), .c(n_29922), .d(FE_OCP_RBN4168_n_29553), .o(n_30401) );
ao22s01 g750026 ( .a(n_29869), .b(n_29083), .c(n_29896), .d(n_29113), .o(n_30447) );
in01s01 g750027 ( .a(n_30367), .o(n_30368) );
oa22s01 g750028 ( .a(n_29869), .b(n_29485), .c(n_29896), .d(n_29507), .o(n_30367) );
oa22s01 g750029 ( .a(FE_OCPN1298_n_30134), .b(n_29059), .c(n_29922), .d(n_29913), .o(n_30485) );
in01s01 g750030 ( .a(n_31038), .o(n_31039) );
oa12s01 g750031 ( .a(n_30953), .b(n_30952), .c(n_30951), .o(n_31038) );
in01s01 g750032 ( .a(n_30970), .o(n_30971) );
ao12s01 g750033 ( .a(n_30903), .b(n_30925), .c(n_30902), .o(n_30970) );
in01s01 g750034 ( .a(n_30139), .o(n_30140) );
na02s01 g750035 ( .a(n_30007), .b(n_30049), .o(n_30139) );
oa22s01 g750037 ( .a(FE_OCPN1298_n_30134), .b(FE_OCP_RBN2650_n_29470), .c(n_29922), .d(n_45489), .o(n_30385) );
in01s01 g750038 ( .a(n_30347), .o(n_30348) );
oa22s01 g750039 ( .a(n_29896), .b(n_29501), .c(n_29869), .d(n_29530), .o(n_30347) );
oa22s01 g750041 ( .a(n_29869), .b(FE_OCPN4853_n_29502), .c(n_29896), .d(n_29523), .o(n_30345) );
na02f01 g750043 ( .a(n_29809), .b(n_28830), .o(n_29901) );
in01s01 g750044 ( .a(n_29897), .o(n_29965) );
no02s02 g750045 ( .a(n_29869), .b(n_28892), .o(n_29897) );
in01s01 g750046 ( .a(n_29899), .o(n_29870) );
no02s02 g750047 ( .a(n_29846), .b(FE_OCPN7083_n_28891), .o(n_29899) );
no02s02 g750048 ( .a(n_29869), .b(n_29898), .o(n_29928) );
na02s01 g750049 ( .a(n_29896), .b(n_30364), .o(n_30423) );
in01s01 g750050 ( .a(n_30383), .o(n_30384) );
no02s01 g750051 ( .a(n_29896), .b(n_30364), .o(n_30383) );
in01s01 g750053 ( .a(n_29960), .o(n_29982) );
no02s06 g750054 ( .a(n_29869), .b(n_29082), .o(n_29960) );
no02s04 g750055 ( .a(n_29896), .b(FE_OCPN5132_n_29081), .o(n_30018) );
in01s01 g750056 ( .a(n_29958), .o(n_29959) );
no02s02 g750057 ( .a(n_29869), .b(FE_OCP_DRV_N6263_FE_OCP_RBN5603_n_29056), .o(n_29958) );
in01m01 g750058 ( .a(n_30010), .o(n_30011) );
no02m01 g750059 ( .a(n_29869), .b(n_29057), .o(n_30010) );
na02m01 g750060 ( .a(n_29869), .b(n_29057), .o(n_30120) );
na02s02 g750061 ( .a(n_29896), .b(FE_OCP_RBN2583_n_29091), .o(n_30114) );
na02s02 g750062 ( .a(n_29869), .b(FE_OCP_RBN2584_n_29091), .o(n_30053) );
in01s01 g750063 ( .a(n_30172), .o(n_30138) );
no02s02 g750064 ( .a(n_29869), .b(n_29161), .o(n_30172) );
in01s02 g750065 ( .a(n_30077), .o(n_30171) );
na02s03 g750066 ( .a(n_29869), .b(n_29161), .o(n_30077) );
na02s01 g750067 ( .a(n_29869), .b(n_46960), .o(n_30113) );
na02s01 g750068 ( .a(n_29896), .b(n_29327), .o(n_30196) );
in01s01 g750069 ( .a(n_30244), .o(n_30217) );
no02s01 g750070 ( .a(n_29896), .b(FE_OCP_RBN7131_n_29262), .o(n_30244) );
no02s01 g750071 ( .a(n_29869), .b(FE_OCP_RBN7130_n_29262), .o(n_30577) );
no02s01 g750072 ( .a(n_29869), .b(n_30111), .o(n_30173) );
no02s01 g750073 ( .a(n_29896), .b(n_29477), .o(n_30194) );
no02s01 g750074 ( .a(n_29896), .b(n_30192), .o(n_30262) );
in01s01 g750075 ( .a(n_30216), .o(n_30261) );
na02s01 g750076 ( .a(n_29896), .b(n_30192), .o(n_30216) );
na02s01 g750077 ( .a(n_29869), .b(n_30214), .o(n_30215) );
na02s01 g750078 ( .a(n_29896), .b(n_29472), .o(n_30245) );
no02m01 g750079 ( .a(n_29869), .b(n_29417), .o(n_30294) );
no02s01 g750080 ( .a(n_29896), .b(n_29442), .o(n_30318) );
na02s01 g750081 ( .a(n_29896), .b(n_29501), .o(n_30272) );
na02s01 g750082 ( .a(n_30952), .b(n_30951), .o(n_30953) );
in01s01 g750083 ( .a(n_30969), .o(n_31065) );
na02s02 g750084 ( .a(n_30896), .b(n_30234), .o(n_30969) );
in01s01 g750086 ( .a(n_29956), .o(n_29957) );
na02s10 g750087 ( .a(n_29922), .b(FE_OCP_RBN5023_n_29080), .o(n_29956) );
in01s01 g750088 ( .a(n_29894), .o(n_29895) );
na02m04 g750089 ( .a(n_29841), .b(FE_OCPN5298_n_29866), .o(n_29894) );
na02s06 g750090 ( .a(n_29841), .b(FE_OCPN5298_n_29866), .o(n_29868) );
in01s01 g750091 ( .a(n_29864), .o(n_29865) );
in01s01 g750094 ( .a(n_29893), .o(n_29920) );
in01s01 g750096 ( .a(n_29918), .o(n_29919) );
no02s06 g750097 ( .a(n_29857), .b(FE_OCP_DRV_N5304_n_29892), .o(n_29918) );
no02s06 g750098 ( .a(n_29857), .b(n_28889), .o(n_29986) );
na02s06 g750099 ( .a(n_29857), .b(n_29031), .o(n_29985) );
in01s01 g750102 ( .a(n_30051), .o(n_30076) );
na02s04 g750103 ( .a(n_29857), .b(FE_OCP_RBN5026_n_29053), .o(n_30051) );
no02s01 g750104 ( .a(FE_OCP_RBN5026_n_29053), .b(n_29857), .o(n_30356) );
in01s01 g750105 ( .a(n_30213), .o(n_30277) );
na02s01 g750106 ( .a(n_30134), .b(n_30191), .o(n_30213) );
no02s01 g750107 ( .a(n_30134), .b(n_29260), .o(n_30198) );
no02s01 g750108 ( .a(n_29857), .b(n_30136), .o(n_30470) );
no02s01 g750109 ( .a(n_29857), .b(n_29167), .o(n_30195) );
no02s02 g750113 ( .a(n_29857), .b(n_29292), .o(n_30050) );
no02s02 g750114 ( .a(n_29922), .b(FE_OCP_RBN4070_n_29292), .o(n_30116) );
no02s01 g750115 ( .a(n_30134), .b(n_29398), .o(n_30279) );
no02s02 g750116 ( .a(n_30134), .b(n_30191), .o(n_30278) );
na02s01 g750117 ( .a(FE_OCPN1298_n_30134), .b(n_45758), .o(n_30371) );
na02m01 g750118 ( .a(n_29922), .b(FE_OCP_RBN2635_n_29371), .o(n_30349) );
na02s01 g750120 ( .a(n_30134), .b(FE_OCPN1300_n_30136), .o(n_30170) );
no02s01 g750121 ( .a(n_29922), .b(n_29231), .o(n_30212) );
na02s01 g750122 ( .a(n_29922), .b(FE_OCP_RBN3710_n_29055), .o(n_30049) );
na02s01 g750123 ( .a(n_29857), .b(n_29055), .o(n_30007) );
no02s01 g750124 ( .a(n_29922), .b(n_29160), .o(n_30108) );
no02s01 g750125 ( .a(n_29922), .b(FE_OCP_RBN4156_n_29378), .o(n_30258) );
na02s01 g750126 ( .a(FE_OCPN1298_n_30134), .b(n_30310), .o(n_30372) );
in01s01 g750127 ( .a(n_30343), .o(n_30344) );
no02m01 g750128 ( .a(n_30134), .b(n_30310), .o(n_30343) );
in01s01 g750129 ( .a(n_30421), .o(n_30422) );
na02s01 g750130 ( .a(FE_OCPN1298_n_30134), .b(n_30399), .o(n_30421) );
no02s01 g750131 ( .a(FE_OCPN1298_n_30134), .b(n_30399), .o(n_30443) );
in01s01 g750134 ( .a(n_29890), .o(n_29916) );
na02f02 g750135 ( .a(n_29839), .b(FE_OCP_DRV_N1468_n_28775), .o(n_29890) );
na02s01 g750136 ( .a(n_29815), .b(n_29814), .o(n_29904) );
in01s01 g750137 ( .a(n_29832), .o(n_29833) );
no02f06 g750138 ( .a(n_29813), .b(FE_OCPUNCON3476_n_29812), .o(n_29832) );
na02m04 g750139 ( .a(n_29813), .b(FE_OCPUNCON3476_n_29812), .o(n_29872) );
na02f02 g750140 ( .a(n_29845), .b(FE_OCPUNCON3478_n_29844), .o(n_29925) );
in01s01 g750141 ( .a(n_29862), .o(n_29863) );
no02s04 g750142 ( .a(n_29845), .b(FE_OCPUNCON3478_n_29844), .o(n_29862) );
na02s01 g750143 ( .a(n_29955), .b(n_29889), .o(n_30025) );
no02s01 g750144 ( .a(n_30925), .b(n_30902), .o(n_30903) );
in01s01 g750145 ( .a(n_29954), .o(n_30019) );
no03f04 TIMEBOOST_cell_8349 ( .a(n_9763), .b(n_9663), .c(n_9928), .o(TIMEBOOST_net_673) );
no02s06 g750147 ( .a(n_29869), .b(n_29112), .o(n_29915) );
na02m01 g750149 ( .a(n_29869), .b(n_29211), .o(n_30071) );
oa12m01 g750150 ( .a(n_29869), .b(n_30111), .c(FE_OCP_RBN7130_n_29262), .o(n_30295) );
na03s03 TIMEBOOST_cell_759 ( .a(n_27659), .b(n_27465), .c(n_27709), .o(n_27771) );
ao12s01 g750152 ( .a(n_30096), .b(n_30923), .c(n_30431), .o(n_30973) );
in01s01 g750153 ( .a(n_30921), .o(n_30922) );
oa12s01 g750154 ( .a(n_30128), .b(n_30835), .c(n_30091), .o(n_30921) );
in01s01 g750155 ( .a(n_29952), .o(n_29953) );
in01s01 g750157 ( .a(n_29951), .o(n_30016) );
ao12s02 g750158 ( .a(n_29841), .b(n_29913), .c(n_28996), .o(n_29951) );
in01s01 g750159 ( .a(n_30210), .o(n_30211) );
oa12f01 g750160 ( .a(n_30134), .b(n_29260), .c(FE_OCPN1300_n_30136), .o(n_30210) );
na02s02 g750161 ( .a(n_29922), .b(n_29139), .o(n_30046) );
in01s01 g750162 ( .a(n_29816), .o(n_29780) );
no02f08 g750163 ( .a(n_29740), .b(n_29738), .o(n_29816) );
ao12s01 g750164 ( .a(n_29794), .b(n_29793), .c(n_29792), .o(n_31303) );
in01s01 g750165 ( .a(n_29795), .o(n_29796) );
oa12f08 g750166 ( .a(n_29764), .b(n_29755), .c(n_29728), .o(n_29795) );
in01s01 g750167 ( .a(n_29842), .o(n_29843) );
ao12s01 g750168 ( .a(n_29791), .b(n_29790), .c(n_29789), .o(n_29842) );
ao12s01 g750169 ( .a(n_30899), .b(n_30898), .c(n_30897), .o(n_31275) );
oa12s01 g750170 ( .a(n_30901), .b(n_30923), .c(n_30900), .o(n_31371) );
no02s02 g750171 ( .a(n_30836), .b(n_30127), .o(n_30952) );
na02s01 g750172 ( .a(n_30923), .b(n_30900), .o(n_30901) );
no02s01 g750173 ( .a(n_30898), .b(n_30897), .o(n_30899) );
na02m06 g750174 ( .a(n_29861), .b(FE_OCP_DRV_N1466_n_29860), .o(n_29955) );
ao12f04 g750175 ( .a(n_29739), .b(n_29736), .c(n_29611), .o(n_29740) );
in01s01 g750176 ( .a(n_29888), .o(n_29889) );
no02m06 g750177 ( .a(n_29861), .b(FE_OCP_DRV_N1466_n_29860), .o(n_29888) );
no02s01 g750178 ( .a(n_29793), .b(n_29792), .o(n_29794) );
no02s01 g750179 ( .a(n_29810), .b(n_29848), .o(n_29811) );
na02m06 g750180 ( .a(n_29754), .b(n_28657), .o(n_29815) );
na02f04 g750181 ( .a(n_29753), .b(FE_OCPN1256_n_28656), .o(n_29814) );
no02s01 g750182 ( .a(n_29859), .b(n_29787), .o(n_29930) );
no02s01 g750183 ( .a(n_29790), .b(n_29789), .o(n_29791) );
in01s10 g750217 ( .a(n_29869), .o(n_29896) );
in01m10 g750218 ( .a(n_29846), .o(n_29869) );
in01m08 g750219 ( .a(n_29809), .o(n_29846) );
ao12m08 g750220 ( .a(FE_RN_522_0), .b(n_29788), .c(n_29671), .o(n_29809) );
in01s02 g750242 ( .a(n_29922), .o(n_30134) );
in01s10 g750251 ( .a(n_29857), .o(n_29922) );
in01s10 g750253 ( .a(n_29841), .o(n_29857) );
in01m08 g750254 ( .a(n_29831), .o(n_29841) );
oa12m08 g750256 ( .a(FE_OCPN1364_n_29615), .b(n_29808), .c(FE_OCP_RBN5720_n_29624), .o(n_29831) );
in01s01 g750257 ( .a(n_30895), .o(n_30896) );
no02f08 g750258 ( .a(n_30840), .b(n_30232), .o(n_30895) );
ao12f04 g750259 ( .a(n_29737), .b(n_29736), .c(n_29602), .o(n_29738) );
in01s01 g750264 ( .a(n_30920), .o(n_31277) );
oa12s01 g750265 ( .a(n_30839), .b(n_30838), .c(n_30837), .o(n_30920) );
in01s01 g750266 ( .a(n_31213), .o(n_30968) );
ao12s01 g750267 ( .a(n_30894), .b(n_30893), .c(n_30892), .o(n_31213) );
ao12s01 g750268 ( .a(n_30253), .b(n_30812), .c(n_30125), .o(n_30925) );
in01s01 g750269 ( .a(n_30840), .o(n_30923) );
no02f08 g750270 ( .a(n_30812), .b(n_30230), .o(n_30840) );
no02s01 g750271 ( .a(n_30893), .b(n_30892), .o(n_30894) );
na02s01 g750272 ( .a(n_30838), .b(n_30837), .o(n_30839) );
no02f06 g750273 ( .a(FE_OCP_RBN5213_n_29773), .b(n_28655), .o(n_29859) );
no02m04 g750276 ( .a(n_29773), .b(FE_OCPUNCON3470_n_28654), .o(n_29787) );
no02f06 g750277 ( .a(n_29751), .b(FE_OCP_DRV_N6275_n_28582), .o(n_29810) );
no02f06 g750278 ( .a(n_29752), .b(n_28583), .o(n_29848) );
na02s01 g750279 ( .a(n_29785), .b(n_29828), .o(n_29873) );
in01s01 g750280 ( .a(n_29826), .o(n_29827) );
na02s01 g750281 ( .a(n_29807), .b(n_29776), .o(n_29826) );
in01s01 g750282 ( .a(n_30835), .o(n_30836) );
ao12s01 g750283 ( .a(n_30811), .b(n_30756), .c(n_30159), .o(n_30835) );
na02m06 g750284 ( .a(n_29779), .b(n_29786), .o(n_29861) );
in01s01 g750285 ( .a(n_29755), .o(n_29792) );
oa12f08 g750286 ( .a(n_29698), .b(n_29735), .c(n_29660), .o(n_29755) );
ao12s01 g750287 ( .a(n_29734), .b(n_29733), .c(n_29735), .o(n_31206) );
in01m02 g750288 ( .a(n_29753), .o(n_29754) );
ao12s01 g750290 ( .a(n_29641), .b(n_29720), .c(n_29602), .o(n_29790) );
ao12s02 g750291 ( .a(n_29707), .b(n_29720), .c(n_29706), .o(n_31327) );
ao12s01 g750292 ( .a(n_30722), .b(n_30721), .c(n_30720), .o(n_31216) );
ao12s01 g750293 ( .a(n_30787), .b(n_30786), .c(n_30785), .o(n_31214) );
oa12s01 g750294 ( .a(n_30167), .b(n_30783), .c(n_30094), .o(n_30898) );
na02s06 TIMEBOOST_cell_2842 ( .a(n_7117), .b(FE_RN_2833_0), .o(TIMEBOOST_net_712) );
na02m04 g750296 ( .a(n_29762), .b(n_29502), .o(n_29786) );
no02s01 g750297 ( .a(n_30756), .b(n_30811), .o(n_30893) );
no02s01 g750298 ( .a(n_30786), .b(n_30785), .o(n_30787) );
na02f06 g750299 ( .a(n_29778), .b(FE_OCP_DRV_N1462_n_29777), .o(n_29828) );
in01s01 g750300 ( .a(n_29784), .o(n_29785) );
no02f08 g750301 ( .a(n_29778), .b(FE_OCP_DRV_N1462_n_29777), .o(n_29784) );
na02f06 g750302 ( .a(n_29766), .b(FE_OCP_DRV_N5147_n_29765), .o(n_29807) );
na02f06 g750303 ( .a(n_29674), .b(n_29589), .o(n_29736) );
in01s01 g750304 ( .a(n_29775), .o(n_29776) );
no02f06 g750305 ( .a(n_29766), .b(FE_OCP_DRV_N5147_n_29765), .o(n_29775) );
na02s01 g750306 ( .a(n_29764), .b(n_29729), .o(n_29793) );
no02s01 g750307 ( .a(n_29733), .b(n_29735), .o(n_29734) );
oa12m02 g750308 ( .a(n_29657), .b(n_29648), .c(n_29702), .o(n_29719) );
no02m04 g750309 ( .a(FE_OCP_RBN2732_n_29657), .b(n_29703), .o(n_29732) );
no02s01 g750310 ( .a(n_29720), .b(n_29706), .o(n_29707) );
no02s01 g750311 ( .a(n_30721), .b(n_30720), .o(n_30722) );
in01m02 g750312 ( .a(n_29788), .o(n_29763) );
na02f10 g750313 ( .a(n_29696), .b(n_29718), .o(n_29788) );
no02f06 g750314 ( .a(n_30719), .b(n_30160), .o(n_30812) );
ao12s01 g750315 ( .a(n_30101), .b(n_30688), .c(n_30126), .o(n_30838) );
in01m02 g750318 ( .a(n_29751), .o(n_29752) );
no02s06 TIMEBOOST_cell_2059 ( .a(n_24268), .b(n_23925), .o(TIMEBOOST_net_644) );
ao12s01 g750320 ( .a(n_30691), .b(n_30690), .c(n_30689), .o(n_31288) );
na02m02 TIMEBOOST_cell_8788 ( .a(n_9239), .b(n_9264), .o(TIMEBOOST_net_2881) );
in01m02 g750323 ( .a(n_29689), .o(n_29690) );
na02m04 g750324 ( .a(n_29648), .b(n_29604), .o(n_29689) );
na02m08 g750325 ( .a(FE_OCP_RBN5047_n_29648), .b(n_29631), .o(n_29718) );
na02s01 TIMEBOOST_cell_6183 ( .a(n_42962), .b(FE_OCPN878_n_43022), .o(TIMEBOOST_net_1943) );
no03s03 TIMEBOOST_cell_8362 ( .a(n_3678), .b(FE_OCP_RBN6761_n_3705), .c(TIMEBOOST_net_1303), .o(n_4113) );
in01s01 TIMEBOOST_cell_5916 ( .a(TIMEBOOST_net_1804), .o(TIMEBOOST_net_1805) );
na02m02 g750329 ( .a(FE_OCP_RBN2723_FE_RN_522_0), .b(n_29671), .o(n_29704) );
no02m02 g750330 ( .a(n_29681), .b(FE_RN_522_0), .o(n_29717) );
no02s01 g750331 ( .a(n_30690), .b(n_30689), .o(n_30691) );
na02s01 g750332 ( .a(n_30687), .b(n_30100), .o(n_30786) );
na02f06 g750333 ( .a(n_29716), .b(FE_OCPN5109_n_29715), .o(n_29764) );
in01s01 g750334 ( .a(n_29728), .o(n_29729) );
no02f06 g750335 ( .a(n_29716), .b(FE_OCPN5109_n_29715), .o(n_29728) );
no02s02 g750336 ( .a(n_29648), .b(n_29702), .o(n_29703) );
no02s02 g750337 ( .a(n_29730), .b(n_29551), .o(n_29762) );
na02s06 TIMEBOOST_cell_2841 ( .a(n_7456), .b(TIMEBOOST_net_711), .o(n_7507) );
in01s01 g750340 ( .a(n_30756), .o(n_30783) );
in01s01 g750341 ( .a(n_30719), .o(n_30756) );
na02f08 g750342 ( .a(n_30662), .b(n_30158), .o(n_30719) );
oa12s01 g750343 ( .a(n_29943), .b(n_30663), .c(n_30380), .o(n_30721) );
na02f08 g750344 ( .a(n_29714), .b(n_29700), .o(n_29778) );
na02s02 TIMEBOOST_cell_5531 ( .a(TIMEBOOST_net_1713), .b(n_6143), .o(n_6243) );
in01s01 g750346 ( .a(n_29674), .o(n_29720) );
oa12f04 g750347 ( .a(n_29592), .b(n_29666), .c(n_29632), .o(n_29674) );
oa12f08 g750348 ( .a(n_29587), .b(n_29687), .c(n_29622), .o(n_29735) );
ao12s01 g750349 ( .a(n_29670), .b(n_29687), .c(n_29669), .o(n_31164) );
oa12s01 g750350 ( .a(n_29727), .b(n_29739), .c(n_29737), .o(n_29789) );
oa12s01 g750351 ( .a(n_29668), .b(n_29667), .c(n_29666), .o(n_31264) );
in01s01 g750352 ( .a(n_31210), .o(n_30718) );
ao12s01 g750353 ( .a(n_30636), .b(n_30663), .c(n_30635), .o(n_31210) );
in01s02 g750354 ( .a(n_29672), .o(n_29673) );
no02f04 g750356 ( .a(n_29658), .b(n_29663), .o(n_29686) );
no02s06 TIMEBOOST_cell_4150 ( .a(TIMEBOOST_net_1165), .b(FE_OCP_RBN6877_n_16920), .o(n_17283) );
na02m06 g750358 ( .a(n_29676), .b(n_29442), .o(n_29714) );
na02s04 g750359 ( .a(n_29697), .b(n_29417), .o(n_29700) );
in01s01 g750364 ( .a(n_29671), .o(n_29681) );
na02m08 g750365 ( .a(n_29628), .b(n_25859), .o(n_29671) );
in01s01 g750366 ( .a(n_30687), .o(n_30688) );
in01s01 g750367 ( .a(n_30662), .o(n_30687) );
no02f08 g750368 ( .a(n_30663), .b(n_30084), .o(n_30662) );
no02s01 g750369 ( .a(n_30663), .b(n_30635), .o(n_30636) );
na02s01 g750370 ( .a(n_29661), .b(n_29698), .o(n_29733) );
no02s01 g750371 ( .a(n_29687), .b(n_29669), .o(n_29670) );
na02s01 g750372 ( .a(n_29739), .b(n_29737), .o(n_29727) );
na02s01 g750373 ( .a(n_29666), .b(n_29667), .o(n_29668) );
in01m04 g750380 ( .a(n_29730), .o(n_29749) );
no02m04 TIMEBOOST_cell_2067 ( .a(n_8694), .b(n_7601), .o(TIMEBOOST_net_648) );
ao12s01 g750383 ( .a(n_30090), .b(n_30634), .c(n_29976), .o(n_30690) );
no02s02 TIMEBOOST_cell_2838 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_13_), .b(n_33015), .o(TIMEBOOST_net_710) );
in01s01 g750385 ( .a(FE_OFN4733_n_29677), .o(n_29678) );
ao22s01 g750386 ( .a(n_29610), .b(n_29633), .c(n_29584), .d(n_29565), .o(n_29677) );
oa12s01 g750387 ( .a(n_30591), .b(n_30590), .c(n_30589), .o(n_31251) );
oa12s01 g750388 ( .a(n_30617), .b(n_30634), .c(n_30616), .o(n_31184) );
na02f06 g750390 ( .a(n_29634), .b(n_29612), .o(n_29635) );
no02s01 TIMEBOOST_cell_3919 ( .a(n_37945), .b(n_37575), .o(TIMEBOOST_net_1050) );
in01m02 g750392 ( .a(n_29697), .o(n_29676) );
no02f08 g750393 ( .a(n_29663), .b(n_29643), .o(n_29697) );
na02s01 g750396 ( .a(n_30590), .b(n_30589), .o(n_30591) );
na02s01 g750397 ( .a(n_30634), .b(n_30616), .o(n_30617) );
na02m06 g750398 ( .a(n_29645), .b(FE_OCPUNCON3468_n_29644), .o(n_29698) );
in01s01 g750399 ( .a(n_29660), .o(n_29661) );
no02f06 g750400 ( .a(n_29645), .b(FE_OCPUNCON3468_n_29644), .o(n_29660) );
na02f08 g750401 ( .a(n_29609), .b(n_29633), .o(n_29687) );
no02s01 g750402 ( .a(n_29632), .b(n_29593), .o(n_29667) );
in01f02 g750403 ( .a(n_29658), .o(n_29659) );
no02s04 TIMEBOOST_cell_4145 ( .a(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n_36607), .o(TIMEBOOST_net_1163) );
oa12m04 g750407 ( .a(n_29630), .b(n_29594), .c(n_29545), .o(n_29631) );
na02m04 TIMEBOOST_cell_8617 ( .a(TIMEBOOST_net_2795), .b(FE_OCP_RBN3261_n_21360), .o(n_21586) );
ao12f04 g750409 ( .a(n_29525), .b(n_29606), .c(n_29570), .o(n_29666) );
na02f04 g750410 ( .a(n_29656), .b(n_29642), .o(n_29739) );
na02m08 g750412 ( .a(n_29579), .b(n_29554), .o(n_29628) );
ao12s01 g750413 ( .a(n_29608), .b(n_29607), .c(n_29606), .o(n_31197) );
na02s04 g750416 ( .a(n_29568), .b(n_29630), .o(n_29615) );
no02f04 g750417 ( .a(n_29566), .b(FE_RN_1384_0), .o(n_29643) );
na02f08 g750420 ( .a(FE_OCP_RBN5702_n_29568), .b(n_25859), .o(n_29624) );
na02f02 g750422 ( .a(n_29620), .b(n_29494), .o(n_29642) );
na02f04 g750423 ( .a(n_29621), .b(FE_OCP_RBN6652_n_29494), .o(n_29656) );
in01s04 g750424 ( .a(n_29612), .o(n_29613) );
na02f06 g750425 ( .a(n_29596), .b(n_29549), .o(n_29612) );
no02f06 TIMEBOOST_cell_5519 ( .a(TIMEBOOST_net_1707), .b(FE_RN_1932_0), .o(n_46996) );
no02m04 g750427 ( .a(n_29562), .b(n_25859), .o(n_29702) );
na02m06 g750428 ( .a(FE_OCP_RBN4169_n_29553), .b(n_29630), .o(n_29579) );
na02s04 g750429 ( .a(n_29553), .b(n_25859), .o(n_29554) );
na02f06 TIMEBOOST_cell_2019 ( .a(FE_OCP_RBN4067_n_18829), .b(n_18371), .o(TIMEBOOST_net_624) );
no02s01 g750431 ( .a(n_30519), .b(n_30034), .o(n_30634) );
in01s01 g750432 ( .a(n_29592), .o(n_29593) );
na02f04 g750433 ( .a(n_29577), .b(n_29576), .o(n_29592) );
no02f04 g750434 ( .a(n_29577), .b(n_29576), .o(n_29632) );
no02f04 g750435 ( .a(n_29590), .b(n_28476), .o(n_29611) );
in01s01 g750436 ( .a(n_29609), .o(n_29610) );
na02f08 g750437 ( .a(n_29583), .b(n_29564), .o(n_29609) );
no02s01 g750438 ( .a(n_29588), .b(n_29622), .o(n_29669) );
no02s01 g750439 ( .a(n_29641), .b(n_29590), .o(n_29706) );
no02s01 g750440 ( .a(n_29607), .b(n_29606), .o(n_29608) );
in01m02 g750441 ( .a(n_29634), .o(n_29591) );
na02f08 g750442 ( .a(n_29529), .b(n_29532), .o(n_29634) );
in01f02 g750443 ( .a(n_29663), .o(n_29640) );
in01m02 g750446 ( .a(n_29604), .o(n_29605) );
na02s10 TIMEBOOST_cell_6590 ( .a(FE_RN_199_0), .b(TIMEBOOST_net_2052), .o(n_37252) );
oa12s01 g750448 ( .a(n_30000), .b(n_30552), .c(n_30381), .o(n_30590) );
na02m02 TIMEBOOST_cell_7982 ( .a(n_5114), .b(n_4497), .o(TIMEBOOST_net_2622) );
in01s01 g750451 ( .a(n_31223), .o(n_30615) );
oa12s01 g750452 ( .a(n_30550), .b(n_30549), .c(n_30548), .o(n_31223) );
oa12s01 g750453 ( .a(n_30521), .b(n_30552), .c(n_30520), .o(n_31253) );
na02s02 TIMEBOOST_cell_2033 ( .a(n_29488), .b(n_29023), .o(TIMEBOOST_net_631) );
na02s01 TIMEBOOST_cell_7659 ( .a(TIMEBOOST_net_2460), .b(n_34509), .o(n_34568) );
in01s02 g750458 ( .a(n_29550), .o(n_29551) );
na02s06 g750459 ( .a(n_29530), .b(n_29630), .o(n_29550) );
in01f02 g750460 ( .a(n_29620), .o(n_29621) );
na02f02 g750461 ( .a(n_29585), .b(n_29603), .o(n_29620) );
na02s06 g750462 ( .a(n_29500), .b(n_25738), .o(n_29596) );
na02f04 g750463 ( .a(FE_OCP_RBN2669_n_29500), .b(FE_OFN775_n_25834), .o(n_29549) );
na02m08 g750464 ( .a(FE_OCP_RBN2668_n_29500), .b(FE_OFN775_n_25834), .o(n_29616) );
na02s01 g750465 ( .a(n_30552), .b(n_30520), .o(n_30521) );
in01s01 g750466 ( .a(n_30518), .o(n_30519) );
na02f06 g750467 ( .a(n_30475), .b(n_29990), .o(n_30518) );
na02s01 g750468 ( .a(n_30549), .b(n_30548), .o(n_30550) );
in01m02 g750471 ( .a(n_29590), .o(n_29602) );
no02m04 g750472 ( .a(n_29574), .b(FE_OCPN1366_n_29573), .o(n_29590) );
in01s01 g750473 ( .a(n_29589), .o(n_29641) );
na02f04 g750474 ( .a(n_29574), .b(FE_OCPN1366_n_29573), .o(n_29589) );
no02m06 g750475 ( .a(n_29572), .b(FE_OCPN1918_n_29571), .o(n_29622) );
in01s01 g750476 ( .a(n_29587), .o(n_29588) );
na02m06 g750477 ( .a(n_29572), .b(FE_OCPN1918_n_29571), .o(n_29587) );
na03m04 TIMEBOOST_cell_8322 ( .a(FE_OCP_RBN3090_n_4872), .b(n_4879), .c(n_4898), .o(n_5085) );
na02s01 g750479 ( .a(n_29570), .b(n_29526), .o(n_29607) );
na02s01 TIMEBOOST_cell_2832 ( .a(n_7036), .b(n_7037), .o(TIMEBOOST_net_707) );
no03s20 TIMEBOOST_cell_2192 ( .a(FE_RN_1956_0), .b(FE_OCPN4520_n_32820), .c(FE_OCP_RBN3990_n_32772), .o(n_32856) );
oa12f06 g750486 ( .a(n_29444), .b(n_29542), .c(n_29498), .o(n_29606) );
in01s01 g750487 ( .a(n_29564), .o(n_29565) );
ao12f06 g750488 ( .a(n_29466), .b(n_29558), .c(n_29516), .o(n_29564) );
oa12s01 g750489 ( .a(n_29560), .b(n_29559), .c(n_29558), .o(n_31012) );
oa12s01 g750492 ( .a(n_29544), .b(n_29543), .c(n_29542), .o(n_31125) );
ao12s01 g750493 ( .a(n_30481), .b(n_30480), .c(n_30479), .o(n_31171) );
in01s01 g750494 ( .a(n_31256), .o(n_31211) );
oa12s01 g750495 ( .a(n_30478), .b(n_30477), .c(n_30476), .o(n_31256) );
in01m02 g750497 ( .a(n_29545), .o(n_29562) );
no02m08 TIMEBOOST_cell_5129 ( .a(TIMEBOOST_net_1512), .b(n_34225), .o(n_34289) );
na02s06 TIMEBOOST_cell_8689 ( .a(TIMEBOOST_net_2831), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_36983) );
in01f04 g750502 ( .a(n_29585), .o(n_29586) );
na02f06 g750504 ( .a(n_29518), .b(FE_OFN774_n_25834), .o(n_29603) );
na02m08 TIMEBOOST_cell_2831 ( .a(n_7222), .b(TIMEBOOST_net_706), .o(n_7284) );
no03f06 TIMEBOOST_cell_8329 ( .a(n_14711), .b(n_14819), .c(n_14858), .o(n_14978) );
no02s01 g750509 ( .a(n_30480), .b(n_30479), .o(n_30481) );
na02f02 g750510 ( .a(n_29505), .b(n_29504), .o(n_29570) );
in01s01 g750511 ( .a(n_29525), .o(n_29526) );
no02f02 g750512 ( .a(n_29505), .b(n_29504), .o(n_29525) );
na02s01 g750513 ( .a(n_29558), .b(n_29559), .o(n_29560) );
na02s01 g750514 ( .a(n_29542), .b(n_29543), .o(n_29544) );
na02s01 g750515 ( .a(n_30477), .b(n_30476), .o(n_30478) );
na02f06 TIMEBOOST_cell_2034 ( .a(TIMEBOOST_net_631), .b(n_29487), .o(n_29489) );
in01s01 g750519 ( .a(n_30475), .o(n_30552) );
oa12f06 g750520 ( .a(n_30002), .b(n_30441), .c(n_29998), .o(n_30475) );
na02s06 TIMEBOOST_cell_1933 ( .a(n_32433), .b(n_32577), .o(TIMEBOOST_net_581) );
in01s01 g750526 ( .a(n_29502), .o(n_29523) );
in01s02 g750527 ( .a(n_29480), .o(n_29502) );
ao22m04 g750528 ( .a(n_29386), .b(n_28803), .c(n_29385), .d(n_28802), .o(n_29480) );
in01s02 g750529 ( .a(n_29530), .o(n_29501) );
in01s04 g750532 ( .a(n_29479), .o(n_29530) );
na03f08 TIMEBOOST_cell_8282 ( .a(n_44872), .b(n_38209), .c(n_37944), .o(n_38034) );
no02f06 TIMEBOOST_cell_4141 ( .a(n_35576), .b(n_35575), .o(TIMEBOOST_net_1161) );
na02m06 g750538 ( .a(n_29453), .b(n_29476), .o(n_29572) );
in01s01 g750539 ( .a(n_29555), .o(n_29556) );
oa12s01 g750540 ( .a(n_29497), .b(n_29496), .c(n_29495), .o(n_29555) );
no02f04 g750544 ( .a(n_29399), .b(n_47251), .o(n_29428) );
no02s04 TIMEBOOST_cell_4140 ( .a(TIMEBOOST_net_1160), .b(n_11458), .o(n_11604) );
na02s06 g750546 ( .a(n_29378), .b(n_29379), .o(n_29406) );
no02s01 g750547 ( .a(n_30441), .b(n_29937), .o(n_30442) );
na02s01 g750548 ( .a(n_30441), .b(n_29910), .o(n_30480) );
na02m02 g750549 ( .a(n_29422), .b(n_30111), .o(n_29454) );
no03m08 TIMEBOOST_cell_8281 ( .a(n_33882), .b(FE_RN_2846_0), .c(FE_RN_2845_0), .o(n_33969) );
na02m04 g750551 ( .a(n_29419), .b(n_29260), .o(n_29476) );
na02s03 g750552 ( .a(n_29418), .b(n_29231), .o(n_29453) );
na02s01 g750553 ( .a(n_29583), .b(n_29633), .o(n_29584) );
no02s01 g750554 ( .a(n_29498), .b(n_29445), .o(n_29543) );
na02s01 g750555 ( .a(n_29496), .b(n_29495), .o(n_29497) );
na02m04 TIMEBOOST_cell_2001 ( .a(n_33609), .b(n_33216), .o(TIMEBOOST_net_615) );
na02f06 g750562 ( .a(n_29381), .b(n_29270), .o(n_29451) );
in01s04 g750564 ( .a(n_29481), .o(n_29473) );
na02s08 g750565 ( .a(n_29401), .b(n_29241), .o(n_29481) );
oa12s01 g750566 ( .a(n_29884), .b(n_30440), .c(n_30332), .o(n_30477) );
in01f02 g750567 ( .a(n_29485), .o(n_29507) );
no02f08 g750570 ( .a(n_29446), .b(n_29424), .o(n_29518) );
in01s01 g750571 ( .a(n_30214), .o(n_29472) );
in01s01 g750572 ( .a(n_29450), .o(n_30214) );
ao12f06 g750575 ( .a(n_29443), .b(n_29396), .c(n_29322), .o(n_29542) );
na02f02 g750576 ( .a(n_29403), .b(n_29382), .o(n_29505) );
oa12f06 g750577 ( .a(n_29413), .b(n_29513), .c(n_29465), .o(n_29558) );
ao12s01 g750578 ( .a(n_29515), .b(n_29514), .c(n_29513), .o(n_30917) );
in01s01 g750579 ( .a(FE_OCP_RBN2652_n_29448), .o(n_30310) );
no02s02 TIMEBOOST_cell_2005 ( .a(n_7943), .b(n_7415), .o(TIMEBOOST_net_617) );
in01s01 g750590 ( .a(n_31172), .o(n_30474) );
ao12s01 g750591 ( .a(n_30434), .b(n_30440), .c(n_30433), .o(n_31172) );
no02s04 TIMEBOOST_cell_6106 ( .a(TIMEBOOST_net_1904), .b(n_3300), .o(n_3403) );
no02s02 g750593 ( .a(n_29329), .b(n_28848), .o(n_29405) );
na02f08 TIMEBOOST_cell_2004 ( .a(n_616), .b(TIMEBOOST_net_616), .o(n_628) );
na02s06 TIMEBOOST_cell_7395 ( .a(TIMEBOOST_net_2328), .b(n_17159), .o(n_17367) );
no02f08 g750596 ( .a(n_29395), .b(n_25738), .o(n_29446) );
no02f06 g750597 ( .a(n_30192), .b(FE_OFN774_n_25834), .o(n_29424) );
na02s01 TIMEBOOST_cell_5032 ( .a(n_41605), .b(FE_OCP_RBN6592_n_41491), .o(TIMEBOOST_net_1464) );
no02m08 TIMEBOOST_cell_6182 ( .a(TIMEBOOST_net_1942), .b(n_10507), .o(n_10599) );
na02f08 g750600 ( .a(n_30394), .b(n_29936), .o(n_30441) );
no02s01 g750601 ( .a(n_30440), .b(n_30433), .o(n_30434) );
in01m04 g750602 ( .a(n_29385), .o(n_29386) );
ao12m06 g750603 ( .a(n_28761), .b(n_29353), .c(n_28742), .o(n_29385) );
in01s02 g750604 ( .a(n_29383), .o(n_29384) );
oa12s04 g750605 ( .a(n_28784), .b(n_29353), .c(n_28828), .o(n_29383) );
in01m04 g750606 ( .a(n_29422), .o(n_29475) );
no02m06 g750607 ( .a(FE_OCP_RBN2060_n_29380), .b(n_29328), .o(n_29422) );
no02f06 g750608 ( .a(n_29421), .b(FE_OCPUNCON1745_n_29420), .o(n_29498) );
in01s01 g750609 ( .a(n_29444), .o(n_29445) );
na02f06 g750610 ( .a(n_29421), .b(FE_OCPUNCON1745_n_29420), .o(n_29444) );
na02m02 g750611 ( .a(n_29380), .b(n_46960), .o(n_29382) );
na02f02 g750612 ( .a(FE_OCP_RBN2059_n_29380), .b(n_29327), .o(n_29403) );
na02m06 g750613 ( .a(n_29491), .b(FE_OCP_DRV_N5145_n_28349), .o(n_29583) );
na02m08 g750614 ( .a(n_29492), .b(n_28350), .o(n_29633) );
na02s01 g750615 ( .a(n_29516), .b(n_29467), .o(n_29559) );
no02s01 g750616 ( .a(n_29513), .b(n_29514), .o(n_29515) );
no02s01 g750617 ( .a(n_29443), .b(n_29397), .o(n_29496) );
na02f04 g750618 ( .a(n_29380), .b(n_29239), .o(n_29381) );
in01m02 g750619 ( .a(n_29418), .o(n_29419) );
in01m04 g750620 ( .a(n_29401), .o(n_29418) );
no02m06 TIMEBOOST_cell_8747 ( .a(TIMEBOOST_net_2860), .b(n_14539), .o(TIMEBOOST_net_2224) );
ao12m06 g750622 ( .a(FE_OFN773_n_25834), .b(n_29272), .c(n_29160), .o(n_29407) );
in01s01 g750625 ( .a(n_29417), .o(n_29442) );
na02s06 g750626 ( .a(n_29330), .b(n_29352), .o(n_29417) );
oa12s01 g750627 ( .a(n_29438), .b(n_29437), .c(n_29436), .o(n_30859) );
in01s01 g750628 ( .a(n_29441), .o(n_31045) );
ao12s01 g750629 ( .a(n_29374), .b(n_29373), .c(n_29372), .o(n_29441) );
ao12s01 g750630 ( .a(n_30420), .b(n_30419), .c(n_30418), .o(n_31189) );
in01m02 g750631 ( .a(n_29399), .o(n_29400) );
in01s01 g750633 ( .a(FE_OCP_RBN4156_n_29378), .o(n_29398) );
na02s02 g750637 ( .a(n_29303), .b(n_28850), .o(n_29352) );
na02s02 g750638 ( .a(n_29353), .b(n_28849), .o(n_29330) );
na02m08 TIMEBOOST_cell_2845 ( .a(n_7560), .b(TIMEBOOST_net_713), .o(n_7659) );
no02s01 g750641 ( .a(n_30419), .b(n_30418), .o(n_30420) );
no02f06 TIMEBOOST_cell_8847 ( .a(TIMEBOOST_net_2910), .b(TIMEBOOST_net_659), .o(n_30619) );
no02f04 g750644 ( .a(n_29376), .b(FE_OCPN1288_n_29375), .o(n_29443) );
in01s01 g750645 ( .a(n_29396), .o(n_29397) );
na02f04 g750646 ( .a(n_29376), .b(FE_OCPN1288_n_29375), .o(n_29396) );
in01s01 g750647 ( .a(n_29466), .o(n_29467) );
no02s01 g750650 ( .a(n_29465), .b(n_29414), .o(n_29514) );
na02s01 g750651 ( .a(n_29436), .b(n_29437), .o(n_29438) );
no02m08 g750653 ( .a(n_29280), .b(n_28801), .o(n_29347) );
no02s01 g750654 ( .a(n_29373), .b(n_29372), .o(n_29374) );
na02s01 g750655 ( .a(n_31145), .b(n_30393), .o(n_30432) );
in01s02 g750657 ( .a(n_29329), .o(n_29345) );
oa12m06 g750658 ( .a(n_28798), .b(n_29279), .c(n_28804), .o(n_29329) );
ao12m04 g750661 ( .a(n_25738), .b(n_29327), .c(n_29262), .o(n_29328) );
in01s01 g750662 ( .a(n_30394), .o(n_30440) );
ao12f06 g750663 ( .a(n_30304), .b(n_30337), .c(n_29887), .o(n_30394) );
in01m02 g750664 ( .a(n_29343), .o(n_29344) );
oa12m04 g750665 ( .a(n_28789), .b(FE_OCP_RBN5645_n_29236), .c(n_28787), .o(n_29343) );
in01f04 g750666 ( .a(n_30192), .o(n_29395) );
no02m02 TIMEBOOST_cell_1922 ( .a(n_22476), .b(TIMEBOOST_net_575), .o(n_22593) );
na02s02 TIMEBOOST_cell_4063 ( .a(n_4547), .b(n_4366), .o(TIMEBOOST_net_1122) );
in01s03 g750669 ( .a(n_29491), .o(n_29492) );
na02m08 g750670 ( .a(n_29415), .b(n_29393), .o(n_29491) );
ao12f06 g750671 ( .a(n_29340), .b(n_29389), .c(n_29436), .o(n_29513) );
in01s01 g750678 ( .a(n_30703), .o(n_30832) );
na02m06 TIMEBOOST_cell_6008 ( .a(TIMEBOOST_net_1855), .b(n_28893), .o(TIMEBOOST_net_248) );
no02f02 TIMEBOOST_cell_8797 ( .a(TIMEBOOST_net_2885), .b(n_14571), .o(TIMEBOOST_net_2127) );
in01s01 g750681 ( .a(n_30416), .o(n_30417) );
oa12s01 g750682 ( .a(n_30360), .b(n_30359), .c(n_30358), .o(n_30416) );
in01s01 g750683 ( .a(n_29353), .o(n_29303) );
no02s08 g750684 ( .a(n_29236), .b(n_28788), .o(n_29353) );
no02s02 TIMEBOOST_cell_7927 ( .a(TIMEBOOST_net_2594), .b(n_4974), .o(TIMEBOOST_net_908) );
no02m08 g750686 ( .a(n_29279), .b(FE_OCP_RBN2500_n_28773), .o(n_29280) );
na02s01 g750687 ( .a(n_30359), .b(n_30358), .o(n_30360) );
no02f04 g750689 ( .a(n_29265), .b(n_29143), .o(n_29302) );
no03m06 TIMEBOOST_cell_8252 ( .a(n_14506), .b(n_14505), .c(n_14607), .o(TIMEBOOST_net_1546) );
na02s02 g750691 ( .a(n_29217), .b(FE_OFN773_n_25834), .o(n_29241) );
na02s06 g750694 ( .a(n_29368), .b(n_30136), .o(n_29393) );
na02m08 g750695 ( .a(n_29369), .b(FE_OCP_RBN2567_n_29163), .o(n_29415) );
no02s01 g750696 ( .a(n_30338), .b(n_29886), .o(n_30419) );
no02f08 g750697 ( .a(n_29263), .b(n_28740), .o(n_29301) );
no02s01 TIMEBOOST_cell_8506 ( .a(n_37856), .b(n_37857), .o(TIMEBOOST_net_2740) );
no02f04 g750699 ( .a(n_29392), .b(FE_OCPUNCON3466_n_29391), .o(n_29465) );
in01s01 g750700 ( .a(n_29413), .o(n_29414) );
na02m04 g750701 ( .a(n_29392), .b(FE_OCPUNCON3466_n_29391), .o(n_29413) );
no02s04 TIMEBOOST_cell_6656 ( .a(TIMEBOOST_net_2085), .b(n_25142), .o(n_25223) );
na02s02 TIMEBOOST_cell_4136 ( .a(TIMEBOOST_net_1158), .b(n_10861), .o(n_10959) );
na02s01 g750706 ( .a(n_29389), .b(n_29341), .o(n_29437) );
no02s01 TIMEBOOST_cell_1991 ( .a(n_19014), .b(n_18280), .o(TIMEBOOST_net_610) );
in01s01 TIMEBOOST_cell_5921 ( .a(FE_OFN1_n_43918), .o(TIMEBOOST_net_1810) );
in01m02 g750710 ( .a(n_29477), .o(n_30111) );
no02s08 TIMEBOOST_cell_1919 ( .a(n_31993), .b(n_32106), .o(TIMEBOOST_net_574) );
na02f04 g750712 ( .a(n_29269), .b(n_29235), .o(n_29376) );
in01s01 g750713 ( .a(n_29322), .o(n_29495) );
oa12f06 g750714 ( .a(n_29189), .b(n_29299), .c(n_29190), .o(n_29322) );
in01s02 g750715 ( .a(FE_OCP_RBN2611_n_29298), .o(n_30191) );
na02f06 g750719 ( .a(n_29198), .b(n_29219), .o(n_29298) );
na02s02 TIMEBOOST_cell_5190 ( .a(FE_OCP_RBN6633_n_2633), .b(n_3058), .o(TIMEBOOST_net_1543) );
ao12s01 g750721 ( .a(n_29268), .b(n_29299), .c(n_29267), .o(n_29373) );
ao12s01 g750722 ( .a(n_30341), .b(n_30340), .c(n_30339), .o(n_31145) );
in01m02 g750723 ( .a(n_29271), .o(n_29272) );
no02s06 TIMEBOOST_cell_8145 ( .a(TIMEBOOST_net_2703), .b(n_13839), .o(n_14018) );
no02m04 g750726 ( .a(n_29194), .b(n_28766), .o(n_29240) );
na02m02 g750727 ( .a(n_29196), .b(n_28769), .o(n_29198) );
na02m04 g750728 ( .a(n_29169), .b(n_28768), .o(n_29219) );
na02s04 TIMEBOOST_cell_6642 ( .a(TIMEBOOST_net_2078), .b(n_41502), .o(n_41672) );
no02s01 g750730 ( .a(n_30340), .b(n_30339), .o(n_30341) );
na02m06 g750731 ( .a(n_29327), .b(n_25738), .o(n_29270) );
na02f04 g750732 ( .a(n_46960), .b(FE_OFN774_n_25834), .o(n_29239) );
in01s01 g750733 ( .a(n_30337), .o(n_30338) );
ao12f06 g750734 ( .a(n_30307), .b(n_30306), .c(n_29882), .o(n_30337) );
no02m04 g750736 ( .a(n_28725), .b(n_29218), .o(n_29236) );
na02f02 g750737 ( .a(n_29215), .b(FE_OCP_RBN2582_n_29091), .o(n_29235) );
na02f04 g750738 ( .a(n_29216), .b(FE_OCP_RBN2583_n_29091), .o(n_29269) );
na02f08 TIMEBOOST_cell_5189 ( .a(TIMEBOOST_net_1542), .b(n_15628), .o(n_15765) );
no02s04 g750740 ( .a(n_29316), .b(n_29167), .o(n_29319) );
in01s01 g750741 ( .a(n_29340), .o(n_29341) );
no02s01 g750744 ( .a(n_29299), .b(n_29267), .o(n_29268) );
na02m10 g750746 ( .a(n_29165), .b(n_28851), .o(n_29279) );
ao12s01 g750747 ( .a(n_30307), .b(n_30306), .c(n_29850), .o(n_30359) );
in01f02 g750748 ( .a(n_29265), .o(n_29266) );
in01f04 g750749 ( .a(n_29233), .o(n_29265) );
no02s01 TIMEBOOST_cell_6824 ( .a(TIMEBOOST_net_2169), .b(FE_OCP_RBN3402_n_43775), .o(FE_RN_1622_0) );
in01s06 g750751 ( .a(n_29368), .o(n_29369) );
in01m06 g750752 ( .a(n_29339), .o(n_29368) );
in01f04 g750755 ( .a(n_29232), .o(n_29263) );
na02m04 TIMEBOOST_cell_2850 ( .a(n_37368), .b(n_37142), .o(TIMEBOOST_net_716) );
in01s01 g750768 ( .a(n_29231), .o(n_29260) );
in01m03 g750769 ( .a(n_29217), .o(n_29231) );
oa12f06 g750771 ( .a(n_29156), .b(n_29313), .c(n_29158), .o(n_29436) );
in01s01 g750773 ( .a(n_29364), .o(n_29365) );
oa12s01 g750774 ( .a(n_29291), .b(n_29313), .c(n_29290), .o(n_29364) );
na02f10 g750775 ( .a(n_29164), .b(n_28734), .o(n_29218) );
in01m02 g750776 ( .a(n_29196), .o(n_29169) );
na02m08 g750777 ( .a(n_29120), .b(n_28805), .o(n_29196) );
no02s01 g750778 ( .a(n_30306), .b(n_30290), .o(n_30340) );
no02f06 TIMEBOOST_cell_4435 ( .a(n_16052), .b(n_14452), .o(TIMEBOOST_net_1308) );
no02s02 TIMEBOOST_cell_1908 ( .a(n_31476), .b(TIMEBOOST_net_568), .o(n_31607) );
na02m08 g750784 ( .a(n_29121), .b(n_28724), .o(n_29165) );
na02s01 g750785 ( .a(n_29313), .b(n_29290), .o(n_29291) );
in01m02 g750786 ( .a(n_29193), .o(n_29194) );
no02m02 g750787 ( .a(n_29164), .b(n_28746), .o(n_29193) );
in01f02 g750788 ( .a(n_29215), .o(n_29216) );
in01f02 g750789 ( .a(n_29192), .o(n_29215) );
ao12f06 g750790 ( .a(n_29379), .b(n_29115), .c(n_29033), .o(n_29192) );
na02s06 TIMEBOOST_cell_8710 ( .a(FE_RN_1375_0), .b(FE_RN_1374_0), .o(TIMEBOOST_net_2842) );
in01m06 g750795 ( .a(n_46960), .o(n_29327) );
in01s02 g750800 ( .a(FE_OCP_RBN2567_n_29163), .o(n_30136) );
na02m04 g750802 ( .a(n_29097), .b(n_29065), .o(n_29163) );
na02s01 TIMEBOOST_cell_6859 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_0_), .o(TIMEBOOST_net_2188) );
in01s01 g750804 ( .a(n_31116), .o(n_30393) );
oa12s01 g750805 ( .a(n_30336), .b(n_30335), .c(n_30334), .o(n_31116) );
no02f10 g750806 ( .a(n_29118), .b(n_28645), .o(n_29164) );
na02m04 g750808 ( .a(n_29092), .b(n_28701), .o(n_29122) );
no02s01 TIMEBOOST_cell_4043 ( .a(n_20081), .b(n_20022), .o(TIMEBOOST_net_1112) );
no02s01 TIMEBOOST_cell_8662 ( .a(FE_OCP_RBN6872_n_31520), .b(n_31017), .o(TIMEBOOST_net_2818) );
in01m03 g750811 ( .a(n_29120), .o(n_29121) );
na02m08 g750812 ( .a(n_29095), .b(n_28718), .o(n_29120) );
no02f08 g750813 ( .a(n_30335), .b(n_30256), .o(n_30306) );
na02s01 g750814 ( .a(n_30335), .b(n_30334), .o(n_30336) );
na02s06 TIMEBOOST_cell_1937 ( .a(n_1467), .b(n_1455), .o(TIMEBOOST_net_583) );
na02s02 TIMEBOOST_cell_1973 ( .a(n_18477), .b(n_18440), .o(TIMEBOOST_net_601) );
in01s02 g750817 ( .a(n_29144), .o(n_29145) );
na02m04 g750818 ( .a(n_29118), .b(n_28770), .o(n_29144) );
no02f04 g750819 ( .a(n_29188), .b(n_29187), .o(n_29190) );
na02f04 g750820 ( .a(n_29188), .b(n_29187), .o(n_29189) );
no02m06 TIMEBOOST_cell_8561 ( .a(TIMEBOOST_net_2767), .b(n_29605), .o(n_29657) );
no02f08 TIMEBOOST_cell_5183 ( .a(TIMEBOOST_net_1539), .b(n_15356), .o(n_15510) );
na02s01 g750823 ( .a(FE_OCP_RBN2583_n_29091), .b(n_29058), .o(n_29211) );
in01s02 g750824 ( .a(n_29116), .o(n_29117) );
no02m02 g750825 ( .a(n_29095), .b(n_28774), .o(n_29116) );
na02m10 g750827 ( .a(n_29210), .b(n_29094), .o(n_29258) );
in01s04 g750832 ( .a(n_29143), .o(n_29161) );
in01s06 g750838 ( .a(n_29167), .o(n_29160) );
na02m08 g750839 ( .a(n_29064), .b(n_29038), .o(n_29167) );
no02f06 g750840 ( .a(n_29180), .b(n_29159), .o(n_29313) );
in01s01 g750841 ( .a(n_29228), .o(n_29229) );
ao22s01 g750842 ( .a(FE_OCP_RBN2049_n_29056), .b(FE_OCP_DRV_N3502_n_29140), .c(FE_OCP_DRV_N6263_FE_OCP_RBN5603_n_29056), .d(n_27961), .o(n_29228) );
na02f10 g750843 ( .a(n_29063), .b(n_28567), .o(n_29118) );
no02m08 g750844 ( .a(n_29039), .b(n_28678), .o(n_29095) );
na02m06 TIMEBOOST_cell_8138 ( .a(FE_OCP_RBN5552_n_23328), .b(n_23178), .o(TIMEBOOST_net_2700) );
no02s02 TIMEBOOST_cell_4042 ( .a(n_16104), .b(TIMEBOOST_net_1111), .o(n_16263) );
in01f02 g750849 ( .a(n_29115), .o(n_29141) );
na02f06 g750850 ( .a(n_29056), .b(FE_OFN774_n_25834), .o(n_29115) );
na02m08 g750851 ( .a(n_29055), .b(FE_OFN773_n_25834), .o(n_29094) );
no02f04 g750852 ( .a(FE_OCP_RBN2564_n_29110), .b(n_29053), .o(n_29159) );
no02f04 g750853 ( .a(n_29137), .b(FE_OCP_RBN5025_n_29053), .o(n_29180) );
no02s02 g750854 ( .a(n_30235), .b(n_30233), .o(n_30267) );
in01s01 g750855 ( .a(n_29188), .o(n_29372) );
na02f06 g750856 ( .a(FE_OCP_RBN5604_n_29056), .b(FE_OCP_DRV_N3502_n_29140), .o(n_29188) );
no02m04 g750857 ( .a(n_29157), .b(FE_OCPN1268_n_29155), .o(n_29158) );
na02m04 g750858 ( .a(n_29157), .b(FE_OCPN1268_n_29155), .o(n_29156) );
na02s01 g750859 ( .a(n_29055), .b(FE_OCP_RBN5026_n_29053), .o(n_29139) );
no02s01 g750861 ( .a(n_29113), .b(n_30364), .o(n_29112) );
no02f04 g750863 ( .a(n_29063), .b(n_28683), .o(n_29092) );
no02f06 g750864 ( .a(n_30168), .b(n_30040), .o(n_30335) );
in01m08 g750865 ( .a(n_29154), .o(n_29210) );
oa22s01 g750874 ( .a(FE_OCP_RBN5022_n_29080), .b(n_29109), .c(FE_OCP_RBN5023_n_29080), .d(n_27914), .o(n_30671) );
in01m02 g750877 ( .a(n_29062), .o(n_29292) );
no02f08 g750879 ( .a(n_29020), .b(n_28605), .o(n_29063) );
in01f02 g750882 ( .a(FE_OCP_RBN2565_n_29110), .o(n_29137) );
na02f06 g750884 ( .a(n_29054), .b(FE_OFN773_n_25834), .o(n_29110) );
na02f04 g750886 ( .a(n_29020), .b(n_28682), .o(n_29034) );
na02s01 g750887 ( .a(n_29059), .b(n_30399), .o(n_29060) );
no04s02 TIMEBOOST_cell_6562 ( .a(n_5546), .b(n_5212), .c(n_5213), .d(n_5545), .o(n_5746) );
in01s01 g750889 ( .a(n_29157), .o(n_29135) );
no02m04 g750890 ( .a(n_29080), .b(n_29109), .o(n_29157) );
in01s01 TIMEBOOST_cell_5909 ( .a(FE_OFN1_n_43918), .o(TIMEBOOST_net_1798) );
ao12s02 g750892 ( .a(n_30156), .b(n_30183), .c(n_29852), .o(n_30235) );
in01f02 g750893 ( .a(n_29057), .o(n_29058) );
in01f02 g750896 ( .a(n_29033), .o(n_29057) );
in01s01 g750910 ( .a(n_29113), .o(n_29083) );
ao12s01 g750911 ( .a(n_29016), .b(n_29015), .c(FE_OFN5079_n_29014), .o(n_29113) );
in01s01 g750912 ( .a(FE_OCPN5132_n_29081), .o(n_29082) );
ao12s01 g750913 ( .a(n_29013), .b(n_29012), .c(n_29011), .o(n_29081) );
in01s01 g750914 ( .a(n_31294), .o(n_30392) );
no02s02 g750915 ( .a(n_30333), .b(n_30305), .o(n_31294) );
na02f08 g750916 ( .a(n_28976), .b(n_28600), .o(n_29020) );
in01s02 g750917 ( .a(n_28979), .o(n_29018) );
no02m08 g750918 ( .a(n_28952), .b(n_28627), .o(n_28979) );
in01s02 g750919 ( .a(n_28977), .o(n_28978) );
na02s04 g750920 ( .a(n_28952), .b(n_28726), .o(n_28977) );
no02s01 g750921 ( .a(n_29015), .b(FE_OFN5079_n_29014), .o(n_29016) );
no02s01 g750922 ( .a(n_29012), .b(n_29011), .o(n_29013) );
no02m04 TIMEBOOST_cell_8524 ( .a(n_33675), .b(n_34037), .o(TIMEBOOST_net_2749) );
no02s01 g750924 ( .a(n_30068), .b(n_30289), .o(n_30333) );
no02s01 g750925 ( .a(n_30105), .b(n_30288), .o(n_30305) );
no02s02 g750926 ( .a(n_30185), .b(n_30254), .o(n_30255) );
na02s01 g750927 ( .a(n_30229), .b(n_30208), .o(n_30253) );
in01s01 g750928 ( .a(n_30233), .o(n_30234) );
oa12s02 g750929 ( .a(n_30208), .b(n_30130), .c(n_29944), .o(n_30233) );
in01f02 g750930 ( .a(n_28997), .o(n_28998) );
oa12s01 g750933 ( .a(n_28975), .b(n_28974), .c(n_28973), .o(n_29031) );
in01s01 g750934 ( .a(n_29059), .o(n_29913) );
oa12s01 g750935 ( .a(n_28972), .b(n_28971), .c(n_28970), .o(n_29059) );
in01m01 g750940 ( .a(n_29054), .o(n_29080) );
in01f01 g750944 ( .a(n_29030), .o(n_29053) );
na02s01 g750947 ( .a(n_28974), .b(n_28973), .o(n_28975) );
na02s01 g750948 ( .a(n_28971), .b(n_28970), .o(n_28972) );
no02s03 TIMEBOOST_cell_1791 ( .a(n_5946), .b(n_4875), .o(TIMEBOOST_net_510) );
in01s01 g750950 ( .a(n_30105), .o(n_30068) );
na02f04 g750951 ( .a(n_30039), .b(n_29821), .o(n_30105) );
no02s02 g750952 ( .a(n_30039), .b(n_30038), .o(n_30040) );
no02s01 g750953 ( .a(n_30811), .b(n_30089), .o(n_30167) );
in01f02 g750954 ( .a(n_28950), .o(n_28951) );
na02f04 g750955 ( .a(n_28935), .b(n_28652), .o(n_28950) );
ao12f04 g750957 ( .a(n_28526), .b(n_28871), .c(n_28530), .o(n_28968) );
oa12s01 g750958 ( .a(n_28815), .b(n_28967), .c(n_28867), .o(n_29015) );
oa12s01 g750959 ( .a(n_28509), .b(n_28967), .c(n_28510), .o(n_29012) );
in01f04 g750960 ( .a(n_28965), .o(n_28966) );
oa12f06 g750961 ( .a(n_28681), .b(n_28934), .c(n_28568), .o(n_28965) );
na02s02 g750962 ( .a(n_30231), .b(n_30162), .o(n_30232) );
oa12s01 g750963 ( .a(n_30231), .b(n_30182), .c(n_30156), .o(n_30975) );
in01s02 g750964 ( .a(n_30229), .o(n_30230) );
no02s02 g750965 ( .a(n_30811), .b(n_30163), .o(n_30229) );
in01s01 g750966 ( .a(n_30185), .o(n_30186) );
ao12s01 g750967 ( .a(n_30097), .b(n_30166), .c(n_30165), .o(n_30185) );
in01s01 g750968 ( .a(n_30183), .o(n_30184) );
oa12s02 g750969 ( .a(n_30097), .b(n_30164), .c(n_30166), .o(n_30183) );
ao22s01 g750970 ( .a(n_28871), .b(n_28886), .c(n_28967), .d(n_28885), .o(n_30364) );
in01s01 g750971 ( .a(n_30102), .o(n_30103) );
oa12s01 g750972 ( .a(n_30005), .b(n_30004), .c(n_30003), .o(n_30102) );
oa22s01 g750973 ( .a(n_30166), .b(n_30303), .c(n_29883), .d(n_30156), .o(n_31119) );
oa22s01 g750974 ( .a(FE_OCPUNCON3480_n_28872), .b(n_28865), .c(FE_OCPUNCON3479_n_28872), .d(n_28866), .o(n_29898) );
in01f02 g750975 ( .a(n_28948), .o(n_28949) );
na02f06 g750976 ( .a(n_28934), .b(FE_OCP_RBN4035_n_28651), .o(n_28948) );
na02f06 g750977 ( .a(n_29947), .b(n_29820), .o(n_30039) );
na02s01 g750978 ( .a(n_30004), .b(n_30003), .o(n_30005) );
no02s01 g750979 ( .a(n_30129), .b(n_29856), .o(n_30130) );
na02s01 g750980 ( .a(n_30182), .b(n_29944), .o(n_30231) );
na02s01 g750981 ( .a(n_30100), .b(n_30099), .o(n_30101) );
no02s01 g750982 ( .a(n_30127), .b(n_30088), .o(n_30128) );
oa12s01 g750983 ( .a(n_28632), .b(n_28933), .c(n_28485), .o(n_28974) );
oa12s01 g750984 ( .a(n_28887), .b(n_28933), .c(n_28842), .o(n_28971) );
oa12s01 g750985 ( .a(n_30067), .b(n_30064), .c(n_29944), .o(n_30163) );
na02s01 g750986 ( .a(n_30100), .b(n_30036), .o(n_30811) );
oa12s02 g750987 ( .a(n_30035), .b(n_29996), .c(n_29944), .o(n_30098) );
no02s02 g750988 ( .a(n_30001), .b(n_29946), .o(n_30002) );
ao12s01 g750989 ( .a(n_30254), .b(n_30207), .c(n_30303), .o(n_31090) );
in01s01 g750991 ( .a(n_30399), .o(n_28996) );
oa22s01 g750992 ( .a(n_28890), .b(n_28914), .c(n_28933), .d(n_28915), .o(n_30399) );
ao22s01 g750995 ( .a(n_29880), .b(n_179), .c(n_29879), .d(n_186), .o(n_31043) );
in01s01 g750996 ( .a(FE_OCP_DRV_N5304_n_29892), .o(n_28995) );
oa22s01 g750997 ( .a(n_28869), .b(n_28913), .c(n_28870), .d(n_28912), .o(n_29892) );
no02s01 g750999 ( .a(n_30161), .b(n_30124), .o(n_30162) );
no02s01 g751000 ( .a(n_30161), .b(n_30129), .o(n_30902) );
no02s01 g751001 ( .a(n_30207), .b(n_30097), .o(n_30254) );
no02s01 g751002 ( .a(n_30438), .b(n_30164), .o(n_31041) );
ao12s01 g751004 ( .a(n_28505), .b(n_28853), .c(n_28474), .o(n_28872) );
in01s01 g751006 ( .a(n_28871), .o(n_28967) );
ao12f08 g751011 ( .a(n_28529), .b(n_28853), .c(n_28511), .o(n_28871) );
in01s01 g751012 ( .a(n_29947), .o(n_30004) );
in01s01 TIMEBOOST_cell_8896 ( .a(n_1142), .o(TIMEBOOST_net_2940) );
na02s02 g751014 ( .a(n_30093), .b(n_30159), .o(n_30160) );
oa12s01 g751015 ( .a(n_29907), .b(n_29886), .c(n_29818), .o(n_29887) );
in01s01 g751016 ( .a(n_30067), .o(n_30127) );
oa12s01 g751017 ( .a(n_29932), .b(n_30089), .c(n_30030), .o(n_30067) );
oa12s01 g751018 ( .a(n_29909), .b(n_30037), .c(n_30083), .o(n_30100) );
oa12s01 g751019 ( .a(n_29909), .b(n_29977), .c(n_30086), .o(n_30036) );
in01s01 g751020 ( .a(n_30034), .o(n_30035) );
ao12s02 g751021 ( .a(n_29944), .b(n_30000), .c(n_29999), .o(n_30034) );
in01s01 g751022 ( .a(n_30001), .o(n_29910) );
ao12s01 g751023 ( .a(n_29837), .b(n_29884), .c(n_29935), .o(n_30001) );
ao12s01 g751024 ( .a(n_29837), .b(n_29945), .c(n_29938), .o(n_29946) );
oa12s01 g751025 ( .a(n_30097), .b(n_30096), .c(n_30095), .o(n_30208) );
na02f08 g751026 ( .a(n_28894), .b(n_28893), .o(n_28934) );
in01s01 g751027 ( .a(n_28891), .o(n_28892) );
ao12s01 g751028 ( .a(n_28833), .b(n_28853), .c(n_28832), .o(n_28891) );
in01s01 g751029 ( .a(n_30166), .o(n_29883) );
oa12s01 g751030 ( .a(n_29825), .b(n_29824), .c(n_29823), .o(n_30166) );
in01s01 g751031 ( .a(n_29856), .o(n_30182) );
oa12s01 g751032 ( .a(n_29806), .b(n_29805), .c(n_29804), .o(n_29856) );
no02s01 g751033 ( .a(n_28853), .b(n_28832), .o(n_28833) );
no02m20 TIMEBOOST_cell_2953 ( .a(n_2151), .b(TIMEBOOST_net_767), .o(n_45903) );
na02s01 g751035 ( .a(n_29805), .b(n_29804), .o(n_29806) );
na02s01 g751036 ( .a(n_29824), .b(n_29823), .o(n_29825) );
no02s01 g751037 ( .a(n_30059), .b(n_30094), .o(n_30159) );
no02s01 g751038 ( .a(n_30092), .b(n_30091), .o(n_30093) );
no02s01 g751039 ( .a(n_30085), .b(n_30157), .o(n_30158) );
na02s01 g751040 ( .a(n_30028), .b(n_30065), .o(n_30066) );
no02s02 g751041 ( .a(n_29881), .b(n_29878), .o(n_29882) );
na02s01 g751042 ( .a(n_29997), .b(n_29974), .o(n_29998) );
na02s01 g751043 ( .a(n_29997), .b(n_29945), .o(n_30479) );
na02s01 g751044 ( .a(n_30126), .b(n_30099), .o(n_30785) );
no02s01 g751045 ( .a(n_30090), .b(n_29995), .o(n_30616) );
no02s01 g751046 ( .a(n_29822), .b(n_29819), .o(n_30003) );
in01s01 g751047 ( .a(n_29879), .o(n_29880) );
na02s01 g751048 ( .a(n_29854), .b(n_29853), .o(n_29879) );
no02s01 g751049 ( .a(n_30290), .b(n_30256), .o(n_30334) );
no02s01 g751050 ( .a(n_30094), .b(n_30089), .o(n_30892) );
no02s01 g751051 ( .a(n_30097), .b(n_30033), .o(n_30161) );
no02s01 g751052 ( .a(n_30088), .b(n_30063), .o(n_30064) );
no02s01 g751053 ( .a(n_29995), .b(n_29600), .o(n_29996) );
in01s01 g751054 ( .a(n_30062), .o(n_30129) );
na02s01 g751055 ( .a(n_29932), .b(n_30033), .o(n_30062) );
in01s01 g751056 ( .a(n_30061), .o(n_30164) );
na02s01 g751057 ( .a(n_30165), .b(n_29909), .o(n_30061) );
no02s01 g751058 ( .a(n_29886), .b(n_29878), .o(n_30358) );
no02s01 g751059 ( .a(n_30332), .b(n_29836), .o(n_30433) );
no02s01 g751060 ( .a(n_30381), .b(n_29939), .o(n_30520) );
no02s01 g751061 ( .a(n_30380), .b(n_30037), .o(n_30635) );
no02s01 g751062 ( .a(n_30303), .b(n_30165), .o(n_30438) );
na02s01 g751063 ( .a(n_30431), .b(n_30029), .o(n_30900) );
no02s01 g751064 ( .a(n_30091), .b(n_30088), .o(n_30951) );
in01s01 g751065 ( .a(n_28869), .o(n_28870) );
ao12s01 g751066 ( .a(n_28501), .b(n_28852), .c(n_28547), .o(n_28869) );
ao12s01 g751067 ( .a(n_30304), .b(n_30303), .c(n_29907), .o(n_30418) );
ao12s01 g751068 ( .a(n_29881), .b(n_30156), .c(n_29838), .o(n_30339) );
ao12s01 g751069 ( .a(n_29975), .b(n_30303), .c(n_29534), .o(n_30548) );
oa12s01 g751070 ( .a(n_30065), .b(n_30156), .c(n_29992), .o(n_30689) );
ao12s01 g751071 ( .a(n_30157), .b(n_30303), .c(n_30086), .o(n_30837) );
oa12s01 g751072 ( .a(n_30060), .b(n_30156), .c(n_29781), .o(n_30897) );
in01s01 g751073 ( .a(n_30412), .o(n_30413) );
ao12s01 g751074 ( .a(n_30092), .b(n_30303), .c(n_30063), .o(n_30412) );
in01s01 g751075 ( .a(n_30124), .o(n_30125) );
ao12s01 g751076 ( .a(n_29909), .b(n_30095), .c(n_29756), .o(n_30124) );
in01s01 g751078 ( .a(n_28933), .o(n_28890) );
in01s01 g751079 ( .a(n_28894), .o(n_28933) );
ao12f08 g751080 ( .a(n_28507), .b(n_28852), .c(n_28532), .o(n_28894) );
in01s01 g751081 ( .a(n_28888), .o(n_28889) );
ao22s01 g751082 ( .a(n_28852), .b(n_28570), .c(n_28807), .d(n_28569), .o(n_28888) );
in01s01 g751083 ( .a(n_29852), .o(n_30207) );
ao12s01 g751084 ( .a(n_29803), .b(n_29802), .c(n_29801), .o(n_29852) );
in01s01 g751085 ( .a(n_30288), .o(n_30289) );
oa22s01 g751086 ( .a(n_30097), .b(n_30038), .c(n_30156), .d(n_30104), .o(n_30288) );
oa22s01 g751087 ( .a(n_30303), .b(n_29490), .c(n_30156), .d(n_29935), .o(n_30476) );
oa22s01 g751088 ( .a(n_30303), .b(n_29535), .c(n_30156), .d(n_29999), .o(n_30589) );
oa22s01 g751089 ( .a(n_30303), .b(n_30083), .c(n_30156), .d(n_29691), .o(n_30720) );
ao22s01 g751090 ( .a(n_30156), .b(n_29797), .c(n_30303), .d(n_30095), .o(n_30972) );
in01s01 g751115 ( .a(n_30546), .o(n_30614) );
in01s02 g751122 ( .a(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_30588) );
in01s04 g751124 ( .a(FE_OFN5087_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_30546) );
in01s01 g751126 ( .a(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_30504) );
in01s02 g751138 ( .a(n_30587), .o(n_30612) );
in01s01 g751139 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_30587) );
in01s02 g751145 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_30545) );
no02s01 g751151 ( .a(n_29802), .b(n_29801), .o(n_29803) );
no02s01 g751152 ( .a(n_30097), .b(n_29817), .o(n_30332) );
in01s01 g751153 ( .a(n_30059), .o(n_30060) );
no02s01 g751154 ( .a(n_29932), .b(n_30030), .o(n_30059) );
in01s01 g751155 ( .a(n_29821), .o(n_29822) );
na02s02 g751156 ( .a(n_29800), .b(n_29799), .o(n_29821) );
no02s01 g751157 ( .a(n_29932), .b(n_29768), .o(n_30091) );
na02s01 g751158 ( .a(n_30156), .b(n_29993), .o(n_30431) );
no02s01 g751159 ( .a(n_30097), .b(n_29335), .o(n_30290) );
no02s01 g751160 ( .a(n_30303), .b(n_30082), .o(n_30380) );
in01s01 g751161 ( .a(n_30096), .o(n_30029) );
no02s01 g751162 ( .a(n_29944), .b(n_29993), .o(n_30096) );
no02s01 g751163 ( .a(n_30303), .b(n_29908), .o(n_30381) );
no02s01 g751164 ( .a(n_29944), .b(n_29709), .o(n_30089) );
no02s01 g751165 ( .a(n_29944), .b(n_29767), .o(n_30088) );
in01s01 g751166 ( .a(n_29943), .o(n_30037) );
na02s01 g751167 ( .a(n_29909), .b(n_30082), .o(n_29943) );
in01s01 g751168 ( .a(n_29977), .o(n_30099) );
no02s01 g751169 ( .a(n_29944), .b(n_29942), .o(n_29977) );
no02s01 g751170 ( .a(n_29932), .b(n_29710), .o(n_30094) );
no02s01 g751171 ( .a(n_29932), .b(n_30063), .o(n_30092) );
no02s01 g751172 ( .a(n_29909), .b(n_30086), .o(n_30157) );
in01s01 g751173 ( .a(n_30126), .o(n_30085) );
na02s01 g751174 ( .a(n_29944), .b(n_29942), .o(n_30126) );
in01s01 g751175 ( .a(n_29995), .o(n_29976) );
no02s01 g751176 ( .a(n_29837), .b(n_29940), .o(n_29995) );
in01s01 g751177 ( .a(n_30000), .o(n_29939) );
na02s01 g751178 ( .a(n_29909), .b(n_29908), .o(n_30000) );
na02s01 g751179 ( .a(n_29944), .b(n_29992), .o(n_30065) );
in01s01 g751180 ( .a(n_30028), .o(n_30090) );
na02s01 g751181 ( .a(n_29944), .b(n_29940), .o(n_30028) );
in01s01 g751182 ( .a(n_29945), .o(n_29877) );
na02s01 g751183 ( .a(n_29818), .b(n_29851), .o(n_29945) );
in01s01 g751184 ( .a(n_29881), .o(n_29850) );
no02s02 g751185 ( .a(n_29837), .b(n_29838), .o(n_29881) );
no02s02 g751186 ( .a(n_29837), .b(n_29312), .o(n_29878) );
na02f04 g751187 ( .a(n_29800), .b(n_28928), .o(n_29854) );
na02s06 g751188 ( .a(FE_OCP_RBN2860_n_29800), .b(n_28929), .o(n_29853) );
in01s02 g751189 ( .a(n_29819), .o(n_29820) );
no02s02 g751190 ( .a(n_29800), .b(n_29799), .o(n_29819) );
no02s02 g751191 ( .a(n_29837), .b(n_29359), .o(n_30256) );
no02s02 g751192 ( .a(n_29818), .b(n_29311), .o(n_29886) );
no02s02 g751193 ( .a(n_29818), .b(n_29907), .o(n_30304) );
in01s01 g751194 ( .a(n_29974), .o(n_29975) );
na02s01 g751195 ( .a(n_29837), .b(n_29938), .o(n_29974) );
in01s01 g751196 ( .a(n_29937), .o(n_29997) );
no02s01 g751197 ( .a(n_29909), .b(n_29851), .o(n_29937) );
in01s01 g751198 ( .a(n_29884), .o(n_29836) );
na02s01 g751199 ( .a(n_29818), .b(n_29817), .o(n_29884) );
ao12f08 g751200 ( .a(n_28468), .b(n_28791), .c(n_28504), .o(n_28853) );
ao12s01 g751201 ( .a(n_29128), .b(n_29771), .c(n_29124), .o(n_29805) );
oa12s01 g751202 ( .a(n_29334), .b(n_29783), .c(n_29310), .o(n_29824) );
ao12s01 g751203 ( .a(n_29909), .b(n_30083), .c(n_30082), .o(n_30084) );
oa12s01 g751204 ( .a(n_29944), .b(n_29999), .c(n_29509), .o(n_29990) );
no02s02 g751205 ( .a(n_29818), .b(n_29360), .o(n_30307) );
oa12s01 g751206 ( .a(n_29837), .b(n_29935), .c(n_29408), .o(n_29936) );
oa12s01 g751208 ( .a(n_28780), .b(n_28791), .c(n_28779), .o(n_28830) );
oa12s01 g751209 ( .a(n_29770), .b(n_29783), .c(n_29769), .o(n_30165) );
oa12s01 g751210 ( .a(n_29761), .b(n_29771), .c(n_29760), .o(n_30033) );
na02s01 g751211 ( .a(n_28791), .b(n_28779), .o(n_28780) );
na02s01 g751212 ( .a(n_29771), .b(n_29760), .o(n_29761) );
na02s01 g751213 ( .a(n_29783), .b(n_29769), .o(n_29770) );
in01s01 g751214 ( .a(n_28852), .o(n_28807) );
oa12f08 g751215 ( .a(FE_OCPN896_n_28506), .b(n_28790), .c(FE_OCPN894_n_28471), .o(n_28852) );
in01s06 g751216 ( .a(n_29818), .o(n_29837) );
in01s02 g751229 ( .a(n_30156), .o(n_30303) );
in01s02 g751236 ( .a(n_30097), .o(n_30156) );
in01s01 g751240 ( .a(n_29944), .o(n_30097) );
in01s01 g751252 ( .a(n_29944), .o(n_29932) );
in01s03 g751253 ( .a(n_29909), .o(n_29944) );
in01s04 g751254 ( .a(n_29837), .o(n_29909) );
in01s04 g751259 ( .a(n_29800), .o(n_29818) );
no02s06 TIMEBOOST_cell_2952 ( .a(FE_RN_2560_0), .b(FE_RN_2555_0), .o(TIMEBOOST_net_767) );
in01s01 g751262 ( .a(FE_OCP_DRV_N6884_n_28829), .o(n_29866) );
oa12s01 g751263 ( .a(n_28778), .b(n_28790), .c(n_28777), .o(n_28829) );
ao12s01 g751264 ( .a(n_29250), .b(n_29722), .c(n_29203), .o(n_29802) );
in01s01 g751265 ( .a(n_30095), .o(n_29797) );
oa12s01 g751266 ( .a(n_29759), .b(n_29758), .c(n_29757), .o(n_30095) );
oa12s01 g751267 ( .a(n_29748), .b(n_29747), .c(n_29746), .o(n_30063) );
in01s01 g751268 ( .a(n_29767), .o(n_29768) );
ao12s01 g751269 ( .a(n_29725), .b(n_29724), .c(n_29723), .o(n_29767) );
na02s01 g751270 ( .a(n_28790), .b(n_28777), .o(n_28778) );
na02s01 g751271 ( .a(n_29758), .b(n_29757), .o(n_29759) );
na02s01 g751272 ( .a(n_29747), .b(n_29746), .o(n_29748) );
na02s01 g751273 ( .a(n_29744), .b(n_29249), .o(n_29783) );
no02s01 g751274 ( .a(n_29724), .b(n_29723), .o(n_29725) );
oa12f08 g751275 ( .a(n_28448), .b(n_28748), .c(n_28423), .o(n_28791) );
ao12s01 g751276 ( .a(n_29205), .b(n_29721), .c(n_29150), .o(n_29771) );
no02m02 TIMEBOOST_cell_4009 ( .a(n_35221), .b(n_35253), .o(TIMEBOOST_net_1095) );
oa22s01 g751278 ( .a(n_28708), .b(n_28463), .c(n_28748), .d(n_28464), .o(n_29844) );
in01s01 g751279 ( .a(n_29993), .o(n_29756) );
ao12s01 g751280 ( .a(n_29713), .b(n_29712), .c(n_29711), .o(n_29993) );
in01s01 g751281 ( .a(n_30030), .o(n_29781) );
oa12s01 g751282 ( .a(n_29743), .b(n_29742), .c(n_29741), .o(n_30030) );
oa12s01 g751283 ( .a(n_29694), .b(n_29693), .c(n_29692), .o(n_30086) );
na02s01 g751284 ( .a(n_29742), .b(n_29741), .o(n_29743) );
na02s01 g751285 ( .a(n_29693), .b(n_29692), .o(n_29694) );
no02s01 g751286 ( .a(n_29712), .b(n_29711), .o(n_29713) );
oa12f08 g751287 ( .a(n_28465), .b(n_28747), .c(n_28439), .o(n_28790) );
in01s01 g751288 ( .a(n_29744), .o(n_29722) );
na02f08 g751289 ( .a(n_29721), .b(n_29202), .o(n_29744) );
no02s01 TIMEBOOST_cell_1875 ( .a(FE_OCP_RBN3222_n_21242), .b(FE_OCP_RBN3251_n_21312), .o(TIMEBOOST_net_552) );
ao12s01 g751291 ( .a(n_29051), .b(n_29708), .c(n_29072), .o(n_29747) );
oa12s01 g751292 ( .a(n_29050), .b(n_29649), .c(n_29308), .o(n_29724) );
oa22s01 g751294 ( .a(n_28747), .b(n_28487), .c(n_28707), .d(n_28486), .o(n_28775) );
in01s01 g751295 ( .a(n_29709), .o(n_29710) );
ao12s01 g751296 ( .a(n_29652), .b(n_29651), .c(n_29650), .o(n_29709) );
in01s01 g751297 ( .a(n_30083), .o(n_29691) );
oa12s01 g751298 ( .a(n_29639), .b(n_29638), .c(n_29637), .o(n_30083) );
ao12s01 g751299 ( .a(n_29655), .b(n_29654), .c(n_29653), .o(n_29942) );
no02s01 g751300 ( .a(n_29654), .b(n_29653), .o(n_29655) );
no02f08 g751301 ( .a(n_29675), .b(n_29098), .o(n_29721) );
na02s01 g751302 ( .a(n_29638), .b(n_29637), .o(n_29639) );
na02s01 g751303 ( .a(n_29675), .b(n_29132), .o(n_29712) );
no02s01 g751304 ( .a(n_29651), .b(n_29650), .o(n_29652) );
in01s01 g751305 ( .a(n_28748), .o(n_28708) );
oa12f08 g751306 ( .a(n_28420), .b(n_28685), .c(n_28389), .o(n_28748) );
ao12s01 g751307 ( .a(n_29333), .b(n_29599), .c(n_29043), .o(n_29693) );
no02m01 TIMEBOOST_cell_1855 ( .a(n_21490), .b(n_21521), .o(TIMEBOOST_net_542) );
ao12s01 g751309 ( .a(n_28661), .b(n_28685), .c(n_28660), .o(n_29812) );
no02s01 g751310 ( .a(n_28685), .b(n_28660), .o(n_28661) );
na02s01 g751311 ( .a(n_29598), .b(n_29332), .o(n_29654) );
na02f08 g751312 ( .a(n_29130), .b(n_29636), .o(n_29675) );
in01s01 g751313 ( .a(n_29649), .o(n_29708) );
na02s01 g751314 ( .a(n_29636), .b(n_29045), .o(n_29649) );
na02s01 g751315 ( .a(n_29597), .b(n_28961), .o(n_29651) );
in01s01 g751316 ( .a(n_28747), .o(n_28707) );
oa12f08 g751317 ( .a(n_28421), .b(n_28684), .c(n_28387), .o(n_28747) );
ao12s01 g751318 ( .a(n_29243), .b(n_29601), .c(n_29285), .o(n_29638) );
ao12s01 g751319 ( .a(n_28659), .b(n_28684), .c(n_28658), .o(n_29860) );
oa12s01 g751320 ( .a(n_29582), .b(n_29601), .c(n_29581), .o(n_30082) );
in01s01 g751321 ( .a(n_29600), .o(n_29992) );
oa12s01 g751322 ( .a(n_29538), .b(n_29537), .c(n_29536), .o(n_29600) );
no02s01 g751323 ( .a(n_28684), .b(n_28658), .o(n_28659) );
in01s01 g751324 ( .a(n_29598), .o(n_29599) );
na02s01 g751325 ( .a(n_29601), .b(n_29074), .o(n_29598) );
na02s01 g751326 ( .a(n_29537), .b(n_29536), .o(n_29538) );
na02s01 g751327 ( .a(n_29601), .b(n_29581), .o(n_29582) );
oa12f08 g751328 ( .a(n_28403), .b(n_28612), .c(n_28357), .o(n_28685) );
in01f04 g751329 ( .a(n_29597), .o(n_29636) );
na02f06 g751330 ( .a(n_29601), .b(n_29102), .o(n_29597) );
in01s01 g751331 ( .a(FE_OCPN1256_n_28656), .o(n_28657) );
ao22s01 g751332 ( .a(n_28612), .b(n_28416), .c(n_28552), .d(n_28415), .o(n_28656) );
ao12s01 g751333 ( .a(n_29512), .b(n_29511), .c(n_29510), .o(n_29940) );
in01s01 g751334 ( .a(n_29999), .o(n_29535) );
ao12s01 g751335 ( .a(n_29461), .b(n_29460), .c(n_29459), .o(n_29999) );
in01s01 g751336 ( .a(n_29938), .o(n_29534) );
ao12s01 g751337 ( .a(n_29464), .b(n_29463), .c(n_29462), .o(n_29938) );
no02s06 g751338 ( .a(n_28806), .b(n_28744), .o(n_28851) );
no02s01 g751339 ( .a(n_29463), .b(n_29462), .o(n_29464) );
no02s01 g751340 ( .a(n_29460), .b(n_29459), .o(n_29461) );
no02s01 g751341 ( .a(n_29511), .b(n_29510), .o(n_29512) );
oa12f08 g751342 ( .a(n_28404), .b(n_28611), .c(n_28355), .o(n_28684) );
na02f06 g751343 ( .a(n_29489), .b(n_29048), .o(n_29601) );
in01s01 g751344 ( .a(FE_OCPUNCON3470_n_28654), .o(n_28655) );
ao22s01 g751345 ( .a(n_28611), .b(n_28418), .c(n_28551), .d(n_28417), .o(n_28654) );
ao12s01 g751346 ( .a(n_29079), .b(n_29487), .c(n_29488), .o(n_29537) );
in01s01 g751347 ( .a(n_29908), .o(n_29509) );
oa12s01 g751348 ( .a(n_29433), .b(n_29432), .c(n_29431), .o(n_29908) );
in01s01 g751349 ( .a(n_29935), .o(n_29490) );
ao12s01 g751350 ( .a(n_29411), .b(n_29410), .c(n_29409), .o(n_29935) );
oa12s01 g751351 ( .a(n_29458), .b(n_29457), .c(n_29456), .o(n_29851) );
na02m01 g751352 ( .a(n_29036), .b(FE_OCP_RBN2499_FE_RN_1553_0), .o(n_28774) );
in01m02 g751353 ( .a(n_28805), .o(n_28806) );
no02f06 TIMEBOOST_cell_1854 ( .a(TIMEBOOST_net_541), .b(n_26846), .o(n_26847) );
no02s01 g751355 ( .a(n_29410), .b(n_29409), .o(n_29411) );
na02s01 g751356 ( .a(n_29457), .b(n_29456), .o(n_29458) );
no02s01 g751357 ( .a(n_29487), .b(n_29047), .o(n_29511) );
na02s01 g751358 ( .a(n_29432), .b(n_29431), .o(n_29433) );
no02s02 g751359 ( .a(n_28788), .b(n_28743), .o(n_28789) );
in01s01 g751360 ( .a(n_28612), .o(n_28552) );
ao12f08 g751361 ( .a(n_28320), .b(n_28536), .c(n_28344), .o(n_28612) );
no02s01 TIMEBOOST_cell_6339 ( .a(n_39600), .b(FE_OCP_RBN6159_n_39816), .o(TIMEBOOST_net_2021) );
ao12s01 g751363 ( .a(n_28908), .b(n_29361), .c(n_28991), .o(n_29463) );
ao12s01 g751364 ( .a(n_29010), .b(n_29388), .c(n_29006), .o(n_29460) );
in01s01 g751365 ( .a(FE_OCP_DRV_N6275_n_28582), .o(n_28583) );
ao12s01 g751366 ( .a(n_28515), .b(n_28536), .c(n_28514), .o(n_28582) );
no02s04 g751367 ( .a(n_28745), .b(n_28626), .o(n_29017) );
na02s02 g751368 ( .a(n_28770), .b(n_28631), .o(n_28746) );
in01s02 g751369 ( .a(n_29036), .o(n_28771) );
no02m08 g751370 ( .a(n_28745), .b(n_28607), .o(n_29036) );
no02s01 g751371 ( .a(n_28536), .b(n_28514), .o(n_28515) );
na02s01 g751372 ( .a(n_29362), .b(n_28946), .o(n_29457) );
no02s01 g751373 ( .a(n_29388), .b(n_28960), .o(n_29432) );
no02f04 TIMEBOOST_cell_3197 ( .a(TIMEBOOST_net_889), .b(n_9867), .o(n_10023) );
in01s01 g751376 ( .a(n_28611), .o(n_28551) );
oa12f08 g751377 ( .a(n_28402), .b(n_28535), .c(n_28353), .o(n_28611) );
oa12s01 g751378 ( .a(n_29171), .b(n_29363), .c(n_29200), .o(n_29410) );
no02f06 g751379 ( .a(n_29358), .b(n_29007), .o(n_29487) );
ao12s01 g751380 ( .a(n_28513), .b(n_28535), .c(n_28512), .o(n_29777) );
in01s01 g751381 ( .a(n_29817), .o(n_29408) );
oa12s01 g751382 ( .a(n_29337), .b(n_29363), .c(n_29336), .o(n_29817) );
na02s02 g751383 ( .a(n_28682), .b(n_28522), .o(n_28683) );
no02s01 g751384 ( .a(n_28535), .b(n_28512), .o(n_28513) );
in01s02 g751385 ( .a(n_28745), .o(n_28726) );
na02s08 g751386 ( .a(FE_OCP_RBN4036_n_28651), .b(n_28579), .o(n_28745) );
no02m02 g751387 ( .a(n_28651), .b(n_28577), .o(n_28681) );
in01s01 g751388 ( .a(n_29361), .o(n_29362) );
no02s01 g751389 ( .a(n_29363), .b(n_28927), .o(n_29361) );
na02s01 g751390 ( .a(n_29363), .b(n_29336), .o(n_29337) );
in01m02 g751391 ( .a(n_28705), .o(n_28770) );
no02s01 g751393 ( .a(n_29838), .b(n_29359), .o(n_29360) );
oa12f08 g751394 ( .a(n_28318), .b(n_28478), .c(n_28288), .o(n_28536) );
in01f04 g751395 ( .a(n_29388), .o(n_29358) );
no02f06 g751396 ( .a(n_29363), .b(n_28992), .o(n_29388) );
oa22s01 g751397 ( .a(n_28441), .b(n_28329), .c(n_28478), .d(n_28330), .o(n_29715) );
in01s01 g751398 ( .a(n_29311), .o(n_29312) );
ao12s01 g751399 ( .a(n_29227), .b(n_29226), .c(n_29225), .o(n_29311) );
oa12s01 g751400 ( .a(n_29288), .b(n_29287), .c(n_29286), .o(n_29907) );
in01s01 TIMEBOOST_cell_7378 ( .a(TIMEBOOST_net_2314), .o(TIMEBOOST_net_2313) );
na02s01 g751404 ( .a(n_29287), .b(n_29286), .o(n_29288) );
no02s01 g751405 ( .a(n_29226), .b(n_29225), .o(n_29227) );
no02m04 g751406 ( .a(n_28610), .b(n_28534), .o(n_28682) );
oa12f08 g751407 ( .a(n_28316), .b(n_28477), .c(n_28341), .o(n_28535) );
no02f06 g751408 ( .a(n_29224), .b(n_28959), .o(n_29363) );
oa12s01 g751409 ( .a(n_28455), .b(n_28477), .c(n_28454), .o(n_29765) );
oa12s01 g751410 ( .a(n_29256), .b(n_29255), .c(n_29254), .o(n_29838) );
in01m04 g751412 ( .a(n_28610), .o(n_28652) );
na02s08 g751413 ( .a(n_28527), .b(n_28520), .o(n_28610) );
no02m08 g751414 ( .a(n_28609), .b(n_28608), .o(n_28893) );
na02s01 g751415 ( .a(n_29255), .b(n_29254), .o(n_29256) );
no02f04 g751416 ( .a(n_29176), .b(n_29223), .o(n_29224) );
na02s01 g751417 ( .a(n_28477), .b(n_28454), .o(n_28455) );
in01s01 g751418 ( .a(n_28478), .o(n_28441) );
oa12f08 g751419 ( .a(n_28284), .b(n_28428), .c(n_28252), .o(n_28478) );
na02s02 TIMEBOOST_cell_7031 ( .a(n_3853), .b(n_3760), .o(TIMEBOOST_net_2274) );
oa12s01 g751421 ( .a(n_28958), .b(n_29177), .c(n_28878), .o(n_29226) );
na02s06 g751422 ( .a(n_28475), .b(n_28467), .o(n_28511) );
in01s01 g751424 ( .a(n_28649), .o(n_28650) );
ao12m01 g751425 ( .a(n_28460), .b(n_28631), .c(n_28630), .o(n_28649) );
na02m06 g751426 ( .a(n_28437), .b(n_28496), .o(n_28532) );
in01s01 g751427 ( .a(n_28476), .o(n_29737) );
oa12s01 g751428 ( .a(n_28427), .b(FE_OCP_DRV_N5143_n_28426), .c(n_28425), .o(n_28476) );
in01s01 TIMEBOOST_cell_7377 ( .a(TIMEBOOST_net_2313), .o(TIMEBOOST_net_2312) );
oa12s02 g751430 ( .a(n_28458), .b(n_28577), .c(delay_sub_ln21_0_unr17_stage7_stallmux_q_21_), .o(n_28579) );
ao12s01 g751433 ( .a(n_28407), .b(n_28428), .c(n_28406), .o(n_29644) );
ao12s01 g751434 ( .a(FE_OCP_RBN6555_n_28458), .b(n_28698), .c(n_27807), .o(n_28744) );
ao12s01 g751435 ( .a(FE_OCP_RBN5587_FE_RN_1367_0), .b(n_28773), .c(n_28795), .o(n_28804) );
na02s01 g751436 ( .a(n_28786), .b(n_28762), .o(n_28787) );
na02s01 g751437 ( .a(n_28719), .b(n_28721), .o(n_28725) );
no02s08 g751439 ( .a(n_28510), .b(n_28494), .o(n_28530) );
na02m10 g751440 ( .a(n_28493), .b(n_28528), .o(n_28529) );
in01s04 g751441 ( .a(n_28526), .o(n_28527) );
na02s08 g751442 ( .a(n_28509), .b(n_28508), .o(n_28526) );
na02s01 g751443 ( .a(n_28742), .b(n_28741), .o(n_28743) );
na02s06 g751444 ( .a(n_28491), .b(n_28489), .o(n_28507) );
na02m08 g751445 ( .a(n_28484), .b(n_28549), .o(n_28609) );
no02s01 g751447 ( .a(n_28736), .b(n_28723), .o(n_28724) );
na02s06 g751448 ( .a(n_28474), .b(n_28473), .o(n_28475) );
no02s01 g751449 ( .a(n_28574), .b(delay_add_ln22_unr17_stage7_stallmux_q_23_), .o(n_28575) );
in01s01 g751450 ( .a(n_28802), .o(n_28803) );
na02s01 g751451 ( .a(n_28786), .b(n_28741), .o(n_28802) );
in01s01 g751452 ( .a(n_28739), .o(n_28740) );
na02s01 g751453 ( .a(n_28722), .b(n_28721), .o(n_28739) );
no02s01 g751455 ( .a(n_28574), .b(n_28605), .o(n_28628) );
in01s02 g751456 ( .a(n_28572), .o(n_28573) );
no02s02 g751457 ( .a(n_28492), .b(n_28550), .o(n_28572) );
in01s02 g751458 ( .a(n_28603), .o(n_28604) );
no02s04 g751459 ( .a(n_28521), .b(n_28571), .o(n_28603) );
in01s01 g751460 ( .a(n_28679), .o(n_28680) );
no02s01 g751461 ( .a(n_28565), .b(n_28645), .o(n_28679) );
na02s02 g751463 ( .a(n_28720), .b(n_28719), .o(n_28737) );
in01s01 g751464 ( .a(n_28849), .o(n_28850) );
no02s01 g751465 ( .a(n_28785), .b(n_28828), .o(n_28849) );
na02s06 g751466 ( .a(n_28547), .b(n_28466), .o(n_28496) );
na02s01 g751467 ( .a(n_28549), .b(n_28548), .o(n_28973) );
in01s01 g751468 ( .a(n_28914), .o(n_28915) );
na02s01 g751469 ( .a(n_28843), .b(n_28887), .o(n_28914) );
na02s01 g751470 ( .a(n_28426), .b(n_28425), .o(n_28427) );
na02s01 g751471 ( .a(FE_OCPN896_n_28506), .b(n_28472), .o(n_28777) );
in01s01 g751472 ( .a(n_28569), .o(n_28570) );
na02s01 g751473 ( .a(n_28491), .b(n_28547), .o(n_28569) );
in01s01 g751474 ( .a(n_28601), .o(n_28602) );
no02s02 g751475 ( .a(n_28568), .b(n_28577), .o(n_28601) );
na02s06 g751476 ( .a(n_28548), .b(n_27654), .o(n_28525) );
in01s01 g751477 ( .a(n_28643), .o(n_28644) );
no02s02 g751478 ( .a(n_28627), .b(n_28626), .o(n_28643) );
in01s02 g751479 ( .a(n_28703), .o(n_28704) );
no02s06 g751480 ( .a(FE_RN_1553_0), .b(n_28678), .o(n_28703) );
in01s01 g751481 ( .a(n_28768), .o(n_28769) );
no02s01 g751482 ( .a(n_28736), .b(n_28735), .o(n_28768) );
no02s01 g751483 ( .a(n_28428), .b(n_28406), .o(n_28407) );
no02s01 g751485 ( .a(n_28801), .b(FE_OCP_RBN2500_n_28773), .o(n_28826) );
na02s01 g751486 ( .a(n_28798), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_30_), .o(n_28799) );
no02s01 g751487 ( .a(n_28505), .b(n_28451), .o(n_28832) );
in01s01 g751488 ( .a(n_28885), .o(n_28886) );
no02s01 g751489 ( .a(n_28816), .b(n_28867), .o(n_28885) );
na02s01 g751490 ( .a(n_28508), .b(n_28495), .o(n_29011) );
na02s01 g751491 ( .a(n_29177), .b(n_29201), .o(n_29255) );
in01s01 g751492 ( .a(n_28766), .o(n_28767) );
oa12s02 g751493 ( .a(n_28734), .b(FE_OCPN6917_n_28460), .c(n_28630), .o(n_28766) );
in01s01 g751494 ( .a(n_28624), .o(n_28625) );
na02s02 g751495 ( .a(n_28600), .b(n_28545), .o(n_28624) );
ao12s01 g751497 ( .a(n_28566), .b(n_28467), .c(delay_add_ln22_unr17_stage7_stallmux_q_23_), .o(n_28701) );
oa12f08 g751498 ( .a(n_28286), .b(n_28372), .c(n_28294), .o(n_28477) );
in01s01 g751499 ( .a(n_28676), .o(n_28677) );
ao12s02 g751500 ( .a(n_28608), .b(n_28458), .c(delay_sub_ln21_0_unr17_stage7_stallmux_q_19_), .o(n_28676) );
in01s01 g751501 ( .a(n_28912), .o(n_28913) );
ao12s01 g751502 ( .a(n_28490), .b(n_28817), .c(delay_sub_ln21_0_unr17_stage7_stallmux_q_15_), .o(n_28912) );
in01s01 g751503 ( .a(n_28732), .o(n_28733) );
oa12s01 g751504 ( .a(n_28718), .b(FE_OCP_RBN6555_n_28458), .c(n_28646), .o(n_28732) );
in01s02 g751505 ( .a(n_28674), .o(n_28675) );
ao22s04 g751506 ( .a(FE_OCP_RBN4031_n_28458), .b(n_28541), .c(FE_OCP_RBN4030_n_28458), .d(delay_sub_ln21_0_unr17_stage7_stallmux_q_21_), .o(n_28674) );
ao12s01 g751510 ( .a(n_28723), .b(FE_OCP_RBN2490_FE_RN_1367_0), .c(delay_sub_ln21_0_unr17_stage7_stallmux_q_27_), .o(n_28764) );
na02s01 g751511 ( .a(n_28469), .b(n_28504), .o(n_28779) );
in01s01 g751512 ( .a(n_28865), .o(n_28866) );
oa12s01 g751513 ( .a(n_28528), .b(FE_OCPN4849_n_28460), .c(n_28473), .o(n_28865) );
in01f02 g751514 ( .a(n_29175), .o(n_29176) );
no02m04 g751515 ( .a(n_29177), .b(n_28906), .o(n_29175) );
in01s01 g751516 ( .a(n_28824), .o(n_28825) );
oa22s01 g751517 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_31_), .c(n_28460), .d(n_27824), .o(n_28824) );
in01s01 g751518 ( .a(n_28822), .o(n_28823) );
ao22s01 g751519 ( .a(FE_OCPN6917_n_28460), .b(n_27834), .c(n_28467), .d(delay_add_ln22_unr17_stage7_stallmux_q_29_), .o(n_28822) );
oa22s01 g751520 ( .a(n_28817), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_), .c(FE_OCP_RBN5591_FE_RN_1367_0), .d(n_27623), .o(n_28970) );
oa22s01 g751522 ( .a(FE_OCP_RBN2490_FE_RN_1367_0), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_29_), .c(FE_OCP_RBN5590_FE_RN_1367_0), .d(n_28795), .o(n_28820) );
in01s01 g751523 ( .a(n_28847), .o(n_28848) );
oa22s01 g751524 ( .a(FE_OCP_RBN2490_FE_RN_1367_0), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_30_), .c(FE_OCP_RBN5590_FE_RN_1367_0), .d(n_27806), .o(n_28847) );
in01s01 g751525 ( .a(n_28845), .o(n_28846) );
oa22s01 g751526 ( .a(FE_OCP_RBN2490_FE_RN_1367_0), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_31_), .c(FE_OCP_RBN5590_FE_RN_1367_0), .d(n_27803), .o(n_28845) );
oa22s01 g751527 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_17_), .c(FE_OCPN4849_n_28460), .d(n_27712), .o(n_29014) );
in01s01 g751528 ( .a(n_29359), .o(n_29335) );
oa12s01 g751529 ( .a(n_29253), .b(n_29252), .c(n_29251), .o(n_29359) );
in01s01 g751531 ( .a(FE_OCPN894_n_28471), .o(n_28472) );
na02s01 g751533 ( .a(FE_OCPN6917_n_28460), .b(n_27833), .o(n_28786) );
in01s01 g751534 ( .a(n_28673), .o(n_28721) );
no02s01 g751535 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_26_), .o(n_28673) );
na02s01 g751536 ( .a(FE_OCPN6917_n_28460), .b(n_27860), .o(n_28719) );
na02s06 g751537 ( .a(FE_OCPN6917_n_28460), .b(n_28630), .o(n_28734) );
no02m02 g751538 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_24_), .o(n_28645) );
no02s02 g751539 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_22_), .o(n_28605) );
in01s01 g751540 ( .a(n_28494), .o(n_28495) );
no02s06 g751541 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_18_), .o(n_28494) );
no02s06 g751542 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_19_), .o(n_28571) );
in01s08 g751543 ( .a(n_28505), .o(n_28493) );
no02s10 g751544 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_14_), .o(n_28505) );
na02s06 g751545 ( .a(n_28438), .b(n_28473), .o(n_28528) );
in01s01 g751546 ( .a(n_28474), .o(n_28451) );
na02s06 g751547 ( .a(n_28419), .b(delay_add_ln22_unr17_stage7_stallmux_q_14_), .o(n_28474) );
in01s01 g751548 ( .a(n_28468), .o(n_28469) );
no02m08 g751549 ( .a(n_28450), .b(n_28449), .o(n_28468) );
na02m08 g751550 ( .a(n_28450), .b(n_28449), .o(n_28504) );
no02s02 g751551 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_20_), .o(n_28550) );
na02s06 g751552 ( .a(n_28460), .b(n_28523), .o(n_28600) );
in01s01 g751553 ( .a(n_28566), .o(n_28567) );
no02s01 g751554 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_23_), .o(n_28566) );
in01s01 g751555 ( .a(n_28522), .o(n_28574) );
na02m01 g751556 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_22_), .o(n_28522) );
na02s06 g751557 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_18_), .o(n_28508) );
in01s01 g751558 ( .a(n_28520), .o(n_28521) );
na02s03 g751559 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_19_), .o(n_28520) );
in01s01 g751560 ( .a(n_28533), .o(n_28492) );
na02s02 g751561 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_20_), .o(n_28533) );
in01s01 g751562 ( .a(n_28722), .o(n_28672) );
na02s01 g751563 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_26_), .o(n_28722) );
na02s01 g751564 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_27_), .o(n_28720) );
in01s01 g751565 ( .a(n_28631), .o(n_28565) );
na02f01 g751566 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_24_), .o(n_28631) );
na02s01 g751567 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_30_), .o(n_28741) );
in01s01 g751568 ( .a(n_28784), .o(n_28785) );
na02s01 g751569 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_28_), .o(n_28784) );
no02s01 g751570 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_28_), .o(n_28828) );
na02s01 g751571 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_21_), .o(n_28545) );
na02s08 g751572 ( .a(n_28437), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_14_), .o(n_28547) );
in01s01 g751574 ( .a(n_28491), .o(n_28501) );
in01s01 g751576 ( .a(n_28489), .o(n_28490) );
na02s06 g751577 ( .a(n_28447), .b(n_28466), .o(n_28489) );
na02s04 g751578 ( .a(n_28437), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_18_), .o(n_28548) );
na02s06 g751579 ( .a(n_28447), .b(n_27637), .o(n_28549) );
na02s01 g751580 ( .a(n_28817), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_), .o(n_28887) );
in01s01 g751581 ( .a(n_28842), .o(n_28843) );
no02s01 g751582 ( .a(n_28817), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_), .o(n_28842) );
no02s06 g751583 ( .a(n_28458), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_19_), .o(n_28608) );
in01s01 g751584 ( .a(n_28486), .o(n_28487) );
na02s01 g751585 ( .a(n_28440), .b(n_28465), .o(n_28486) );
no02s06 g751586 ( .a(n_28447), .b(n_27669), .o(n_28577) );
in01s06 g751587 ( .a(n_28568), .o(n_28544) );
no02s10 g751588 ( .a(n_28458), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_20_), .o(n_28568) );
na02s03 g751589 ( .a(FE_OCP_RBN6555_n_28458), .b(n_28646), .o(n_28718) );
in01s01 g751590 ( .a(n_28543), .o(n_28626) );
na02s02 g751591 ( .a(n_28458), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_22_), .o(n_28543) );
na02s06 g751593 ( .a(FE_OCP_RBN6553_n_28458), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_24_), .o(n_28647) );
no02s06 g751594 ( .a(FE_OCP_RBN6553_n_28458), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_24_), .o(n_28678) );
no02s02 g751596 ( .a(n_28458), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_22_), .o(n_28627) );
na02s06 g751597 ( .a(n_28447), .b(n_28541), .o(n_28542) );
in01s02 g751598 ( .a(n_28698), .o(n_28735) );
na02s02 g751599 ( .a(FE_OCP_RBN2490_FE_RN_1367_0), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_26_), .o(n_28698) );
no02s01 g751600 ( .a(FE_OCP_RBN2491_FE_RN_1367_0), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_26_), .o(n_28736) );
no02s01 g751601 ( .a(FE_OCP_RBN2490_FE_RN_1367_0), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_27_), .o(n_28723) );
na02s01 g751603 ( .a(FE_OCP_RBN2490_FE_RN_1367_0), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_28_), .o(n_28773) );
no02m01 g751604 ( .a(FE_OCP_RBN2490_FE_RN_1367_0), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_28_), .o(n_28801) );
in01s01 g751605 ( .a(n_28463), .o(n_28464) );
na02s01 g751606 ( .a(n_28448), .b(n_28424), .o(n_28463) );
in01s01 g751607 ( .a(n_28815), .o(n_28816) );
na02s01 g751608 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_16_), .o(n_28815) );
no02s01 g751609 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_16_), .o(n_28867) );
na02f04 g751610 ( .a(n_29252), .b(n_29105), .o(n_29177) );
na02s01 g751611 ( .a(n_29252), .b(n_29251), .o(n_29253) );
na02s01 g751612 ( .a(n_29249), .b(n_29103), .o(n_29250) );
in01s01 g751613 ( .a(n_28761), .o(n_28762) );
ao12m01 g751614 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_28_), .c(delay_add_ln22_unr17_stage7_stallmux_q_29_), .o(n_28761) );
na02s06 g751616 ( .a(n_28467), .b(n_27711), .o(n_28509) );
oa12m01 g751617 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_28_), .c(delay_add_ln22_unr17_stage7_stallmux_q_29_), .o(n_28742) );
in01s01 g751618 ( .a(n_28484), .o(n_28485) );
na02s06 g751619 ( .a(n_28447), .b(n_27642), .o(n_28484) );
ao12s01 g751621 ( .a(n_28371), .b(n_28391), .c(n_28293), .o(n_28426) );
oa12s06 g751622 ( .a(FE_OCP_RBN5590_FE_RN_1367_0), .b(n_28795), .c(n_27778), .o(n_28798) );
na02m04 g751623 ( .a(n_29249), .b(n_29174), .o(n_29248) );
oa12f08 g751624 ( .a(n_28250), .b(n_28373), .c(n_28210), .o(n_28428) );
ao12s01 g751625 ( .a(n_28370), .b(n_28391), .c(n_28369), .o(n_29573) );
oa22s01 g751626 ( .a(n_28335), .b(n_28265), .c(n_28373), .d(n_28266), .o(n_29571) );
in01s01 g751627 ( .a(n_28423), .o(n_28424) );
no02m06 g751628 ( .a(n_28405), .b(delay_add_ln22_unr17_stage7_stallmux_q_12_), .o(n_28423) );
na02m06 g751629 ( .a(n_28405), .b(delay_add_ln22_unr17_stage7_stallmux_q_12_), .o(n_28448) );
no02f08 g751630 ( .a(n_28391), .b(n_28371), .o(n_28372) );
in01s01 g751631 ( .a(n_28439), .o(n_28440) );
no02s08 g751632 ( .a(n_28422), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_12_), .o(n_28439) );
na02m06 g751633 ( .a(n_28422), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_12_), .o(n_28465) );
na02s01 g751634 ( .a(n_28421), .b(n_28388), .o(n_28658) );
na02s01 g751635 ( .a(n_28390), .b(n_28420), .o(n_28660) );
in01s02 g751655 ( .a(n_28467), .o(n_28460) );
in01f20 g751656 ( .a(n_28438), .o(n_28467) );
in01f10 g751658 ( .a(n_28419), .o(n_28438) );
na02f10 g751659 ( .a(n_28383), .b(n_28360), .o(n_28419) );
in01s01 g751669 ( .a(FE_OCP_RBN5591_FE_RN_1367_0), .o(n_28817) );
in01m20 g751691 ( .a(n_28447), .o(n_28458) );
in01m20 g751692 ( .a(n_28437), .o(n_28447) );
no02m04 TIMEBOOST_cell_8595 ( .a(TIMEBOOST_net_2784), .b(n_19755), .o(n_19886) );
no02m08 g751694 ( .a(n_28384), .b(n_28361), .o(n_28450) );
no02s01 g751696 ( .a(n_28369), .b(n_28391), .o(n_28370) );
ao12s04 g751697 ( .a(n_29205), .b(n_29125), .c(n_28919), .o(n_29249) );
oa12f04 g751698 ( .a(n_28962), .b(n_28994), .c(n_28793), .o(n_29252) );
oa12s01 g751699 ( .a(n_28364), .b(n_28363), .c(n_28362), .o(n_29576) );
na02f06 g751700 ( .a(n_28368), .b(n_28367), .o(n_28420) );
in01s01 g751701 ( .a(n_28389), .o(n_28390) );
no02m08 g751702 ( .a(n_28368), .b(n_28367), .o(n_28389) );
na02s06 g751703 ( .a(n_28366), .b(n_28365), .o(n_28421) );
oa12f08 g751704 ( .a(n_28247), .b(n_28303), .c(n_28223), .o(n_28391) );
in01s01 g751705 ( .a(n_28387), .o(n_28388) );
no02m08 g751706 ( .a(n_28366), .b(n_28365), .o(n_28387) );
in01s01 g751707 ( .a(n_28417), .o(n_28418) );
na02s01 g751708 ( .a(n_28356), .b(n_28404), .o(n_28417) );
na02s01 g751709 ( .a(n_28363), .b(n_28362), .o(n_28364) );
in01s01 g751710 ( .a(n_28415), .o(n_28416) );
na02s01 g751711 ( .a(n_28403), .b(n_28358), .o(n_28415) );
ao12s04 g751712 ( .a(n_28359), .b(n_27976), .c(n_28360), .o(n_28361) );
in01s04 g751714 ( .a(n_28383), .o(n_28384) );
na02s03 TIMEBOOST_cell_4307 ( .a(n_8187), .b(FE_OCP_RBN5609_n_7730), .o(TIMEBOOST_net_1244) );
na02s04 g751717 ( .a(n_29132), .b(n_29028), .o(n_29205) );
in01s01 g751718 ( .a(n_28373), .o(n_28335) );
ao12f08 g751719 ( .a(n_28147), .b(n_28322), .c(n_28187), .o(n_28373) );
no02s02 TIMEBOOST_cell_6792 ( .a(TIMEBOOST_net_2153), .b(n_4925), .o(TIMEBOOST_net_1314) );
in01s01 g751722 ( .a(FE_OCP_DRV_N5145_n_28349), .o(n_28350) );
oa12s01 g751723 ( .a(n_28312), .b(n_28322), .c(n_28311), .o(n_28349) );
in01s01 g751724 ( .a(n_30038), .o(n_30104) );
ao12s01 g751725 ( .a(n_29247), .b(n_29246), .c(n_29245), .o(n_30038) );
na02m10 g751726 ( .a(FE_OCPN3548_n_28043), .b(n_28334), .o(n_28359) );
na02f08 g751727 ( .a(n_28348), .b(delay_add_ln22_unr17_stage7_stallmux_q_10_), .o(n_28403) );
in01s01 g751728 ( .a(n_28357), .o(n_28358) );
no02f08 g751729 ( .a(n_28348), .b(delay_add_ln22_unr17_stage7_stallmux_q_10_), .o(n_28357) );
na02s03 g751730 ( .a(n_28334), .b(n_28332), .o(n_28333) );
na02s06 g751732 ( .a(n_28347), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_10_), .o(n_28404) );
in01s01 g751733 ( .a(n_28355), .o(n_28356) );
no02s06 g751734 ( .a(n_28347), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_10_), .o(n_28355) );
no02s01 TIMEBOOST_cell_6791 ( .a(FE_OCP_RBN2964_n_4046), .b(n_4316), .o(TIMEBOOST_net_2153) );
no02s06 g751736 ( .a(n_28319), .b(n_28091), .o(n_28331) );
na02s01 g751737 ( .a(n_28402), .b(n_28354), .o(n_28512) );
na02s01 g751738 ( .a(n_28222), .b(n_28304), .o(n_28363) );
na02s01 g751739 ( .a(n_28322), .b(n_28311), .o(n_28312) );
na02s01 g751740 ( .a(n_28321), .b(n_28344), .o(n_28514) );
no02m04 g751741 ( .a(n_29246), .b(n_28993), .o(n_28994) );
no02s01 g751742 ( .a(n_29246), .b(n_29245), .o(n_29247) );
na02s01 g751743 ( .a(n_29050), .b(n_29049), .o(n_29051) );
na02s01 g751744 ( .a(n_29029), .b(n_28988), .o(n_29079) );
in01s02 g751745 ( .a(n_29078), .o(n_29132) );
na02s02 g751746 ( .a(n_29050), .b(n_28990), .o(n_29078) );
ao12s02 g751747 ( .a(n_29047), .b(n_28989), .c(n_28919), .o(n_29048) );
oa12s01 g751748 ( .a(n_28919), .b(n_29104), .c(n_29172), .o(n_29174) );
na02m08 g751750 ( .a(n_28307), .b(n_28295), .o(n_28366) );
ao12s01 g751751 ( .a(n_28302), .b(FE_OCP_RBN2040_n_28268), .c(n_28300), .o(n_29504) );
no02m06 g751752 ( .a(n_28309), .b(n_28308), .o(n_28310) );
na02m10 TIMEBOOST_cell_8609 ( .a(TIMEBOOST_net_2791), .b(n_26147), .o(n_26318) );
no02s10 g751755 ( .a(n_28309), .b(n_28015), .o(n_28334) );
na02m08 g751756 ( .a(n_28306), .b(n_28305), .o(n_28344) );
in01s01 g751757 ( .a(n_28320), .o(n_28321) );
no02m08 g751758 ( .a(n_28306), .b(n_28305), .o(n_28320) );
na02m08 g751761 ( .a(n_28343), .b(n_28342), .o(n_28402) );
in01s01 g751762 ( .a(n_28353), .o(n_28354) );
no02m08 g751763 ( .a(n_28343), .b(n_28342), .o(n_28353) );
in01s01 g751764 ( .a(n_28303), .o(n_28304) );
no02f08 g751765 ( .a(n_28268), .b(n_28166), .o(n_28303) );
no02s01 g751766 ( .a(n_28341), .b(n_28317), .o(n_28454) );
no02s01 g751767 ( .a(FE_OCP_RBN2040_n_28268), .b(n_28300), .o(n_28302) );
in01s01 g751768 ( .a(n_28329), .o(n_28330) );
na02s01 g751769 ( .a(n_28318), .b(n_28289), .o(n_28329) );
na02m04 g751770 ( .a(n_28930), .b(n_28841), .o(n_29246) );
na02s03 g751771 ( .a(n_28931), .b(n_28993), .o(n_28962) );
na02s01 g751772 ( .a(n_29203), .b(n_29149), .o(n_29204) );
na02s01 g751773 ( .a(n_29008), .b(n_28898), .o(n_29010) );
ao12s02 g751774 ( .a(n_44045), .b(n_28941), .c(n_28793), .o(n_29050) );
in01s01 g751775 ( .a(n_29047), .o(n_29029) );
na02s02 g751776 ( .a(n_28945), .b(n_29008), .o(n_29047) );
ao12s01 g751778 ( .a(n_28233), .b(n_28232), .c(n_28234), .o(n_29439) );
oa12s01 g751779 ( .a(n_28910), .b(n_28911), .c(n_28909), .o(n_29799) );
no02s06 TIMEBOOST_cell_1767 ( .a(n_39553), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(TIMEBOOST_net_498) );
na02f08 g751782 ( .a(n_28293), .b(n_28285), .o(n_28294) );
na02s10 g751783 ( .a(n_27917), .b(n_28254), .o(n_28309) );
na02f06 g751784 ( .a(n_28291), .b(n_28290), .o(n_28292) );
in01s01 g751785 ( .a(n_28288), .o(n_28289) );
no02f08 g751786 ( .a(n_28273), .b(delay_add_ln22_unr17_stage7_stallmux_q_8_), .o(n_28288) );
na02f08 g751788 ( .a(n_28273), .b(delay_add_ln22_unr17_stage7_stallmux_q_8_), .o(n_28318) );
no03s02 TIMEBOOST_cell_8229 ( .a(n_28799), .b(FE_OCP_RBN2490_FE_RN_1367_0), .c(FE_OCP_RBN5593_FE_RN_1367_0), .o(TIMEBOOST_net_2435) );
na02s06 TIMEBOOST_cell_8042 ( .a(FE_OCPN5122_n_44438), .b(n_31783), .o(TIMEBOOST_net_2652) );
no02s01 TIMEBOOST_cell_6779 ( .a(FE_OCP_RBN4302_n_44579), .b(FE_OCP_RBN6731_n_44579), .o(TIMEBOOST_net_2147) );
in01s01 g751792 ( .a(n_28316), .o(n_28317) );
na02m08 g751793 ( .a(n_28299), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_8_), .o(n_28316) );
no02m08 g751794 ( .a(n_28299), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_8_), .o(n_28341) );
na02s01 g751795 ( .a(n_28286), .b(n_28285), .o(n_28425) );
na02s01 g751796 ( .a(n_28253), .b(n_28284), .o(n_28406) );
no02s01 g751797 ( .a(n_28234), .b(n_28232), .o(n_28233) );
in01s02 g751798 ( .a(n_28930), .o(n_28931) );
na02m06 g751799 ( .a(n_28911), .b(n_28840), .o(n_28930) );
na02s01 g751800 ( .a(n_28911), .b(n_28909), .o(n_28910) );
no02s01 g751801 ( .a(n_29131), .b(n_29101), .o(n_29203) );
in01s01 g751802 ( .a(n_44045), .o(n_28961) );
in01s01 g751804 ( .a(n_28960), .o(n_29008) );
oa12s02 g751805 ( .a(n_28946), .b(n_28882), .c(n_28836), .o(n_28960) );
oa12s02 g751806 ( .a(n_28958), .b(n_28903), .c(n_28793), .o(n_28959) );
oa12f08 g751808 ( .a(n_28181), .b(n_28255), .c(n_28139), .o(n_28268) );
no02s01 g751809 ( .a(n_29127), .b(n_29151), .o(n_29202) );
ao12s01 g751810 ( .a(n_29131), .b(n_29077), .c(n_28919), .o(n_29823) );
ao12s01 g751811 ( .a(n_29148), .b(n_29172), .c(n_28919), .o(n_29801) );
oa12s01 g751812 ( .a(n_29126), .b(n_29123), .c(n_28897), .o(n_29804) );
in01s01 g751813 ( .a(n_29103), .o(n_29104) );
oa12s01 g751814 ( .a(n_28919), .b(n_29077), .c(n_29076), .o(n_29103) );
no04m06 TIMEBOOST_cell_7364 ( .a(FE_RN_259_0), .b(FE_OCPN1906_n_23322), .c(n_23326), .d(FE_OCP_RBN2448_n_23246), .o(FE_RN_260_0) );
oa12s01 g751817 ( .a(n_28225), .b(n_28255), .c(n_28224), .o(n_29420) );
in01s01 g751818 ( .a(n_28928), .o(n_28929) );
oa22s01 g751819 ( .a(n_28838), .b(n_179), .c(n_28839), .d(n_186), .o(n_28928) );
no04s20 TIMEBOOST_cell_6420 ( .a(n_32830), .b(n_32651), .c(n_32851), .d(n_32652), .o(n_32953) );
no02s06 g751821 ( .a(n_28230), .b(n_28229), .o(n_28231) );
no03s02 TIMEBOOST_cell_7363 ( .a(n_18051), .b(n_18052), .c(n_18003), .o(TIMEBOOST_net_2066) );
na02m10 g751823 ( .a(n_28282), .b(n_28088), .o(n_28283) );
in01m08 g751824 ( .a(n_28254), .o(n_28291) );
no02m10 g751825 ( .a(n_28230), .b(n_28014), .o(n_28254) );
na02f06 g751826 ( .a(n_28228), .b(n_28227), .o(n_28284) );
in01s01 g751827 ( .a(n_28252), .o(n_28253) );
no02m08 g751828 ( .a(n_28228), .b(n_28227), .o(n_28252) );
in01s06 g751829 ( .a(n_28271), .o(n_28251) );
na02m08 g751831 ( .a(n_28208), .b(n_26972), .o(n_28286) );
na02f06 g751832 ( .a(n_28207), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_7_), .o(n_28285) );
no02s01 g751833 ( .a(n_28264), .b(n_28371), .o(n_28369) );
na02s01 g751834 ( .a(n_28255), .b(n_28224), .o(n_28225) );
in01s01 g751835 ( .a(n_28265), .o(n_28266) );
na02s01 g751836 ( .a(n_28250), .b(n_28211), .o(n_28265) );
na02s01 g751838 ( .a(n_29150), .b(n_29070), .o(n_29151) );
na02s01 g751839 ( .a(n_29334), .b(n_29309), .o(n_29769) );
no02s01 g751840 ( .a(n_29128), .b(n_29069), .o(n_29760) );
in01s01 g751841 ( .a(n_29126), .o(n_29127) );
na02s01 g751842 ( .a(n_29123), .b(n_28897), .o(n_29126) );
na02s01 g751843 ( .a(n_29124), .b(n_29123), .o(n_29125) );
in01s01 g751844 ( .a(n_29148), .o(n_29149) );
no02s01 g751845 ( .a(n_29172), .b(n_28919), .o(n_29148) );
no02s01 g751846 ( .a(n_29077), .b(n_28919), .o(n_29131) );
ao12f08 g751847 ( .a(n_28093), .b(n_28192), .c(n_28142), .o(n_28234) );
na02m06 g751848 ( .a(n_28813), .b(n_28812), .o(n_28911) );
ao12s01 g751849 ( .a(n_29129), .b(n_28919), .c(n_29026), .o(n_29746) );
no02s04 TIMEBOOST_cell_1796 ( .a(TIMEBOOST_net_512), .b(n_10833), .o(n_10896) );
no02s02 g751851 ( .a(n_29073), .b(n_29044), .o(n_29102) );
ao12s01 g751852 ( .a(n_29100), .b(n_28919), .c(n_29068), .o(n_29757) );
oa12s01 g751853 ( .a(n_28793), .b(n_28943), .c(n_28942), .o(n_28945) );
oa12s01 g751854 ( .a(n_28919), .b(n_28921), .c(n_29026), .o(n_28990) );
oa12s01 g751855 ( .a(n_28919), .b(n_29068), .c(n_29067), .o(n_29028) );
no02m08 g751857 ( .a(n_28209), .b(n_28218), .o(n_28299) );
oa22s01 g751858 ( .a(n_28161), .b(n_28146), .c(n_28162), .d(n_28192), .o(n_29391) );
oa12f08 g751859 ( .a(n_28222), .b(n_28221), .c(n_28220), .o(n_28223) );
na02m10 g751860 ( .a(n_28191), .b(n_27971), .o(n_28230) );
na02s06 g751861 ( .a(n_28191), .b(n_28189), .o(n_28190) );
in01s01 g751862 ( .a(n_28210), .o(n_28211) );
no02m06 g751863 ( .a(n_28188), .b(delay_add_ln22_unr17_stage7_stallmux_q_6_), .o(n_28210) );
na02f06 g751864 ( .a(n_28188), .b(delay_add_ln22_unr17_stage7_stallmux_q_6_), .o(n_28250) );
in01m10 g751865 ( .a(n_28249), .o(n_28282) );
no02m10 g751866 ( .a(n_28217), .b(n_28219), .o(n_28249) );
no02s06 g751867 ( .a(n_28217), .b(n_28056), .o(n_28218) );
ao12m06 g751868 ( .a(n_28057), .b(n_28123), .c(FE_OCP_RBN5523_n_28058), .o(n_28209) );
no02m08 g751869 ( .a(n_28248), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_6_), .o(n_28371) );
in01s01 g751870 ( .a(n_28293), .o(n_28264) );
na02f06 g751871 ( .a(n_28248), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_6_), .o(n_28293) );
oa12s01 g751872 ( .a(n_28247), .b(n_28221), .c(n_28220), .o(n_28362) );
na02s01 g751873 ( .a(n_28187), .b(n_28148), .o(n_28311) );
oa22f08 g751874 ( .a(n_28066), .b(delay_xor_ln21_unr18_stage7_stallmux_q_13_), .c(n_28070), .d(FE_OCP_RBN2039_n_44722), .o(n_28381) );
na02m06 g751875 ( .a(n_28811), .b(n_179), .o(n_28813) );
na02s01 g751876 ( .a(n_28946), .b(n_28907), .o(n_28908) );
na02s01 g751877 ( .a(n_29045), .b(n_29025), .o(n_29046) );
na02s01 g751878 ( .a(n_28905), .b(n_28904), .o(n_28906) );
in01s01 g751879 ( .a(n_28926), .o(n_28927) );
no02s01 g751880 ( .a(n_28859), .b(n_29200), .o(n_28926) );
na02s01 g751881 ( .a(n_29006), .b(n_28956), .o(n_29007) );
na02s01 g751882 ( .a(n_29003), .b(n_29043), .o(n_29044) );
in01s01 g751883 ( .a(n_29073), .o(n_29074) );
na02s01 g751884 ( .a(n_29001), .b(n_29285), .o(n_29073) );
no02s01 g751885 ( .a(n_29308), .b(n_29071), .o(n_29072) );
na02s01 g751886 ( .a(n_29332), .b(n_29042), .o(n_29333) );
na02s01 g751888 ( .a(n_29045), .b(n_28940), .o(n_29650) );
na02s01 g751889 ( .a(n_29201), .b(n_29105), .o(n_29251) );
na02s01 g751890 ( .a(n_28841), .b(n_28840), .o(n_28909) );
in01s01 g751891 ( .a(n_28838), .o(n_28839) );
na02s01 g751892 ( .a(n_28812), .b(n_28811), .o(n_28838) );
na02s01 g751893 ( .a(n_29043), .b(n_29042), .o(n_29653) );
in01s01 g751894 ( .a(n_29101), .o(n_29334) );
no02s01 g751895 ( .a(n_29076), .b(n_28919), .o(n_29101) );
na02s01 g751896 ( .a(n_29040), .b(n_29049), .o(n_29723) );
in01s01 g751897 ( .a(n_29070), .o(n_29128) );
na02s01 g751898 ( .a(n_28897), .b(n_29041), .o(n_29070) );
na02s01 g751899 ( .a(n_28991), .b(n_28907), .o(n_29456) );
no02s01 g751900 ( .a(n_28986), .b(n_28943), .o(n_29431) );
no02s01 g751901 ( .a(n_29004), .b(n_28957), .o(n_29510) );
na02s01 g751902 ( .a(n_29285), .b(n_29242), .o(n_29581) );
no02s02 g751903 ( .a(n_28864), .b(n_28984), .o(n_28883) );
na02s01 g751904 ( .a(n_28940), .b(n_28939), .o(n_28941) );
in01s01 g751905 ( .a(n_29069), .o(n_29124) );
no02s01 g751906 ( .a(n_29041), .b(n_28897), .o(n_29069) );
in01s01 g751907 ( .a(n_29100), .o(n_29150) );
no02s01 g751908 ( .a(n_28919), .b(n_29068), .o(n_29100) );
no02s01 g751909 ( .a(n_28919), .b(n_29026), .o(n_29129) );
no02s02 g751910 ( .a(n_28863), .b(n_28901), .o(n_28882) );
na02s01 g751911 ( .a(n_28988), .b(n_28987), .o(n_28989) );
na02s01 g751912 ( .a(n_28881), .b(n_28904), .o(n_29225) );
no02s01 g751913 ( .a(n_28902), .b(n_28923), .o(n_28903) );
in01s01 g751914 ( .a(n_29309), .o(n_29310) );
na02s01 g751915 ( .a(n_28919), .b(n_29076), .o(n_29309) );
na02s01 g751916 ( .a(n_29099), .b(n_29305), .o(n_29711) );
no02s01 g751917 ( .a(n_29170), .b(n_29200), .o(n_29336) );
oa12f08 g751918 ( .a(n_28160), .b(n_28186), .c(n_28112), .o(n_28255) );
ao12s01 g751919 ( .a(n_29308), .b(n_28919), .c(n_28689), .o(n_29741) );
ao12s01 g751920 ( .a(n_29000), .b(n_28919), .c(n_28982), .o(n_29637) );
ao12s01 g751921 ( .a(n_29002), .b(n_28919), .c(n_28984), .o(n_29692) );
ao12s01 g751922 ( .a(n_29024), .b(n_28919), .c(n_28557), .o(n_29536) );
ao12s01 g751923 ( .a(n_28955), .b(n_28919), .c(n_28942), .o(n_29459) );
oa12s01 g751924 ( .a(n_28905), .b(n_28919), .c(n_28862), .o(n_29254) );
ao12s01 g751925 ( .a(n_29223), .b(n_28897), .c(n_28923), .o(n_29286) );
oa12s01 g751926 ( .a(n_28858), .b(n_28897), .c(n_28834), .o(n_29409) );
ao12s01 g751927 ( .a(n_28924), .b(n_28919), .c(n_28901), .o(n_29462) );
no02s02 TIMEBOOST_cell_3987 ( .a(n_24344), .b(n_24230), .o(TIMEBOOST_net_1084) );
in01s04 g751929 ( .a(n_28207), .o(n_28208) );
ao22s01 g751931 ( .a(n_28186), .b(n_28180), .c(FE_OCP_RBN5374_n_28186), .d(n_28179), .o(n_29375) );
oa12s01 g751932 ( .a(n_28758), .b(n_28757), .c(n_28756), .o(n_29172) );
oa12s01 g751933 ( .a(n_28755), .b(n_28754), .c(n_28753), .o(n_29077) );
ao12s01 g751934 ( .a(n_28752), .b(n_28751), .c(n_28750), .o(n_29123) );
oa22s01 g751935 ( .a(n_28919), .b(n_28134), .c(n_28897), .d(n_28993), .o(n_29245) );
in01s40 g751936 ( .a(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_34037) );
no02s01 TIMEBOOST_cell_3986 ( .a(TIMEBOOST_net_1083), .b(n_42467), .o(n_42492) );
no02s06 g751939 ( .a(n_28149), .b(n_28040), .o(n_28150) );
no02m10 g751940 ( .a(n_28149), .b(n_28010), .o(n_28191) );
na02f08 g751941 ( .a(n_28125), .b(n_28124), .o(n_28187) );
in01s01 g751942 ( .a(n_28147), .o(n_28148) );
no02f08 g751943 ( .a(n_28125), .b(n_28124), .o(n_28147) );
na02s10 g751944 ( .a(FE_OCP_RBN5523_n_28058), .b(n_28123), .o(n_28217) );
na02s06 g751945 ( .a(n_28221), .b(n_28220), .o(n_28247) );
na02s01 g751946 ( .a(n_28222), .b(FE_OCP_RBN7019_n_28166), .o(n_28300) );
na02s01 g751947 ( .a(n_28183), .b(n_28182), .o(n_28232) );
na02s01 g751948 ( .a(n_28757), .b(n_28756), .o(n_28758) );
na02s01 g751949 ( .a(n_28754), .b(n_28753), .o(n_28755) );
no02s01 g751950 ( .a(n_28751), .b(n_28750), .o(n_28752) );
in01s01 g751951 ( .a(n_28924), .o(n_28925) );
no02s01 g751952 ( .a(n_28793), .b(n_28901), .o(n_28924) );
no02s01 g751953 ( .a(n_28836), .b(n_28923), .o(n_29223) );
in01s01 g751954 ( .a(n_28902), .o(n_28881) );
no02s01 g751955 ( .a(n_28793), .b(n_28860), .o(n_28902) );
in01s01 g751956 ( .a(n_29242), .o(n_29243) );
na02s01 g751957 ( .a(n_28919), .b(n_28669), .o(n_29242) );
in01s01 g751958 ( .a(n_29071), .o(n_29040) );
no02s01 g751959 ( .a(n_28919), .b(n_28899), .o(n_29071) );
in01s01 g751960 ( .a(n_29305), .o(n_29306) );
na02s01 g751961 ( .a(n_28919), .b(n_29067), .o(n_29305) );
in01s01 g751962 ( .a(n_29006), .o(n_28986) );
na02s01 g751963 ( .a(n_28897), .b(n_28879), .o(n_29006) );
in01s01 g751964 ( .a(n_28864), .o(n_29042) );
no02s01 g751965 ( .a(n_28836), .b(n_28837), .o(n_28864) );
in01s01 g751966 ( .a(n_28940), .o(n_28922) );
na02s01 g751967 ( .a(n_28793), .b(n_28664), .o(n_28940) );
in01s01 g751968 ( .a(n_29049), .o(n_28921) );
na02s01 g751969 ( .a(n_28793), .b(n_28899), .o(n_29049) );
in01s01 g751970 ( .a(n_29025), .o(n_29308) );
na02s01 g751971 ( .a(n_28897), .b(n_28939), .o(n_29025) );
na02s01 g751972 ( .a(n_28897), .b(n_28665), .o(n_29045) );
in01s01 g751973 ( .a(n_28943), .o(n_28898) );
no02s01 g751974 ( .a(n_28836), .b(n_28879), .o(n_28943) );
in01s01 g751975 ( .a(n_28863), .o(n_28907) );
no02s01 g751976 ( .a(n_28836), .b(n_28835), .o(n_28863) );
in01s01 g751977 ( .a(n_28988), .o(n_28957) );
na02s01 g751978 ( .a(n_28793), .b(n_28937), .o(n_28988) );
in01s01 g751979 ( .a(n_29170), .o(n_29171) );
no02s01 g751980 ( .a(n_28897), .b(n_28327), .o(n_29170) );
na02s02 g751981 ( .a(n_28749), .b(n_27957), .o(n_28812) );
na02m06 g751982 ( .a(FE_OCP_RBN2524_n_28749), .b(n_27958), .o(n_28811) );
na02s02 g751983 ( .a(FE_OCP_RBN2524_n_28749), .b(n_27994), .o(n_28840) );
na02s02 g751984 ( .a(n_28781), .b(n_27995), .o(n_28841) );
na02s01 g751985 ( .a(n_28793), .b(n_28856), .o(n_29105) );
in01s01 g751986 ( .a(n_28905), .o(n_28878) );
na02s01 g751987 ( .a(n_28793), .b(n_28862), .o(n_28905) );
na02s01 g751988 ( .a(n_28793), .b(n_28860), .o(n_28904) );
na02s01 g751989 ( .a(n_28781), .b(n_28835), .o(n_28991) );
no02s01 g751990 ( .a(n_28793), .b(n_28810), .o(n_29200) );
in01s01 g751991 ( .a(n_28858), .o(n_28859) );
na02s01 g751992 ( .a(n_28781), .b(n_28834), .o(n_28858) );
in01s01 g751993 ( .a(n_28955), .o(n_28956) );
no02s01 g751994 ( .a(n_28793), .b(n_28942), .o(n_28955) );
in01s01 g751995 ( .a(n_29004), .o(n_29488) );
no02s01 g751996 ( .a(n_28919), .b(n_28937), .o(n_29004) );
in01s01 g751997 ( .a(n_29023), .o(n_29024) );
na02s01 g751998 ( .a(n_28897), .b(n_28987), .o(n_29023) );
na02s01 g751999 ( .a(n_28897), .b(n_28837), .o(n_29043) );
in01s01 g752000 ( .a(n_29002), .o(n_29003) );
no02s01 g752001 ( .a(n_28919), .b(n_28984), .o(n_29002) );
in01s01 g752002 ( .a(n_29000), .o(n_29001) );
no02s01 g752003 ( .a(n_28919), .b(n_28982), .o(n_29000) );
na02s01 g752004 ( .a(n_28897), .b(n_28555), .o(n_29285) );
in01s01 g752005 ( .a(n_29098), .o(n_29099) );
no02s02 g752006 ( .a(n_28919), .b(n_29067), .o(n_29098) );
na02s01 g752007 ( .a(n_28897), .b(n_28203), .o(n_29201) );
in01s01 g752009 ( .a(n_28192), .o(n_28146) );
na02s01 g752011 ( .a(n_28919), .b(n_28691), .o(n_29332) );
oa12s01 g752012 ( .a(n_28793), .b(n_28396), .c(n_28810), .o(n_28946) );
in01s01 g752013 ( .a(n_28877), .o(n_28958) );
ao12s01 g752014 ( .a(n_28793), .b(n_28862), .c(n_28856), .o(n_28877) );
in01s01 g752015 ( .a(n_29187), .o(n_29267) );
oa12s02 g752016 ( .a(n_28165), .b(FE_OCP_DRV_N1880_n_28164), .c(n_28163), .o(n_29187) );
ao12s01 g752017 ( .a(n_28122), .b(n_28121), .c(n_28120), .o(n_29317) );
in01s01 g752018 ( .a(FE_OCPN1268_n_29155), .o(n_29290) );
oa12s01 g752019 ( .a(n_28100), .b(n_28099), .c(n_28098), .o(n_29155) );
oa12s01 g752020 ( .a(n_28730), .b(n_28729), .c(n_28728), .o(n_29076) );
oa12s01 g752021 ( .a(n_28694), .b(n_28693), .c(n_28692), .o(n_29026) );
oa12s01 g752022 ( .a(n_28715), .b(n_28714), .c(n_28713), .o(n_29068) );
ao12s01 g752023 ( .a(n_28712), .b(n_28711), .c(n_28710), .o(n_29041) );
na03f08 TIMEBOOST_cell_7125 ( .a(FE_RN_1246_0), .b(n_40798), .c(n_40915), .o(n_40997) );
na02s01 TIMEBOOST_cell_4881 ( .a(TIMEBOOST_net_1388), .b(FE_RN_739_0), .o(FE_RN_741_0) );
in01m08 g752026 ( .a(n_28102), .o(n_28149) );
no02m10 g752027 ( .a(n_28071), .b(n_27968), .o(n_28102) );
na02s06 g752028 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_4_), .b(n_28086), .o(n_28183) );
na03f08 TIMEBOOST_cell_4731 ( .a(n_24231), .b(FE_OFN743_delay_sub_ln23_0_unr15_stage6_stallmux_q), .c(n_24269), .o(n_24320) );
na02m04 g752032 ( .a(n_28071), .b(n_28002), .o(n_28072) );
no02s02 TIMEBOOST_cell_6152 ( .a(TIMEBOOST_net_1927), .b(n_15319), .o(TIMEBOOST_net_1541) );
no02m06 TIMEBOOST_cell_7489 ( .a(TIMEBOOST_net_2375), .b(n_12505), .o(n_12584) );
na02f08 g752039 ( .a(n_28143), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_4_), .o(n_28222) );
no02m06 g752041 ( .a(n_28143), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_4_), .o(n_28166) );
na02s01 g752042 ( .a(n_28140), .b(n_28181), .o(n_28224) );
na02s01 g752043 ( .a(n_28164), .b(n_28163), .o(n_28165) );
na02s01 g752044 ( .a(n_28099), .b(n_28098), .o(n_28100) );
in01s01 g752045 ( .a(n_28161), .o(n_28162) );
na02s01 g752046 ( .a(n_28142), .b(n_28094), .o(n_28161) );
na02s01 g752047 ( .a(n_28729), .b(n_28728), .o(n_28730) );
na02s01 g752048 ( .a(n_28693), .b(n_28692), .o(n_28694) );
na02s01 g752049 ( .a(n_28714), .b(n_28713), .o(n_28715) );
no02s01 g752050 ( .a(n_28711), .b(n_28710), .o(n_28712) );
na02m06 g752051 ( .a(n_28044), .b(n_28043), .o(n_28332) );
ao12f10 g752053 ( .a(n_28015), .b(FE_OCP_RBN2414_n_44722), .c(delay_xor_ln22_unr18_stage7_stallmux_q_11_), .o(n_28308) );
ao12m10 g752054 ( .a(n_28014), .b(FE_OCP_RBN2414_n_44722), .c(delay_xor_ln22_unr18_stage7_stallmux_q_9_), .o(n_28229) );
no04m03 g752055 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_11_), .b(delay_xor_ln21_unr18_stage7_stallmux_q_9_), .c(n_28032), .d(delay_xor_ln21_unr18_stage7_stallmux_q_10_), .o(n_28070) );
ao12f08 g752057 ( .a(n_28114), .b(n_28059), .c(n_27910), .o(n_28186) );
no02s01 g752058 ( .a(n_28120), .b(n_28121), .o(n_28122) );
in01s01 g752059 ( .a(n_28690), .o(n_28691) );
no02s02 g752060 ( .a(n_28982), .b(n_28669), .o(n_28690) );
ao12s01 g752061 ( .a(n_28263), .b(n_28709), .c(n_28214), .o(n_28757) );
in01s04 g752092 ( .a(n_28897), .o(n_28919) );
in01s03 g752100 ( .a(n_28793), .o(n_28897) );
in01s02 g752107 ( .a(n_28793), .o(n_28836) );
in01s06 g752109 ( .a(n_28781), .o(n_28793) );
in01s04 g752110 ( .a(FE_OCP_RBN2524_n_28749), .o(n_28781) );
ao12s01 g752113 ( .a(n_28157), .b(n_28636), .c(n_28174), .o(n_28751) );
ao12s01 g752114 ( .a(n_28262), .b(n_28709), .c(n_28173), .o(n_28754) );
na02m10 g752116 ( .a(n_28097), .b(n_28119), .o(n_28221) );
oa12s01 g752117 ( .a(n_28621), .b(n_28620), .c(n_28619), .o(n_28984) );
in01s01 g752118 ( .a(n_28939), .o(n_28689) );
ao12s01 g752119 ( .a(n_28618), .b(n_28617), .c(n_28616), .o(n_28939) );
oa12s01 g752120 ( .a(n_28639), .b(n_28638), .c(n_28637), .o(n_28899) );
oa12s01 g752121 ( .a(n_28668), .b(n_28667), .c(n_28666), .o(n_29067) );
no02m08 TIMEBOOST_cell_3978 ( .a(TIMEBOOST_net_1079), .b(n_9095), .o(n_9313) );
na02m10 g752123 ( .a(n_27965), .b(n_28061), .o(n_28119) );
oa12s10 g752124 ( .a(n_27964), .b(n_28096), .c(FE_OCP_RBN3982_n_27911), .o(n_28097) );
no02s01 g752125 ( .a(n_28709), .b(n_28216), .o(n_28729) );
na02s20 g752126 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_12_), .b(FE_OCP_RBN2414_n_44722), .o(n_28044) );
no02f40 g752127 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_11_), .b(FE_OCP_RBN2414_n_44722), .o(n_28015) );
no02s40 g752128 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_9_), .b(FE_OCP_RBN2415_n_44722), .o(n_28014) );
in01s02 g752129 ( .a(n_28071), .o(n_28042) );
na02m10 g752130 ( .a(n_28012), .b(n_27872), .o(n_28071) );
na02m10 g752131 ( .a(n_27922), .b(FE_OCP_RBN2039_n_44722), .o(n_28043) );
in01s01 g752132 ( .a(n_28093), .o(n_28094) );
no02f08 g752133 ( .a(n_46961), .b(delay_add_ln22_unr17_stage7_stallmux_q_3_), .o(n_28093) );
na02f08 g752134 ( .a(n_46961), .b(delay_add_ln22_unr17_stage7_stallmux_q_3_), .o(n_28142) );
in01s06 g752135 ( .a(n_28117), .o(n_28118) );
no02s02 TIMEBOOST_cell_3069 ( .a(TIMEBOOST_net_825), .b(n_8863), .o(n_8910) );
na02s08 g752137 ( .a(n_28116), .b(n_28115), .o(n_28181) );
in01s01 g752138 ( .a(n_28139), .o(n_28140) );
no02m08 g752139 ( .a(n_28116), .b(n_28115), .o(n_28139) );
in01s01 g752140 ( .a(n_28179), .o(n_28180) );
na02s01 g752141 ( .a(n_28113), .b(n_28160), .o(n_28179) );
no02s01 g752142 ( .a(n_28114), .b(n_28060), .o(n_28164) );
no02s01 g752143 ( .a(n_28067), .b(n_28068), .o(n_28121) );
na02s01 g752144 ( .a(n_28638), .b(n_28637), .o(n_28639) );
na02s01 g752145 ( .a(n_28620), .b(n_28619), .o(n_28621) );
no02s01 g752146 ( .a(n_28617), .b(n_28616), .o(n_28618) );
na02s01 g752147 ( .a(n_28635), .b(n_28202), .o(n_28711) );
no02m10 g752148 ( .a(n_28064), .b(FE_OCP_RBN2039_n_44722), .o(n_28066) );
in01s04 g752149 ( .a(n_28090), .o(n_28091) );
no02s10 g752150 ( .a(n_28064), .b(n_28065), .o(n_28090) );
na02s01 g752151 ( .a(n_28667), .b(n_28666), .o(n_28668) );
in01m06 g752152 ( .a(n_28040), .o(n_28041) );
ao12m10 g752153 ( .a(n_28010), .b(FE_OCP_RBN2037_n_44722), .c(delay_xor_ln22_unr18_stage7_stallmux_q_7_), .o(n_28040) );
in01s06 g752154 ( .a(n_28062), .o(n_28063) );
ao12s10 g752155 ( .a(n_28039), .b(FE_OCP_RBN2415_n_44722), .c(delay_xor_ln21_unr18_stage7_stallmux_q_11_), .o(n_28062) );
in01m03 g752156 ( .a(n_28088), .o(n_28089) );
ao12s06 g752157 ( .a(n_28226), .b(FE_OCP_RBN2415_n_44722), .c(delay_xor_ln21_unr18_stage7_stallmux_q_9_), .o(n_28088) );
na02m08 TIMEBOOST_cell_7411 ( .a(n_1551), .b(TIMEBOOST_net_2336), .o(n_1635) );
ao12s01 g752161 ( .a(n_27973), .b(n_28009), .c(delay_add_ln22_unr17_stage7_stallmux_q_1_), .o(n_28099) );
oa12s01 g752162 ( .a(n_28560), .b(n_28559), .c(n_28558), .o(n_28982) );
ao12s01 g752163 ( .a(n_28587), .b(n_28586), .c(n_28585), .o(n_28837) );
in01s01 g752164 ( .a(n_28664), .o(n_28665) );
oa12s01 g752165 ( .a(n_28590), .b(n_28589), .c(n_28588), .o(n_28664) );
no02s02 TIMEBOOST_cell_1763 ( .a(FE_OCP_RBN4352_FE_OCPN1263_n_20971), .b(FE_OCP_RBN5962_n_20459), .o(TIMEBOOST_net_496) );
no02s01 TIMEBOOST_cell_4875 ( .a(TIMEBOOST_net_1385), .b(n_1377), .o(n_1669) );
ao12f08 g752169 ( .a(n_28038), .b(n_28037), .c(n_28036), .o(n_28143) );
in01s20 g752170 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_12_), .o(n_27922) );
no02s02 TIMEBOOST_cell_1837 ( .a(FE_RN_2880_0), .b(n_47273), .o(TIMEBOOST_net_533) );
na02s01 g752175 ( .a(n_28592), .b(n_28054), .o(n_28638) );
no02s01 g752176 ( .a(n_44826), .b(n_28106), .o(n_28591) );
no02m40 g752177 ( .a(FE_OCP_RBN2037_n_44722), .b(delay_xor_ln22_unr18_stage7_stallmux_q_7_), .o(n_28010) );
na02s06 g752179 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_13_), .b(FE_OCP_RBN2414_n_44722), .o(n_28360) );
na02s02 g752180 ( .a(n_27921), .b(FE_OCP_RBN2039_n_44722), .o(n_27976) );
na02f10 g752181 ( .a(FE_OCP_RBN5531_n_27941), .b(n_27895), .o(n_28008) );
no02f06 TIMEBOOST_cell_4920 ( .a(n_21785), .b(n_23175), .o(TIMEBOOST_net_1408) );
no02f10 g752183 ( .a(n_27940), .b(n_26566), .o(n_28068) );
no02f08 g752184 ( .a(n_27939), .b(delay_add_ln22_unr17_stage7_stallmux_q_2_), .o(n_28067) );
no02m20 g752185 ( .a(n_27944), .b(FE_OCP_RBN2039_n_44722), .o(n_28064) );
no02s40 g752186 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_11_), .b(FE_OCP_RBN2415_n_44722), .o(n_28039) );
no02m10 g752187 ( .a(n_28096), .b(FE_OCPN1400_n_28095), .o(n_28061) );
no02f06 g752188 ( .a(FE_OCP_RBN2416_n_44722), .b(delay_xor_ln21_unr18_stage7_stallmux_q_9_), .o(n_28226) );
no02s20 g752189 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_12_), .b(FE_OCP_RBN2415_n_44722), .o(n_28065) );
no02m08 g752190 ( .a(n_28037), .b(n_28036), .o(n_28038) );
na02f08 g752191 ( .a(n_28085), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_2_), .o(n_28160) );
in01s01 g752192 ( .a(n_28112), .o(n_28113) );
no02f08 g752193 ( .a(n_28085), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_2_), .o(n_28112) );
in01s01 g752194 ( .a(n_28059), .o(n_28060) );
na02f08 g752195 ( .a(n_28034), .b(n_28035), .o(n_28059) );
no02f08 g752196 ( .a(n_28035), .b(n_28034), .o(n_28114) );
no02s01 g752197 ( .a(n_28009), .b(delay_add_ln22_unr17_stage7_stallmux_q_1_), .o(n_27973) );
no02s01 g752198 ( .a(n_44825), .b(n_28615), .o(n_28667) );
na02s01 g752199 ( .a(n_28559), .b(n_28558), .o(n_28560) );
na02s01 g752200 ( .a(n_28589), .b(n_28588), .o(n_28590) );
in01s01 g752201 ( .a(n_28635), .o(n_28636) );
na02s01 g752202 ( .a(n_44825), .b(n_28130), .o(n_28635) );
na02m10 g752203 ( .a(n_27971), .b(n_27972), .o(n_28189) );
no02s01 g752204 ( .a(n_28586), .b(n_28585), .o(n_28587) );
ao12m10 g752205 ( .a(n_27916), .b(FE_OCP_RBN2414_n_44722), .c(delay_xor_ln22_unr18_stage7_stallmux_q_10_), .o(n_28290) );
oa22f10 g752206 ( .a(n_27871), .b(FE_OCP_RBN7127_n_44722), .c(n_44723), .d(delay_xor_ln22_unr18_stage7_stallmux_q_5_), .o(n_28011) );
in01f08 g752208 ( .a(n_28083), .o(n_28084) );
no02s04 TIMEBOOST_cell_3935 ( .a(n_29271), .b(n_29379), .o(TIMEBOOST_net_1058) );
in01s01 g752210 ( .a(n_28634), .o(n_28709) );
na02m06 g752211 ( .a(n_44827), .b(n_28201), .o(n_28634) );
ao12s01 g752212 ( .a(n_28027), .b(n_28539), .c(n_27950), .o(n_28617) );
ao12s01 g752215 ( .a(n_28238), .b(n_28538), .c(n_28154), .o(n_28620) );
in01s01 g752216 ( .a(n_28987), .o(n_28557) );
ao22s01 g752217 ( .a(n_28479), .b(n_28315), .c(n_28480), .d(n_28314), .o(n_28987) );
in01s01 g752218 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_13_), .o(n_27921) );
in01m20 g752223 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_12_), .o(n_27944) );
na02f10 g752226 ( .a(n_27839), .b(n_27919), .o(n_27920) );
na02s01 g752227 ( .a(n_28539), .b(n_28079), .o(n_28592) );
no02s01 g752228 ( .a(n_28539), .b(n_44046), .o(n_28589) );
na02s20 g752229 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_8_), .b(FE_OCP_RBN2415_n_44722), .o(n_27972) );
no02f20 g752231 ( .a(n_27919), .b(n_27918), .o(n_27941) );
na02m10 g752232 ( .a(n_27871), .b(FE_OCP_RBN7127_n_44722), .o(n_27872) );
na02m40 g752233 ( .a(n_27869), .b(FE_OCP_RBN2039_n_44722), .o(n_27971) );
in01s06 g752234 ( .a(n_27916), .o(n_27917) );
no02s40 g752235 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_10_), .b(FE_OCP_RBN2414_n_44722), .o(n_27916) );
no02m40 g752237 ( .a(n_44723), .b(delay_xor_ln21_unr18_stage7_stallmux_q_7_), .o(n_28058) );
in01s20 g752238 ( .a(n_28037), .o(n_28096) );
in01s03 g752240 ( .a(n_28005), .o(n_28006) );
na02s40 g752241 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_13_), .b(FE_OCP_RBN2414_n_44722), .o(n_28005) );
na02s01 TIMEBOOST_cell_8778 ( .a(n_11154), .b(n_10239), .o(TIMEBOOST_net_2876) );
no02s01 g752243 ( .a(n_28538), .b(n_28195), .o(n_28586) );
in01m08 g752244 ( .a(n_28056), .o(n_28057) );
no02s20 g752245 ( .a(n_28032), .b(n_28219), .o(n_28056) );
in01s06 g752246 ( .a(n_28002), .o(n_28003) );
in01s06 g752248 ( .a(n_28030), .o(n_28031) );
ao12m06 g752249 ( .a(n_28001), .b(FE_OCP_RBN2415_n_44722), .c(delay_xor_ln21_unr18_stage7_stallmux_q_10_), .o(n_28030) );
oa12s01 g752250 ( .a(n_28212), .b(FE_OCP_RBN2481_FE_RN_734_0), .c(n_28259), .o(n_28559) );
na02m06 g752252 ( .a(n_28539), .b(n_28177), .o(n_28556) );
in01s01 g752258 ( .a(n_28669), .o(n_28555) );
oa12s01 g752259 ( .a(n_28499), .b(FE_OCP_RBN2481_FE_RN_734_0), .c(n_28498), .o(n_28669) );
in01f08 g752260 ( .a(n_27939), .o(n_27940) );
in01m40 g752264 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_8_), .o(n_27869) );
in01m40 g752266 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_5_), .o(n_27871) );
in01s20 g752269 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_7_), .o(n_27938) );
in01s01 g752271 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_27_), .o(n_27807) );
in01s01 g752273 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_29_), .o(n_28795) );
in01s01 g752275 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_30_), .o(n_27806) );
no02m40 g752279 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_6_), .b(FE_OCP_RBN2038_n_44722), .o(n_27968) );
in01m01 g752283 ( .a(n_28001), .o(n_28270) );
no02s40 g752284 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_10_), .b(FE_OCP_RBN2416_n_44722), .o(n_28001) );
no02s20 g752286 ( .a(n_27970), .b(n_27937), .o(n_27966) );
no02s40 g752287 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_8_), .b(FE_OCP_RBN2416_n_44722), .o(n_28219) );
no02s01 g752288 ( .a(FE_OCP_RBN2480_FE_RN_734_0), .b(n_28109), .o(n_28538) );
na02s01 g752289 ( .a(FE_OCP_RBN2481_FE_RN_734_0), .b(n_28498), .o(n_28499) );
in01f10 g752290 ( .a(n_27895), .o(n_27896) );
ao12f20 g752291 ( .a(n_27864), .b(n_44723), .c(delay_xor_ln22_unr18_stage7_stallmux_q_4_), .o(n_27895) );
in01f08 g752294 ( .a(n_28028), .o(n_28029) );
in01s06 g752297 ( .a(n_27964), .o(n_27965) );
no02s06 TIMEBOOST_cell_8855 ( .a(TIMEBOOST_net_2914), .b(n_16407), .o(n_16499) );
no02m20 g752300 ( .a(n_27889), .b(n_27936), .o(n_27962) );
in01s01 g752302 ( .a(n_28479), .o(n_28480) );
ao12s01 g752303 ( .a(n_28050), .b(n_28457), .c(n_27949), .o(n_28479) );
in01s01 g752309 ( .a(FE_OCP_DRV_N3502_n_29140), .o(n_27961) );
oa12s01 g752310 ( .a(n_27887), .b(n_27888), .c(delay_sub_ln21_0_unr17_stage7_stallmux_q_0_), .o(n_29140) );
in01s01 g752311 ( .a(n_29109), .o(n_27914) );
ao12s01 g752312 ( .a(n_27830), .b(FE_OCP_RBN6369_n_27773), .c(delay_add_ln22_unr17_stage7_stallmux_q_0_), .o(n_29109) );
oa12s01 g752313 ( .a(n_28436), .b(n_28435), .c(n_28434), .o(n_28942) );
oa12s01 g752314 ( .a(n_28446), .b(n_28457), .c(n_28445), .o(n_28937) );
in01s01 g752315 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_27_), .o(n_27860) );
in01s01 g752317 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_29_), .o(n_27834) );
in01s01 g752319 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_30_), .o(n_27833) );
in01s01 g752325 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_25_), .o(n_28646) );
in01s01 g752327 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_31_), .o(n_27803) );
in01f08 g752329 ( .a(n_27831), .o(n_27832) );
na02f40 g752330 ( .a(n_27868), .b(n_27802), .o(n_27831) );
in01s10 g752331 ( .a(n_27970), .o(n_27912) );
na02s80 g752332 ( .a(n_27893), .b(n_27885), .o(n_27970) );
no02f80 g752333 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_4_), .b(n_44723), .o(n_27864) );
no02f80 g752334 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_3_), .b(n_44761), .o(n_27918) );
na02f10 g752335 ( .a(n_27773), .b(delay_add_ln22_unr17_stage7_stallmux_q_0_), .o(n_28098) );
no02m40 g752336 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_6_), .b(n_44723), .o(n_27999) );
na02m40 g752338 ( .a(n_45200), .b(FE_OCP_RBN7128_n_44722), .o(n_27911) );
no02s80 g752339 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_3_), .b(n_44761), .o(n_27936) );
no02s40 g752340 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_5_), .b(n_44723), .o(n_28092) );
no02s01 TIMEBOOST_cell_5096 ( .a(n_29365), .b(n_29135), .o(TIMEBOOST_net_1496) );
no02s20 g752342 ( .a(n_27823), .b(FE_OCP_RBN7128_n_44722), .o(n_27889) );
in01s01 g752343 ( .a(n_27910), .o(n_28163) );
na02s01 g752345 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_0_), .b(n_27888), .o(n_27887) );
no02s01 g752346 ( .a(FE_OCP_RBN6369_n_27773), .b(delay_add_ln22_unr17_stage7_stallmux_q_0_), .o(n_27830) );
na02s01 g752347 ( .a(n_28435), .b(n_28434), .o(n_28436) );
na02s01 g752348 ( .a(n_28457), .b(n_28445), .o(n_28446) );
na02s10 g752352 ( .a(n_27802), .b(n_27738), .o(n_27825) );
no02f08 TIMEBOOST_cell_5115 ( .a(TIMEBOOST_net_1505), .b(n_29730), .o(n_29808) );
in01s01 g752363 ( .a(n_27785), .o(n_27758) );
in01s01 g752365 ( .a(n_27784), .o(n_27757) );
in01s01 g752367 ( .a(n_27783), .o(n_27756) );
oa22s01 g752369 ( .a(n_28397), .b(n_28277), .c(n_28398), .d(n_28276), .o(n_28901) );
in01s01 g752370 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_25_), .o(n_28630) );
in01s01 g752372 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_31_), .o(n_27824) );
in01s20 g752379 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_3_), .o(n_27823) );
in01s20 g752381 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_5_), .o(n_27822) );
in01s01 g752383 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_23_), .o(n_28606) );
in01s01 g752386 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_28_), .o(n_27778) );
na03s08 TIMEBOOST_cell_5704 ( .a(n_17480), .b(n_17395), .c(n_17442), .o(n_17620) );
na02s80 g752389 ( .a(n_27732), .b(FE_OCP_RBN7127_n_44722), .o(n_27802) );
in01s20 g752391 ( .a(n_27884), .o(n_27937) );
na02m40 g752392 ( .a(n_27794), .b(FE_OCP_RBN7128_n_44722), .o(n_27884) );
na02f80 g752393 ( .a(n_44420), .b(FE_OCP_RBN7128_n_44722), .o(n_27885) );
na02m04 TIMEBOOST_cell_3890 ( .a(TIMEBOOST_net_1035), .b(n_41191), .o(n_41256) );
no02s01 g752396 ( .a(n_28399), .b(FE_RN_728_0), .o(n_28457) );
oa12s01 g752397 ( .a(n_28256), .b(n_28401), .c(n_28297), .o(n_28435) );
in01m02 g752401 ( .a(n_27835), .o(n_27795) );
ao22f10 g752408 ( .a(n_44759), .b(n_27719), .c(FE_OCP_RBN7127_n_44722), .d(delay_xor_ln22_unr18_stage7_stallmux_q_0_), .o(n_27773) );
in01s01 g752413 ( .a(n_27781), .o(n_27752) );
ao12s01 g752415 ( .a(n_28380), .b(n_28401), .c(n_28379), .o(n_28879) );
in01f40 g752418 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_2_), .o(n_27776) );
in01s80 g752420 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_1_), .o(n_27732) );
in01m40 g752422 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_2_), .o(n_27794) );
in01f08 g752428 ( .a(n_27868), .o(n_27751) );
na02f80 g752429 ( .a(n_27719), .b(FE_OCP_RBN7127_n_44722), .o(n_27868) );
na02f80 g752431 ( .a(n_44696), .b(FE_OCP_RBN7128_n_44722), .o(n_27893) );
no02s01 g752434 ( .a(n_28401), .b(n_28379), .o(n_28380) );
in01s01 g752435 ( .a(n_28397), .o(n_28398) );
oa12s01 g752436 ( .a(n_27848), .b(n_28378), .c(n_27903), .o(n_28397) );
in01s02 g752443 ( .a(n_27800), .o(n_27767) );
in01s01 g752445 ( .a(n_27799), .o(n_27766) );
in01s02 g752447 ( .a(n_27720), .o(n_27698) );
in01s01 g752449 ( .a(n_27739), .o(n_27730) );
oa22s02 g752450 ( .a(n_27639), .b(n_27423), .c(FE_OCP_RBN4495_n_27639), .d(n_27424), .o(n_27739) );
oa12s02 g752451 ( .a(n_27395), .b(n_27639), .c(n_27254), .o(n_27675) );
ao12s02 g752452 ( .a(n_27294), .b(FE_OCP_RBN4496_n_27639), .c(FE_OCPN1396_n_27211), .o(n_27697) );
in01s01 g752453 ( .a(n_27729), .o(n_27755) );
oa12s01 g752455 ( .a(n_27461), .b(n_27672), .c(n_27336), .o(n_27674) );
ao12s02 g752456 ( .a(n_27411), .b(n_27648), .c(n_27337), .o(n_27696) );
oa12s02 g752457 ( .a(n_27469), .b(n_27648), .c(n_27371), .o(n_27695) );
ao12s01 g752458 ( .a(n_27507), .b(n_27672), .c(n_27326), .o(n_27673) );
ao12s01 g752459 ( .a(n_28352), .b(n_28378), .c(n_28351), .o(n_28835) );
in01s01 g752460 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_21_), .o(n_28523) );
in01f80 g752465 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_0_), .o(n_27719) );
in01s01 g752471 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_21_), .o(n_28541) );
no02s01 g752474 ( .a(n_28378), .b(n_28351), .o(n_28352) );
ao12m04 g752475 ( .a(n_28052), .b(n_28328), .c(n_27905), .o(n_28401) );
oa22f02 g752478 ( .a(n_27643), .b(n_24350), .c(n_27619), .d(n_27845), .o(n_27671) );
in01s02 g752479 ( .a(n_27772), .o(n_27745) );
ao12m06 g752482 ( .a(n_27223), .b(n_27661), .c(n_27144), .o(n_27723) );
in01s01 g752483 ( .a(n_27771), .o(n_27744) );
no02s02 TIMEBOOST_cell_1520 ( .a(TIMEBOOST_net_374), .b(n_30116), .o(n_30175) );
oa12s01 g752485 ( .a(n_27418), .b(n_27691), .c(FE_OCPN5134_n_27667), .o(n_27692) );
no02s02 g752486 ( .a(n_27668), .b(n_27384), .o(n_27717) );
oa12m01 g752488 ( .a(n_27302), .b(n_27691), .c(n_27401), .o(n_27715) );
in01s02 g752489 ( .a(n_27736), .o(n_27768) );
ao22s04 g752490 ( .a(n_44265), .b(n_27503), .c(n_27620), .d(n_27502), .o(n_27736) );
oa12s04 g752491 ( .a(n_27463), .b(n_44265), .c(n_27415), .o(n_27670) );
no02m08 TIMEBOOST_cell_1542 ( .a(n_14478), .b(TIMEBOOST_net_385), .o(n_14515) );
oa22m02 g752495 ( .a(n_27653), .b(n_24350), .c(n_27635), .d(n_27796), .o(n_27687) );
in01s01 g752496 ( .a(n_28834), .o(n_28396) );
ao12s01 g752497 ( .a(n_28340), .b(n_28339), .c(n_28338), .o(n_28834) );
in01s01 g752500 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_19_), .o(n_27654) );
in01s01 g752502 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_20_), .o(n_27669) );
na02s01 g752505 ( .a(n_27712), .b(n_27710), .o(n_27711) );
na02s01 g752506 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_), .o(n_27642) );
no02s01 g752507 ( .a(n_28328), .b(n_27955), .o(n_28378) );
no02s01 g752508 ( .a(n_28339), .b(n_28338), .o(n_28340) );
na02s02 g752509 ( .a(n_27691), .b(n_27466), .o(n_27709) );
no02s01 TIMEBOOST_cell_1519 ( .a(n_29167), .b(n_29922), .o(TIMEBOOST_net_374) );
no02s01 g752511 ( .a(n_27691), .b(FE_OCPN5134_n_27667), .o(n_27668) );
oa22f02 g752512 ( .a(n_27665), .b(n_24350), .c(n_27644), .d(n_27796), .o(n_27708) );
oa22s02 g752513 ( .a(n_27622), .b(n_24350), .c(n_27607), .d(n_27845), .o(n_27652) );
in01f02 g752514 ( .a(n_27728), .o(n_27706) );
in01m02 g752516 ( .a(n_27727), .o(n_27705) );
oa12s06 g752522 ( .a(n_27426), .b(n_27645), .c(n_27343), .o(n_27684) );
ao12s04 g752523 ( .a(n_27388), .b(n_27634), .c(n_27425), .o(n_27703) );
in01s02 g752524 ( .a(n_27701), .o(n_27702) );
na02s04 g752525 ( .a(n_27646), .b(n_27531), .o(n_27701) );
in01m02 g752526 ( .a(n_27655), .o(n_27641) );
in01s02 g752528 ( .a(n_27693), .o(n_27666) );
na02s01 TIMEBOOST_cell_2884 ( .a(n_18090), .b(n_17944), .o(TIMEBOOST_net_733) );
oa12s02 g752530 ( .a(n_27256), .b(n_27602), .c(n_27601), .o(n_27610) );
no02s03 g752531 ( .a(n_27603), .b(n_27295), .o(n_27624) );
na02s06 g752535 ( .a(n_27600), .b(n_27551), .o(n_27639) );
in01s06 g752536 ( .a(n_27672), .o(n_27648) );
in01s02 g752537 ( .a(n_27648), .o(n_27649) );
na02s06 g752539 ( .a(n_27599), .b(n_27550), .o(n_27672) );
no02m04 TIMEBOOST_cell_1541 ( .a(n_14321), .b(n_13514), .o(TIMEBOOST_net_385) );
in01s01 g752541 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_17_), .o(n_27712) );
in01s01 g752544 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_), .o(n_27623) );
in01s01 g752546 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_18_), .o(n_27637) );
no02f02 TIMEBOOST_cell_8740 ( .a(FE_OCPN5128_n_22280), .b(n_24891), .o(TIMEBOOST_net_2857) );
na02s02 g752550 ( .a(n_27602), .b(n_27397), .o(n_27621) );
na02f06 TIMEBOOST_cell_2883 ( .a(TIMEBOOST_net_732), .b(n_18433), .o(n_18645) );
no02s03 g752552 ( .a(n_27602), .b(n_27601), .o(n_27603) );
na02s02 g752558 ( .a(n_27598), .b(n_27297), .o(n_27600) );
na02s02 g752559 ( .a(n_27598), .b(n_27427), .o(n_27599) );
in01f02 g752560 ( .a(n_27686), .o(n_27662) );
in01f02 g752562 ( .a(n_27714), .o(n_27683) );
in01s02 g752564 ( .a(n_27681), .o(n_27682) );
in01s03 g752565 ( .a(n_27661), .o(n_27681) );
no02f04 TIMEBOOST_cell_1514 ( .a(TIMEBOOST_net_371), .b(n_25239), .o(n_25401) );
in01s01 g752568 ( .a(n_27691), .o(n_27659) );
na02s06 g752569 ( .a(n_27608), .b(n_27471), .o(n_27691) );
na02s02 g752570 ( .a(n_27634), .b(n_27429), .o(n_27646) );
in01f02 g752571 ( .a(n_27643), .o(n_27619) );
oa22f02 g752572 ( .a(n_27569), .b(n_27457), .c(n_27570), .d(n_27458), .o(n_27643) );
in01s02 g752573 ( .a(n_27653), .o(n_27635) );
no02s01 TIMEBOOST_cell_1496 ( .a(TIMEBOOST_net_362), .b(FE_OCP_RBN2769_n_3238), .o(n_3324) );
in01s01 g752575 ( .a(n_28810), .o(n_28327) );
oa12s01 g752576 ( .a(n_28279), .b(n_28298), .c(n_28278), .o(n_28810) );
no03s03 TIMEBOOST_cell_7145 ( .a(n_41654), .b(FE_OCP_RBN6589_n_41491), .c(n_41688), .o(n_41742) );
na02s01 g752578 ( .a(n_28298), .b(n_28278), .o(n_28279) );
in01s06 g752582 ( .a(n_27634), .o(n_27645) );
na02s10 g752583 ( .a(FE_OCP_RBN1176_n_27593), .b(n_27433), .o(n_27634) );
no02s01 TIMEBOOST_cell_1513 ( .a(n_24217), .b(n_25181), .o(TIMEBOOST_net_371) );
na02s06 g752585 ( .a(n_27593), .b(n_27353), .o(n_27608) );
na02m04 g752586 ( .a(n_27571), .b(FE_OCP_RBN6233_n_27504), .o(n_27585) );
no02s01 TIMEBOOST_cell_1495 ( .a(n_3286), .b(n_2437), .o(TIMEBOOST_net_362) );
in01s01 g752589 ( .a(n_27602), .o(n_27595) );
na02s06 g752590 ( .a(n_27573), .b(n_27512), .o(n_27602) );
oa22s01 g752591 ( .a(n_27578), .b(n_27544), .c(n_27579), .d(n_27545), .o(n_27617) );
in01f02 g752592 ( .a(n_27665), .o(n_27644) );
oa22m04 g752593 ( .a(FE_OCP_RBN3418_n_27590), .b(n_27270), .c(n_27590), .d(n_27271), .o(n_27665) );
oa22s01 g752600 ( .a(n_27555), .b(n_27542), .c(FE_OCP_RBN4494_n_27555), .d(n_27543), .o(n_27584) );
in01s02 g752601 ( .a(n_27622), .o(n_27607) );
oa22s02 g752602 ( .a(n_27565), .b(n_27348), .c(n_27566), .d(n_27349), .o(n_27622) );
oa12m04 g752604 ( .a(n_27511), .b(n_27567), .c(n_27213), .o(n_27582) );
no02s06 g752606 ( .a(n_27573), .b(n_27300), .o(n_27598) );
ao12s01 g752607 ( .a(n_28246), .b(n_28245), .c(n_28244), .o(n_28860) );
oa22s01 g752608 ( .a(n_28239), .b(n_28024), .c(n_28240), .d(n_28023), .o(n_28923) );
in01s01 g752609 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_16_), .o(n_27710) );
no02s01 g752612 ( .a(n_28245), .b(n_28244), .o(n_28246) );
in01f04 g752613 ( .a(n_27614), .o(n_27615) );
na02f08 g752614 ( .a(n_27568), .b(n_27403), .o(n_27614) );
in01s02 g752615 ( .a(n_27571), .o(n_27572) );
na02s06 g752616 ( .a(n_27567), .b(n_27430), .o(n_27571) );
no03m02 TIMEBOOST_cell_3589 ( .a(n_9582), .b(n_9461), .c(FE_OCP_RBN5919_n_9456), .o(n_9675) );
in01f02 g752618 ( .a(n_27604), .o(n_27605) );
ao12f04 g752619 ( .a(n_27269), .b(n_27554), .c(n_27233), .o(n_27604) );
in01f02 g752623 ( .a(n_27569), .o(n_27570) );
oa12f02 g752624 ( .a(n_27301), .b(n_27476), .c(n_27219), .o(n_27569) );
na02s08 g752625 ( .a(n_27535), .b(n_27264), .o(n_27573) );
ao12s01 g752626 ( .a(n_28243), .b(n_28242), .c(n_28241), .o(n_28862) );
in01s01 g752627 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_15_), .o(n_28473) );
in01s01 g752629 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_15_), .o(n_28466) );
no02s01 g752631 ( .a(n_28242), .b(n_28241), .o(n_28243) );
in01s01 TIMEBOOST_cell_8904 ( .a(n_1304), .o(TIMEBOOST_net_2948) );
no02m04 g752634 ( .a(n_27554), .b(n_27168), .o(n_27590) );
in01s01 g752635 ( .a(n_27565), .o(n_27566) );
na02s02 g752636 ( .a(n_27476), .b(n_27206), .o(n_27565) );
in01s01 g752637 ( .a(n_28239), .o(n_28240) );
no02s02 TIMEBOOST_cell_1630 ( .a(TIMEBOOST_net_429), .b(n_3846), .o(n_3853) );
oa12s01 g752639 ( .a(n_28204), .b(n_28158), .c(n_27990), .o(n_28245) );
oa22s01 g752640 ( .a(n_27533), .b(n_27529), .c(n_27532), .d(n_27528), .o(n_27580) );
in01s01 g752641 ( .a(n_27578), .o(n_27579) );
oa12s01 g752642 ( .a(n_27506), .b(n_27533), .c(n_27422), .o(n_27578) );
oa22s01 g752647 ( .a(n_27473), .b(n_27546), .c(n_27442), .d(n_27547), .o(n_27576) );
oa12s01 g752649 ( .a(n_27527), .b(n_27442), .c(n_27454), .o(n_27555) );
in01s04 g752650 ( .a(n_27535), .o(n_27567) );
no02s01 g752652 ( .a(n_28159), .b(n_27987), .o(n_28242) );
oa22s01 g752662 ( .a(n_27441), .b(n_27191), .c(n_27440), .d(n_27190), .o(n_27534) );
oa22s01 g752663 ( .a(n_27314), .b(n_27225), .c(n_27313), .d(n_27224), .o(n_27443) );
in01s01 g752664 ( .a(n_28856), .o(n_28203) );
ao12s01 g752665 ( .a(n_28137), .b(n_28136), .c(n_28135), .o(n_28856) );
in01s01 g752667 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_13_), .o(n_28452) );
na02s01 g752671 ( .a(n_28261), .b(FE_RN_739_0), .o(n_28263) );
na02s01 g752672 ( .a(n_28261), .b(n_28132), .o(n_28262) );
in01s01 g752674 ( .a(n_28158), .o(n_28159) );
in01s01 g752675 ( .a(n_28138), .o(n_28158) );
no02s04 g752676 ( .a(n_28082), .b(n_27876), .o(n_28138) );
no02s01 g752677 ( .a(n_28136), .b(n_28135), .o(n_28137) );
in01s01 g752680 ( .a(n_27532), .o(n_27533) );
in01s01 g752681 ( .a(n_27514), .o(n_27532) );
oa12f08 g752682 ( .a(n_27157), .b(n_27363), .c(n_27127), .o(n_27514) );
in01s01 g752684 ( .a(n_27442), .o(n_27473) );
in01s01 g752685 ( .a(n_27404), .o(n_27442) );
ao12f08 g752686 ( .a(n_27183), .b(n_27245), .c(n_27153), .o(n_27404) );
in01s01 g752687 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_13_), .o(n_28449) );
na02s01 g752689 ( .a(n_28202), .b(n_28156), .o(n_28157) );
in01s04 g752690 ( .a(n_28216), .o(n_28261) );
oa12s04 g752691 ( .a(n_28202), .b(n_28129), .c(n_27923), .o(n_28216) );
in01s01 g752692 ( .a(n_28082), .o(n_28136) );
no02s04 g752693 ( .a(n_27998), .b(n_27933), .o(n_28082) );
oa22s01 g752694 ( .a(n_27358), .b(n_27101), .c(n_27359), .d(n_27102), .o(n_27472) );
in01s01 g752695 ( .a(n_27440), .o(n_27441) );
ao12s01 g752696 ( .a(n_27361), .b(n_27362), .c(n_27125), .o(n_27440) );
oa22s01 g752697 ( .a(n_27240), .b(n_27071), .c(n_27239), .d(n_27072), .o(n_27365) );
oa22s01 g752698 ( .a(n_27242), .b(n_27214), .c(n_27241), .d(n_27215), .o(n_27364) );
in01s01 g752699 ( .a(n_27313), .o(n_27314) );
oa12s01 g752700 ( .a(n_27243), .b(n_27244), .c(n_27151), .o(n_27313) );
ao12s04 g752702 ( .a(n_28615), .b(n_27993), .c(n_27899), .o(n_28202) );
no02f08 g752703 ( .a(n_27362), .b(n_27361), .o(n_27363) );
na02f08 g752704 ( .a(n_27244), .b(n_27243), .o(n_27245) );
ao12s04 g752705 ( .a(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .b(n_27997), .c(n_27988), .o(n_27998) );
oa22s01 g752706 ( .a(n_27238), .b(n_27043), .c(n_27237), .d(n_27042), .o(n_27360) );
in01s01 g752707 ( .a(n_28993), .o(n_28134) );
oa22s02 g752708 ( .a(n_27932), .b(n_28021), .c(n_27997), .d(n_28022), .o(n_28993) );
na02s01 g752710 ( .a(n_28054), .b(n_28053), .o(n_28055) );
oa12s04 g752711 ( .a(n_28054), .b(n_27954), .c(n_27923), .o(n_28615) );
in01s01 g752712 ( .a(n_27358), .o(n_27359) );
in01s01 g752713 ( .a(n_27362), .o(n_27358) );
na02f08 g752714 ( .a(n_27194), .b(n_27026), .o(n_27362) );
in01s01 g752715 ( .a(n_27241), .o(n_27242) );
in01s01 g752716 ( .a(n_27244), .o(n_27241) );
oa22s01 g752718 ( .a(n_27161), .b(n_27082), .c(n_27128), .d(n_27081), .o(n_27279) );
in01s01 g752719 ( .a(n_27239), .o(n_27240) );
oa12s01 g752720 ( .a(n_27068), .b(n_27128), .c(n_27073), .o(n_27239) );
in01s01 g752721 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_11_), .o(n_28365) );
na02s01 g752723 ( .a(n_27960), .b(n_27813), .o(n_28027) );
no02s02 g752724 ( .a(n_27883), .b(n_27988), .o(n_27933) );
in01s01 g752725 ( .a(n_27997), .o(n_27932) );
ao12s06 g752726 ( .a(n_27787), .b(n_27909), .c(n_27882), .o(n_27997) );
ao12s04 g752727 ( .a(n_44046), .b(n_27814), .c(n_27899), .o(n_28054) );
no02s02 g752728 ( .a(n_27549), .b(n_27292), .o(n_27551) );
no02s02 g752729 ( .a(n_27549), .b(n_27548), .o(n_27550) );
ao12s02 g752730 ( .a(n_27906), .b(n_27956), .c(n_27928), .o(n_28052) );
oa22s01 g752731 ( .a(n_27159), .b(n_27021), .c(n_27158), .d(n_27022), .o(n_27278) );
in01s01 g752732 ( .a(n_27237), .o(n_27238) );
ao12s01 g752733 ( .a(n_27192), .b(n_27193), .c(n_26958), .o(n_27237) );
oa12f06 g752734 ( .a(n_27011), .b(n_27193), .c(n_27192), .o(n_27194) );
in01s01 g752735 ( .a(n_27994), .o(n_27995) );
ao12s01 g752736 ( .a(n_27908), .b(n_27909), .c(n_27907), .o(n_27994) );
in01s01 g752737 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_11_), .o(n_28367) );
na02s02 g752740 ( .a(n_27909), .b(n_27882), .o(n_27883) );
no02s01 g752741 ( .a(n_27909), .b(n_27907), .o(n_27908) );
in01s01 g752742 ( .a(n_44046), .o(n_27960) );
oa12s02 g752745 ( .a(n_28204), .b(n_27880), .c(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n_27959) );
na02m08 g752746 ( .a(n_27355), .b(n_27433), .o(n_27513) );
no02s02 g752747 ( .a(n_27434), .b(n_27470), .o(n_27471) );
na02s08 g752750 ( .a(n_27512), .b(n_27352), .o(n_27549) );
ao12s02 g752751 ( .a(n_27548), .b(n_27510), .c(FE_OCPN945_n_27287), .o(n_27561) );
oa22s01 g752752 ( .a(n_27077), .b(n_27037), .c(n_27076), .d(n_27038), .o(n_27129) );
in01s01 g752754 ( .a(n_27128), .o(n_27161) );
in01s01 g752755 ( .a(n_27104), .o(n_27128) );
oa12f08 g752756 ( .a(n_27020), .b(n_27058), .c(n_26980), .o(n_27104) );
in01s01 g752757 ( .a(n_27957), .o(n_27958) );
oa22s01 g752758 ( .a(n_27851), .b(n_186), .c(n_27852), .d(n_179), .o(n_27957) );
no02m04 g752760 ( .a(n_27437), .b(n_27121), .o(n_27439) );
no02s04 g752761 ( .a(n_27437), .b(n_27276), .o(n_27438) );
no02s08 g752762 ( .a(n_27402), .b(n_27307), .o(n_27512) );
no02m02 g752763 ( .a(n_27402), .b(n_27464), .o(n_27511) );
oa12s06 g752765 ( .a(n_27812), .b(n_27763), .c(n_179), .o(n_27909) );
in01s01 g752766 ( .a(n_27955), .o(n_27956) );
ao12s02 g752767 ( .a(n_27929), .b(n_27875), .c(n_27791), .o(n_27955) );
na02s01 TIMEBOOST_cell_7658 ( .a(FE_OCP_RBN4920_n_33691), .b(FE_OCP_RBN6668_n_34297), .o(TIMEBOOST_net_2460) );
na02s06 TIMEBOOST_cell_8619 ( .a(TIMEBOOST_net_2796), .b(TIMEBOOST_net_1153), .o(n_10991) );
ao12s01 g752771 ( .a(n_27923), .b(n_28132), .c(n_27721), .o(n_28152) );
oa12s02 g752772 ( .a(n_27899), .b(n_27902), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_11_), .o(n_27928) );
oa22s01 g752773 ( .a(n_27089), .b(n_26984), .c(n_27088), .d(n_26983), .o(n_27160) );
in01s01 g752774 ( .a(n_27158), .o(n_27159) );
in01s01 g752775 ( .a(n_27193), .o(n_27158) );
oa12f08 g752776 ( .a(n_26875), .b(n_27075), .c(n_26960), .o(n_27193) );
no02m02 g752777 ( .a(n_27437), .b(n_27356), .o(n_27436) );
in01s06 g752779 ( .a(n_27434), .o(n_27433) );
na02m06 g752780 ( .a(n_27357), .b(n_27312), .o(n_27434) );
na02s01 g752782 ( .a(n_28196), .b(n_27790), .o(n_28238) );
in01s01 g752784 ( .a(n_27905), .o(n_27906) );
no02s02 g752785 ( .a(n_27881), .b(n_27903), .o(n_27905) );
in01s01 g752788 ( .a(n_28079), .o(n_28080) );
no02s01 g752789 ( .a(n_28051), .b(n_27992), .o(n_28079) );
in01s01 g752790 ( .a(n_28130), .o(n_28131) );
no02s01 g752791 ( .a(n_28107), .b(n_28106), .o(n_28130) );
no02s01 g752793 ( .a(n_28199), .b(n_28198), .o(n_28214) );
no02s01 g752794 ( .a(n_28077), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_27_), .o(n_28129) );
na02s02 g752795 ( .a(n_27813), .b(n_27453), .o(n_27814) );
no02s06 g752796 ( .a(n_27853), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_19_), .o(n_27854) );
no02s02 g752797 ( .a(n_27901), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_23_), .o(n_27954) );
na02s01 g752798 ( .a(n_27951), .b(n_27575), .o(n_27993) );
no02s02 g752800 ( .a(n_27810), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_7_), .o(n_27880) );
no02s01 g752801 ( .a(n_28076), .b(n_27853), .o(n_28585) );
no02s01 g752802 ( .a(n_28106), .b(n_28105), .o(n_28666) );
na02s01 g752803 ( .a(n_28053), .b(n_28075), .o(n_28637) );
no02s01 g752804 ( .a(n_28050), .b(n_28025), .o(n_28445) );
no02s01 g752805 ( .a(n_27992), .b(n_27789), .o(n_28588) );
no02s01 g752806 ( .a(n_28297), .b(n_28257), .o(n_28379) );
no02s01 g752807 ( .a(n_28259), .b(n_28213), .o(n_28498) );
na02s01 g752808 ( .a(n_28156), .b(n_28174), .o(n_28710) );
no02s01 g752809 ( .a(n_28198), .b(n_28078), .o(n_28728) );
no02s01 g752810 ( .a(n_27792), .b(n_27929), .o(n_28338) );
no02s01 g752811 ( .a(n_27903), .b(n_27902), .o(n_28351) );
na02s01 g752812 ( .a(n_27879), .b(n_27926), .o(n_28244) );
na02s01 g752813 ( .a(n_27788), .b(n_27882), .o(n_27907) );
in01s01 g752814 ( .a(n_27851), .o(n_27852) );
na02s01 g752815 ( .a(n_27764), .b(n_27812), .o(n_27851) );
no02s01 g752816 ( .a(n_28280), .b(n_27953), .o(n_28278) );
na02s01 g752817 ( .a(n_27986), .b(n_27877), .o(n_28135) );
in01m02 g752818 ( .a(n_27437), .o(n_27403) );
in01m06 g752819 ( .a(n_27357), .o(n_27437) );
no02s02 TIMEBOOST_cell_8606 ( .a(n_39095), .b(n_39089), .o(TIMEBOOST_net_2790) );
na02m02 g752821 ( .a(n_27310), .b(n_27230), .o(n_27356) );
no02m04 g752822 ( .a(n_27276), .b(n_27234), .o(n_27312) );
na02s02 g752823 ( .a(n_27273), .b(n_27355), .o(n_27470) );
no02f08 TIMEBOOST_cell_7054 ( .a(TIMEBOOST_net_2285), .b(n_39709), .o(n_39748) );
in01s02 g752826 ( .a(n_27402), .o(n_27430) );
na02m06 g752827 ( .a(n_27206), .b(n_27272), .o(n_27402) );
na02s01 g752828 ( .a(n_27351), .b(n_27291), .o(n_27548) );
na02s02 g752829 ( .a(n_27469), .b(FE_OCPN6927_n_26464), .o(n_27510) );
ao12s01 g752830 ( .a(n_28199), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_29_), .o(n_28753) );
ao12s01 g752831 ( .a(n_28108), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_19_), .o(n_28619) );
ao12s01 g752832 ( .a(n_28326), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_30_), .o(n_28756) );
ao12s01 g752833 ( .a(n_28051), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_21_), .o(n_28616) );
ao12s01 g752834 ( .a(n_28175), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_23_), .o(n_28692) );
ao12s01 g752835 ( .a(n_28107), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_25_), .o(n_28713) );
ao12s01 g752836 ( .a(n_28200), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_27_), .o(n_28750) );
in01s01 g752837 ( .a(n_28276), .o(n_28277) );
ao12s01 g752838 ( .a(n_27881), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_11_), .o(n_28276) );
in01s01 g752839 ( .a(n_28314), .o(n_28315) );
ao12s01 g752840 ( .a(n_28018), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_15_), .o(n_28314) );
in01s01 g752841 ( .a(n_28023), .o(n_28024) );
ao12s01 g752842 ( .a(n_27991), .b(n_27762), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_7_), .o(n_28023) );
ao12s01 g752843 ( .a(n_27990), .b(n_27762), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_5_), .o(n_28241) );
no02s02 g752844 ( .a(n_27354), .b(n_27304), .o(n_27429) );
oa22s01 g752845 ( .a(n_27047), .b(n_27005), .c(n_27013), .d(n_27004), .o(n_27059) );
in01s01 g752846 ( .a(n_27076), .o(n_27077) );
in01s01 g752847 ( .a(n_27058), .o(n_27076) );
oa12f08 g752848 ( .a(n_26982), .b(n_27047), .c(n_26913), .o(n_27058) );
no02s01 g752849 ( .a(n_27428), .b(n_27394), .o(n_27509) );
oa22s01 g752850 ( .a(n_27285), .b(n_27923), .c(n_27948), .d(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .o(n_28558) );
oa22s01 g752851 ( .a(n_27164), .b(n_27923), .c(n_27948), .d(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_), .o(n_28434) );
in01s01 g752852 ( .a(n_28021), .o(n_28022) );
oa22s01 g752853 ( .a(n_27988), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .c(n_27762), .d(delay_sub_ln23_0_unr20_stage7_stallmux_q_3_), .o(n_28021) );
in01s01 g752854 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_9_), .o(n_28305) );
in01s01 g752856 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_9_), .o(n_28342) );
na02s06 g752903 ( .a(n_27050), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n_27882) );
in01s01 g752904 ( .a(n_28132), .o(n_28078) );
na02s01 g752905 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_28_), .o(n_28132) );
no02s02 g752906 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_10_), .o(n_27903) );
no02s01 g752907 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_7_), .o(n_27991) );
in01s01 g752908 ( .a(n_27986), .o(n_27987) );
na02s01 g752909 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_4_), .o(n_27986) );
in01s01 g752910 ( .a(n_27791), .o(n_27792) );
na02s02 g752911 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_9_), .o(n_27791) );
no02s01 g752912 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_29_), .o(n_28199) );
no02s01 g752913 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_), .o(n_28297) );
in01s01 g752914 ( .a(n_28128), .o(n_28174) );
no02s01 g752915 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_26_), .o(n_28128) );
in01s01 g752916 ( .a(n_27951), .o(n_28105) );
na02s01 g752917 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_24_), .b(n_27899), .o(n_27951) );
in01s03 g752918 ( .a(n_27790), .o(n_27853) );
na02s06 g752919 ( .a(n_27733), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_18_), .o(n_27790) );
na02s06 g752920 ( .a(FE_OCP_RBN2282_delay_sub_ln23_unr21_stage7_stallmux_q_1_), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_1_), .o(n_27812) );
in01s01 g752921 ( .a(n_27992), .o(n_27950) );
no02s01 g752922 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_20_), .o(n_27992) );
in01s01 g752923 ( .a(n_27813), .o(n_27789) );
na02s01 g752924 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_20_), .o(n_27813) );
in01s01 g752925 ( .a(n_28156), .o(n_28077) );
na02s01 g752926 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_26_), .b(n_27899), .o(n_28156) );
in01s01 g752927 ( .a(n_28212), .o(n_28213) );
na02s01 g752928 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .o(n_28212) );
in01s01 g752929 ( .a(n_28053), .o(n_27901) );
na02s01 g752930 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_22_), .o(n_28053) );
no02s01 g752931 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_19_), .o(n_28108) );
in01s01 g752932 ( .a(n_28076), .o(n_28154) );
no02s01 g752933 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_18_), .b(n_27899), .o(n_28076) );
in01s01 g752934 ( .a(n_27949), .o(n_28025) );
na02s01 g752935 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_14_), .b(n_27899), .o(n_27949) );
no02s02 g752936 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_11_), .o(n_27881) );
no02s02 g752937 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_9_), .b(n_27765), .o(n_27929) );
no02s01 g752938 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_5_), .o(n_27990) );
in01s01 g752939 ( .a(n_27878), .o(n_27879) );
no02s01 g752940 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_6_), .o(n_27878) );
in01s01 g752941 ( .a(n_27876), .o(n_27877) );
no02s01 g752942 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_4_), .o(n_27876) );
in01s01 g752943 ( .a(n_27763), .o(n_27764) );
no02s06 g752944 ( .a(FE_OCP_RBN2282_delay_sub_ln23_unr21_stage7_stallmux_q_1_), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_1_), .o(n_27763) );
in01s01 g752945 ( .a(n_27787), .o(n_27788) );
no02s02 g752946 ( .a(n_27050), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n_27787) );
in01s01 g752947 ( .a(n_27926), .o(n_27810) );
na02s02 g752948 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_6_), .o(n_27926) );
no02s01 g752949 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_8_), .o(n_28280) );
in01s01 g752950 ( .a(n_27848), .o(n_27902) );
na02s02 g752951 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_10_), .o(n_27848) );
in01s01 g752952 ( .a(n_27875), .o(n_27953) );
na02s01 g752953 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_8_), .o(n_27875) );
no02s01 g752955 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_14_), .b(n_27899), .o(n_28050) );
no02s01 g752957 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_15_), .b(n_27899), .o(n_28018) );
no02s01 g752958 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_21_), .o(n_28051) );
in01s01 g752959 ( .a(n_28176), .o(n_28075) );
no02s01 g752960 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_22_), .o(n_28176) );
no02s01 g752961 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_23_), .o(n_28175) );
no02s01 g752962 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_25_), .o(n_28107) );
no02s01 g752963 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_24_), .o(n_28106) );
no02s01 g752964 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_27_), .o(n_28200) );
in01s01 g752965 ( .a(n_28198), .o(n_28173) );
no02s01 g752966 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_28_), .o(n_28198) );
no02s01 g752967 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_30_), .o(n_28326) );
no02s01 g752968 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .o(n_28259) );
in01s01 g752969 ( .a(n_28256), .o(n_28257) );
na02s01 g752970 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_), .o(n_28256) );
na02s02 g752971 ( .a(n_27274), .b(FE_OCP_RBN4486_n_27145), .o(n_27277) );
oa12s01 g752972 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_5_), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_4_), .o(n_28204) );
ao12s01 g752973 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .o(n_28109) );
in01s01 g752974 ( .a(n_28195), .o(n_28196) );
no02s01 g752975 ( .a(n_27931), .b(n_27923), .o(n_28195) );
oa12s01 g752977 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_), .o(n_28016) );
oa22s01 g752979 ( .a(n_27044), .b(n_26915), .c(n_27045), .d(n_26916), .o(n_27090) );
in01s01 g752980 ( .a(n_27088), .o(n_27089) );
in01s01 g752981 ( .a(n_27075), .o(n_27088) );
oa12f08 g752982 ( .a(n_26877), .b(n_27028), .c(n_26822), .o(n_27075) );
no02s06 TIMEBOOST_cell_1442 ( .a(TIMEBOOST_net_335), .b(n_24370), .o(n_24626) );
in01s01 g752985 ( .a(n_27276), .o(n_27310) );
no02f04 TIMEBOOST_cell_1444 ( .a(TIMEBOOST_net_336), .b(FE_OCP_RBN7030_n_44259), .o(n_33784) );
in01s01 g752989 ( .a(n_27353), .o(n_27354) );
no02s08 TIMEBOOST_cell_8685 ( .a(TIMEBOOST_net_2829), .b(n_21268), .o(n_21461) );
in01s01 g752992 ( .a(n_27400), .o(n_27401) );
na02s02 g752994 ( .a(n_27263), .b(FE_OCP_RBN6217_n_27110), .o(n_27352) );
na02s02 g752995 ( .a(n_27184), .b(n_27098), .o(n_27272) );
no02s02 g752996 ( .a(n_27226), .b(n_27110), .o(n_27307) );
no03s40 TIMEBOOST_cell_3452 ( .a(n_22889), .b(FE_RN_1592_0), .c(FE_RN_1591_0), .o(n_23066) );
in01s01 g752998 ( .a(n_27427), .o(n_27428) );
no02s02 g752999 ( .a(n_27299), .b(n_27294), .o(n_27427) );
in01s01 g753001 ( .a(n_27469), .o(n_27507) );
na02s02 g753002 ( .a(n_27347), .b(FE_OCP_RBN6222_n_27110), .o(n_27469) );
in01m01 g753012 ( .a(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n_27762) );
in01s01 g753017 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_29_), .o(n_27721) );
in01s03 g753024 ( .a(n_27923), .o(n_27899) );
in01s02 g753028 ( .a(FE_OFN622_n_28336), .o(n_32287) );
in01s01 g753035 ( .a(FE_OFN622_n_28336), .o(n_32566) );
in01f01 g753037 ( .a(n_27948), .o(n_28336) );
in01s03 g753061 ( .a(n_27923), .o(n_27948) );
in01s06 g753073 ( .a(n_27923), .o(n_27765) );
in01s10 g753074 ( .a(n_27923), .o(n_27733) );
in01s01 g753076 ( .a(n_27190), .o(n_27191) );
na02s01 g753077 ( .a(n_27126), .b(n_27157), .o(n_27190) );
in01s01 g753078 ( .a(n_27528), .o(n_27529) );
na02s01 g753079 ( .a(n_27506), .b(n_27421), .o(n_27528) );
na02m08 g753080 ( .a(n_27126), .b(n_27125), .o(n_27127) );
in01s02 g753081 ( .a(n_27270), .o(n_27271) );
na02s04 g753082 ( .a(n_27233), .b(n_27232), .o(n_27270) );
na02m04 g753083 ( .a(n_27208), .b(n_27232), .o(n_27269) );
in01s01 g753084 ( .a(n_27305), .o(n_27306) );
no02s02 g753085 ( .a(n_27146), .b(n_27121), .o(n_27305) );
no02s10 g753086 ( .a(n_27123), .b(n_27150), .o(n_27189) );
no02s02 TIMEBOOST_cell_1441 ( .a(n_24322), .b(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(TIMEBOOST_net_335) );
in01s01 g753088 ( .a(n_27267), .o(n_27268) );
na02s02 g753089 ( .a(FE_OCP_RBN4486_n_27145), .b(n_27230), .o(n_27267) );
in01s01 g753090 ( .a(n_27274), .o(n_27229) );
no02s06 g753091 ( .a(n_27146), .b(n_27188), .o(n_27274) );
in01s01 g753093 ( .a(n_27467), .o(n_27468) );
na02s02 g753094 ( .a(n_27425), .b(n_27426), .o(n_27467) );
no02f04 TIMEBOOST_cell_1443 ( .a(FE_OCP_RBN4921_n_33691), .b(n_33782), .o(TIMEBOOST_net_336) );
in01s01 g753097 ( .a(n_27398), .o(n_27399) );
no02s02 g753098 ( .a(n_27223), .b(n_27178), .o(n_27398) );
no03s02 TIMEBOOST_cell_3465 ( .a(FE_RN_2077_0), .b(FE_RN_2076_0), .c(n_1673), .o(TIMEBOOST_net_723) );
in01s01 g753100 ( .a(n_27465), .o(n_27466) );
no02s01 g753101 ( .a(n_27384), .b(n_27667), .o(n_27465) );
na02s01 g753103 ( .a(n_27302), .b(n_27303), .o(n_27304) );
in01s01 g753104 ( .a(n_27396), .o(n_27397) );
no02m01 g753105 ( .a(n_27295), .b(n_27601), .o(n_27396) );
no02m04 g753107 ( .a(n_27250), .b(n_27173), .o(n_27301) );
na02s02 g753108 ( .a(n_27143), .b(FE_OCP_RBN1015_n_25826), .o(n_27184) );
in01s01 g753109 ( .a(n_27546), .o(n_27547) );
na02s01 g753110 ( .a(n_27455), .b(n_27527), .o(n_27546) );
no02f08 TIMEBOOST_cell_8171 ( .a(n_21705), .b(TIMEBOOST_net_2716), .o(FE_RN_1184_0) );
in01s01 g753113 ( .a(n_27224), .o(n_27225) );
no02s01 g753114 ( .a(n_27152), .b(n_27183), .o(n_27224) );
no02f06 g753115 ( .a(n_27152), .b(n_27151), .o(n_27153) );
in01s01 g753116 ( .a(n_27348), .o(n_27349) );
na02s01 g753117 ( .a(n_27175), .b(n_27143), .o(n_27348) );
no02s06 g753119 ( .a(n_27213), .b(n_27464), .o(n_27504) );
no02s06 g753120 ( .a(n_27213), .b(n_27172), .o(n_27264) );
na02s02 g753121 ( .a(n_27256), .b(n_27218), .o(n_27300) );
na02s02 g753122 ( .a(n_27216), .b(n_27217), .o(n_27263) );
in01s01 g753123 ( .a(n_27502), .o(n_27503) );
na02s01 g753124 ( .a(n_27463), .b(n_27462), .o(n_27502) );
in01s01 g753125 ( .a(n_27423), .o(n_27424) );
na02s01 g753126 ( .a(n_27211), .b(n_27395), .o(n_27423) );
in01s01 g753127 ( .a(n_27500), .o(n_27501) );
na02s01 g753128 ( .a(n_27461), .b(n_27337), .o(n_27500) );
na02s02 g753129 ( .a(n_27298), .b(n_27297), .o(n_27299) );
na02s01 g753130 ( .a(n_27296), .b(n_26398), .o(n_27347) );
na02s01 g753131 ( .a(n_27326), .b(n_27393), .o(n_27394) );
in01f02 g753132 ( .a(n_27498), .o(n_27499) );
na03f06 TIMEBOOST_cell_7229 ( .a(n_15006), .b(n_14919), .c(n_15040), .o(n_15224) );
in01s02 g753134 ( .a(n_27496), .o(n_27497) );
no02s02 g753135 ( .a(n_27391), .b(n_27188), .o(n_27496) );
no02f08 TIMEBOOST_cell_6378 ( .a(TIMEBOOST_net_2040), .b(n_21119), .o(n_21266) );
in01s01 g753138 ( .a(n_27492), .o(n_27493) );
no02s01 g753139 ( .a(n_27309), .b(n_27386), .o(n_27492) );
in01s01 g753140 ( .a(n_27459), .o(n_27460) );
na02s01 g753141 ( .a(n_27303), .b(n_27339), .o(n_27459) );
in01s01 g753142 ( .a(n_27490), .o(n_27491) );
na02s01 g753143 ( .a(n_27338), .b(n_27382), .o(n_27490) );
oa22s01 g753144 ( .a(n_26991), .b(n_26840), .c(n_26992), .d(n_26839), .o(n_27046) );
in01s01 g753145 ( .a(n_27047), .o(n_27013) );
oa12f08 g753146 ( .a(n_26912), .b(n_26993), .c(n_26837), .o(n_27047) );
in01f02 g753147 ( .a(n_27457), .o(n_27458) );
na02m02 g753148 ( .a(n_27334), .b(n_27227), .o(n_27457) );
in01s01 g753149 ( .a(n_27488), .o(n_27489) );
na02s06 TIMEBOOST_cell_2830 ( .a(n_7082), .b(n_7081), .o(TIMEBOOST_net_706) );
in01s01 g753151 ( .a(n_27486), .o(n_27487) );
na02s02 g753152 ( .a(n_27380), .b(n_27329), .o(n_27486) );
in01s01 g753153 ( .a(n_27525), .o(n_27526) );
na02s01 g753154 ( .a(n_27298), .b(n_27413), .o(n_27525) );
in01s01 g753155 ( .a(n_27523), .o(n_27524) );
no02m02 TIMEBOOST_cell_8730 ( .a(n_12614), .b(n_12497), .o(TIMEBOOST_net_2852) );
in01s01 g753157 ( .a(n_27484), .o(n_27485) );
no02m04 TIMEBOOST_cell_8585 ( .a(TIMEBOOST_net_2779), .b(n_35118), .o(n_35139) );
oa22s01 g753159 ( .a(n_26993), .b(n_26954), .c(n_26922), .d(n_26955), .o(n_27029) );
in01s01 g753160 ( .a(n_27544), .o(n_27545) );
na02s01 g753161 ( .a(n_27420), .b(n_27456), .o(n_27544) );
in01s01 g753162 ( .a(n_27482), .o(n_27483) );
na02s02 g753163 ( .a(n_27342), .b(n_27387), .o(n_27482) );
in01s01 g753164 ( .a(n_27480), .o(n_27481) );
na02s01 g753165 ( .a(n_27340), .b(n_27383), .o(n_27480) );
in01s01 g753166 ( .a(n_27542), .o(n_27543) );
oa22s01 g753167 ( .a(FE_OCPN945_n_27287), .b(n_25781), .c(FE_OCP_RBN6218_n_27110), .d(n_25810), .o(n_27542) );
in01s01 g753168 ( .a(n_27521), .o(n_27522) );
na02s01 g753169 ( .a(n_27414), .b(n_27381), .o(n_27521) );
in01s01 g753170 ( .a(n_27519), .o(n_27520) );
na02s01 g753171 ( .a(n_27410), .b(n_27376), .o(n_27519) );
na02s06 g753174 ( .a(n_27070), .b(FE_OCPN5120_n_25595), .o(n_27126) );
na02s01 g753176 ( .a(n_27204), .b(n_25822), .o(n_27506) );
in01s01 g753177 ( .a(n_27421), .o(n_27422) );
na02s01 g753178 ( .a(n_27207), .b(n_25789), .o(n_27421) );
na02s01 g753179 ( .a(n_27204), .b(n_25777), .o(n_27420) );
na02s01 g753180 ( .a(FE_OCPN1236_n_27207), .b(n_25757), .o(n_27456) );
in01m01 g753181 ( .a(n_27124), .o(n_27232) );
no02m04 g753182 ( .a(FE_OCP_RBN5203_n_25729), .b(n_27103), .o(n_27124) );
in01s03 g753183 ( .a(n_27150), .o(n_27233) );
no02f01 g753185 ( .a(n_25816), .b(FE_OCPN1236_n_27207), .o(n_27392) );
no02s06 g753186 ( .a(n_27120), .b(FE_OCP_RBN3078_n_25816), .o(n_27123) );
na02m06 TIMEBOOST_cell_3003 ( .a(TIMEBOOST_net_792), .b(n_41962), .o(n_42030) );
no02m06 g753191 ( .a(n_27103), .b(FE_OCP_RBN5199_n_25893), .o(n_27121) );
no02s06 g753195 ( .a(n_27120), .b(FE_OCP_RBN5198_n_25893), .o(n_27146) );
no02s01 g753196 ( .a(n_27207), .b(n_25962), .o(n_27391) );
no02s06 g753197 ( .a(FE_OCP_RBN6213_n_27086), .b(n_25963), .o(n_27188) );
in01s01 g753198 ( .a(n_27119), .o(n_27230) );
no02s02 g753199 ( .a(n_27103), .b(FE_OCP_RBN6034_n_46962), .o(n_27119) );
no02s04 g753201 ( .a(FE_OCP_RBN6214_n_27086), .b(FE_OCP_RBN3152_n_46962), .o(n_27145) );
no02s01 g753202 ( .a(FE_OCPN1236_n_27207), .b(n_25999), .o(n_27390) );
na03m06 TIMEBOOST_cell_8357 ( .a(n_9524), .b(n_9439), .c(n_9549), .o(n_9791) );
in01s01 g753205 ( .a(n_27426), .o(n_27388) );
na02s02 g753206 ( .a(n_27204), .b(n_25928), .o(n_27426) );
in01s01 g753207 ( .a(n_27425), .o(n_27343) );
na02s02 g753208 ( .a(n_27207), .b(FE_OCP_RBN6029_n_25928), .o(n_27425) );
na02s01 g753209 ( .a(n_27204), .b(n_26107), .o(n_27342) );
na02s01 g753210 ( .a(n_27207), .b(n_26114), .o(n_27387) );
in01s01 g753212 ( .a(n_27144), .o(n_27178) );
na02s02 g753213 ( .a(FE_OCP_RBN6214_n_27086), .b(n_26011), .o(n_27144) );
no02s02 g753217 ( .a(n_27120), .b(n_26011), .o(n_27223) );
no02s01 g753218 ( .a(n_27207), .b(FE_OCP_RBN6031_n_25997), .o(n_27386) );
no02s01 g753219 ( .a(n_27120), .b(FE_OCP_RBN6819_n_25997), .o(n_27309) );
in01s01 g753220 ( .a(n_27222), .o(n_27667) );
na02s01 g753221 ( .a(n_27120), .b(FE_OCPN6935_FE_OCP_RBN6066_n_26081), .o(n_27222) );
in01s01 g753223 ( .a(n_27384), .o(n_27418) );
no02s01 g753224 ( .a(n_27204), .b(FE_OCPN6935_FE_OCP_RBN6066_n_26081), .o(n_27384) );
na02s01 g753225 ( .a(n_27204), .b(n_26200), .o(n_27340) );
na02s01 g753226 ( .a(n_27207), .b(n_26171), .o(n_27383) );
na02s01 g753227 ( .a(n_27204), .b(n_26169), .o(n_27339) );
na02s01 g753228 ( .a(n_27207), .b(FE_OCP_RBN3247_n_26169), .o(n_27303) );
na02s01 g753229 ( .a(n_27204), .b(n_26146), .o(n_27338) );
na02s01 g753230 ( .a(n_27207), .b(FE_OCP_RBN4392_n_26146), .o(n_27382) );
in01s01 g753231 ( .a(n_27336), .o(n_27337) );
in01s01 g753233 ( .a(n_27296), .o(n_27336) );
na02s01 g753234 ( .a(FE_OCP_RBN3253_n_26276), .b(n_27167), .o(n_27296) );
na02s01 g753235 ( .a(FE_OCP_RBN6218_n_27110), .b(n_26201), .o(n_27381) );
in01s02 g753237 ( .a(n_27175), .o(n_27219) );
na02s03 g753238 ( .a(n_27110), .b(FE_OCP_RBN1038_n_45533), .o(n_27175) );
na02s01 g753239 ( .a(n_27110), .b(n_27217), .o(n_27218) );
na02s01 g753240 ( .a(FE_OCP_RBN6218_n_27110), .b(n_27217), .o(n_27380) );
in01s01 g753241 ( .a(n_27216), .o(n_27601) );
na02s06 g753242 ( .a(n_27167), .b(FE_OCP_RBN4367_n_25889), .o(n_27216) );
in01s01 g753243 ( .a(n_27214), .o(n_27215) );
na02s01 g753244 ( .a(n_27113), .b(n_27243), .o(n_27214) );
no02f02 g753245 ( .a(n_27083), .b(n_25598), .o(n_27152) );
in01s01 g753247 ( .a(n_27454), .o(n_27455) );
no02s01 g753248 ( .a(FE_OCPN945_n_27287), .b(n_27416), .o(n_27454) );
na02s01 g753249 ( .a(FE_OCPN945_n_27287), .b(n_27416), .o(n_27527) );
in01s01 g753251 ( .a(n_27143), .o(n_27173) );
na02s02 g753252 ( .a(n_27098), .b(FE_OCP_RBN1039_n_45533), .o(n_27143) );
na02f06 g753253 ( .a(FE_OCPN945_n_27287), .b(FE_OCP_RBN1014_n_25826), .o(n_27334) );
na02s02 g753254 ( .a(n_27110), .b(FE_OCP_RBN1015_n_25826), .o(n_27227) );
no02s04 TIMEBOOST_cell_1399 ( .a(n_42122), .b(n_42196), .o(TIMEBOOST_net_314) );
no02m03 g753260 ( .a(n_27167), .b(FE_OCP_RBN1032_n_25844), .o(n_27213) );
no02s01 g753261 ( .a(FE_OCP_RBN6218_n_27110), .b(n_25915), .o(n_27378) );
no02s06 g753262 ( .a(n_27167), .b(n_27170), .o(n_27172) );
na02f08 TIMEBOOST_cell_2829 ( .a(TIMEBOOST_net_705), .b(n_7270), .o(n_7332) );
in01s01 g753266 ( .a(n_27256), .o(n_27295) );
na02s02 g753267 ( .a(n_27110), .b(FE_OCP_RBN1166_n_25889), .o(n_27256) );
na02s02 g753268 ( .a(FE_OCPN945_n_27287), .b(n_25980), .o(n_27329) );
in01s01 g753269 ( .a(n_27462), .o(n_27415) );
na02s01 g753270 ( .a(FE_OCP_RBN6218_n_27110), .b(n_26110), .o(n_27462) );
na02s01 g753271 ( .a(FE_OCPN945_n_27287), .b(n_26174), .o(n_27414) );
in01s01 g753274 ( .a(n_27211), .o(n_27254) );
na02s01 g753275 ( .a(FE_OCP_RBN4390_n_26173), .b(n_27167), .o(n_27211) );
in01s01 g753277 ( .a(n_27294), .o(n_27395) );
no02m01 g753278 ( .a(n_27167), .b(FE_OCP_RBN4390_n_26173), .o(n_27294) );
na02s01 g753279 ( .a(FE_OCPN945_n_27287), .b(n_26323), .o(n_27413) );
na02s02 g753280 ( .a(FE_OCP_RBN6221_n_27110), .b(FE_OCPN1683_n_27210), .o(n_27298) );
in01s01 g753281 ( .a(n_27461), .o(n_27411) );
na02s01 g753282 ( .a(FE_OCP_RBN6218_n_27110), .b(n_26276), .o(n_27461) );
na02s01 g753283 ( .a(FE_OCPN945_n_27287), .b(FE_OCP_RBN6120_n_26398), .o(n_27410) );
na02s01 g753284 ( .a(FE_OCP_RBN6221_n_27110), .b(n_26398), .o(n_27376) );
na03s01 TIMEBOOST_cell_8256 ( .a(n_977), .b(n_951), .c(n_865), .o(n_943) );
na02s01 g753286 ( .a(FE_OCP_RBN6221_n_27110), .b(FE_OCPN6927_n_26464), .o(n_27393) );
no02s01 TIMEBOOST_cell_6392 ( .a(TIMEBOOST_net_2047), .b(n_22438), .o(n_22457) );
na02s01 g753288 ( .a(FE_OCP_RBN6221_n_27110), .b(n_26652), .o(n_27375) );
in01s01 g753289 ( .a(n_27463), .o(n_27373) );
na02s06 g753290 ( .a(FE_OCPN945_n_27287), .b(n_26048), .o(n_27463) );
in01s01 g753291 ( .a(n_27677), .o(n_27678) );
oa12f02 g753292 ( .a(n_27627), .b(n_27657), .c(n_26896), .o(n_27677) );
in01s01 g753293 ( .a(n_27044), .o(n_27045) );
in01s01 g753294 ( .a(n_27028), .o(n_27044) );
no02f08 g753295 ( .a(n_26971), .b(n_26847), .o(n_27028) );
in01s01 g753298 ( .a(n_27168), .o(n_27208) );
no02s06 g753299 ( .a(n_27086), .b(n_25823), .o(n_27168) );
no02s03 g753300 ( .a(n_27120), .b(n_26116), .o(n_27308) );
na02s02 g753301 ( .a(n_26115), .b(n_27120), .o(n_27355) );
na02s01 g753302 ( .a(n_27207), .b(n_26250), .o(n_27302) );
in01m02 g753305 ( .a(n_27206), .o(n_27250) );
in01s01 g753308 ( .a(n_27291), .o(n_27292) );
na02s01 g753309 ( .a(n_27167), .b(n_26247), .o(n_27291) );
na02s01 g753310 ( .a(n_27110), .b(n_26213), .o(n_27297) );
in01s01 g753312 ( .a(n_27326), .o(n_27371) );
na02s01 g753313 ( .a(FE_OCP_RBN6221_n_27110), .b(n_26471), .o(n_27326) );
oa22s01 g753314 ( .a(n_27611), .b(n_26869), .c(n_27612), .d(n_26870), .o(n_27656) );
oa22s01 g753315 ( .a(n_27626), .b(n_26935), .c(n_27657), .d(n_26936), .o(n_27676) );
in01s01 g753316 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_7_), .o(n_28227) );
in01s01 g753318 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_7_), .o(n_26972) );
no02f06 g753321 ( .a(n_26970), .b(n_26846), .o(n_26971) );
in01s01 g753322 ( .a(n_27101), .o(n_27102) );
na02s01 g753323 ( .a(n_27125), .b(n_27055), .o(n_27101) );
in01s01 g753324 ( .a(n_26991), .o(n_26992) );
na02s01 g753325 ( .a(n_26970), .b(n_26755), .o(n_26991) );
in01s01 g753326 ( .a(n_27151), .o(n_27113) );
no02f06 g753327 ( .a(n_27100), .b(n_27099), .o(n_27151) );
in01s01 g753328 ( .a(n_27071), .o(n_27072) );
na02s01 g753329 ( .a(n_27057), .b(n_27025), .o(n_27071) );
na02f06 g753331 ( .a(n_27100), .b(n_27099), .o(n_27243) );
oa12f02 g753332 ( .a(n_26907), .b(n_27613), .c(FE_OCP_RBN4435_n_26160), .o(n_27627) );
in01s08 g753339 ( .a(n_27070), .o(n_27086) );
in01s06 g753344 ( .a(n_27207), .o(n_27204) );
in01m10 g753352 ( .a(n_27120), .o(n_27207) );
in01f10 g753356 ( .a(n_27103), .o(n_27120) );
in01m08 g753357 ( .a(n_27070), .o(n_27103) );
na02f10 g753359 ( .a(n_27012), .b(n_27027), .o(n_27070) );
oa22s01 g753360 ( .a(n_26882), .b(n_26776), .c(n_26852), .d(n_26777), .o(n_26969) );
in01s01 g753361 ( .a(n_26993), .o(n_26922) );
oa12f08 g753362 ( .a(n_26819), .b(n_26883), .c(n_26774), .o(n_26993) );
in01s10 g753379 ( .a(n_27110), .o(n_27167) );
in01m10 g753380 ( .a(n_27098), .o(n_27110) );
in01m08 g753387 ( .a(n_27083), .o(n_27098) );
oa22s01 g753389 ( .a(n_26883), .b(n_26836), .c(n_26828), .d(n_26835), .o(n_26968) );
na02f08 g753391 ( .a(n_26988), .b(n_26963), .o(n_27027) );
na02f06 g753392 ( .a(n_46422), .b(n_26961), .o(n_27012) );
na02f06 g753393 ( .a(n_26882), .b(n_26754), .o(n_26970) );
in01s01 g753394 ( .a(n_27042), .o(n_27043) );
na02s01 g753395 ( .a(n_26990), .b(n_27026), .o(n_27042) );
no02f06 g753396 ( .a(n_26989), .b(n_26918), .o(n_27011) );
na02m04 g753397 ( .a(n_27041), .b(n_27040), .o(n_27125) );
in01s01 g753398 ( .a(n_27361), .o(n_27055) );
no02m04 g753399 ( .a(n_27041), .b(n_27040), .o(n_27361) );
in01s01 g753400 ( .a(n_27081), .o(n_27082) );
na02s01 g753401 ( .a(n_27068), .b(n_27036), .o(n_27081) );
na02f04 g753402 ( .a(n_27010), .b(FE_OCPN1737_n_27009), .o(n_27057) );
in01s01 g753403 ( .a(n_27024), .o(n_27025) );
no02s04 g753404 ( .a(n_27010), .b(n_27009), .o(n_27024) );
in01s01 g753405 ( .a(n_27657), .o(n_27626) );
no02f04 g753406 ( .a(n_27613), .b(n_26833), .o(n_27657) );
in01s01 g753407 ( .a(n_27611), .o(n_27612) );
ao12s01 g753408 ( .a(n_26769), .b(n_27589), .c(n_26832), .o(n_27611) );
oa22s01 g753409 ( .a(n_26809), .b(n_26719), .c(n_26808), .d(n_26718), .o(n_26881) );
na02f06 g753410 ( .a(n_27039), .b(n_27023), .o(n_27100) );
oa22s01 g753411 ( .a(FE_OCP_DRV_N1514_n_26786), .b(n_26750), .c(n_26787), .d(n_26751), .o(n_26853) );
oa22s01 g753412 ( .a(n_27586), .b(n_26829), .c(n_27587), .d(n_26830), .o(n_27625) );
na02f04 g753416 ( .a(n_27007), .b(n_26487), .o(n_27039) );
na02s04 g753417 ( .a(n_27006), .b(n_26456), .o(n_27023) );
in01s01 g753418 ( .a(n_26882), .o(n_26852) );
ao12f06 g753419 ( .a(n_26691), .b(n_26765), .c(n_26660), .o(n_26882) );
in01s01 g753420 ( .a(n_27021), .o(n_27022) );
no02s01 g753421 ( .a(n_27192), .b(n_26918), .o(n_27021) );
in01s01 g753422 ( .a(n_26989), .o(n_26990) );
no02f04 g753423 ( .a(n_26967), .b(n_26966), .o(n_26989) );
na02s02 g753424 ( .a(n_26967), .b(n_26966), .o(n_27026) );
in01s01 g753425 ( .a(n_26883), .o(n_26828) );
na02f08 g753426 ( .a(n_26768), .b(n_26723), .o(n_26883) );
in01s01 g753427 ( .a(n_27037), .o(n_27038) );
na02s01 g753428 ( .a(n_27020), .b(n_26981), .o(n_27037) );
na02f04 g753429 ( .a(n_27019), .b(FE_OCPN5234_n_27018), .o(n_27068) );
in01s01 g753430 ( .a(n_27073), .o(n_27036) );
no02f04 g753431 ( .a(n_27019), .b(FE_OCPN5234_n_27018), .o(n_27073) );
no02f06 g753433 ( .a(n_46422), .b(n_26871), .o(n_26988) );
oa12f08 g753434 ( .a(n_26387), .b(n_26987), .c(n_26985), .o(n_27008) );
no03s06 TIMEBOOST_cell_7141 ( .a(n_13286), .b(n_13349), .c(n_13700), .o(n_13353) );
no02f06 g753436 ( .a(n_27589), .b(n_26817), .o(n_27613) );
no02f08 TIMEBOOST_cell_8647 ( .a(TIMEBOOST_net_2810), .b(n_39607), .o(FE_RN_1874_0) );
oa22s01 g753439 ( .a(n_27559), .b(n_26906), .c(n_27560), .d(n_26905), .o(n_27588) );
in01s01 g753440 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_25_), .o(n_27575) );
no02f08 TIMEBOOST_cell_7584 ( .a(n_24419), .b(n_24441), .o(TIMEBOOST_net_2423) );
na02s04 g753443 ( .a(n_26879), .b(n_26961), .o(n_26962) );
in01f02 g753445 ( .a(n_27006), .o(n_27007) );
no02m06 g753446 ( .a(n_26987), .b(n_26537), .o(n_27006) );
no02s02 TIMEBOOST_cell_5275 ( .a(TIMEBOOST_net_1585), .b(n_3914), .o(n_4229) );
in01s01 g753448 ( .a(n_26983), .o(n_26984) );
no02s01 g753449 ( .a(n_26960), .b(n_26876), .o(n_26983) );
in01s01 g753451 ( .a(n_26918), .o(n_26958) );
no02f04 g753452 ( .a(n_26844), .b(n_25363), .o(n_26918) );
in01s01 g753454 ( .a(n_27004), .o(n_27005) );
na02s01 g753455 ( .a(n_26914), .b(n_26982), .o(n_27004) );
na02m04 g753456 ( .a(n_26957), .b(n_26956), .o(n_27020) );
in01s01 g753457 ( .a(n_26980), .o(n_26981) );
no02m04 g753458 ( .a(n_26957), .b(n_26956), .o(n_26980) );
in01s01 g753459 ( .a(n_27586), .o(n_27587) );
in01s01 g753460 ( .a(n_27589), .o(n_27586) );
no02s04 TIMEBOOST_cell_1234 ( .a(TIMEBOOST_net_231), .b(n_23616), .o(n_23750) );
oa22s01 g753463 ( .a(n_26788), .b(n_26647), .c(n_26732), .d(n_26648), .o(n_26810) );
in01s01 g753464 ( .a(n_26808), .o(n_26809) );
oa12s01 g753465 ( .a(n_26764), .b(n_26788), .c(n_26658), .o(n_26808) );
oa12f06 g753466 ( .a(n_26696), .b(n_26767), .c(n_26766), .o(n_26768) );
na02s04 TIMEBOOST_cell_7842 ( .a(n_15692), .b(n_14452), .o(TIMEBOOST_net_2552) );
oa12s01 g753468 ( .a(n_26763), .b(n_26767), .c(n_26762), .o(n_26807) );
in01s01 g753469 ( .a(FE_OCP_DRV_N1514_n_26786), .o(n_26787) );
ao12s01 g753470 ( .a(n_26766), .b(n_26767), .c(n_26617), .o(n_26786) );
oa22s01 g753471 ( .a(n_27537), .b(n_26790), .c(n_27538), .d(n_26791), .o(n_27574) );
in01s01 g753472 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_5_), .o(n_28124) );
in01s02 g753474 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_5_), .o(n_28220) );
no02s06 TIMEBOOST_cell_7860 ( .a(n_14805), .b(FE_OCP_RBN6057_n_16011), .o(TIMEBOOST_net_2561) );
no02f04 g753478 ( .a(n_26784), .b(n_26749), .o(n_26827) );
in01s02 g753479 ( .a(n_26879), .o(n_26880) );
no02f06 TIMEBOOST_cell_7841 ( .a(TIMEBOOST_net_2551), .b(n_38689), .o(n_38732) );
na02f02 g753482 ( .a(FE_OCP_RBN3355_FE_RN_1058_0), .b(n_26497), .o(n_26878) );
na02s06 TIMEBOOST_cell_7493 ( .a(TIMEBOOST_net_2377), .b(n_23683), .o(n_23737) );
in01s01 g753484 ( .a(n_26915), .o(n_26916) );
na02s01 g753485 ( .a(n_26877), .b(n_26823), .o(n_26915) );
na02f08 g753486 ( .a(n_26788), .b(n_26764), .o(n_26765) );
no02m08 g753487 ( .a(n_26851), .b(FE_OCP_DRV_N1432_n_26850), .o(n_26960) );
in01s01 g753488 ( .a(n_26875), .o(n_26876) );
na02f06 g753489 ( .a(n_26851), .b(FE_OCP_DRV_N1432_n_26850), .o(n_26875) );
in01s01 g753490 ( .a(n_26913), .o(n_26914) );
no02m04 g753491 ( .a(n_26874), .b(n_26873), .o(n_26913) );
na02m04 g753492 ( .a(n_26874), .b(n_26873), .o(n_26982) );
na02s01 g753493 ( .a(n_26762), .b(n_26767), .o(n_26763) );
in01s01 g753494 ( .a(n_26954), .o(n_26955) );
na02s01 g753495 ( .a(n_26912), .b(n_26838), .o(n_26954) );
no02m06 g753497 ( .a(n_26871), .b(n_26824), .o(n_26961) );
ao12f04 g753499 ( .a(n_23564), .b(n_26804), .c(n_26797), .o(n_26919) );
in01m02 g753500 ( .a(n_26848), .o(n_26849) );
ao12f04 g753501 ( .a(n_26581), .b(n_26781), .c(n_26473), .o(n_26848) );
in01s01 g753502 ( .a(n_27559), .o(n_27560) );
na02s01 g753503 ( .a(n_27540), .b(n_26771), .o(n_27559) );
no03f08 TIMEBOOST_cell_8230 ( .a(FE_RN_1673_0), .b(n_23542), .c(n_23600), .o(TIMEBOOST_net_2397) );
na02m06 g753507 ( .a(n_26805), .b(n_26826), .o(n_26957) );
oa22s01 g753508 ( .a(n_27451), .b(n_26895), .c(n_27452), .d(n_26894), .o(n_27539) );
na02m04 g753511 ( .a(n_26778), .b(n_26422), .o(n_26805) );
na02m04 g753512 ( .a(FE_OCP_RBN6132_n_26778), .b(n_26421), .o(n_26826) );
in01s04 g753513 ( .a(n_26872), .o(n_26871) );
na02m06 g753514 ( .a(n_26804), .b(n_23564), .o(n_26872) );
no02s06 g753516 ( .a(n_26804), .b(n_23564), .o(n_26824) );
in01s01 g753520 ( .a(n_27537), .o(n_27538) );
na02s01 g753521 ( .a(n_27450), .b(n_26793), .o(n_27537) );
na02f04 g753522 ( .a(n_27449), .b(n_26770), .o(n_27540) );
in01s01 g753524 ( .a(n_26822), .o(n_26823) );
no02m06 g753525 ( .a(n_26802), .b(FE_OCPN1934_n_26801), .o(n_26822) );
no02s01 TIMEBOOST_cell_1215 ( .a(FE_RN_743_0), .b(n_28326), .o(TIMEBOOST_net_222) );
in01s01 g753527 ( .a(n_26839), .o(n_26840) );
no02s01 g753528 ( .a(n_26846), .b(n_26799), .o(n_26839) );
na02f04 g753529 ( .a(n_26821), .b(n_26820), .o(n_26912) );
in01s01 g753530 ( .a(n_26837), .o(n_26838) );
no02f04 g753531 ( .a(n_26821), .b(n_26820), .o(n_26837) );
in01f02 g753533 ( .a(n_26783), .o(n_26784) );
ao12f04 g753534 ( .a(n_26704), .b(n_26729), .c(FE_OCP_RBN6870_FE_RN_2289_0), .o(n_26783) );
in01s01 g753535 ( .a(n_26788), .o(n_26732) );
ao12f08 g753536 ( .a(n_26586), .b(n_26705), .c(n_26532), .o(n_26788) );
na03m20 TIMEBOOST_cell_3446 ( .a(n_27884), .b(delay_xor_ln21_unr18_stage7_stallmux_q_2_), .c(n_44759), .o(n_27934) );
oa12s01 g753538 ( .a(n_26675), .b(n_26674), .c(n_26705), .o(n_26731) );
na02s03 TIMEBOOST_cell_8814 ( .a(n_44855), .b(n_44498), .o(TIMEBOOST_net_2894) );
oa12f06 g753540 ( .a(n_26616), .b(n_26701), .c(n_26557), .o(n_26767) );
oa12s01 g753541 ( .a(n_26703), .b(n_26702), .c(n_26701), .o(n_26761) );
oa22s01 g753542 ( .a(n_27368), .b(n_26924), .c(n_27367), .d(n_26925), .o(n_27479) );
in01s01 g753546 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_21_), .o(n_27453) );
no02m06 g753548 ( .a(n_26695), .b(n_26614), .o(n_26759) );
na03f02 TIMEBOOST_cell_7186 ( .a(FE_RN_982_0), .b(n_2535), .c(n_2753), .o(FE_RN_984_0) );
na02f04 g753550 ( .a(n_26670), .b(n_26620), .o(n_26704) );
in01m02 g753551 ( .a(n_26785), .o(n_26758) );
no02m08 g753552 ( .a(n_26729), .b(n_26671), .o(n_26785) );
no02f08 g753554 ( .a(n_26756), .b(n_26389), .o(n_26781) );
in01s01 g753555 ( .a(n_27451), .o(n_27452) );
na02s01 g753556 ( .a(n_27406), .b(n_26897), .o(n_27451) );
in01s01 g753557 ( .a(n_27449), .o(n_27450) );
no02f04 g753558 ( .a(n_27406), .b(n_26860), .o(n_27449) );
no02m08 g753559 ( .a(n_26722), .b(n_25101), .o(n_26846) );
no02f04 g753560 ( .a(n_26721), .b(FE_OCP_DRV_N5157_n_25100), .o(n_26799) );
na02s01 g753561 ( .a(n_26674), .b(n_26705), .o(n_26675) );
no02s01 TIMEBOOST_cell_7049 ( .a(n_10305), .b(n_10306), .o(TIMEBOOST_net_2283) );
no02s01 TIMEBOOST_cell_8539 ( .a(TIMEBOOST_net_2756), .b(FE_RN_888_0), .o(TIMEBOOST_net_1511) );
na02s01 g753564 ( .a(n_26702), .b(n_26701), .o(n_26703) );
in01s01 g753565 ( .a(n_26835), .o(n_26836) );
na02s01 g753566 ( .a(n_26775), .b(n_26819), .o(n_26835) );
na02m04 g753568 ( .a(n_26756), .b(n_26520), .o(n_26778) );
na02m06 g753569 ( .a(n_26698), .b(n_26672), .o(n_26802) );
no02f08 g753570 ( .a(n_26699), .b(n_26673), .o(n_26804) );
na02f04 g753571 ( .a(n_26700), .b(n_26726), .o(n_26821) );
oa22s01 g753572 ( .a(n_27322), .b(n_26736), .c(n_27321), .d(n_26737), .o(n_27448) );
oa22s01 g753573 ( .a(n_27320), .b(n_26928), .c(n_27319), .d(n_26929), .o(n_27447) );
no02s01 g753576 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .o(n_27931) );
na02f02 g753578 ( .a(n_26661), .b(FE_OCP_RBN3283_n_26316), .o(n_26700) );
na02m04 g753579 ( .a(FE_OCP_RBN4412_n_26661), .b(n_26316), .o(n_26726) );
no02f08 g753580 ( .a(n_26669), .b(n_26579), .o(n_26729) );
no02f08 g753581 ( .a(n_26652), .b(n_26663), .o(n_26699) );
no02m04 g753582 ( .a(n_26622), .b(FE_OCP_DRV_N6899_FE_OCPN5276_n_23590), .o(n_26673) );
na02f08 g753583 ( .a(n_26697), .b(n_26301), .o(n_26756) );
na02f04 g753584 ( .a(n_27283), .b(n_26898), .o(n_27406) );
na02s04 g753585 ( .a(n_26629), .b(n_26592), .o(n_26698) );
na02s02 g753586 ( .a(n_26628), .b(n_26590), .o(n_26672) );
in01m04 g753587 ( .a(n_26670), .o(n_26671) );
ao12f04 g753588 ( .a(n_26596), .b(n_26539), .c(n_23590), .o(n_26670) );
in01s01 g753589 ( .a(n_26776), .o(n_26777) );
na02s01 g753590 ( .a(n_26755), .b(n_26754), .o(n_26776) );
in01s02 g753591 ( .a(n_26724), .o(n_26725) );
no02s04 g753592 ( .a(n_26697), .b(n_26519), .o(n_26724) );
na02f06 g753593 ( .a(n_26753), .b(n_26752), .o(n_26819) );
in01s01 g753594 ( .a(n_26774), .o(n_26775) );
no02f06 g753595 ( .a(n_26753), .b(n_26752), .o(n_26774) );
no02f04 g753596 ( .a(n_26584), .b(n_26654), .o(n_26696) );
in01s01 g753597 ( .a(n_26750), .o(n_26751) );
na02s01 g753598 ( .a(n_26723), .b(n_26655), .o(n_26750) );
in01f01 g753599 ( .a(n_26748), .o(n_26749) );
na02s02 TIMEBOOST_cell_3334 ( .a(n_11003), .b(n_11013), .o(TIMEBOOST_net_958) );
in01m02 g753601 ( .a(n_26694), .o(n_26695) );
na02m04 g753602 ( .a(n_26669), .b(n_26563), .o(n_26694) );
no03m08 TIMEBOOST_cell_7126 ( .a(n_23228), .b(n_23039), .c(n_23210), .o(n_23305) );
in01s01 g753605 ( .a(n_27367), .o(n_27368) );
ao12s01 g753606 ( .a(n_26742), .b(n_27284), .c(n_26709), .o(n_27367) );
in01m04 g753607 ( .a(n_26721), .o(n_26722) );
ao12f08 g753609 ( .a(n_26462), .b(n_26599), .c(n_26518), .o(n_26705) );
oa12s01 g753610 ( .a(n_26595), .b(n_26594), .c(n_26599), .o(n_26668) );
oa12f06 g753611 ( .a(n_26495), .b(n_26623), .c(n_26559), .o(n_26701) );
oa12s01 g753612 ( .a(n_26625), .b(n_26624), .c(n_26623), .o(n_26693) );
oa22s01 g753613 ( .a(n_27202), .b(n_26889), .c(n_27201), .d(n_26888), .o(n_27323) );
in01s01 g753615 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_3_), .o(n_28115) );
in01s01 g753617 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .o(n_27285) );
na02f08 g753622 ( .a(n_26597), .b(FE_OCP_RBN3279_FE_RN_1496_0), .o(n_26669) );
in01s02 g753623 ( .a(n_46934), .o(n_26747) );
no02s03 g753626 ( .a(n_26583), .b(FE_OCPN5276_n_23590), .o(n_26666) );
na02f10 TIMEBOOST_cell_3333 ( .a(n_36108), .b(TIMEBOOST_net_957), .o(n_36272) );
no02m06 TIMEBOOST_cell_7076 ( .a(TIMEBOOST_net_2296), .b(FE_OCP_RBN6853_n_39793), .o(n_39966) );
no02f08 g753629 ( .a(n_26630), .b(n_26277), .o(n_26697) );
na02m04 g753631 ( .a(n_26630), .b(n_26319), .o(n_26661) );
in01s01 g753632 ( .a(n_27321), .o(n_27322) );
no02s01 g753633 ( .a(n_27284), .b(n_26714), .o(n_27321) );
in01s02 g753634 ( .a(n_26628), .o(n_26629) );
no02m04 g753635 ( .a(n_26597), .b(n_26596), .o(n_26628) );
no02f04 g753636 ( .a(n_26659), .b(n_26658), .o(n_26660) );
na02f04 g753637 ( .a(n_26657), .b(FE_OCP_DRV_N1490_n_26656), .o(n_26754) );
in01s01 g753638 ( .a(n_26692), .o(n_26755) );
no02m04 g753639 ( .a(n_26657), .b(FE_OCP_DRV_N1490_n_26656), .o(n_26692) );
na02s01 g753640 ( .a(n_26594), .b(n_26599), .o(n_26595) );
in01s01 g753641 ( .a(n_26718), .o(n_26719) );
no02s01 g753642 ( .a(n_26659), .b(n_26691), .o(n_26718) );
in01s01 g753643 ( .a(n_26654), .o(n_26655) );
no02f04 g753644 ( .a(n_26627), .b(n_26626), .o(n_26654) );
na02s02 g753645 ( .a(n_26627), .b(n_26626), .o(n_26723) );
na02s01 g753646 ( .a(n_26624), .b(n_26623), .o(n_26625) );
no02s01 g753647 ( .a(n_26584), .b(n_26766), .o(n_26762) );
no02s02 TIMEBOOST_cell_5676 ( .a(FE_RN_1535_0), .b(FE_OCP_RBN6214_n_27086), .o(TIMEBOOST_net_1786) );
in01s01 g753649 ( .a(n_27319), .o(n_27320) );
in01s01 g753650 ( .a(n_27283), .o(n_27319) );
oa12f04 g753651 ( .a(n_26715), .b(n_27203), .c(n_26792), .o(n_27283) );
in01s01 g753652 ( .a(n_26652), .o(n_26653) );
in01f04 g753653 ( .a(n_26622), .o(n_26652) );
oa22s01 g753657 ( .a(n_27132), .b(n_26926), .c(n_27133), .d(n_26927), .o(n_27247) );
oa22s01 g753658 ( .a(n_27198), .b(n_26681), .c(n_27199), .d(n_26682), .o(n_27318) );
in01s01 g753659 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_2_), .o(n_26566) );
na02s02 g753662 ( .a(FE_OCP_RBN3279_FE_RN_1496_0), .b(n_26504), .o(n_26592) );
no02s02 g753663 ( .a(FE_OCP_RBN6850_n_26504), .b(FE_RN_1496_0), .o(n_26590) );
no02m06 g753664 ( .a(n_26540), .b(n_26434), .o(n_26597) );
na02f06 g753666 ( .a(n_26540), .b(FE_OCP_RBN1867_n_26407), .o(n_26564) );
no02s02 g753667 ( .a(FE_OCP_RBN6850_n_26504), .b(n_26596), .o(n_26563) );
na02f02 g753668 ( .a(n_26504), .b(n_26424), .o(n_26539) );
na02s06 g753673 ( .a(n_26553), .b(n_23509), .o(n_26620) );
na02f08 g753674 ( .a(n_26524), .b(n_26363), .o(n_26630) );
no02s01 g753675 ( .a(n_27203), .b(n_26738), .o(n_27284) );
no02f02 g753676 ( .a(n_26588), .b(n_26587), .o(n_26659) );
in01m02 g753677 ( .a(n_26589), .o(n_26691) );
na02s02 g753678 ( .a(n_26588), .b(n_26587), .o(n_26589) );
no02s01 g753679 ( .a(n_26586), .b(n_26533), .o(n_26674) );
in01s01 g753680 ( .a(n_26647), .o(n_26648) );
na02s01 g753681 ( .a(n_26560), .b(n_26764), .o(n_26647) );
no02f04 TIMEBOOST_cell_8781 ( .a(TIMEBOOST_net_2877), .b(n_14855), .o(n_14979) );
in01s01 g753686 ( .a(n_26584), .o(n_26617) );
no02f02 g753687 ( .a(n_26522), .b(n_25013), .o(n_26584) );
na02s01 g753689 ( .a(n_26558), .b(n_26616), .o(n_26702) );
in01s01 g753690 ( .a(n_27201), .o(n_27202) );
ao12s01 g753691 ( .a(n_26815), .b(n_27135), .c(n_26710), .o(n_27201) );
oa12f08 g753692 ( .a(n_26325), .b(n_26506), .c(n_26403), .o(n_26599) );
in01m02 g753694 ( .a(n_26583), .o(n_26664) );
oa12s01 g753696 ( .a(n_26480), .b(n_26479), .c(n_26506), .o(n_26536) );
oa12f06 g753698 ( .a(n_26461), .b(n_26392), .c(n_26525), .o(n_26623) );
oa12s01 g753699 ( .a(n_26527), .b(n_26526), .c(n_26525), .o(n_26582) );
oa22s01 g753700 ( .a(n_27096), .b(n_26891), .c(n_27095), .d(n_26890), .o(n_27165) );
oa22s01 g753701 ( .a(n_27108), .b(n_26683), .c(n_27109), .d(n_26684), .o(n_27200) );
in01m01 g753702 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_1_), .o(n_27865) );
na02m04 g753708 ( .a(n_26580), .b(n_26478), .o(n_26581) );
na02f02 g753713 ( .a(n_26442), .b(FE_RN_1641_0), .o(n_26504) );
na02f06 g753714 ( .a(n_26444), .b(n_26409), .o(n_26540) );
in01s01 g753715 ( .a(n_27198), .o(n_27199) );
in01s01 g753716 ( .a(n_27203), .o(n_27198) );
no02f06 g753717 ( .a(n_27135), .b(n_26772), .o(n_27203) );
in01s01 g753718 ( .a(n_26658), .o(n_26560) );
no02f04 g753719 ( .a(n_26531), .b(FE_OCPN1352_n_26530), .o(n_26658) );
in01s01 g753720 ( .a(n_26532), .o(n_26533) );
na02m06 g753724 ( .a(n_26531), .b(FE_OCPN1352_n_26530), .o(n_26764) );
na02s01 g753725 ( .a(n_26479), .b(n_26506), .o(n_26480) );
no02s01 g753726 ( .a(n_26496), .b(n_26559), .o(n_26624) );
in01s01 g753727 ( .a(n_26557), .o(n_26558) );
no02f04 g753728 ( .a(n_26529), .b(n_26528), .o(n_26557) );
na02f04 g753729 ( .a(n_26529), .b(n_26528), .o(n_26616) );
na02s01 g753730 ( .a(n_26526), .b(n_26525), .o(n_26527) );
in01m04 g753731 ( .a(n_26502), .o(n_26503) );
oa12m06 g753732 ( .a(n_26335), .b(n_26377), .c(FE_OCPN1088_n_25481), .o(n_26502) );
in01m02 g753733 ( .a(n_26614), .o(n_26615) );
no02s03 g753734 ( .a(n_26579), .b(n_26521), .o(n_26614) );
na02m06 TIMEBOOST_cell_1066 ( .a(n_37353), .b(TIMEBOOST_net_147), .o(n_37373) );
in01m02 g753737 ( .a(n_26524), .o(n_26555) );
na02m06 TIMEBOOST_cell_3416 ( .a(n_11599), .b(n_11569), .o(TIMEBOOST_net_999) );
ao12m04 g753739 ( .a(n_26663), .b(n_26478), .c(FE_OCP_RBN6090_n_26322), .o(n_26537) );
oa12s01 g753741 ( .a(n_26414), .b(n_26413), .c(n_26412), .o(n_26477) );
oa22s01 g753744 ( .a(n_27080), .b(n_26893), .c(n_27079), .d(n_26892), .o(n_27134) );
in01s01 g753745 ( .a(n_27132), .o(n_27133) );
oa12s01 g753746 ( .a(n_26711), .b(n_27097), .c(n_26571), .o(n_27132) );
na02m08 g753748 ( .a(n_26448), .b(n_26472), .o(n_26553) );
in01m01 g753749 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_1_), .o(n_28034) );
in01s01 g753752 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_), .o(n_27164) );
na02s02 TIMEBOOST_cell_3415 ( .a(n_27620), .b(TIMEBOOST_net_998), .o(n_27688) );
na02s04 TIMEBOOST_cell_1065 ( .a(n_37357), .b(n_37366), .o(TIMEBOOST_net_147) );
na02m02 g753760 ( .a(n_26409), .b(FE_OCP_RBN1866_n_26407), .o(n_26501) );
no02m02 g753761 ( .a(n_26407), .b(n_26437), .o(n_26500) );
no02s06 g753762 ( .a(n_26458), .b(n_23509), .o(n_26579) );
no02s02 g753763 ( .a(n_26424), .b(n_23564), .o(n_26521) );
na02s03 g753764 ( .a(n_26398), .b(n_23353), .o(n_26448) );
na02m06 g753765 ( .a(FE_OCP_RBN6121_n_26398), .b(n_23509), .o(n_26472) );
no02m02 g753766 ( .a(n_26519), .b(n_26219), .o(n_26520) );
in01s01 g753767 ( .a(n_26497), .o(n_26498) );
na02s04 g753768 ( .a(n_26478), .b(n_26473), .o(n_26497) );
in01s01 g753769 ( .a(n_27108), .o(n_27109) );
na02s01 g753770 ( .a(n_27097), .b(n_26741), .o(n_27108) );
na02s01 g753771 ( .a(n_26412), .b(n_26413), .o(n_26414) );
na02s01 g753772 ( .a(n_26463), .b(n_26518), .o(n_26594) );
na02s01 g753773 ( .a(FE_OCP_RBN6120_n_26398), .b(FE_OCP_RBN3253_n_26276), .o(n_26471) );
no02f04 g753774 ( .a(n_26366), .b(n_26367), .o(n_26447) );
in01s01 g753775 ( .a(n_26495), .o(n_26496) );
na02s04 g753776 ( .a(n_26469), .b(n_26468), .o(n_26495) );
na02s01 TIMEBOOST_cell_3138 ( .a(n_35765), .b(FE_OCP_RBN3290_n_35539), .o(TIMEBOOST_net_860) );
na03s02 TIMEBOOST_cell_8220 ( .a(n_23943), .b(n_23944), .c(n_24498), .o(TIMEBOOST_net_1468) );
in01s02 g753783 ( .a(n_26493), .o(n_26494) );
na02s04 g753784 ( .a(n_26467), .b(n_26372), .o(n_26493) );
in01s02 g753785 ( .a(n_26465), .o(n_26466) );
in01s02 g753786 ( .a(n_26444), .o(n_26465) );
oa12f06 g753787 ( .a(n_26340), .b(n_26368), .c(n_26359), .o(n_26444) );
in01s01 g753788 ( .a(n_27095), .o(n_27096) );
ao12s01 g753789 ( .a(n_26861), .b(n_27067), .c(n_26547), .o(n_27095) );
no02f06 g753790 ( .a(n_27097), .b(n_26642), .o(n_27135) );
na02s01 TIMEBOOST_cell_8661 ( .a(TIMEBOOST_net_2817), .b(n_31682), .o(n_31796) );
oa12s01 g753801 ( .a(n_26371), .b(n_26370), .c(n_26369), .o(n_26439) );
oa12f06 g753802 ( .a(n_26278), .b(n_26425), .c(n_26362), .o(n_26525) );
na02f04 g753803 ( .a(n_26410), .b(n_26374), .o(n_26529) );
oa12s01 g753804 ( .a(n_26427), .b(n_26426), .c(n_26425), .o(n_26491) );
oa22s01 g753805 ( .a(n_27064), .b(n_26900), .c(n_27063), .d(n_26899), .o(n_27107) );
no02m06 g753806 ( .a(n_26376), .b(FE_OCPN1081_n_24819), .o(n_26377) );
no02s01 TIMEBOOST_cell_5606 ( .a(n_31730), .b(n_31599), .o(TIMEBOOST_net_1751) );
no02s01 TIMEBOOST_cell_7039 ( .a(FE_OCP_RBN2966_n_4046), .b(FE_OCP_RBN2962_n_4046), .o(TIMEBOOST_net_2278) );
na02m02 g753809 ( .a(n_26329), .b(n_26245), .o(n_26374) );
na02f04 g753810 ( .a(n_26330), .b(n_26246), .o(n_26410) );
in01m01 g753812 ( .a(n_26409), .o(n_26437) );
na02f02 g753813 ( .a(n_26373), .b(n_23414), .o(n_26409) );
na03f20 TIMEBOOST_cell_8185 ( .a(FE_OCP_RBN2416_n_44722), .b(delay_xor_ln21_unr18_stage7_stallmux_q_6_), .c(FE_RN_2514_0), .o(FE_RN_2515_0) );
no02m06 g753815 ( .a(FE_OCP_RBN6849_n_26358), .b(n_23509), .o(n_26434) );
no02s04 g753819 ( .a(n_26373), .b(n_23353), .o(n_26407) );
no02f02 g753820 ( .a(n_26358), .b(n_23447), .o(n_26406) );
na02m04 g753823 ( .a(n_26320), .b(FE_OCPN1334_n_23467), .o(n_26478) );
na02s02 g753824 ( .a(n_26322), .b(FE_OCPN1334_n_23467), .o(n_26372) );
na02m06 g753825 ( .a(FE_OCP_RBN6090_n_26322), .b(n_23486), .o(n_26467) );
ao12f04 g753826 ( .a(n_26302), .b(n_26224), .c(FE_RN_1793_0), .o(n_26340) );
in01s01 g753827 ( .a(n_26462), .o(n_26463) );
no02f06 g753828 ( .a(n_26429), .b(FE_OCPN5240_n_26428), .o(n_26462) );
na02f06 g753830 ( .a(n_26429), .b(FE_OCPN5240_n_26428), .o(n_26518) );
na02s01 g753831 ( .a(n_26369), .b(n_26370), .o(n_26371) );
no02s01 g753832 ( .a(n_26337), .b(n_26338), .o(n_26413) );
no02s01 g753833 ( .a(n_26326), .b(n_26403), .o(n_26479) );
na02s01 g753834 ( .a(n_26393), .b(n_26461), .o(n_26526) );
na02s01 g753835 ( .a(n_26426), .b(n_26425), .o(n_26427) );
na02f04 g753837 ( .a(n_26303), .b(n_26368), .o(n_26401) );
na02s10 TIMEBOOST_cell_928 ( .a(FE_OCP_RBN5017_n_12026), .b(TIMEBOOST_net_78), .o(n_12106) );
na02s01 TIMEBOOST_cell_946 ( .a(TIMEBOOST_net_87), .b(n_28205), .o(n_28239) );
in01f02 g753841 ( .a(n_26399), .o(n_26400) );
no02f04 g753842 ( .a(n_26300), .b(n_26367), .o(n_26399) );
ao12f02 g753843 ( .a(n_23414), .b(n_26218), .c(n_26078), .o(n_26366) );
in01s01 g753844 ( .a(n_27079), .o(n_27080) );
oa12s01 g753845 ( .a(n_26508), .b(n_27035), .c(n_26549), .o(n_27079) );
na02f06 g753846 ( .a(n_27067), .b(n_26610), .o(n_27097) );
in01s02 g753848 ( .a(n_26424), .o(n_26458) );
na02s02 TIMEBOOST_cell_6295 ( .a(n_10850), .b(n_10831), .o(TIMEBOOST_net_1999) );
oa12s01 g753857 ( .a(n_26295), .b(n_26294), .c(n_26293), .o(n_26365) );
no02s01 TIMEBOOST_cell_1214 ( .a(TIMEBOOST_net_221), .b(n_38128), .o(n_38174) );
oa22s01 g753860 ( .a(n_27035), .b(n_26575), .c(n_27051), .d(n_26574), .o(n_27092) );
na02s06 g753864 ( .a(n_26264), .b(FE_OCPN1081_n_24819), .o(n_26335) );
na02m04 g753866 ( .a(n_26226), .b(FE_OCP_RBN6067_n_26121), .o(n_26304) );
no02s02 g753867 ( .a(n_26302), .b(n_26179), .o(n_26303) );
no02s02 TIMEBOOST_cell_4438 ( .a(TIMEBOOST_net_1309), .b(FE_OCP_RBN4365_n_4692), .o(n_4936) );
in01m04 g753869 ( .a(n_26332), .o(n_26333) );
na02m08 g753870 ( .a(n_26301), .b(n_26258), .o(n_26332) );
na02s01 TIMEBOOST_cell_945 ( .a(n_28204), .b(n_27926), .o(TIMEBOOST_net_87) );
na02s02 g753872 ( .a(n_26253), .b(n_26218), .o(n_26331) );
no02s02 g753873 ( .a(n_26254), .b(n_26283), .o(n_26364) );
no02f04 g753874 ( .a(n_26298), .b(n_26144), .o(n_26300) );
no02f02 g753875 ( .a(n_26251), .b(n_26221), .o(n_26299) );
in01m02 g753876 ( .a(n_26329), .o(n_26330) );
na02m04 g753877 ( .a(n_26298), .b(n_26216), .o(n_26329) );
na02s10 TIMEBOOST_cell_927 ( .a(FE_RN_2101_0), .b(FE_OCPN4935_n_11993), .o(TIMEBOOST_net_78) );
na02m06 g753880 ( .a(n_26319), .b(n_26363), .o(n_26394) );
na02s02 TIMEBOOST_cell_4553 ( .a(n_40534), .b(n_40223), .o(TIMEBOOST_net_1367) );
no02s01 TIMEBOOST_cell_1213 ( .a(n_38076), .b(n_38093), .o(TIMEBOOST_net_221) );
no02f06 TIMEBOOST_cell_3419 ( .a(n_21959), .b(TIMEBOOST_net_1000), .o(n_22030) );
na02m06 TIMEBOOST_cell_5149 ( .a(TIMEBOOST_net_1522), .b(FE_OCP_RBN4179_n_38592), .o(n_38658) );
in01s02 g753885 ( .a(n_26327), .o(n_26328) );
no02m08 g753887 ( .a(n_26297), .b(FE_OCPN1294_n_26296), .o(n_26403) );
no02f02 g753888 ( .a(n_26184), .b(n_24590), .o(n_26337) );
no02s06 g753889 ( .a(n_24591), .b(n_26185), .o(n_26338) );
in01s01 g753890 ( .a(n_26325), .o(n_26326) );
na02f06 g753891 ( .a(n_26297), .b(FE_OCPN1294_n_26296), .o(n_26325) );
no02s01 g753892 ( .a(n_26279), .b(n_26362), .o(n_26426) );
na02f04 g753893 ( .a(n_26361), .b(n_26360), .o(n_26461) );
in01s01 g753894 ( .a(n_26392), .o(n_26393) );
no02f04 g753895 ( .a(n_26361), .b(n_26360), .o(n_26392) );
na02s01 g753896 ( .a(n_26293), .b(n_26294), .o(n_26295) );
in01m02 g753897 ( .a(n_26376), .o(n_26324) );
na02f08 g753899 ( .a(n_26227), .b(n_26157), .o(n_26368) );
in01s06 g753903 ( .a(n_26456), .o(n_26487) );
no03s02 TIMEBOOST_cell_7926 ( .a(TIMEBOOST_net_1673), .b(n_5147), .c(n_5113), .o(TIMEBOOST_net_2594) );
in01m02 g753906 ( .a(n_26421), .o(n_26422) );
no02f08 TIMEBOOST_cell_930 ( .a(n_40992), .b(TIMEBOOST_net_79), .o(n_41030) );
in01s03 g753908 ( .a(n_26292), .o(n_26367) );
in01s01 g753910 ( .a(n_27063), .o(n_27064) );
in01s01 g753911 ( .a(n_27067), .o(n_27063) );
na02f02 TIMEBOOST_cell_6828 ( .a(TIMEBOOST_net_2171), .b(n_16669), .o(TIMEBOOST_net_1764) );
in01s01 g753913 ( .a(FE_OCPN1683_n_27210), .o(n_26323) );
in01s01 g753914 ( .a(n_26291), .o(n_27210) );
in01m02 g753915 ( .a(n_26291), .o(n_26290) );
na03s20 TIMEBOOST_cell_4569 ( .a(n_11774), .b(n_11696), .c(n_45224), .o(TIMEBOOST_net_16) );
na03f06 TIMEBOOST_cell_4617 ( .a(n_23517), .b(n_23556), .c(n_23631), .o(FE_RN_2375_0) );
ao12s01 g753922 ( .a(n_26215), .b(n_26267), .c(n_26214), .o(n_26370) );
oa22m04 g753925 ( .a(FE_OCP_RBN3246_n_26169), .b(n_23447), .c(n_26169), .d(n_23466), .o(n_26322) );
na02m06 TIMEBOOST_cell_4554 ( .a(TIMEBOOST_net_1367), .b(n_40556), .o(n_40578) );
in01s02 g753930 ( .a(n_26265), .o(n_26266) );
no02m04 g753931 ( .a(n_26228), .b(FE_OCPN1336_n_25673), .o(n_26265) );
in01s02 g753932 ( .a(n_26263), .o(n_26264) );
na02m08 g753933 ( .a(n_26228), .b(n_25694), .o(n_26263) );
in01s02 g753934 ( .a(n_26226), .o(n_26227) );
na02m08 g753935 ( .a(n_26130), .b(n_26178), .o(n_26226) );
no02f04 g753936 ( .a(n_26158), .b(n_26206), .o(n_26262) );
na02f06 TIMEBOOST_cell_8650 ( .a(n_26447), .b(n_26175), .o(TIMEBOOST_net_2812) );
na02m04 g753938 ( .a(n_26220), .b(n_26204), .o(n_26225) );
no02s06 g753939 ( .a(n_26196), .b(FE_OCPN3578_n_23354), .o(n_26359) );
na02m04 g753940 ( .a(n_26167), .b(n_26120), .o(n_26224) );
na02s02 TIMEBOOST_cell_4559 ( .a(FE_RN_2695_0), .b(FE_RN_2697_0), .o(TIMEBOOST_net_1370) );
no02f02 g753942 ( .a(n_26152), .b(n_23414), .o(n_26191) );
no02s02 TIMEBOOST_cell_3325 ( .a(TIMEBOOST_net_953), .b(n_31929), .o(n_32130) );
no02m01 g753944 ( .a(n_26173), .b(n_23414), .o(n_26222) );
na02m06 g753946 ( .a(n_26221), .b(n_26220), .o(n_26298) );
na02s06 g753947 ( .a(n_26190), .b(n_23353), .o(n_26301) );
in01s03 g753949 ( .a(n_26219), .o(n_26258) );
no02f08 g753950 ( .a(n_26190), .b(n_23447), .o(n_26219) );
in01s02 g753952 ( .a(n_26319), .o(n_26355) );
na02m08 g753953 ( .a(n_26195), .b(n_23466), .o(n_26319) );
na02s06 g753954 ( .a(n_26194), .b(n_23447), .o(n_26363) );
in01s01 g753955 ( .a(n_26218), .o(n_26283) );
na02m06 g753959 ( .a(n_26188), .b(n_23466), .o(n_26218) );
in01s02 g753961 ( .a(n_26253), .o(n_26254) );
in01s02 g753962 ( .a(n_26217), .o(n_26253) );
no02f06 g753963 ( .a(n_26188), .b(n_23466), .o(n_26217) );
in01s02 g753964 ( .a(n_26251), .o(n_26252) );
na02f04 g753965 ( .a(n_26220), .b(n_26216), .o(n_26251) );
no02s03 g753966 ( .a(n_26198), .b(n_23466), .o(n_26389) );
no02m08 TIMEBOOST_cell_929 ( .a(n_40716), .b(n_40711), .o(TIMEBOOST_net_79) );
in01s02 g753969 ( .a(n_26354), .o(n_26387) );
no02s06 g753970 ( .a(n_26318), .b(FE_OCP_DRV_N6899_FE_OCPN5276_n_23590), .o(n_26354) );
no03s03 TIMEBOOST_cell_4707 ( .a(n_3198), .b(n_2426), .c(n_3205), .o(n_3498) );
in01s01 g753973 ( .a(n_27035), .o(n_27051) );
na02s02 g753974 ( .a(n_26977), .b(n_26612), .o(n_27035) );
no02s01 g753975 ( .a(n_26267), .b(n_26214), .o(n_26215) );
na02s01 g753976 ( .a(n_26200), .b(FE_OCP_RBN6066_n_26081), .o(n_26250) );
na02s01 g753977 ( .a(n_26174), .b(n_26048), .o(n_26213) );
no02s01 g753978 ( .a(n_26212), .b(n_26186), .o(n_26294) );
in01s01 g753979 ( .a(n_26278), .o(n_26279) );
na02m04 g753980 ( .a(n_26249), .b(n_26248), .o(n_26278) );
no02f04 g753981 ( .a(n_26249), .b(n_26248), .o(n_26362) );
na02s01 g753983 ( .a(n_26201), .b(n_26110), .o(n_26247) );
no03f08 TIMEBOOST_cell_3576 ( .a(n_29659), .b(n_29686), .c(n_29640), .o(n_29766) );
na03m02 TIMEBOOST_cell_8193 ( .a(n_22984), .b(n_23326), .c(n_23246), .o(n_23327) );
in01s01 g753987 ( .a(n_27033), .o(n_27034) );
na02m01 TIMEBOOST_cell_3350 ( .a(FE_OCPN900_n_16923), .b(n_17139), .o(TIMEBOOST_net_966) );
na02s01 TIMEBOOST_cell_1193 ( .a(n_36855), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_), .o(TIMEBOOST_net_211) );
in01s01 g753990 ( .a(n_27031), .o(n_27032) );
no02s02 TIMEBOOST_cell_3418 ( .a(n_21520), .b(n_21480), .o(TIMEBOOST_net_1000) );
na02f04 TIMEBOOST_cell_5542 ( .a(n_36628), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_1719) );
in01s02 g753993 ( .a(n_26184), .o(n_26185) );
na02s01 TIMEBOOST_cell_5285 ( .a(TIMEBOOST_net_1590), .b(n_20708), .o(n_20836) );
oa22s01 g754000 ( .a(n_26974), .b(n_26903), .c(n_26949), .d(n_26904), .o(n_27016) );
oa22s01 g754001 ( .a(n_26978), .b(n_26901), .c(n_26950), .d(n_26902), .o(n_27015) );
oa12s01 g754002 ( .a(n_26953), .b(n_26952), .c(n_26951), .o(n_27002) );
no02m08 g754006 ( .a(n_26112), .b(n_25672), .o(n_26228) );
na02s04 g754007 ( .a(n_26129), .b(n_26083), .o(n_26131) );
no02f04 TIMEBOOST_cell_5541 ( .a(TIMEBOOST_net_1718), .b(n_30988), .o(n_31265) );
no02m06 g754011 ( .a(n_26129), .b(n_26128), .o(n_26130) );
no02s04 g754012 ( .a(n_26129), .b(n_26128), .o(n_26158) );
no02f08 TIMEBOOST_cell_7813 ( .a(TIMEBOOST_net_2537), .b(n_24657), .o(n_24839) );
no02f02 g754014 ( .a(FE_OCP_RBN3173_n_26178), .b(n_26136), .o(n_26181) );
no02m08 TIMEBOOST_cell_4190 ( .a(TIMEBOOST_net_1185), .b(FE_OCP_RBN1175_n_27593), .o(n_27661) );
no02s06 TIMEBOOST_cell_4430 ( .a(TIMEBOOST_net_1305), .b(n_46959), .o(TIMEBOOST_net_1129) );
no02s04 TIMEBOOST_cell_2131 ( .a(n_10141), .b(n_9966), .o(TIMEBOOST_net_680) );
no02s02 g754019 ( .a(n_26179), .b(n_26156), .o(n_26208) );
in01m02 g754020 ( .a(n_26206), .o(n_26207) );
na02f04 g754021 ( .a(n_26178), .b(FE_OCP_RBN6068_n_26121), .o(n_26206) );
na02s04 g754022 ( .a(n_26087), .b(n_23466), .o(n_26216) );
no02s06 g754024 ( .a(n_26176), .b(n_23398), .o(n_26277) );
no02s01 TIMEBOOST_cell_5666 ( .a(FE_OCP_RBN6175_n_16923), .b(FE_OCP_RBN4396_n_16146), .o(TIMEBOOST_net_1781) );
no02f06 TIMEBOOST_cell_3349 ( .a(n_27540), .b(TIMEBOOST_net_965), .o(n_27589) );
na02s01 g754027 ( .a(n_26952), .b(n_26951), .o(n_26953) );
in01s01 g754028 ( .a(n_26976), .o(n_26977) );
no02f06 g754029 ( .a(n_26911), .b(n_26484), .o(n_26976) );
na02m08 TIMEBOOST_cell_3417 ( .a(TIMEBOOST_net_999), .b(n_11603), .o(n_11777) );
no02f04 g754033 ( .a(n_26085), .b(n_24432), .o(n_26186) );
no02m08 g754034 ( .a(n_26086), .b(n_24433), .o(n_26212) );
in01f02 g754035 ( .a(n_26153), .o(n_26154) );
in01s02 g754037 ( .a(n_26245), .o(n_26246) );
na02s03 g754038 ( .a(n_26204), .b(n_26149), .o(n_26245) );
no02s01 TIMEBOOST_cell_8507 ( .a(TIMEBOOST_net_2740), .b(n_37827), .o(n_37878) );
in01m04 g754041 ( .a(n_26221), .o(n_26306) );
na02m08 g754042 ( .a(n_26089), .b(n_26101), .o(n_26221) );
in01s01 g754045 ( .a(n_26174), .o(n_26201) );
in01s02 g754046 ( .a(n_26152), .o(n_26174) );
no02f08 TIMEBOOST_cell_6714 ( .a(TIMEBOOST_net_2114), .b(n_38719), .o(n_38743) );
in01m04 g754056 ( .a(n_26171), .o(n_26200) );
oa22m04 g754062 ( .a(n_26040), .b(n_25720), .c(n_26041), .d(n_25719), .o(n_26169) );
in01s01 g754064 ( .a(n_26198), .o(n_26240) );
oa22m04 g754065 ( .a(n_26081), .b(n_23447), .c(FE_OCP_RBN6065_n_26081), .d(n_23398), .o(n_26198) );
no02s02 TIMEBOOST_cell_3106 ( .a(n_9696), .b(n_9729), .o(TIMEBOOST_net_844) );
na02s06 TIMEBOOST_cell_4417 ( .a(n_20466), .b(n_20429), .o(TIMEBOOST_net_1299) );
no02s01 TIMEBOOST_cell_4419 ( .a(FE_OFN748_n_22641), .b(n_23398), .o(TIMEBOOST_net_1300) );
in01m02 g754069 ( .a(n_26318), .o(n_26272) );
na02m04 TIMEBOOST_cell_4220 ( .a(TIMEBOOST_net_1200), .b(n_12517), .o(n_12565) );
oa12s01 g754071 ( .a(n_26092), .b(n_26091), .c(n_26090), .o(n_26150) );
in01m04 g754073 ( .a(n_26167), .o(n_26196) );
no02s02 TIMEBOOST_cell_4558 ( .a(TIMEBOOST_net_1369), .b(FE_OCP_RBN1026_n_17417), .o(FE_RN_344_0) );
in01s04 g754075 ( .a(n_26194), .o(n_26195) );
na02s08 TIMEBOOST_cell_8755 ( .a(TIMEBOOST_net_2864), .b(n_14402), .o(n_14535) );
no02f08 TIMEBOOST_cell_6713 ( .a(FE_OFN5092_delay_sub_ln23_0_unr25_stage9_stallmux_q), .b(n_38703), .o(TIMEBOOST_net_2114) );
na02s02 TIMEBOOST_cell_4555 ( .a(n_17331), .b(FE_RN_340_0), .o(TIMEBOOST_net_1368) );
in01s02 g754082 ( .a(n_26129), .o(n_26104) );
na02m08 g754083 ( .a(n_26068), .b(FE_OCP_RBN1035_FE_RN_557_0), .o(n_26129) );
no02s10 TIMEBOOST_cell_4213 ( .a(n_32870), .b(n_32717), .o(TIMEBOOST_net_1197) );
no02f04 g754085 ( .a(n_26060), .b(n_26015), .o(n_26124) );
na02s06 TIMEBOOST_cell_4418 ( .a(TIMEBOOST_net_1299), .b(n_20694), .o(n_20777) );
no02s01 TIMEBOOST_cell_8499 ( .a(TIMEBOOST_net_2736), .b(n_37725), .o(n_37773) );
na02m06 g754088 ( .a(n_26027), .b(n_26100), .o(n_26101) );
na02f04 TIMEBOOST_cell_3315 ( .a(TIMEBOOST_net_948), .b(n_39803), .o(n_39895) );
no02m02 g754090 ( .a(n_26097), .b(n_23466), .o(n_26156) );
na02m08 g754092 ( .a(n_26098), .b(n_23317), .o(n_26178) );
no02f08 g754094 ( .a(n_26098), .b(n_23317), .o(n_26121) );
in01s02 g754095 ( .a(n_26120), .o(n_26179) );
na02m04 g754096 ( .a(n_26097), .b(n_23339), .o(n_26120) );
na02s03 g754097 ( .a(n_26079), .b(n_23466), .o(n_26149) );
na02s06 g754098 ( .a(n_26146), .b(FE_OCPN1334_n_23467), .o(n_26147) );
no02s02 TIMEBOOST_cell_6259 ( .a(n_4860), .b(n_4477), .o(TIMEBOOST_net_1981) );
no02s20 TIMEBOOST_cell_8468 ( .a(n_32399), .b(FE_OCP_RBN6527_n_44962), .o(TIMEBOOST_net_2721) );
no02s01 TIMEBOOST_cell_3123 ( .a(TIMEBOOST_net_852), .b(FE_OCP_RBN5947_n_14982), .o(n_15297) );
na02s06 g754102 ( .a(n_25999), .b(FE_OFN748_n_22641), .o(n_26032) );
na02s06 g754103 ( .a(n_26039), .b(n_23353), .o(n_26175) );
in01s01 g754104 ( .a(n_26204), .o(n_26144) );
na02f06 g754105 ( .a(n_26118), .b(n_23353), .o(n_26204) );
na02m06 TIMEBOOST_cell_3131 ( .a(TIMEBOOST_net_856), .b(n_34953), .o(n_35077) );
no02m08 TIMEBOOST_cell_5429 ( .a(TIMEBOOST_net_1662), .b(n_5610), .o(n_5802) );
no02s04 TIMEBOOST_cell_6944 ( .a(TIMEBOOST_net_2230), .b(n_29329), .o(n_29425) );
na02f10 TIMEBOOST_cell_5195 ( .a(n_34570), .b(TIMEBOOST_net_1545), .o(n_34440) );
na02s02 TIMEBOOST_cell_5545 ( .a(TIMEBOOST_net_1720), .b(n_6136), .o(n_6248) );
in01s01 g754111 ( .a(n_26978), .o(n_26950) );
in01s01 g754112 ( .a(n_26911), .o(n_26978) );
na02f04 TIMEBOOST_cell_1088 ( .a(n_37369), .b(TIMEBOOST_net_158), .o(n_37418) );
na02f04 g754114 ( .a(n_26021), .b(n_26090), .o(n_26369) );
no02s01 g754115 ( .a(n_26114), .b(FE_OCP_RBN6029_n_25928), .o(n_26116) );
na02s01 g754116 ( .a(n_26114), .b(FE_OCP_RBN6029_n_25928), .o(n_26115) );
na02s01 g754117 ( .a(n_26091), .b(n_26090), .o(n_26092) );
in01s02 g754118 ( .a(n_26142), .o(n_26143) );
in01m02 g754119 ( .a(n_26112), .o(n_26142) );
no02s01 TIMEBOOST_cell_1048 ( .a(n_23276), .b(TIMEBOOST_net_138), .o(n_23357) );
in01f02 g754121 ( .a(n_26061), .o(n_26062) );
na02f04 g754122 ( .a(n_25947), .b(FE_OCP_RBN1036_FE_RN_557_0), .o(n_26061) );
na02s01 TIMEBOOST_cell_5398 ( .a(n_3884), .b(n_3885), .o(TIMEBOOST_net_1647) );
oa12m06 g754125 ( .a(FE_OCPN1390_n_26054), .b(n_26055), .c(n_26026), .o(n_26089) );
in01s01 g754126 ( .a(n_26974), .o(n_26949) );
na02s01 g754127 ( .a(n_26834), .b(n_26382), .o(n_26974) );
ao12s01 g754128 ( .a(n_26812), .b(n_26947), .c(n_26866), .o(n_26952) );
oa12s01 g754129 ( .a(n_26051), .b(n_25984), .c(n_24219), .o(n_26111) );
in01f02 g754130 ( .a(n_26176), .o(n_26139) );
in01s01 TIMEBOOST_cell_8891 ( .a(TIMEBOOST_net_2934), .o(TIMEBOOST_net_2935) );
na02m04 TIMEBOOST_cell_6896 ( .a(TIMEBOOST_net_2206), .b(n_29479), .o(FE_RN_317_0) );
in01s03 g754134 ( .a(n_26085), .o(n_26086) );
oa12s01 g754136 ( .a(n_26948), .b(n_26947), .c(n_26946), .o(n_27001) );
in01s02 g754138 ( .a(n_26069), .o(n_26029) );
no02f08 g754139 ( .a(n_25966), .b(n_25588), .o(n_26069) );
in01m02 g754140 ( .a(n_26068), .o(n_26028) );
no02f08 g754141 ( .a(n_26004), .b(n_26003), .o(n_26068) );
in01f02 g754142 ( .a(n_26059), .o(n_26060) );
in01f03 g754143 ( .a(n_26027), .o(n_26059) );
no02f06 g754144 ( .a(n_25972), .b(n_26002), .o(n_26027) );
na02m02 g754146 ( .a(n_25920), .b(n_23259), .o(n_25947) );
na02m02 TIMEBOOST_cell_6895 ( .a(n_29480), .b(FE_RN_315_0), .o(TIMEBOOST_net_2206) );
in01f02 g754148 ( .a(n_26057), .o(n_26058) );
no02f06 g754149 ( .a(n_26026), .b(n_26002), .o(n_26057) );
na02f10 TIMEBOOST_cell_3111 ( .a(n_3456), .b(TIMEBOOST_net_846), .o(n_3564) );
na02f02 g754152 ( .a(n_25938), .b(n_23254), .o(n_25976) );
na02m06 g754153 ( .a(n_25982), .b(FE_OFN747_n_22641), .o(n_26100) );
na02s04 g754154 ( .a(n_25986), .b(n_23398), .o(n_26025) );
na02s01 g754155 ( .a(n_26947), .b(n_26452), .o(n_26834) );
in01s01 g754156 ( .a(n_26293), .o(n_26051) );
no02m06 g754157 ( .a(n_25983), .b(n_24218), .o(n_26293) );
na02s01 g754158 ( .a(n_26947), .b(n_26946), .o(n_26948) );
no02s01 TIMEBOOST_cell_1047 ( .a(n_22695), .b(n_22700), .o(TIMEBOOST_net_138) );
ao12s04 g754160 ( .a(n_25540), .b(n_25974), .c(FE_OCPN5111_n_25973), .o(n_26000) );
na02f04 g754161 ( .a(n_25975), .b(n_25506), .o(n_26022) );
in01m02 g754162 ( .a(n_26083), .o(n_26084) );
no02s20 TIMEBOOST_cell_848 ( .a(TIMEBOOST_net_38), .b(n_17245), .o(n_17561) );
no02f04 g754165 ( .a(n_25969), .b(n_26003), .o(n_26049) );
na02s02 g754166 ( .a(n_26076), .b(n_26036), .o(n_26138) );
no03s10 TIMEBOOST_cell_3438 ( .a(FE_OCPN1651_n_11918), .b(n_11919), .c(n_11718), .o(TIMEBOOST_net_55) );
no02s02 TIMEBOOST_cell_5517 ( .a(TIMEBOOST_net_1706), .b(n_36483), .o(TIMEBOOST_net_1176) );
in01s01 g754169 ( .a(n_26021), .o(n_26091) );
no02m06 TIMEBOOST_cell_8648 ( .a(n_39579), .b(n_45840), .o(TIMEBOOST_net_2811) );
in01s01 g754171 ( .a(n_26048), .o(n_26110) );
in01s01 g754174 ( .a(n_26020), .o(n_26048) );
in01s02 g754175 ( .a(n_26020), .o(n_26019) );
no03f08 TIMEBOOST_cell_8064 ( .a(FE_OCP_RBN5327_FE_RN_2034_0), .b(n_19969), .c(n_20093), .o(TIMEBOOST_net_2663) );
in01s01 g754181 ( .a(n_25999), .o(n_27117) );
in01f04 g754182 ( .a(n_25999), .o(n_25998) );
in01s01 g754185 ( .a(n_26114), .o(n_26107) );
in01s01 g754186 ( .a(n_26045), .o(n_26114) );
in01s03 g754187 ( .a(n_26045), .o(n_26044) );
oa22m02 g754192 ( .a(n_25900), .b(n_25616), .c(FE_OCP_RBN6013_n_25900), .d(n_25615), .o(n_25997) );
oa12s08 g754197 ( .a(n_25645), .b(n_26016), .c(n_25614), .o(n_26042) );
in01m02 g754198 ( .a(n_26040), .o(n_26041) );
oa12s02 g754199 ( .a(n_25618), .b(n_26016), .c(n_25749), .o(n_26040) );
no02m08 TIMEBOOST_cell_924 ( .a(TIMEBOOST_net_76), .b(FE_RN_1640_0), .o(n_32740) );
in01s02 g754202 ( .a(n_26118), .o(n_26079) );
no02s01 TIMEBOOST_cell_4465 ( .a(n_43692), .b(n_43412), .o(TIMEBOOST_net_1323) );
oa12s01 g754204 ( .a(n_26745), .b(n_26744), .c(n_26743), .o(n_26796) );
oa12s01 g754205 ( .a(n_26910), .b(n_26909), .c(n_26908), .o(n_26973) );
in01f02 g754206 ( .a(n_26077), .o(n_26078) );
in01f02 g754207 ( .a(n_26039), .o(n_26077) );
na02f04 g754209 ( .a(n_25974), .b(FE_OCPN5111_n_25973), .o(n_25975) );
in01s02 g754211 ( .a(n_25972), .o(n_25994) );
na02f08 g754212 ( .a(n_25939), .b(n_25919), .o(n_25972) );
na02f10 TIMEBOOST_cell_3257 ( .a(n_43528), .b(TIMEBOOST_net_919), .o(n_43638) );
in01f01 g754214 ( .a(n_26004), .o(n_25971) );
no02f04 g754215 ( .a(FE_OCP_RBN1851_n_25898), .b(n_23254), .o(n_26004) );
no02f08 TIMEBOOST_cell_4548 ( .a(FE_RN_154_0), .b(TIMEBOOST_net_1364), .o(n_16646) );
in01s01 g754217 ( .a(n_26136), .o(n_26076) );
in01s01 TIMEBOOST_cell_8908 ( .a(n_1354), .o(TIMEBOOST_net_2952) );
no02m04 g754219 ( .a(n_26037), .b(n_23398), .o(n_26136) );
na02f04 TIMEBOOST_cell_4563 ( .a(n_36505), .b(FE_OCPN1940_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_1372) );
no02s06 g754221 ( .a(n_25916), .b(n_25824), .o(n_26003) );
no02s10 TIMEBOOST_cell_847 ( .a(n_17244), .b(n_17197), .o(TIMEBOOST_net_38) );
no02f02 g754223 ( .a(n_25917), .b(FE_OFN745_n_22641), .o(n_25969) );
no02f04 TIMEBOOST_cell_7762 ( .a(FE_OCP_RBN1139_n_19270), .b(n_19694), .o(TIMEBOOST_net_2512) );
na02s02 g754225 ( .a(n_26037), .b(n_23466), .o(n_26036) );
no02s02 TIMEBOOST_cell_5478 ( .a(n_10944), .b(n_44498), .o(TIMEBOOST_net_1687) );
no02s06 g754227 ( .a(n_25912), .b(n_25829), .o(n_26002) );
no02s02 g754228 ( .a(n_25898), .b(n_23254), .o(n_25922) );
no02f04 g754229 ( .a(n_25931), .b(n_23254), .o(n_26128) );
no02s06 g754230 ( .a(n_46962), .b(n_23259), .o(n_25968) );
in01s02 g754231 ( .a(n_26014), .o(n_26015) );
in01s02 g754232 ( .a(n_26026), .o(n_26014) );
na02s01 g754234 ( .a(n_26744), .b(n_26743), .o(n_26745) );
na02s01 g754235 ( .a(n_26909), .b(n_26908), .o(n_26910) );
na02s03 g754236 ( .a(n_25955), .b(n_25747), .o(n_26013) );
no02s06 TIMEBOOST_cell_923 ( .a(n_32643), .b(FE_OCP_RBN6533_n_32436), .o(TIMEBOOST_net_76) );
in01m04 g754238 ( .a(n_25966), .o(n_25967) );
no02m08 g754239 ( .a(n_25940), .b(n_25565), .o(n_25966) );
na02f04 g754241 ( .a(n_25939), .b(n_25881), .o(n_25964) );
in01s01 g754246 ( .a(n_25962), .o(n_25963) );
in01s01 g754247 ( .a(n_25938), .o(n_25962) );
in01s02 g754248 ( .a(n_25938), .o(n_25937) );
in01s01 g754251 ( .a(n_26010), .o(n_26011) );
in01f02 g754252 ( .a(n_25986), .o(n_26010) );
oa22f04 g754254 ( .a(FE_OCP_RBN6018_n_25895), .b(n_25586), .c(n_25895), .d(n_25585), .o(n_25986) );
in01s01 g754255 ( .a(n_25983), .o(n_25984) );
in01f04 g754257 ( .a(n_25982), .o(n_26055) );
in01s01 g754259 ( .a(n_26795), .o(n_26947) );
na02s02 TIMEBOOST_cell_3314 ( .a(n_40202), .b(n_39894), .o(TIMEBOOST_net_948) );
oa12s01 g754261 ( .a(n_26945), .b(n_26944), .c(n_26943), .o(n_27000) );
in01s02 g754264 ( .a(n_25919), .o(n_25935) );
na02f08 g754265 ( .a(n_25874), .b(FE_OFN747_n_22641), .o(n_25919) );
na02s02 g754266 ( .a(n_25847), .b(n_23254), .o(n_25881) );
na02s01 g754269 ( .a(n_26944), .b(n_26943), .o(n_26945) );
in01m04 g754270 ( .a(n_25940), .o(n_25974) );
in01s04 g754271 ( .a(n_25940), .o(n_25918) );
ao12s01 g754273 ( .a(n_26343), .b(n_26646), .c(n_26690), .o(n_26744) );
no02s01 g754274 ( .a(n_26689), .b(n_26384), .o(n_26909) );
in01s01 g754276 ( .a(n_27217), .o(n_25980) );
in01s01 g754277 ( .a(n_25934), .o(n_27217) );
in01m02 g754278 ( .a(n_25934), .o(n_25933) );
in01s02 g754280 ( .a(n_25931), .o(n_25932) );
no02s01 TIMEBOOST_cell_4545 ( .a(n_21254), .b(n_21295), .o(TIMEBOOST_net_1363) );
in01f01 g754282 ( .a(n_25916), .o(n_25917) );
na02f04 g754283 ( .a(n_25832), .b(n_45532), .o(n_25916) );
in01s01 g754286 ( .a(n_25915), .o(n_27170) );
in01s03 g754287 ( .a(n_25915), .o(n_25914) );
in01s01 g754289 ( .a(n_26037), .o(n_26009) );
no03s03 TIMEBOOST_cell_4585 ( .a(n_6716), .b(n_6745), .c(n_6710), .o(n_6711) );
in01f04 g754295 ( .a(n_25902), .o(n_25903) );
no02m06 g754296 ( .a(n_25828), .b(n_25482), .o(n_25902) );
na02f08 g754301 ( .a(n_25876), .b(n_25854), .o(n_25928) );
na02m08 g754303 ( .a(n_25875), .b(n_25503), .o(n_25925) );
oa12m02 g754305 ( .a(n_25536), .b(n_25819), .c(FE_OCP_RBN4341_n_25500), .o(n_25900) );
in01s01 g754306 ( .a(n_26016), .o(n_25956) );
no02s01 TIMEBOOST_cell_8700 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_1_), .b(n_6669), .o(TIMEBOOST_net_2837) );
in01s02 g754308 ( .a(n_25954), .o(n_25955) );
ao12s03 g754309 ( .a(n_25723), .b(n_25870), .c(n_25751), .o(n_25954) );
na02s06 TIMEBOOST_cell_8688 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_), .o(TIMEBOOST_net_2831) );
no02m04 g754316 ( .a(n_25763), .b(n_25831), .o(n_25793) );
na02m04 g754317 ( .a(n_25889), .b(n_23317), .o(n_25911) );
na03f80 TIMEBOOST_cell_4584 ( .a(n_27868), .b(n_27802), .c(TIMEBOOST_net_1006), .o(n_27919) );
na02f02 g754320 ( .a(n_25817), .b(FE_OFN748_n_22641), .o(n_25856) );
no02s01 TIMEBOOST_cell_7041 ( .a(n_4606), .b(FE_OCP_RBN2964_n_4046), .o(TIMEBOOST_net_2279) );
na02f02 g754322 ( .a(n_45533), .b(n_25831), .o(n_25832) );
no02f06 TIMEBOOST_cell_8513 ( .a(TIMEBOOST_net_2743), .b(n_29302), .o(n_29421) );
na02m08 g754325 ( .a(n_25813), .b(n_25479), .o(n_25855) );
no02m04 g754326 ( .a(n_25783), .b(n_25445), .o(n_25828) );
na02f06 g754327 ( .a(n_25843), .b(n_25537), .o(n_25876) );
na02s04 g754328 ( .a(n_25812), .b(n_25538), .o(n_25854) );
na02s04 g754329 ( .a(n_25843), .b(n_25502), .o(n_25875) );
no02f06 g754331 ( .a(FE_OCP_RBN3105_n_25819), .b(n_25647), .o(n_25895) );
na03m08 TIMEBOOST_cell_4853 ( .a(FE_OCP_RBN6237_n_11853), .b(n_11729), .c(n_11848), .o(n_12027) );
in01s01 g754336 ( .a(n_26688), .o(n_26689) );
na02m06 g754337 ( .a(n_26646), .b(n_26312), .o(n_26688) );
oa12s01 g754338 ( .a(n_26613), .b(FE_OCP_RBN6860_n_26160), .c(n_26855), .o(n_26944) );
na02m08 g754346 ( .a(n_25821), .b(n_25788), .o(n_25893) );
no02f08 g754348 ( .a(n_25764), .b(n_25416), .o(n_25849) );
oa12s01 g754351 ( .a(n_26942), .b(n_26941), .c(n_26940), .o(n_26999) );
in01s02 g754352 ( .a(n_25890), .o(n_25891) );
in01s02 g754353 ( .a(n_25874), .o(n_25890) );
na02f03 TIMEBOOST_cell_5171 ( .a(n_34196), .b(TIMEBOOST_net_1533), .o(FE_RN_706_0) );
no02m06 TIMEBOOST_cell_5381 ( .a(TIMEBOOST_net_1638), .b(n_35444), .o(n_35468) );
no02f10 TIMEBOOST_cell_3009 ( .a(TIMEBOOST_net_795), .b(n_23949), .o(n_24072) );
na02s01 g754358 ( .a(n_26941), .b(n_26940), .o(n_26942) );
no02s01 g754360 ( .a(n_25777), .b(n_25822), .o(n_25823) );
na02m06 g754361 ( .a(n_25758), .b(n_25447), .o(n_25788) );
na02m08 g754362 ( .a(n_25759), .b(n_25446), .o(n_25821) );
no02f08 g754363 ( .a(n_25733), .b(n_25415), .o(n_25764) );
ao12f01 g754365 ( .a(n_25782), .b(n_25704), .c(n_25561), .o(n_25819) );
in01m02 g754366 ( .a(n_25845), .o(n_25846) );
oa12m06 g754367 ( .a(n_25454), .b(n_25727), .c(n_25425), .o(n_25845) );
ao12m06 g754369 ( .a(n_25422), .b(FE_OCP_RBN5996_n_25732), .c(n_25760), .o(n_25785) );
na02m06 g754370 ( .a(n_25761), .b(n_25389), .o(n_25818) );
in01s01 g754371 ( .a(n_26646), .o(n_26613) );
no02m06 g754372 ( .a(n_26941), .b(n_26232), .o(n_26646) );
na02s02 TIMEBOOST_cell_6640 ( .a(TIMEBOOST_net_2077), .b(n_18665), .o(n_18666) );
ao22f02 g754381 ( .a(n_25732), .b(n_25488), .c(FE_OCP_RBN5998_n_25732), .d(n_25487), .o(n_25817) );
na02f08 TIMEBOOST_cell_6726 ( .a(TIMEBOOST_net_2120), .b(n_19700), .o(n_19774) );
in01m04 g754388 ( .a(n_25783), .o(n_25813) );
na02s01 TIMEBOOST_cell_6754 ( .a(TIMEBOOST_net_2134), .b(n_39261), .o(n_39342) );
in01s01 g754390 ( .a(n_25869), .o(n_25870) );
in01s02 g754391 ( .a(n_25843), .o(n_25869) );
in01f04 g754392 ( .a(n_25812), .o(n_25843) );
ao12m04 g754394 ( .a(n_25782), .b(n_25704), .c(n_25504), .o(n_25812) );
in01s01 g754397 ( .a(n_25781), .o(n_25810) );
in01s01 g754398 ( .a(n_25763), .o(n_25781) );
in01s02 g754399 ( .a(n_25763), .o(n_25762) );
in01s01 g754405 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_3_), .o(n_27988) );
na02s04 TIMEBOOST_cell_5636 ( .a(n_27595), .b(n_27396), .o(TIMEBOOST_net_1766) );
no02f04 TIMEBOOST_cell_4546 ( .a(TIMEBOOST_net_1363), .b(n_21699), .o(n_21754) );
na02m04 g754409 ( .a(FE_OCP_RBN5997_n_25732), .b(n_25760), .o(n_25761) );
no02f08 g754412 ( .a(n_25677), .b(n_25378), .o(n_25734) );
na02s02 TIMEBOOST_cell_5619 ( .a(TIMEBOOST_net_1757), .b(n_6276), .o(n_6419) );
in01m06 g754414 ( .a(n_25758), .o(n_25759) );
in01m06 g754415 ( .a(n_25733), .o(n_25758) );
no02f10 g754416 ( .a(n_25704), .b(n_25453), .o(n_25733) );
no02f10 TIMEBOOST_cell_3007 ( .a(FE_RN_2382_0), .b(TIMEBOOST_net_794), .o(n_23949) );
ao12m04 g754419 ( .a(n_26386), .b(n_26420), .c(FE_OCP_RBN6096_n_26160), .o(n_26941) );
in01s01 g754424 ( .a(n_25757), .o(n_25777) );
in01s01 g754425 ( .a(n_25731), .o(n_25757) );
in01f04 g754426 ( .a(n_25731), .o(n_25730) );
no02m08 g754432 ( .a(n_25726), .b(n_25457), .o(n_25727) );
no02f02 g754435 ( .a(n_25635), .b(n_25401), .o(n_25656) );
no02f10 g754439 ( .a(n_25654), .b(n_25353), .o(n_25704) );
ao12m10 g754444 ( .a(n_25457), .b(n_25631), .c(n_25458), .o(n_25732) );
oa12m04 g754445 ( .a(n_25397), .b(FE_OCP_RBN1005_n_25545), .c(n_25331), .o(n_25655) );
ao12m02 g754446 ( .a(n_25239), .b(FE_OCP_RBN1004_n_25545), .c(n_25398), .o(n_25634) );
in01m04 g754447 ( .a(n_25676), .o(n_25677) );
oa22s01 g754450 ( .a(n_25653), .b(n_25427), .c(n_25675), .d(n_25428), .o(n_27416) );
oa12s01 g754451 ( .a(n_26939), .b(n_26938), .c(n_26937), .o(n_26998) );
in01s01 g754453 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_2_), .o(n_27050) );
no02f02 g754456 ( .a(n_25545), .b(n_25272), .o(n_25635) );
na02s01 g754457 ( .a(n_26814), .b(n_26816), .o(n_26817) );
na02s01 g754458 ( .a(n_26831), .b(n_26832), .o(n_26833) );
na02s01 g754459 ( .a(n_26773), .b(n_26639), .o(n_26815) );
in01s01 g754460 ( .a(n_26869), .o(n_26870) );
na02s01 g754461 ( .a(n_26831), .b(n_26816), .o(n_26869) );
na02f04 g754462 ( .a(FE_OCP_RBN2976_n_25295), .b(n_25567), .o(n_25633) );
no02f02 g754463 ( .a(n_25601), .b(n_25295), .o(n_25602) );
na02f10 g754464 ( .a(n_25601), .b(n_25321), .o(n_25654) );
na02m04 g754465 ( .a(n_26938), .b(n_26419), .o(n_26420) );
oa12s01 g754466 ( .a(n_26793), .b(n_26713), .c(n_26541), .o(n_26794) );
na02s01 g754467 ( .a(n_26938), .b(n_26937), .o(n_26939) );
na02s04 TIMEBOOST_cell_1087 ( .a(n_37368), .b(n_37143), .o(TIMEBOOST_net_158) );
in01s01 g754470 ( .a(n_25789), .o(n_25822) );
ao12s01 g754471 ( .a(n_25630), .b(n_25629), .c(n_25628), .o(n_25789) );
oa12f04 g754472 ( .a(n_25323), .b(FE_OCP_RBN5942_n_25544), .c(n_25231), .o(n_25632) );
ao12s04 g754473 ( .a(n_25292), .b(n_25544), .c(n_25206), .o(n_25600) );
ao12s01 g754475 ( .a(n_25519), .b(n_25518), .c(n_25517), .o(n_25598) );
in01s01 g754476 ( .a(n_26935), .o(n_26936) );
oa22s01 g754477 ( .a(n_26907), .b(FE_OCP_RBN4435_n_26160), .c(n_26350), .d(n_26896), .o(n_26935) );
ao12s02 g754478 ( .a(n_26381), .b(n_26418), .c(FE_OCP_RBN6857_n_26160), .o(n_26514) );
na02s01 g754479 ( .a(n_26686), .b(n_26708), .o(n_26742) );
na02s01 g754480 ( .a(n_26352), .b(FE_OCP_RBN4434_n_26160), .o(n_26831) );
no02s03 g754481 ( .a(n_26314), .b(n_26419), .o(n_26386) );
na02s01 g754482 ( .a(n_26351), .b(FE_OCP_RBN4433_n_26160), .o(n_26816) );
in01s01 g754483 ( .a(n_25675), .o(n_25653) );
in01m04 g754484 ( .a(n_25631), .o(n_25675) );
in01m08 g754485 ( .a(FE_OCP_RBN1005_n_25545), .o(n_25631) );
oa12f06 g754488 ( .a(n_25277), .b(n_25433), .c(n_25243), .o(n_25545) );
no02s01 g754489 ( .a(n_25629), .b(n_25628), .o(n_25630) );
no02s01 g754490 ( .a(n_25518), .b(n_25517), .o(n_25519) );
oa12s02 g754491 ( .a(n_26383), .b(n_26349), .c(n_26160), .o(n_26454) );
no02s02 TIMEBOOST_cell_5354 ( .a(n_5009), .b(n_5021), .o(TIMEBOOST_net_1625) );
in01s01 g754493 ( .a(n_26772), .o(n_26773) );
na02s02 g754494 ( .a(n_26687), .b(n_26741), .o(n_26772) );
no02s02 g754495 ( .a(n_26714), .b(n_26644), .o(n_26715) );
in01s01 g754496 ( .a(n_26905), .o(n_26906) );
ao12s01 g754497 ( .a(n_26868), .b(n_26740), .c(FE_OCP_RBN4435_n_26160), .o(n_26905) );
no02m04 g754498 ( .a(n_26313), .b(n_26193), .o(n_26938) );
oa12s01 g754500 ( .a(n_25516), .b(n_25515), .c(n_25514), .o(n_25595) );
in01f02 g754501 ( .a(n_25601), .o(n_25567) );
oa12s01 g754503 ( .a(n_26934), .b(n_26933), .c(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_26997) );
oa12s01 g754504 ( .a(n_26932), .b(n_26931), .c(n_26930), .o(n_26996) );
na02s01 g754505 ( .a(n_26933), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_26934) );
na02s02 g754506 ( .a(n_26452), .b(n_26415), .o(n_26453) );
no02s01 g754507 ( .a(n_26707), .b(n_26712), .o(n_26771) );
in01s01 g754508 ( .a(n_26829), .o(n_26830) );
na02s01 g754509 ( .a(n_26814), .b(n_26832), .o(n_26829) );
no02s01 g754510 ( .a(FE_OCP_RBN4434_n_26160), .b(n_26740), .o(n_26868) );
no02s01 g754511 ( .a(n_26712), .b(n_26740), .o(n_26713) );
na02s01 g754512 ( .a(n_25515), .b(n_25514), .o(n_25516) );
in01s01 g754513 ( .a(FE_OCP_RBN5942_n_25544), .o(n_25629) );
in01f02 g754515 ( .a(n_25513), .o(n_25544) );
na02f08 g754516 ( .a(n_25429), .b(n_25207), .o(n_25513) );
na02s01 g754517 ( .a(n_26931), .b(n_26930), .o(n_26932) );
na02s03 g754518 ( .a(n_26739), .b(n_26685), .o(n_26792) );
in01s02 g754519 ( .a(n_26313), .o(n_26314) );
no02s01 TIMEBOOST_cell_876 ( .a(TIMEBOOST_net_52), .b(n_36925), .o(n_37023) );
in01s01 g754521 ( .a(n_26611), .o(n_26612) );
no02s06 TIMEBOOST_cell_5102 ( .a(n_8700), .b(n_8699), .o(TIMEBOOST_net_1499) );
no02s10 TIMEBOOST_cell_882 ( .a(FE_OCPN1342_n_11927), .b(TIMEBOOST_net_55), .o(n_11998) );
no02s01 TIMEBOOST_cell_5266 ( .a(n_44925), .b(n_38587), .o(TIMEBOOST_net_1581) );
in01s01 g754525 ( .a(n_26714), .o(n_26686) );
no02s01 g754526 ( .a(n_26541), .b(n_26573), .o(n_26714) );
ao12s02 g754527 ( .a(n_26541), .b(n_26708), .c(n_26643), .o(n_26644) );
no02s01 g754528 ( .a(n_25430), .b(n_25466), .o(n_27009) );
ao12s02 g754529 ( .a(n_25465), .b(n_25464), .c(n_25463), .o(n_27099) );
ao12s01 g754530 ( .a(n_25431), .b(n_25432), .c(n_25241), .o(n_25518) );
in01s01 g754531 ( .a(n_26351), .o(n_26352) );
ao12s01 g754532 ( .a(n_26236), .b(n_26235), .c(n_26234), .o(n_26351) );
in01s01 g754533 ( .a(n_26907), .o(n_26350) );
oa12s01 g754534 ( .a(n_26239), .b(n_26238), .c(n_26237), .o(n_26907) );
na02s01 g754535 ( .a(n_26238), .b(n_26237), .o(n_26239) );
no02s01 g754536 ( .a(n_26235), .b(n_26234), .o(n_26236) );
no02s02 g754537 ( .a(n_26551), .b(n_26550), .o(n_26552) );
no02s02 g754538 ( .a(n_26602), .b(n_26636), .o(n_26685) );
no02s02 g754539 ( .a(n_26311), .b(n_26271), .o(n_26312) );
no02s02 g754540 ( .a(n_26385), .b(n_26345), .o(n_26452) );
no02s01 g754541 ( .a(n_26608), .b(n_26609), .o(n_26610) );
no02s01 g754542 ( .a(n_26633), .b(n_26572), .o(n_26711) );
na02s02 g754543 ( .a(n_26641), .b(n_26640), .o(n_26642) );
in01s02 g754544 ( .a(n_26738), .o(n_26739) );
na02s02 g754545 ( .a(n_26710), .b(n_26638), .o(n_26738) );
na02s01 g754546 ( .a(n_26383), .b(n_26346), .o(n_26384) );
na02s01 g754548 ( .a(n_26813), .b(n_26866), .o(n_26946) );
in01s01 g754549 ( .a(n_26903), .o(n_26904) );
na02s01 g754550 ( .a(n_26865), .b(n_26864), .o(n_26903) );
no02s01 g754551 ( .a(n_26308), .b(n_26348), .o(n_26349) );
na02s02 g754552 ( .a(n_26864), .b(n_26417), .o(n_26418) );
in01s01 g754553 ( .a(n_26901), .o(n_26902) );
na02s01 g754554 ( .a(n_26863), .b(n_26862), .o(n_26901) );
no02s01 TIMEBOOST_cell_7067 ( .a(FE_OCPN3592_n_45301), .b(FE_OCP_RBN4483_n_11439), .o(TIMEBOOST_net_2292) );
in01s01 g754556 ( .a(n_26574), .o(n_26575) );
no02s01 g754557 ( .a(n_26550), .b(n_26549), .o(n_26574) );
no02f06 TIMEBOOST_cell_8637 ( .a(TIMEBOOST_net_2805), .b(FE_RN_588_0), .o(n_30727) );
in01s01 g754559 ( .a(n_26899), .o(n_26900) );
no02s01 g754560 ( .a(n_26861), .b(n_26608), .o(n_26899) );
in01s01 g754561 ( .a(n_26683), .o(n_26684) );
na02s01 g754562 ( .a(n_26640), .b(n_26606), .o(n_26683) );
in01s01 g754563 ( .a(n_26681), .o(n_26682) );
na02s01 g754564 ( .a(n_26710), .b(n_26639), .o(n_26681) );
no02s01 g754565 ( .a(n_26548), .b(n_26604), .o(n_26573) );
in01s01 g754566 ( .a(n_26736), .o(n_26737) );
na02s01 g754567 ( .a(n_26709), .b(n_26708), .o(n_26736) );
in01s01 g754568 ( .a(n_26928), .o(n_26929) );
na02s01 g754569 ( .a(n_26898), .b(n_26897), .o(n_26928) );
in01s01 g754570 ( .a(n_26790), .o(n_26791) );
na02s01 g754571 ( .a(n_26770), .b(n_26677), .o(n_26790) );
na02s01 g754572 ( .a(FE_OCP_RBN4434_n_26160), .b(n_26734), .o(n_26832) );
in01s01 g754573 ( .a(n_26769), .o(n_26814) );
no02s01 g754574 ( .a(FE_OCP_RBN4434_n_26160), .b(n_26734), .o(n_26769) );
no02s01 g754575 ( .a(n_26308), .b(n_26311), .o(n_26743) );
no02f08 g754576 ( .a(n_25432), .b(FE_OCPN1310_n_25431), .o(n_25433) );
no02s01 g754577 ( .a(n_25404), .b(n_25212), .o(n_25430) );
no02s01 g754578 ( .a(n_25405), .b(n_25213), .o(n_25466) );
no02s01 g754579 ( .a(n_25464), .b(n_25463), .o(n_25465) );
in01s01 g754580 ( .a(n_26233), .o(n_26930) );
ao12m04 g754581 ( .a(FE_OCPN3580_n_25370), .b(n_26163), .c(n_25372), .o(n_26233) );
in01s01 g754582 ( .a(n_26926), .o(n_26927) );
oa12s01 g754583 ( .a(n_26641), .b(n_26896), .c(n_26605), .o(n_26926) );
ao12s01 g754584 ( .a(n_26716), .b(FE_OCP_RBN4438_n_26160), .c(n_26348), .o(n_26908) );
in01s01 g754585 ( .a(n_26894), .o(n_26895) );
ao12s01 g754586 ( .a(n_26860), .b(FE_OCP_RBN4435_n_26160), .c(n_26680), .o(n_26894) );
in01s01 g754587 ( .a(n_26892), .o(n_26893) );
ao12s01 g754588 ( .a(n_26551), .b(FE_OCP_RBN4435_n_26160), .c(n_26510), .o(n_26892) );
in01s01 g754589 ( .a(n_26890), .o(n_26891) );
ao12s01 g754590 ( .a(n_26609), .b(FE_OCP_RBN4435_n_26160), .c(n_26546), .o(n_26890) );
in01s01 g754591 ( .a(n_26888), .o(n_26889) );
ao12s01 g754592 ( .a(n_26637), .b(FE_OCP_RBN4435_n_26160), .c(n_26604), .o(n_26888) );
in01s01 g754593 ( .a(n_26924), .o(n_26925) );
oa12s01 g754594 ( .a(n_26601), .b(n_26896), .c(n_26643), .o(n_26924) );
oa12s01 g754595 ( .a(n_26690), .b(FE_OCP_RBN6860_n_26160), .c(n_25605), .o(n_26943) );
ao12s01 g754596 ( .a(n_26385), .b(FE_OCP_RBN4438_n_26160), .c(n_26310), .o(n_26951) );
in01s01 g754597 ( .a(n_26793), .o(n_26707) );
oa12s01 g754598 ( .a(FE_OCP_RBN4434_n_26160), .b(n_26680), .c(n_26679), .o(n_26793) );
oa12s01 g754599 ( .a(n_25462), .b(n_25461), .c(n_25460), .o(n_27040) );
oa12s01 g754600 ( .a(n_25203), .b(n_25403), .c(n_25268), .o(n_25515) );
oa12f06 g754601 ( .a(n_25234), .b(n_25365), .c(n_25175), .o(n_25429) );
in01s01 g754602 ( .a(n_26886), .o(n_26887) );
oa22s01 g754603 ( .a(FE_OCP_RBN6857_n_26160), .b(n_25686), .c(FE_OCP_RBN4437_n_26160), .d(n_26417), .o(n_26886) );
in01s01 g754604 ( .a(n_26884), .o(n_26885) );
oa22s01 g754605 ( .a(FE_OCP_RBN6857_n_26160), .b(n_26512), .c(FE_OCP_RBN4437_n_26160), .d(n_25745), .o(n_26884) );
ao22s01 g754606 ( .a(FE_OCP_RBN6860_n_26160), .b(n_25371), .c(FE_OCP_RBN4439_n_26160), .d(n_25342), .o(n_26933) );
oa22s01 g754607 ( .a(n_26133), .b(n_25740), .c(n_26132), .d(n_25739), .o(n_26740) );
oa22s01 g754608 ( .a(FE_OCP_RBN4439_n_26160), .b(n_26162), .c(FE_OCP_RBN4435_n_26160), .d(n_26192), .o(n_26931) );
ao22s01 g754609 ( .a(FE_OCP_RBN4438_n_26160), .b(n_25524), .c(FE_OCP_RBN6860_n_26160), .d(n_26419), .o(n_26937) );
ao22s01 g754610 ( .a(FE_OCP_RBN4435_n_26160), .b(n_26855), .c(FE_OCP_RBN4438_n_26160), .d(n_26307), .o(n_26940) );
in01s01 g754611 ( .a(n_27014), .o(n_27062) );
in01s01 g754617 ( .a(n_27014), .o(n_27130) );
in01s01 g754626 ( .a(n_27366), .o(n_27536) );
in01s01 g754630 ( .a(FE_OCPN1340_n_27246), .o(n_27518) );
in01s04 g754637 ( .a(n_27246), .o(n_27366) );
in01s02 g754641 ( .a(n_27131), .o(n_27246) );
in01s01 g754647 ( .a(n_27131), .o(n_27315) );
in01s02 g754655 ( .a(n_27014), .o(n_27131) );
in01s01 g754656 ( .a(n_27130), .o(n_30823) );
in01s01 g754674 ( .a(FE_OCPN5130_FE_OFN1198_n_27014), .o(n_30584) );
in01s01 g754677 ( .a(n_27014), .o(n_30790) );
in01s02 g754679 ( .a(FE_OFN1199_n_27014), .o(n_30466) );
no02s01 g754684 ( .a(FE_OCP_RBN4434_n_26160), .b(n_26680), .o(n_26860) );
in01s01 g754685 ( .a(n_26606), .o(n_26572) );
na02s01 g754686 ( .a(FE_OCP_RBN6858_n_26160), .b(n_26544), .o(n_26606) );
no02s02 g754687 ( .a(FE_OCP_RBN6097_n_26160), .b(n_26310), .o(n_26385) );
in01s01 g754688 ( .a(n_26486), .o(n_26862) );
no02s01 g754689 ( .a(FE_OCP_RBN6097_n_26160), .b(n_26451), .o(n_26486) );
na02s01 g754690 ( .a(FE_OCP_RBN4435_n_26160), .b(n_26679), .o(n_26897) );
in01s01 g754691 ( .a(n_26548), .o(n_26639) );
no02s01 g754692 ( .a(FE_OCP_RBN3269_n_26160), .b(n_26509), .o(n_26548) );
no02s01 g754693 ( .a(FE_OCP_RBN4433_n_26160), .b(n_26507), .o(n_26861) );
in01s01 g754694 ( .a(n_26812), .o(n_26813) );
no02s01 g754695 ( .a(FE_OCP_RBN6860_n_26160), .b(n_25575), .o(n_26812) );
na02s01 g754696 ( .a(n_26160), .b(n_25685), .o(n_26864) );
na02s01 g754697 ( .a(FE_OCP_RBN4438_n_26160), .b(n_25547), .o(n_26865) );
no02s01 g754698 ( .a(FE_OCP_RBN6096_n_26160), .b(n_26348), .o(n_26716) );
no02s01 TIMEBOOST_cell_875 ( .a(n_37022), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_1_), .o(TIMEBOOST_net_52) );
no02s02 g754700 ( .a(n_26160), .b(n_26192), .o(n_26193) );
no02s02 g754701 ( .a(FE_OCP_RBN6096_n_26160), .b(n_26307), .o(n_26232) );
no02s02 g754702 ( .a(FE_OCP_RBN6096_n_26160), .b(n_25440), .o(n_26311) );
in01s01 g754703 ( .a(n_26271), .o(n_26690) );
no02s02 g754704 ( .a(FE_OCP_RBN6096_n_26160), .b(n_26230), .o(n_26271) );
in01s01 g754706 ( .a(n_26308), .o(n_26346) );
no02s02 g754707 ( .a(n_26160), .b(n_25441), .o(n_26308) );
in01s01 g754708 ( .a(n_26345), .o(n_26866) );
no02s02 g754709 ( .a(FE_OCP_RBN6096_n_26160), .b(n_25683), .o(n_26345) );
na02s01 g754710 ( .a(FE_OCP_RBN4437_n_26160), .b(n_26451), .o(n_26863) );
no02s01 g754711 ( .a(FE_OCP_RBN6097_n_26160), .b(n_25712), .o(n_26549) );
in01s01 g754712 ( .a(n_26550), .o(n_26508) );
no02s02 g754713 ( .a(FE_OCP_RBN6858_n_26160), .b(n_25713), .o(n_26550) );
no02s02 g754714 ( .a(FE_OCP_RBN6858_n_26160), .b(n_26510), .o(n_26551) );
in01s01 g754715 ( .a(n_26547), .o(n_26608) );
na02s01 g754716 ( .a(FE_OCP_RBN6856_n_26160), .b(n_26507), .o(n_26547) );
no02s01 g754717 ( .a(FE_OCP_RBN6858_n_26160), .b(n_26546), .o(n_26609) );
in01s01 g754718 ( .a(n_26571), .o(n_26640) );
no02s01 g754719 ( .a(FE_OCP_RBN6858_n_26160), .b(n_26544), .o(n_26571) );
na02s02 g754720 ( .a(n_26541), .b(n_26605), .o(n_26641) );
na02s02 g754721 ( .a(n_26541), .b(n_26509), .o(n_26710) );
in01s01 g754722 ( .a(n_26637), .o(n_26638) );
no02s01 g754723 ( .a(FE_OCP_RBN4434_n_26160), .b(n_26604), .o(n_26637) );
na02s01 g754724 ( .a(FE_OCP_RBN4434_n_26160), .b(n_26542), .o(n_26708) );
in01s01 g754725 ( .a(n_26636), .o(n_26709) );
no02s01 g754726 ( .a(FE_OCP_RBN4434_n_26160), .b(n_26542), .o(n_26636) );
in01s01 g754727 ( .a(n_26601), .o(n_26602) );
na02s02 g754728 ( .a(n_26541), .b(n_26643), .o(n_26601) );
na02s01 g754729 ( .a(n_26541), .b(n_26033), .o(n_26898) );
in01s01 g754730 ( .a(n_26712), .o(n_26677) );
no02s01 g754731 ( .a(n_26541), .b(n_26634), .o(n_26712) );
na02s01 g754732 ( .a(n_26541), .b(n_26634), .o(n_26770) );
in01s01 g754733 ( .a(n_25432), .o(n_25464) );
na02s01 g754735 ( .a(n_25461), .b(n_25460), .o(n_25462) );
oa12s01 g754736 ( .a(n_25287), .b(n_26161), .c(n_25312), .o(n_26238) );
ao12s01 g754737 ( .a(n_25771), .b(n_26161), .c(n_25736), .o(n_26235) );
in01s01 g754738 ( .a(n_26381), .o(n_26382) );
no02s01 g754739 ( .a(n_26160), .b(n_25684), .o(n_26381) );
in01s01 g754740 ( .a(n_26383), .o(n_26343) );
oa12s02 g754741 ( .a(FE_OCP_RBN6096_n_26160), .b(n_26230), .c(n_26307), .o(n_26383) );
in01s01 g754742 ( .a(n_26415), .o(n_26416) );
na02s01 g754743 ( .a(FE_OCP_RBN6097_n_26160), .b(n_25687), .o(n_26415) );
no02s01 g754744 ( .a(FE_OCP_RBN6857_n_26160), .b(n_25746), .o(n_26484) );
in01s01 g754745 ( .a(n_26741), .o(n_26633) );
na02s01 g754746 ( .a(FE_OCP_RBN6858_n_26160), .b(n_25882), .o(n_26741) );
ao12s01 g754747 ( .a(n_25337), .b(n_25336), .c(n_25335), .o(n_26966) );
ao12s01 g754748 ( .a(n_25334), .b(n_25366), .c(n_25333), .o(n_27018) );
in01s01 g754749 ( .a(n_25404), .o(n_25405) );
oa12s01 g754750 ( .a(n_25209), .b(n_25366), .c(n_25154), .o(n_25404) );
oa12s01 g754751 ( .a(n_26135), .b(n_26161), .c(n_26134), .o(n_26734) );
na02s01 g754753 ( .a(n_26161), .b(n_26134), .o(n_26135) );
no02s01 g754754 ( .a(n_25336), .b(n_25335), .o(n_25337) );
in01s01 g754755 ( .a(n_25403), .o(n_25461) );
in01s01 g754756 ( .a(n_25365), .o(n_25403) );
oa12f08 g754757 ( .a(n_25176), .b(n_25248), .c(n_25146), .o(n_25365) );
no02s01 g754758 ( .a(n_25366), .b(n_25333), .o(n_25334) );
in01s01 g754759 ( .a(n_26132), .o(n_26133) );
oa12s01 g754760 ( .a(n_25306), .b(n_26106), .c(n_25191), .o(n_26132) );
in01s01 g754767 ( .a(FE_OCP_RBN4435_n_26160), .o(n_26896) );
in01s03 g754786 ( .a(FE_OCP_RBN4434_n_26160), .o(n_26541) );
in01m06 g754798 ( .a(n_26163), .o(n_26160) );
na02s10 TIMEBOOST_cell_868 ( .a(n_17561), .b(TIMEBOOST_net_48), .o(n_17683) );
ao22s01 g754800 ( .a(n_25952), .b(n_25709), .c(n_25953), .d(n_25708), .o(n_26643) );
oa22s01 g754801 ( .a(n_26006), .b(n_25710), .c(n_26005), .d(n_25711), .o(n_26680) );
ao12s01 g754802 ( .a(n_26073), .b(n_26106), .c(n_26072), .o(n_26634) );
no02s01 g754805 ( .a(n_26106), .b(n_26072), .o(n_26073) );
no02s01 g754806 ( .a(n_26008), .b(n_25309), .o(n_26161) );
na02m10 g754809 ( .a(n_25361), .b(FE_OCP_RBN2935_n_25401), .o(n_25457) );
in01s01 TIMEBOOST_cell_8905 ( .a(TIMEBOOST_net_2948), .o(TIMEBOOST_net_2949) );
na02m03 TIMEBOOST_cell_867 ( .a(n_17458), .b(n_17560), .o(TIMEBOOST_net_48) );
ao12f08 g754812 ( .a(n_25116), .b(n_25282), .c(n_25069), .o(n_25366) );
ao12s01 g754814 ( .a(n_25281), .b(n_25280), .c(n_25279), .o(n_25363) );
ao12s01 g754815 ( .a(n_25246), .b(n_25247), .c(n_25144), .o(n_25336) );
ao12s01 g754816 ( .a(n_25245), .b(n_25282), .c(n_25244), .o(n_26956) );
na02s01 g754817 ( .a(n_25949), .b(n_25290), .o(n_26106) );
no02s01 g754818 ( .a(n_25280), .b(n_25279), .o(n_25281) );
no02f08 g754819 ( .a(n_25247), .b(n_25246), .o(n_25248) );
na02s02 g754820 ( .a(n_25511), .b(n_25451), .o(n_25782) );
no02s01 g754821 ( .a(n_25282), .b(n_25244), .o(n_25245) );
na02s06 g754825 ( .a(n_25210), .b(n_25303), .o(n_25361) );
no02s06 TIMEBOOST_cell_3154 ( .a(n_42633), .b(n_42593), .o(TIMEBOOST_net_868) );
in01s01 g754827 ( .a(n_26007), .o(n_26008) );
na02f06 g754828 ( .a(n_25948), .b(n_25341), .o(n_26007) );
in01s01 g754829 ( .a(n_26005), .o(n_26006) );
ao12s01 g754830 ( .a(n_25679), .b(n_25977), .c(n_25741), .o(n_26005) );
in01s01 g754831 ( .a(n_25952), .o(n_25953) );
oa12s01 g754832 ( .a(n_25254), .b(n_25923), .c(n_25189), .o(n_25952) );
oa12s01 g754833 ( .a(n_25906), .b(n_25923), .c(n_25905), .o(n_26542) );
in01s01 g754834 ( .a(n_26679), .o(n_26033) );
oa12s01 g754835 ( .a(n_25951), .b(n_25977), .c(n_25950), .o(n_26679) );
na02s01 g754838 ( .a(n_25564), .b(n_25973), .o(n_25565) );
na02m04 TIMEBOOST_cell_3130 ( .a(n_34946), .b(n_30545), .o(TIMEBOOST_net_856) );
na02s01 g754840 ( .a(n_25625), .b(n_25626), .o(n_25627) );
in01s01 g754844 ( .a(n_25487), .o(n_25488) );
na02s02 g754845 ( .a(n_25389), .b(n_25388), .o(n_25487) );
na02s04 g754846 ( .a(n_25275), .b(n_24332), .o(n_25303) );
in01s01 g754847 ( .a(n_25593), .o(n_25594) );
na02s02 g754848 ( .a(n_25506), .b(n_25973), .o(n_25593) );
na02s01 g754850 ( .a(n_25486), .b(n_25424), .o(n_25509) );
in01s01 g754853 ( .a(n_25650), .o(n_25651) );
na02s01 g754854 ( .a(n_25624), .b(n_25625), .o(n_25650) );
in01s01 g754855 ( .a(n_25695), .o(n_25696) );
no02s01 g754856 ( .a(n_25673), .b(n_25672), .o(n_25695) );
no02f06 TIMEBOOST_cell_6258 ( .a(TIMEBOOST_net_1980), .b(FE_OCP_RBN3324_n_5813), .o(n_5946) );
in01s01 g754858 ( .a(n_25724), .o(n_25725) );
na02s01 g754859 ( .a(FE_RN_1509_0), .b(n_25694), .o(n_25724) );
in01s01 g754860 ( .a(n_25427), .o(n_25428) );
na02s01 g754861 ( .a(n_25398), .b(n_25397), .o(n_25427) );
na02s01 g754862 ( .a(n_25977), .b(n_25950), .o(n_25951) );
na02s01 g754863 ( .a(n_25923), .b(n_25905), .o(n_25906) );
na02f06 g754864 ( .a(n_25242), .b(n_25241), .o(n_25243) );
na02s01 g754865 ( .a(n_25668), .b(n_25667), .o(n_25723) );
na02s01 g754866 ( .a(n_25277), .b(n_25242), .o(n_25517) );
in01s01 g754867 ( .a(n_25670), .o(n_25671) );
na02s01 g754868 ( .a(n_25626), .b(n_25591), .o(n_25670) );
no02s01 g754869 ( .a(n_25329), .b(n_25328), .o(n_25396) );
na02s02 g754870 ( .a(n_25301), .b(n_25357), .o(n_25426) );
in01s01 g754871 ( .a(n_25622), .o(n_25623) );
na02s01 g754872 ( .a(n_25564), .b(n_25543), .o(n_25622) );
in01s01 g754873 ( .a(n_25948), .o(n_25949) );
no02f06 g754874 ( .a(n_25904), .b(n_25308), .o(n_25948) );
oa12s01 g754875 ( .a(n_25885), .b(n_25884), .c(n_25883), .o(n_26604) );
ao12f08 g754876 ( .a(n_25046), .b(n_25187), .c(n_25105), .o(n_25282) );
ao12s01 g754877 ( .a(n_25186), .b(n_25185), .c(n_25184), .o(n_26850) );
in01s01 g754878 ( .a(n_25247), .o(n_25280) );
oa12f08 g754879 ( .a(n_25008), .b(n_25128), .c(n_25066), .o(n_25247) );
in01s01 g754880 ( .a(n_25775), .o(n_25776) );
oa22s01 g754881 ( .a(n_25542), .b(n_24857), .c(FE_OCPN1088_n_25481), .d(n_24872), .o(n_25775) );
no02m08 g754882 ( .a(n_25453), .b(n_25382), .o(n_25511) );
oa12s01 g754883 ( .a(n_25158), .b(n_25187), .c(n_25157), .o(n_26873) );
in01s02 g754884 ( .a(n_25394), .o(n_25395) );
na02s02 g754885 ( .a(n_25276), .b(n_25302), .o(n_25394) );
na02s02 g754887 ( .a(n_25485), .b(n_25452), .o(n_25562) );
na02s02 g754889 ( .a(n_25385), .b(n_25421), .o(n_25507) );
in01s01 g754890 ( .a(n_25721), .o(n_25722) );
oa22s01 g754891 ( .a(n_25542), .b(FE_OCPN1081_n_24819), .c(FE_OCP_RBN6797_n_25211), .d(n_24865), .o(n_25721) );
na02s01 g754892 ( .a(FE_OCP_RBN2907_n_25238), .b(n_24458), .o(n_25452) );
in01s01 g754893 ( .a(n_25331), .o(n_25398) );
no02s02 g754894 ( .a(n_25210), .b(FE_OCP_RBN1002_n_24079), .o(n_25331) );
na02s01 g754895 ( .a(n_25210), .b(n_24217), .o(n_25302) );
na02s01 g754896 ( .a(n_25181), .b(FE_OCP_RBN4149_n_24173), .o(n_25276) );
na02s02 g754897 ( .a(FE_OCP_RBN6796_n_25211), .b(n_24632), .o(n_25625) );
in01s01 g754899 ( .a(n_25301), .o(n_25329) );
na02s06 g754900 ( .a(FE_OCP_RBN5922_n_25211), .b(n_24332), .o(n_25301) );
no02s04 g754901 ( .a(n_25210), .b(FE_OCP_RBN1009_n_24175), .o(n_25359) );
na02s02 g754902 ( .a(FE_OCP_RBN5924_n_25211), .b(FE_OCP_RBN2621_n_24175), .o(n_25399) );
in01s01 g754904 ( .a(n_25275), .o(n_25358) );
na02s03 g754905 ( .a(n_25211), .b(FE_OCP_RBN1010_n_24175), .o(n_25275) );
na02s01 g754906 ( .a(FE_OCP_RBN6796_n_25211), .b(n_24518), .o(n_25564) );
na02s01 g754907 ( .a(FE_OCP_RBN2907_n_25238), .b(n_24486), .o(n_25973) );
na02s02 g754908 ( .a(n_25542), .b(n_24612), .o(n_25624) );
na02s01 g754909 ( .a(n_25542), .b(n_24717), .o(n_25591) );
na02s01 g754910 ( .a(FE_OCP_RBN6796_n_25211), .b(n_24794), .o(n_25626) );
na02s02 g754911 ( .a(FE_OCP_RBN5925_n_25211), .b(n_24457), .o(n_25486) );
na02m08 TIMEBOOST_cell_7789 ( .a(TIMEBOOST_net_2525), .b(n_34730), .o(n_34828) );
in01s01 g754913 ( .a(n_25424), .o(n_25425) );
na02m01 g754915 ( .a(n_25327), .b(n_25390), .o(n_25424) );
na02s01 g754916 ( .a(FE_OCP_RBN6793_n_25211), .b(n_24438), .o(n_25485) );
in01s01 g754918 ( .a(n_25389), .o(n_25422) );
na02s02 g754919 ( .a(FE_OCP_RBN5925_n_25211), .b(FE_OCP_RBN5671_n_24288), .o(n_25389) );
na02s01 g754920 ( .a(FE_OCP_RBN5923_n_25211), .b(n_25386), .o(n_25388) );
na02s02 g754921 ( .a(n_25327), .b(n_25386), .o(n_25760) );
na02s01 g754922 ( .a(n_25327), .b(n_24419), .o(n_25385) );
na02s01 g754923 ( .a(FE_OCP_RBN5925_n_25211), .b(n_24305), .o(n_25421) );
na02s01 g754924 ( .a(n_25542), .b(n_24546), .o(n_25543) );
no02s01 g754925 ( .a(FE_OCP_RBN6797_n_25211), .b(n_24680), .o(n_25673) );
no02m01 g754926 ( .a(n_25542), .b(n_24959), .o(n_25672) );
no02s01 g754928 ( .a(FE_OCP_RBN6797_n_25211), .b(n_24774), .o(n_25648) );
na02m01 g754929 ( .a(FE_OCP_RBN6797_n_25211), .b(n_24774), .o(n_25694) );
no02s01 g754930 ( .a(n_25327), .b(n_24332), .o(n_25328) );
na02s01 g754931 ( .a(FE_OCP_RBN4157_n_24222), .b(FE_OCP_RBN4298_n_25238), .o(n_25357) );
in01s01 g754933 ( .a(n_25239), .o(n_25397) );
no02f01 g754934 ( .a(n_25181), .b(FE_OCP_RBN1001_n_24079), .o(n_25239) );
in01s01 g754936 ( .a(n_25506), .o(n_25540) );
na02s02 g754937 ( .a(FE_OCP_RBN6794_n_25211), .b(n_24633), .o(n_25506) );
na02s01 g754938 ( .a(n_25884), .b(n_25883), .o(n_25885) );
na02f04 g754939 ( .a(n_25149), .b(n_24054), .o(n_25242) );
na02m06 g754940 ( .a(n_25150), .b(n_24055), .o(n_25277) );
no02s01 g754941 ( .a(n_25185), .b(n_25184), .o(n_25186) );
no02f02 g754943 ( .a(n_25505), .b(n_25553), .o(n_25561) );
in01s02 g754944 ( .a(n_25668), .o(n_25669) );
ao12s02 g754945 ( .a(n_25647), .b(n_25552), .c(n_25551), .o(n_25668) );
na02s01 g754946 ( .a(n_25187), .b(n_25157), .o(n_25158) );
na02s01 g754947 ( .a(n_25867), .b(n_26507), .o(n_25882) );
na02s02 g754948 ( .a(n_25327), .b(n_24392), .o(n_25455) );
no02s04 g754950 ( .a(n_25210), .b(FE_OCPN5364_n_24221), .o(n_25272) );
in01s01 g754952 ( .a(n_25383), .o(n_25418) );
na02s01 g754953 ( .a(n_25210), .b(n_24420), .o(n_25383) );
in01s01 g754954 ( .a(n_25588), .o(n_25589) );
no02s02 g754955 ( .a(FE_OCP_RBN6796_n_25211), .b(n_24635), .o(n_25588) );
in01s01 g754956 ( .a(n_25904), .o(n_25977) );
oa12s01 g754958 ( .a(n_25288), .b(n_25868), .c(n_25200), .o(n_25923) );
na02s06 TIMEBOOST_cell_8840 ( .a(n_45304), .b(FE_OCPN4845_FE_OFN4779_n_44490), .o(TIMEBOOST_net_2907) );
ao12s01 g754961 ( .a(n_25153), .b(n_25152), .c(n_25151), .o(n_26820) );
ao12s01 g754962 ( .a(n_25804), .b(n_25803), .c(n_25802), .o(n_26605) );
ao12s01 g754963 ( .a(n_25840), .b(n_25868), .c(n_25839), .o(n_26509) );
no02s01 g754964 ( .a(n_25868), .b(n_25839), .o(n_25840) );
no02s01 g754965 ( .a(n_25803), .b(n_25802), .o(n_25804) );
ao12f08 g754967 ( .a(n_25050), .b(n_25076), .c(n_25025), .o(n_25187) );
in01s01 g754969 ( .a(n_25212), .o(n_25213) );
no02s01 g754970 ( .a(n_25182), .b(n_25155), .o(n_25212) );
na02s01 g754971 ( .a(n_25148), .b(n_25241), .o(n_25463) );
no02s01 g754972 ( .a(n_25152), .b(n_25151), .o(n_25153) );
in01m02 g754974 ( .a(n_25149), .o(n_25150) );
oa12s01 g754976 ( .a(n_25108), .b(n_25118), .c(n_25107), .o(n_26801) );
in01s01 g754977 ( .a(n_25128), .o(n_25185) );
oa12f08 g754978 ( .a(n_24983), .b(n_25118), .c(n_25035), .o(n_25128) );
in01f01 g754979 ( .a(n_25504), .o(n_25505) );
no02f04 g754980 ( .a(n_25414), .b(n_25482), .o(n_25504) );
na02s01 g754981 ( .a(n_25381), .b(FE_OCP_RBN4311_n_25178), .o(n_25451) );
na02s02 g754982 ( .a(n_25555), .b(n_25500), .o(n_25750) );
na02s01 g754983 ( .a(n_25619), .b(n_25551), .o(n_25667) );
in01s01 g754984 ( .a(n_25867), .o(n_26546) );
ao12s01 g754985 ( .a(n_25774), .b(n_25773), .c(n_25772), .o(n_25867) );
oa12s01 g754986 ( .a(n_25801), .b(n_25800), .c(n_25799), .o(n_26544) );
oa12s01 g754987 ( .a(n_25344), .b(n_25744), .c(n_25193), .o(n_25884) );
in01s06 g755000 ( .a(FE_OCP_RBN6796_n_25211), .o(n_25542) );
in01s06 g755017 ( .a(n_25181), .o(n_25211) );
in01s06 g755021 ( .a(n_25210), .o(n_25327) );
in01s06 g755025 ( .a(n_25181), .o(n_25210) );
no02f08 g755026 ( .a(n_25117), .b(n_25106), .o(n_25181) );
ao12f06 g755027 ( .a(FE_OCPN1354_n_22484), .b(n_25048), .c(n_24829), .o(n_25117) );
no02f08 g755028 ( .a(n_25743), .b(n_25343), .o(n_25868) );
no02s01 g755029 ( .a(n_25773), .b(n_25772), .o(n_25774) );
na02s01 g755030 ( .a(n_25800), .b(n_25799), .o(n_25801) );
na02s03 g755031 ( .a(n_25127), .b(FE_OCPN1314_n_25126), .o(n_25241) );
no02m08 g755032 ( .a(n_25103), .b(n_23888), .o(n_25182) );
no02m02 g755033 ( .a(n_25102), .b(FE_OCP_DRV_N1476_n_23887), .o(n_25155) );
in01s01 g755034 ( .a(n_25431), .o(n_25148) );
no02m06 g755035 ( .a(n_25127), .b(FE_OCPN1314_n_25126), .o(n_25431) );
na02s01 g755036 ( .a(n_25118), .b(n_25107), .o(n_25108) );
no02s01 g755037 ( .a(n_25233), .b(n_25208), .o(n_25514) );
na02s01 g755038 ( .a(n_25323), .b(n_25206), .o(n_25628) );
no02f06 g755039 ( .a(n_25233), .b(n_25268), .o(n_25234) );
in01f02 g755041 ( .a(n_25355), .o(n_25356) );
na02f06 g755042 ( .a(n_25321), .b(n_25267), .o(n_25355) );
na02s04 TIMEBOOST_cell_2113 ( .a(n_35327), .b(n_30633), .o(TIMEBOOST_net_671) );
in01s02 g755045 ( .a(n_25446), .o(n_25447) );
no02m04 g755046 ( .a(n_25415), .b(n_25416), .o(n_25446) );
na02m04 g755047 ( .a(n_25352), .b(n_25350), .o(n_25382) );
no02s06 g755049 ( .a(n_25445), .b(n_25375), .o(n_25479) );
na02s02 g755050 ( .a(n_25413), .b(n_25412), .o(n_25414) );
na02m01 g755051 ( .a(n_25349), .b(n_24422), .o(n_25381) );
in01s01 g755052 ( .a(n_25537), .o(n_25538) );
na02s02 g755053 ( .a(n_25503), .b(n_25502), .o(n_25537) );
in01s01 g755054 ( .a(n_25585), .o(n_25586) );
no02s01 g755055 ( .a(FE_OCP_RBN4341_n_25500), .b(n_25535), .o(n_25585) );
no02s01 g755056 ( .a(n_25647), .b(n_25535), .o(n_25536) );
in01s01 g755057 ( .a(n_25661), .o(n_25662) );
na02s01 g755058 ( .a(n_25613), .b(n_25645), .o(n_25661) );
no02s01 g755059 ( .a(n_25554), .b(n_25553), .o(n_25555) );
na02s02 g755060 ( .a(n_25499), .b(n_25531), .o(n_25552) );
na02s01 g755061 ( .a(n_25618), .b(FE_OCP_RBN2709_n_24505), .o(n_25619) );
no02s01 g755062 ( .a(n_25077), .b(n_24972), .o(n_25152) );
na02s01 g755063 ( .a(n_25125), .b(n_25209), .o(n_25333) );
oa12s01 g755064 ( .a(n_25196), .b(n_25715), .c(n_25217), .o(n_25803) );
no02s02 g755065 ( .a(n_25319), .b(n_25229), .o(n_25354) );
na02m02 g755066 ( .a(n_25320), .b(n_25205), .o(n_25380) );
in01s04 g755067 ( .a(n_25378), .o(n_25379) );
no02s06 g755068 ( .a(n_25291), .b(n_25353), .o(n_25378) );
in01s02 g755069 ( .a(n_25477), .o(n_25478) );
no02s02 g755070 ( .a(n_25351), .b(n_25377), .o(n_25477) );
in01s01 g755071 ( .a(n_25533), .o(n_25534) );
na02s02 g755072 ( .a(n_25413), .b(n_25444), .o(n_25533) );
in01s01 g755073 ( .a(n_25615), .o(n_25616) );
no02s01 g755074 ( .a(n_25554), .b(n_25532), .o(n_25615) );
in01s01 g755075 ( .a(n_25719), .o(n_25720) );
no02s01 g755076 ( .a(n_25693), .b(n_25644), .o(n_25719) );
in01s01 g755077 ( .a(n_25747), .o(n_25748) );
oa22s01 g755078 ( .a(n_25551), .b(n_24621), .c(n_25373), .d(n_24650), .o(n_25747) );
oa12s02 g755079 ( .a(n_25075), .b(n_25074), .c(n_25073), .o(n_26752) );
oa12s01 g755080 ( .a(n_25718), .b(n_25717), .c(n_25716), .o(n_26510) );
in01s01 g755081 ( .a(n_25583), .o(n_25584) );
na02s02 g755082 ( .a(n_25476), .b(n_25501), .o(n_25583) );
in01s01 g755083 ( .a(n_25691), .o(n_25692) );
na02s02 g755084 ( .a(n_25612), .b(n_25582), .o(n_25691) );
no03s04 TIMEBOOST_cell_8203 ( .a(FE_RN_1903_0), .b(FE_RN_1904_0), .c(n_1713), .o(n_1766) );
na02s01 g755086 ( .a(n_25717), .b(n_25716), .o(n_25718) );
no02s01 g755087 ( .a(n_25688), .b(n_25195), .o(n_25800) );
in01s01 g755088 ( .a(n_25154), .o(n_25125) );
no02s06 g755089 ( .a(n_25098), .b(FE_OCP_DRV_N1474_n_23792), .o(n_25154) );
no02f06 g755090 ( .a(n_25024), .b(n_24972), .o(n_25025) );
in01s01 g755091 ( .a(n_25076), .o(n_25077) );
na02f08 g755092 ( .a(n_25074), .b(n_25018), .o(n_25076) );
in01s01 g755093 ( .a(n_25147), .o(n_25209) );
no02m06 g755094 ( .a(n_25099), .b(n_23793), .o(n_25147) );
no02s01 g755095 ( .a(n_25268), .b(n_25204), .o(n_25460) );
no02f04 g755096 ( .a(n_25180), .b(n_25179), .o(n_25233) );
in01s01 g755097 ( .a(n_25207), .o(n_25208) );
na02s02 g755098 ( .a(n_25180), .b(n_25179), .o(n_25207) );
in01s01 g755100 ( .a(n_25206), .o(n_25231) );
na02m06 g755101 ( .a(n_25178), .b(n_24093), .o(n_25206) );
na02f01 g755102 ( .a(FE_OCP_RBN2911_n_25178), .b(FE_OCPN871_n_24098), .o(n_25323) );
no02s02 g755103 ( .a(FE_OCP_RBN4307_n_25178), .b(n_24093), .o(n_25292) );
in01s02 g755104 ( .a(n_25319), .o(n_25320) );
no02s02 g755105 ( .a(FE_OCP_RBN4309_n_25178), .b(FE_OCP_RBN1022_n_24181), .o(n_25319) );
in01s01 g755107 ( .a(n_25205), .o(n_25229) );
na02m04 g755108 ( .a(n_25178), .b(FE_OCP_RBN1022_n_24181), .o(n_25205) );
na02s10 g755109 ( .a(FE_OCP_RBN4309_n_25178), .b(FE_OCPN1312_FE_OCP_RBN1024_n_24125), .o(n_25321) );
in01m02 g755110 ( .a(FE_OCP_RBN6763_FE_RN_2259_0), .o(n_25267) );
no02s02 g755112 ( .a(FE_OCP_RBN1019_n_24165), .b(FE_OCP_RBN4309_n_25178), .o(n_25291) );
no02m06 g755113 ( .a(FE_OCP_RBN2911_n_25178), .b(n_25265), .o(n_25353) );
in01s02 g755114 ( .a(n_25352), .o(n_25416) );
na02s04 g755115 ( .a(FE_OCPN1096_n_25318), .b(FE_OCP_RBN4311_n_25178), .o(n_25352) );
no02m02 g755116 ( .a(FE_OCP_RBN4311_n_25178), .b(FE_OCPN1096_n_25318), .o(n_25415) );
no02s01 g755117 ( .a(FE_OCP_RBN4311_n_25178), .b(n_25316), .o(n_25377) );
in01s01 g755118 ( .a(n_25350), .o(n_25351) );
na02s02 g755119 ( .a(n_25316), .b(FE_OCP_RBN4311_n_25178), .o(n_25350) );
no02f01 g755120 ( .a(FE_OCP_RBN5901_n_25178), .b(n_24310), .o(n_25482) );
no02s02 g755121 ( .a(FE_OCP_RBN4311_n_25178), .b(n_24310), .o(n_25375) );
in01m01 g755122 ( .a(n_25349), .o(n_25445) );
na02s06 g755123 ( .a(FE_OCP_RBN4311_n_25178), .b(n_24310), .o(n_25349) );
na02s02 g755124 ( .a(FE_OCP_RBN5903_n_25178), .b(n_24422), .o(n_25413) );
na02s01 g755125 ( .a(FE_OCP_RBN4311_n_25178), .b(n_24395), .o(n_25444) );
na02s02 g755126 ( .a(FE_OCP_RBN5901_n_25178), .b(FE_OCP_RBN2666_n_24372), .o(n_25503) );
na02s02 g755127 ( .a(n_25373), .b(n_24529), .o(n_25502) );
na02s01 g755128 ( .a(n_25373), .b(FE_OCP_RBN2695_n_24436), .o(n_25476) );
na02s01 g755129 ( .a(FE_OCP_RBN5901_n_25178), .b(n_24469), .o(n_25501) );
na02s01 g755131 ( .a(n_25373), .b(FE_OCP_RBN5707_n_24451), .o(n_25500) );
in01s01 g755132 ( .a(n_25535), .o(n_25499) );
no02s02 g755133 ( .a(n_25373), .b(FE_OCP_RBN5707_n_24451), .o(n_25535) );
no02s01 g755134 ( .a(FE_OCP_RBN5901_n_25178), .b(FE_OCP_RBN2704_n_24510), .o(n_25554) );
no02s01 g755135 ( .a(n_25373), .b(n_25531), .o(n_25532) );
in01s01 g755136 ( .a(n_25613), .o(n_25614) );
na02s01 g755137 ( .a(n_25373), .b(n_45633), .o(n_25613) );
na02s02 g755138 ( .a(n_25551), .b(FE_OCP_RBN5722_n_24506), .o(n_25645) );
na02s01 g755139 ( .a(n_25373), .b(n_24555), .o(n_25582) );
na02s01 g755140 ( .a(n_25551), .b(FE_OCP_RBN2715_n_24501), .o(n_25612) );
no02s01 g755141 ( .a(n_25551), .b(n_25104), .o(n_25693) );
no02s01 g755142 ( .a(n_25373), .b(FE_OCP_RBN2709_n_24505), .o(n_25644) );
no02s01 g755143 ( .a(n_25050), .b(n_25024), .o(n_25151) );
na02s01 g755144 ( .a(n_25074), .b(n_25073), .o(n_25075) );
no02s01 g755145 ( .a(n_25070), .b(n_25116), .o(n_25244) );
no02s01 g755146 ( .a(n_25745), .b(n_26451), .o(n_25746) );
na02s01 g755147 ( .a(n_25105), .b(n_25047), .o(n_25157) );
in01m02 g755148 ( .a(n_25071), .o(n_25072) );
ao12f04 g755149 ( .a(n_24695), .b(n_24989), .c(n_24690), .o(n_25071) );
in01s01 g755150 ( .a(n_25743), .o(n_25744) );
no02f06 g755151 ( .a(n_25715), .b(n_25198), .o(n_25743) );
oa12s01 g755152 ( .a(n_25571), .b(n_25714), .c(n_25604), .o(n_25773) );
in01s04 g755154 ( .a(n_25102), .o(n_25103) );
oa12f08 g755156 ( .a(n_24961), .b(n_25049), .c(n_24913), .o(n_25118) );
in01s01 g755157 ( .a(FE_OCP_DRV_N5157_n_25100), .o(n_25101) );
ao12s01 g755158 ( .a(n_25021), .b(n_25020), .c(n_25049), .o(n_25100) );
no02m10 g755160 ( .a(FE_OCP_RBN4309_n_25178), .b(n_24201), .o(n_25295) );
na02s06 g755161 ( .a(FE_OCP_RBN5903_n_25178), .b(n_24316), .o(n_25412) );
no02s01 g755162 ( .a(FE_OCP_RBN5901_n_25178), .b(n_24531), .o(n_25553) );
no02s02 g755163 ( .a(n_25373), .b(n_24570), .o(n_25647) );
no02s01 g755164 ( .a(n_25551), .b(n_24642), .o(n_25749) );
na02s01 g755165 ( .a(n_25551), .b(n_24639), .o(n_25618) );
ao12s01 g755166 ( .a(n_25690), .b(n_25714), .c(n_25689), .o(n_26507) );
na02f06 g755167 ( .a(n_25042), .b(n_24694), .o(n_25048) );
no02s01 g755168 ( .a(n_25714), .b(n_25689), .o(n_25690) );
no02m04 g755169 ( .a(n_25045), .b(FE_OCP_DRV_N1472_n_25044), .o(n_25116) );
in01s01 g755170 ( .a(n_25046), .o(n_25047) );
no02m04 g755171 ( .a(n_25023), .b(FE_OCP_DRV_N1470_n_25022), .o(n_25046) );
no02m06 g755172 ( .a(n_24946), .b(n_23628), .o(n_25050) );
no02f04 g755173 ( .a(n_24945), .b(n_23627), .o(n_25024) );
na02s06 g755174 ( .a(n_25023), .b(FE_OCP_DRV_N1470_n_25022), .o(n_25105) );
in01s01 g755175 ( .a(n_25069), .o(n_25070) );
na02s06 g755176 ( .a(n_25045), .b(FE_OCP_DRV_N1472_n_25044), .o(n_25069) );
no02s01 g755177 ( .a(n_25049), .b(n_25020), .o(n_25021) );
na02s01 g755178 ( .a(n_25145), .b(n_25176), .o(n_25335) );
no02f04 g755179 ( .a(n_25114), .b(n_23892), .o(n_25268) );
in01s01 g755180 ( .a(n_25203), .o(n_25204) );
in01s01 g755181 ( .a(n_25175), .o(n_25203) );
na02f08 g755183 ( .a(n_25145), .b(n_25144), .o(n_25146) );
oa12s01 g755185 ( .a(n_25194), .b(n_25660), .c(n_25052), .o(n_25717) );
in01s01 g755186 ( .a(n_25715), .o(n_25688) );
na02f06 g755187 ( .a(n_25640), .b(n_25218), .o(n_25715) );
in01m02 g755188 ( .a(n_25098), .o(n_25099) );
no02s01 TIMEBOOST_cell_3114 ( .a(n_9956), .b(n_9875), .o(TIMEBOOST_net_848) );
no02s04 TIMEBOOST_cell_2970 ( .a(n_24857), .b(n_22207), .o(TIMEBOOST_net_776) );
ao12s01 g755192 ( .a(n_24978), .b(n_24977), .c(n_24976), .o(n_26626) );
in01s01 g755193 ( .a(n_25745), .o(n_26512) );
ao12s01 g755194 ( .a(n_25608), .b(n_25607), .c(n_25606), .o(n_25745) );
in01s01 g755195 ( .a(n_25712), .o(n_25713) );
ao12s01 g755196 ( .a(n_25642), .b(n_25660), .c(n_25641), .o(n_25712) );
in01s02 g755205 ( .a(n_25373), .o(n_25551) );
in01m03 g755207 ( .a(FE_OCP_RBN5901_n_25178), .o(n_25373) );
no02m06 g755230 ( .a(n_24992), .b(FE_OCP_RBN5815_n_24823), .o(n_25042) );
na02s02 TIMEBOOST_cell_6837 ( .a(n_16908), .b(n_16909), .o(TIMEBOOST_net_2176) );
na02m04 g755232 ( .a(n_24992), .b(n_24805), .o(n_24993) );
no02m08 TIMEBOOST_cell_6932 ( .a(TIMEBOOST_net_2224), .b(n_14540), .o(TIMEBOOST_net_1077) );
no02m02 TIMEBOOST_cell_4083 ( .a(FE_RN_2434_0), .b(FE_OCP_RBN3098_n_15561), .o(TIMEBOOST_net_1132) );
oa12m04 g755235 ( .a(n_24691), .b(n_24970), .c(n_24896), .o(n_25041) );
no02s01 g755236 ( .a(n_25607), .b(n_25606), .o(n_25608) );
no02s01 g755237 ( .a(n_25660), .b(n_25641), .o(n_25642) );
na02f06 g755238 ( .a(n_25095), .b(n_23890), .o(n_25145) );
na02m08 g755239 ( .a(n_25096), .b(n_23891), .o(n_25176) );
no02s01 g755240 ( .a(n_24977), .b(n_24976), .o(n_24978) );
na02s01 g755241 ( .a(n_25686), .b(n_25685), .o(n_25687) );
na02s01 g755242 ( .a(n_25018), .b(n_24987), .o(n_25073) );
ao12m06 g755244 ( .a(n_24842), .b(n_24975), .c(n_24803), .o(n_24990) );
in01s01 g755245 ( .a(n_25640), .o(n_25714) );
no02m04 TIMEBOOST_cell_2964 ( .a(n_18870), .b(n_18513), .o(TIMEBOOST_net_773) );
in01s04 g755247 ( .a(n_25016), .o(n_25017) );
in01m04 g755248 ( .a(n_24989), .o(n_25016) );
ao12f06 g755249 ( .a(n_24881), .b(n_24975), .c(n_24823), .o(n_24989) );
oa22m04 g755251 ( .a(n_24899), .b(n_24757), .c(n_24898), .d(n_24756), .o(n_25023) );
in01m02 g755252 ( .a(n_24945), .o(n_24946) );
oa12f08 g755254 ( .a(n_24851), .b(n_24974), .c(n_24892), .o(n_25049) );
ao12s01 g755255 ( .a(n_24942), .b(n_24941), .c(n_24974), .o(n_26656) );
no02f04 g755257 ( .a(n_25040), .b(n_25015), .o(n_25114) );
no02f04 g755260 ( .a(n_25011), .b(n_24799), .o(n_25040) );
no02s03 g755261 ( .a(n_24986), .b(n_24819), .o(n_25015) );
in01s02 g755262 ( .a(n_25038), .o(n_25039) );
oa12f04 g755263 ( .a(n_24966), .b(n_24937), .c(n_24971), .o(n_25038) );
na02s01 g755264 ( .a(n_25120), .b(n_25529), .o(n_25660) );
in01s01 g755266 ( .a(n_24972), .o(n_24987) );
no02s04 g755267 ( .a(n_24944), .b(n_24943), .o(n_24972) );
na02s04 g755268 ( .a(n_24944), .b(n_24943), .o(n_25018) );
no02s01 g755270 ( .a(n_24941), .b(n_24974), .o(n_24942) );
na02s01 g755271 ( .a(n_25144), .b(n_25094), .o(n_25279) );
no02s01 g755272 ( .a(n_26310), .b(n_25683), .o(n_25684) );
no02f01 TIMEBOOST_cell_2963 ( .a(n_19537), .b(TIMEBOOST_net_772), .o(n_19694) );
ao12s01 g755275 ( .a(n_25521), .b(n_25638), .c(n_25548), .o(n_25607) );
in01m04 g755277 ( .a(n_25095), .o(n_25096) );
na02s02 TIMEBOOST_cell_4235 ( .a(n_1730), .b(n_1729), .o(TIMEBOOST_net_1208) );
ao12s01 g755280 ( .a(n_24940), .b(n_24939), .c(n_24938), .o(n_25013) );
oa12s01 g755281 ( .a(n_24859), .b(n_24877), .c(n_24923), .o(n_24977) );
in01s01 g755282 ( .a(n_25686), .o(n_26417) );
oa12s01 g755283 ( .a(n_25581), .b(n_25580), .c(n_25579), .o(n_25686) );
ao12s01 g755284 ( .a(n_25639), .b(n_25638), .c(n_25637), .o(n_26451) );
no02m10 g755285 ( .a(n_24900), .b(n_24808), .o(n_24975) );
in01m02 g755287 ( .a(n_24986), .o(n_25011) );
na02f08 g755288 ( .a(n_24915), .b(n_24971), .o(n_24986) );
na02s01 g755289 ( .a(n_25580), .b(n_25579), .o(n_25581) );
no02s01 g755290 ( .a(n_25638), .b(n_25637), .o(n_25639) );
no02f08 g755291 ( .a(n_24861), .b(n_24887), .o(n_24924) );
no02s01 g755292 ( .a(n_25066), .b(n_24969), .o(n_25184) );
na02m06 g755293 ( .a(n_25065), .b(n_25064), .o(n_25144) );
in01s01 g755294 ( .a(n_25246), .o(n_25094) );
no02m06 g755295 ( .a(n_25065), .b(n_25064), .o(n_25246) );
no02f08 TIMEBOOST_cell_4234 ( .a(n_41083), .b(TIMEBOOST_net_1207), .o(n_41110) );
na02s04 g755297 ( .a(n_24967), .b(n_24774), .o(n_24985) );
no02m04 g755298 ( .a(n_24971), .b(n_24964), .o(n_24970) );
no02s01 g755299 ( .a(n_24939), .b(n_24938), .o(n_24940) );
in01s02 g755300 ( .a(n_24921), .o(n_24922) );
na02s04 g755301 ( .a(n_24900), .b(n_24729), .o(n_24921) );
in01m02 g755302 ( .a(n_24898), .o(n_24899) );
ao12s04 g755303 ( .a(n_24788), .b(n_24787), .c(n_24660), .o(n_24898) );
in01s01 g755304 ( .a(n_25528), .o(n_25529) );
ao12f08 g755307 ( .a(n_24536), .b(n_24787), .c(n_24535), .o(n_24862) );
oa12f08 g755309 ( .a(n_24822), .b(n_24897), .c(n_24776), .o(n_24974) );
ao12s01 g755310 ( .a(n_24884), .b(n_24883), .c(n_24897), .o(n_26587) );
in01m02 g755311 ( .a(n_25036), .o(n_25037) );
ao12s01 g755313 ( .a(n_24882), .b(n_24920), .c(FE_RN_2389_0), .o(n_24976) );
ao12s01 g755314 ( .a(n_24880), .b(n_24879), .c(n_24878), .o(n_26528) );
in01s01 g755315 ( .a(n_25685), .o(n_25547) );
oa12s01 g755316 ( .a(n_25473), .b(n_25472), .c(n_25471), .o(n_25685) );
oa12s01 g755317 ( .a(n_25578), .b(n_25577), .c(n_25576), .o(n_26310) );
na02s01 g755318 ( .a(n_25472), .b(n_25471), .o(n_25473) );
na02s01 g755319 ( .a(n_25577), .b(n_25576), .o(n_25578) );
na02m06 g755320 ( .a(n_24810), .b(n_24754), .o(n_24842) );
in01s01 g755321 ( .a(n_25470), .o(n_25638) );
ao12f04 g755322 ( .a(n_25223), .b(n_25410), .c(n_25084), .o(n_25470) );
no02s01 g755324 ( .a(n_24984), .b(n_25035), .o(n_25107) );
no02s01 g755325 ( .a(n_24897), .b(n_24883), .o(n_24884) );
no02m06 g755326 ( .a(n_24935), .b(n_23669), .o(n_25066) );
in01s04 g755328 ( .a(n_24969), .o(n_25008) );
no02m04 g755329 ( .a(n_24934), .b(FE_OCP_DRV_N1900_n_23668), .o(n_24969) );
na02m08 g755330 ( .a(n_24918), .b(n_24876), .o(n_24971) );
no02s01 g755331 ( .a(n_24887), .b(n_24923), .o(n_24939) );
no02s01 g755332 ( .a(n_24920), .b(FE_RN_2389_0), .o(n_24882) );
na02f04 g755333 ( .a(n_24810), .b(n_24829), .o(n_24881) );
no02s01 g755334 ( .a(n_24879), .b(n_24878), .o(n_24880) );
na02m08 g755335 ( .a(n_24787), .b(n_24705), .o(n_24900) );
in01m02 g755336 ( .a(n_24967), .o(n_24968) );
na02s01 TIMEBOOST_cell_6099 ( .a(FE_OCP_RBN4146_n_7743), .b(FE_OCP_RBN2599_n_7743), .o(TIMEBOOST_net_1901) );
in01s01 g755339 ( .a(n_24877), .o(n_24938) );
in01s01 g755340 ( .a(n_24861), .o(n_24877) );
ao12f06 g755341 ( .a(n_24837), .b(n_24760), .c(n_24784), .o(n_24861) );
no02f02 TIMEBOOST_cell_8605 ( .a(TIMEBOOST_net_2789), .b(n_20508), .o(n_20597) );
no02s02 TIMEBOOST_cell_8819 ( .a(TIMEBOOST_net_2896), .b(n_5242), .o(TIMEBOOST_net_1637) );
no02s01 g755344 ( .a(n_25410), .b(n_25142), .o(n_25472) );
na02s01 g755345 ( .a(n_25410), .b(n_24997), .o(n_25409) );
na02s02 TIMEBOOST_cell_6989 ( .a(n_19238), .b(n_20375), .o(TIMEBOOST_net_2253) );
no02s04 g755347 ( .a(n_24910), .b(n_24620), .o(n_24937) );
ao12m08 g755351 ( .a(n_24788), .b(n_24699), .c(n_22207), .o(n_24810) );
in01s03 g755352 ( .a(n_24860), .o(n_24923) );
na02f06 g755353 ( .a(n_24839), .b(n_24838), .o(n_24860) );
in01s01 g755354 ( .a(n_24887), .o(n_24859) );
no02f06 g755355 ( .a(n_24839), .b(n_24838), .o(n_24887) );
in01s01 g755356 ( .a(n_24983), .o(n_24984) );
na02m06 g755357 ( .a(n_24963), .b(FE_OCPN1922_n_24962), .o(n_24983) );
no02s08 g755358 ( .a(n_24963), .b(FE_OCPN1922_n_24962), .o(n_25035) );
na02s01 g755359 ( .a(n_24914), .b(n_24961), .o(n_25020) );
na02m04 g755360 ( .a(n_24911), .b(n_24680), .o(n_24936) );
no02s01 g755362 ( .a(n_24785), .b(n_24837), .o(n_24879) );
oa12s01 g755363 ( .a(n_25031), .b(n_25494), .c(n_25436), .o(n_25577) );
in01s02 g755365 ( .a(n_24787), .o(n_24836) );
na02f10 g755368 ( .a(n_24703), .b(n_24702), .o(n_24787) );
oa12m04 g755369 ( .a(n_22393), .b(n_24875), .c(n_24874), .o(n_24876) );
in01s02 g755371 ( .a(n_24896), .o(n_24915) );
ao12f04 g755372 ( .a(FE_OCPN5128_n_22280), .b(n_24875), .c(n_24874), .o(n_24896) );
na02m04 g755373 ( .a(n_24829), .b(n_24692), .o(n_24895) );
na02s06 g755374 ( .a(n_24766), .b(n_46963), .o(n_24920) );
oa12f08 g755375 ( .a(n_24711), .b(n_24834), .c(n_24775), .o(n_24897) );
ao12s01 g755376 ( .a(n_24833), .b(n_24832), .c(n_24834), .o(n_26530) );
in01m02 g755377 ( .a(n_24934), .o(n_24935) );
in01f04 g755379 ( .a(n_24932), .o(n_24933) );
no03f04 TIMEBOOST_cell_374 ( .a(n_45134), .b(n_15271), .c(n_15559), .o(n_15706) );
oa12s01 g755382 ( .a(n_24763), .b(n_24762), .c(n_24761), .o(n_26468) );
oa12s01 g755383 ( .a(n_25574), .b(n_25573), .c(n_25572), .o(n_26348) );
in01s01 g755384 ( .a(n_25683), .o(n_25575) );
oa12s01 g755385 ( .a(n_25495), .b(n_25494), .c(n_25493), .o(n_25683) );
no02f04 g755386 ( .a(n_25494), .b(n_24996), .o(n_25410) );
na02s01 g755387 ( .a(n_25494), .b(n_25493), .o(n_25495) );
no02s02 TIMEBOOST_cell_4369 ( .a(n_8696), .b(FE_OCP_RBN4138_n_7743), .o(TIMEBOOST_net_1275) );
no02m06 g755390 ( .a(n_24704), .b(n_24659), .o(n_24705) );
oa12m08 g755391 ( .a(n_22111), .b(n_24701), .c(n_24507), .o(n_24703) );
no02s02 g755392 ( .a(n_24788), .b(n_24726), .o(n_24729) );
no02s02 TIMEBOOST_cell_5612 ( .a(FE_OCPN945_n_27287), .b(n_27170), .o(TIMEBOOST_net_1754) );
no02f04 g755394 ( .a(n_24872), .b(n_22393), .o(n_24873) );
na02s01 g755395 ( .a(n_25573), .b(n_25572), .o(n_25574) );
no02f04 g755396 ( .a(n_24765), .b(n_24764), .o(n_24837) );
in01s01 g755397 ( .a(n_24784), .o(n_24785) );
na02f04 g755398 ( .a(n_24765), .b(n_24764), .o(n_24784) );
na02m06 g755399 ( .a(n_24894), .b(n_24893), .o(n_24961) );
in01s01 g755400 ( .a(n_24913), .o(n_24914) );
no02s08 g755401 ( .a(n_24894), .b(n_24893), .o(n_24913) );
no02s01 g755402 ( .a(n_24832), .b(n_24834), .o(n_24833) );
no02s01 g755403 ( .a(n_24852), .b(n_24892), .o(n_24941) );
na02s01 g755404 ( .a(n_24762), .b(n_24761), .o(n_24763) );
ao12m08 g755405 ( .a(n_24626), .b(n_24701), .c(n_24466), .o(n_24702) );
in01s02 g755406 ( .a(n_24830), .o(n_24831) );
no02s01 TIMEBOOST_cell_4199 ( .a(n_37085), .b(n_36929), .o(TIMEBOOST_net_1190) );
in01s02 g755408 ( .a(n_24911), .o(n_24912) );
in01s02 g755409 ( .a(n_24918), .o(n_24911) );
na02f04 TIMEBOOST_cell_3186 ( .a(n_15704), .b(n_15408), .o(TIMEBOOST_net_884) );
in01m02 g755415 ( .a(n_24868), .o(n_24869) );
no02f04 TIMEBOOST_cell_8870 ( .a(n_39642), .b(n_45188), .o(TIMEBOOST_net_2922) );
no02s06 TIMEBOOST_cell_3094 ( .a(n_29248), .b(n_29204), .o(TIMEBOOST_net_838) );
in01s01 g755418 ( .a(n_24760), .o(n_24878) );
na02m08 g755420 ( .a(n_24867), .b(n_24853), .o(n_24963) );
in01s01 g755421 ( .a(n_25440), .o(n_25441) );
oa12s01 g755422 ( .a(n_25348), .b(n_25347), .c(n_25346), .o(n_25440) );
in01s01 g755423 ( .a(n_26230), .o(n_25605) );
oa12s01 g755424 ( .a(n_25527), .b(n_25526), .c(n_25525), .o(n_26230) );
in01s06 g755425 ( .a(n_24910), .o(n_24964) );
in01s06 g755426 ( .a(n_24891), .o(n_24910) );
na02s01 g755428 ( .a(n_25347), .b(n_25346), .o(n_25348) );
na02s01 g755429 ( .a(n_25526), .b(n_25525), .o(n_25527) );
no02m04 TIMEBOOST_cell_4264 ( .a(TIMEBOOST_net_1222), .b(n_19390), .o(TIMEBOOST_net_1046) );
no02m06 TIMEBOOST_cell_5365 ( .a(TIMEBOOST_net_1630), .b(FE_OCP_RBN6804_n_9742), .o(n_9992) );
no02s10 g755432 ( .a(n_22207), .b(n_24687), .o(n_24808) );
na02m06 g755433 ( .a(n_24655), .b(n_24652), .o(n_24699) );
na03f08 TIMEBOOST_cell_8359 ( .a(n_35424), .b(n_35358), .c(n_35447), .o(n_35501) );
no02s02 g755435 ( .a(n_24802), .b(n_24752), .o(n_24805) );
na02s06 g755436 ( .a(n_24754), .b(n_24803), .o(n_24804) );
no02f20 TIMEBOOST_cell_4198 ( .a(n_40664), .b(TIMEBOOST_net_1189), .o(FE_RN_107_0) );
in01s02 g755438 ( .a(n_24756), .o(n_24757) );
no02s02 g755439 ( .a(n_24704), .b(n_24726), .o(n_24756) );
na02m04 g755440 ( .a(n_24874), .b(FE_OCPN5128_n_22280), .o(n_24828) );
no02s02 TIMEBOOST_cell_5518 ( .a(n_5677), .b(n_5911), .o(TIMEBOOST_net_1707) );
na02s02 g755442 ( .a(n_24750), .b(n_24691), .o(n_24783) );
ao12f04 g755443 ( .a(n_25111), .b(n_25224), .c(n_25057), .o(n_25494) );
na02s06 g755445 ( .a(n_24820), .b(n_24632), .o(n_24853) );
na02m06 g755446 ( .a(n_24821), .b(n_24612), .o(n_24867) );
in01s01 g755447 ( .a(n_24851), .o(n_24852) );
na02m04 g755448 ( .a(n_24826), .b(n_24825), .o(n_24851) );
no02m04 g755449 ( .a(n_24826), .b(n_24825), .o(n_24892) );
na02s01 g755450 ( .a(n_24698), .b(n_24661), .o(n_24762) );
in01s02 g755453 ( .a(n_24659), .o(n_24660) );
ao12m08 g755454 ( .a(n_24624), .b(n_24602), .c(n_24601), .o(n_24659) );
no02m04 TIMEBOOST_cell_4562 ( .a(TIMEBOOST_net_1371), .b(n_36545), .o(TIMEBOOST_net_1177) );
na02f04 TIMEBOOST_cell_8803 ( .a(TIMEBOOST_net_2888), .b(n_15476), .o(n_15652) );
in01s02 g755458 ( .a(n_24870), .o(n_24850) );
ao12s01 g755460 ( .a(n_25113), .b(n_25262), .c(n_25088), .o(n_25573) );
oa12f08 g755461 ( .a(n_24713), .b(n_24779), .c(n_24636), .o(n_24834) );
na02m04 TIMEBOOST_cell_4349 ( .a(n_42100), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(TIMEBOOST_net_1265) );
na03f06 TIMEBOOST_cell_8291 ( .a(FE_OCP_RBN2642_n_13667), .b(FE_RN_145_0), .c(n_13851), .o(n_46984) );
ao12s01 g755465 ( .a(n_24781), .b(n_24780), .c(n_24779), .o(n_24848) );
in01f02 g755466 ( .a(n_24857), .o(n_24872) );
na02s01 g755469 ( .a(n_25261), .b(n_25112), .o(n_25347) );
in01s03 g755470 ( .a(n_24656), .o(n_24657) );
no02f06 g755471 ( .a(n_24579), .b(n_24626), .o(n_24656) );
in01s01 TIMEBOOST_cell_7388 ( .a(n_36750), .o(TIMEBOOST_net_2324) );
na02s02 g755473 ( .a(n_24581), .b(n_24267), .o(n_24604) );
in01s02 g755474 ( .a(n_24655), .o(n_24726) );
na02m06 g755475 ( .a(n_24623), .b(n_24624), .o(n_24655) );
no02s06 TIMEBOOST_cell_3180 ( .a(n_35005), .b(n_30612), .o(TIMEBOOST_net_881) );
in01s06 g755477 ( .a(n_24803), .o(n_24802) );
na02m10 g755478 ( .a(FE_OCP_RBN6681_n_24648), .b(FE_OCPN1920_n_22393), .o(n_24803) );
no02s02 g755479 ( .a(n_24694), .b(FE_OCPN1354_n_22484), .o(n_24695) );
no02s04 g755480 ( .a(n_24778), .b(n_24518), .o(n_24782) );
na02s02 TIMEBOOST_cell_8853 ( .a(TIMEBOOST_net_2913), .b(n_5783), .o(FE_RN_2283_0) );
no02m04 g755483 ( .a(n_24694), .b(n_24691), .o(n_24692) );
na02s02 g755484 ( .a(n_24694), .b(FE_OCPN1354_n_22484), .o(n_24690) );
in01s01 g755486 ( .a(n_24754), .o(n_24752) );
na02s08 g755487 ( .a(n_24648), .b(n_24620), .o(n_24754) );
no02s06 g755488 ( .a(n_24623), .b(n_24624), .o(n_24704) );
na02s06 g755490 ( .a(n_24577), .b(n_23360), .o(n_24698) );
na02f02 g755491 ( .a(n_24576), .b(n_23359), .o(n_24661) );
na02s01 g755492 ( .a(n_24777), .b(n_24822), .o(n_24883) );
no02s01 g755493 ( .a(n_24779), .b(n_24780), .o(n_24781) );
ao12s01 g755494 ( .a(n_24982), .b(n_25468), .c(n_25407), .o(n_25526) );
in01s01 g755496 ( .a(n_24701), .o(n_24653) );
no02m10 g755497 ( .a(n_24578), .b(n_24318), .o(n_24701) );
in01m04 g755498 ( .a(n_24820), .o(n_24821) );
in01m04 g755499 ( .a(n_24800), .o(n_24820) );
in01s02 g755501 ( .a(n_24687), .o(n_24688) );
in01s06 g755502 ( .a(n_24652), .o(n_24687) );
no02m08 g755503 ( .a(n_24539), .b(n_24580), .o(n_24652) );
in01s01 g755508 ( .a(FE_OCPN1081_n_24819), .o(n_24865) );
in01s01 g755511 ( .a(n_24799), .o(n_24819) );
in01f06 g755512 ( .a(n_24799), .o(n_24798) );
no02s06 TIMEBOOST_cell_1949 ( .a(FE_OCPN1653_n_23078), .b(n_23044), .o(TIMEBOOST_net_589) );
in01m02 g755514 ( .a(n_24750), .o(n_24751) );
na02s02 TIMEBOOST_cell_7922 ( .a(n_4995), .b(n_4596), .o(TIMEBOOST_net_2592) );
in01s01 g755517 ( .a(n_26307), .o(n_26855) );
oa12s01 g755518 ( .a(n_25469), .b(n_25468), .c(n_25467), .o(n_26307) );
in01s02 g755519 ( .a(n_24874), .o(n_24797) );
no02m08 g755520 ( .a(n_24722), .b(n_24685), .o(n_24874) );
na02s01 g755521 ( .a(n_25468), .b(n_25467), .o(n_25469) );
in01s01 g755522 ( .a(n_25261), .o(n_25262) );
in01s01 g755523 ( .a(n_25224), .o(n_25261) );
no02f04 g755524 ( .a(n_25172), .b(n_24995), .o(n_25224) );
na02m04 TIMEBOOST_cell_8016 ( .a(n_5636), .b(n_6265), .o(TIMEBOOST_net_2639) );
in01m02 g755527 ( .a(n_24581), .o(n_24582) );
no02s02 TIMEBOOST_cell_2041 ( .a(n_3120), .b(n_2451), .o(TIMEBOOST_net_635) );
no02s04 g755529 ( .a(n_24510), .b(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24539) );
no02m08 g755530 ( .a(FE_OCP_RBN2704_n_24510), .b(FE_OCPN1916_n_22111), .o(n_24580) );
no02s02 TIMEBOOST_cell_4001 ( .a(n_4194), .b(n_4200), .o(TIMEBOOST_net_1091) );
na02m04 TIMEBOOST_cell_2038 ( .a(TIMEBOOST_net_633), .b(FE_OCP_RBN2668_n_29500), .o(n_29604) );
no02s04 g755533 ( .a(n_24638), .b(n_22207), .o(n_24685) );
no02m08 g755534 ( .a(n_24680), .b(FE_OFN742_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24722) );
na02m06 g755535 ( .a(n_24748), .b(FE_OCP_DRV_N1420_n_24747), .o(n_24822) );
in01s01 g755536 ( .a(n_24776), .o(n_24777) );
no02s08 g755537 ( .a(n_24748), .b(FE_OCP_DRV_N1420_n_24747), .o(n_24776) );
no02s01 g755538 ( .a(n_24712), .b(n_24775), .o(n_24832) );
in01f02 g755539 ( .a(n_24720), .o(n_24721) );
no02s04 TIMEBOOST_cell_2042 ( .a(TIMEBOOST_net_635), .b(n_3141), .o(n_4336) );
in01m02 g755541 ( .a(n_24578), .o(n_24579) );
in01s02 g755543 ( .a(n_24778), .o(n_24746) );
na02m08 g755544 ( .a(n_24719), .b(n_24497), .o(n_24778) );
na02s01 TIMEBOOST_cell_2840 ( .a(FE_RN_2566_0), .b(n_7093), .o(TIMEBOOST_net_711) );
in01s02 g755546 ( .a(n_24576), .o(n_24577) );
oa22f02 g755547 ( .a(FE_OCP_RBN1822_n_24473), .b(n_25318), .c(n_24473), .d(n_24204), .o(n_24576) );
na02f06 g755548 ( .a(n_24508), .b(n_24472), .o(n_24761) );
ao12s01 g755550 ( .a(n_24716), .b(n_24715), .c(n_24714), .o(n_26428) );
in01s01 g755553 ( .a(FE_OCP_RBN5718_n_24718), .o(n_24774) );
no02s20 TIMEBOOST_cell_5948 ( .a(TIMEBOOST_net_1825), .b(FE_OCP_RBN5530_n_1541), .o(n_1614) );
ao12s01 g755556 ( .a(n_24569), .b(n_24568), .c(FE_OCP_RBN1163_n_24471), .o(n_26360) );
no02s01 TIMEBOOST_cell_6051 ( .a(n_13463), .b(n_13464), .o(TIMEBOOST_net_1877) );
na02m06 g755559 ( .a(n_24573), .b(n_24537), .o(n_24694) );
na02m10 g755560 ( .a(n_24477), .b(n_24452), .o(n_24602) );
in01s01 g755564 ( .a(n_24717), .o(n_24794) );
in01s02 g755568 ( .a(n_24684), .o(n_24717) );
na02s02 TIMEBOOST_cell_7966 ( .a(FE_OCP_RBN4457_n_43103), .b(n_43199), .o(TIMEBOOST_net_2614) );
na02m06 TIMEBOOST_cell_7078 ( .a(TIMEBOOST_net_2297), .b(n_10988), .o(n_11058) );
no02m02 TIMEBOOST_cell_2016 ( .a(TIMEBOOST_net_622), .b(n_14163), .o(n_14279) );
no02s02 g755575 ( .a(n_24626), .b(n_24368), .o(n_24574) );
na02s06 g755576 ( .a(n_24436), .b(FE_OCPN1916_n_22111), .o(n_24452) );
na02s04 g755577 ( .a(FE_OCP_RBN2708_n_24505), .b(FE_OCPN1920_n_22393), .o(n_24573) );
na02f02 g755578 ( .a(n_24505), .b(n_24620), .o(n_24537) );
no02s02 g755579 ( .a(n_24534), .b(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24536) );
na02s02 g755580 ( .a(n_24534), .b(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24535) );
na02s06 g755582 ( .a(n_24506), .b(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24532) );
na02m08 g755583 ( .a(FE_OCP_RBN2694_n_24436), .b(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24477) );
no02s06 TIMEBOOST_cell_8839 ( .a(TIMEBOOST_net_2906), .b(n_35751), .o(FE_RN_2668_0) );
no02s02 TIMEBOOST_cell_2839 ( .a(TIMEBOOST_net_710), .b(n_33061), .o(n_33143) );
na02m04 g755586 ( .a(n_24451), .b(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24476) );
no02m08 g755588 ( .a(n_24683), .b(FE_OCPN1318_n_24682), .o(n_24775) );
no02s01 g755589 ( .a(n_24715), .b(n_24714), .o(n_24716) );
na02s01 g755590 ( .a(n_24637), .b(n_24713), .o(n_24780) );
no02s01 g755591 ( .a(FE_OCP_RBN2695_n_24436), .b(n_24529), .o(n_24531) );
no02s01 g755592 ( .a(n_24469), .b(FE_OCP_RBN2666_n_24372), .o(n_24570) );
no02s01 g755593 ( .a(n_24555), .b(n_45633), .o(n_24642) );
na02s01 g755594 ( .a(n_24555), .b(n_45633), .o(n_24639) );
no02s01 g755595 ( .a(n_24568), .b(FE_OCP_RBN1163_n_24471), .o(n_24569) );
in01s01 g755596 ( .a(n_24711), .o(n_24712) );
na02f06 g755597 ( .a(n_24683), .b(FE_OCPN1318_n_24682), .o(n_24711) );
na02s02 g755598 ( .a(n_25310), .b(n_25345), .o(n_25408) );
in01s01 g755599 ( .a(n_25172), .o(n_25468) );
ao12f02 g755600 ( .a(n_25062), .b(n_25093), .c(n_24953), .o(n_25172) );
na02f06 TIMEBOOST_cell_8074 ( .a(n_45010), .b(FE_OCP_RBN1843_n_20640), .o(TIMEBOOST_net_2668) );
na02s02 TIMEBOOST_cell_2834 ( .a(n_7048), .b(n_7049), .o(TIMEBOOST_net_708) );
in01s01 g755604 ( .a(FE_OCP_RBN2704_n_24510), .o(n_25531) );
na02s06 TIMEBOOST_cell_4169 ( .a(FE_RN_2887_0), .b(FE_RN_2884_0), .o(TIMEBOOST_net_1175) );
in01s02 g755612 ( .a(n_24680), .o(n_24959) );
in01m06 g755613 ( .a(n_24638), .o(n_24680) );
na02s06 TIMEBOOST_cell_4236 ( .a(n_1847), .b(TIMEBOOST_net_1208), .o(n_1921) );
in01s02 g755615 ( .a(n_24621), .o(n_24650) );
oa22m02 g755616 ( .a(FE_OCP_RBN4184_n_24467), .b(n_24048), .c(n_24467), .d(n_24049), .o(n_24621) );
in01m04 g755617 ( .a(n_24598), .o(n_24646) );
na02s04 TIMEBOOST_cell_2037 ( .a(n_29527), .b(n_25859), .o(TIMEBOOST_net_633) );
na03m02 TIMEBOOST_cell_3526 ( .a(n_19030), .b(FE_OCP_RBN1130_n_18918), .c(n_18978), .o(n_19139) );
na02m06 g755621 ( .a(n_24465), .b(n_24367), .o(n_24507) );
na02s06 TIMEBOOST_cell_2833 ( .a(n_7258), .b(TIMEBOOST_net_707), .o(n_7335) );
na02s08 TIMEBOOST_cell_4168 ( .a(TIMEBOOST_net_1174), .b(n_40538), .o(n_40561) );
na02s04 g755626 ( .a(n_24471), .b(n_24502), .o(n_24472) );
in01s01 g755627 ( .a(n_24636), .o(n_24637) );
no02m08 g755628 ( .a(n_24614), .b(n_24613), .o(n_24636) );
na02f06 g755629 ( .a(n_24614), .b(n_24613), .o(n_24713) );
in01s04 g755630 ( .a(n_24562), .o(n_24563) );
ao12m06 g755631 ( .a(n_23850), .b(n_24463), .c(n_23708), .o(n_24562) );
no02s01 g755632 ( .a(n_24593), .b(n_24554), .o(n_24715) );
no02s01 g755633 ( .a(n_24546), .b(n_24633), .o(n_24635) );
no02m04 g755634 ( .a(n_24566), .b(n_24560), .o(n_24561) );
na02m02 TIMEBOOST_cell_2052 ( .a(TIMEBOOST_net_640), .b(FE_OCP_RBN6640_n_24268), .o(n_24405) );
oa12s01 g755636 ( .a(n_25188), .b(n_25286), .c(n_24979), .o(n_25345) );
in01s01 g755649 ( .a(FE_OCP_RBN2695_n_24436), .o(n_24469) );
in01s01 g755653 ( .a(FE_OCP_RBN2709_n_24505), .o(n_25104) );
oa22m02 g755656 ( .a(n_24406), .b(n_24051), .c(n_24405), .d(n_24050), .o(n_24505) );
in01s02 g755660 ( .a(n_24612), .o(n_24632) );
in01s01 g755662 ( .a(n_24556), .o(n_24714) );
oa12f04 g755663 ( .a(n_24443), .b(n_24549), .c(n_24494), .o(n_24556) );
na02s01 TIMEBOOST_cell_5224 ( .a(n_34748), .b(n_34705), .o(TIMEBOOST_net_1560) );
oa12s01 g755665 ( .a(n_24551), .b(n_24550), .c(n_24549), .o(n_26296) );
oa12s01 g755666 ( .a(n_24448), .b(n_24447), .c(n_24446), .o(n_26248) );
in01s01 g755667 ( .a(n_26419), .o(n_25524) );
ao12s02 g755668 ( .a(n_25439), .b(n_25438), .c(n_25437), .o(n_26419) );
ao12s01 g755669 ( .a(n_24449), .b(n_24503), .c(n_24502), .o(n_24568) );
in01s01 g755673 ( .a(FE_OCP_RBN2715_n_24501), .o(n_24555) );
in01s06 g755676 ( .a(n_24534), .o(n_24601) );
no02s03 TIMEBOOST_cell_2992 ( .a(n_14194), .b(n_13257), .o(TIMEBOOST_net_787) );
ao12f06 g755679 ( .a(n_24321), .b(n_24347), .c(n_21975), .o(n_24473) );
no02f08 g755680 ( .a(n_24500), .b(n_23921), .o(n_24566) );
na02f02 g755681 ( .a(n_25063), .b(n_25092), .o(n_25093) );
no02s01 g755682 ( .a(n_25438), .b(n_25437), .o(n_25439) );
na02s01 g755683 ( .a(n_25371), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_25372) );
no02s01 g755684 ( .a(n_25371), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_25370) );
na02m02 g755685 ( .a(n_24500), .b(n_24498), .o(n_24499) );
na02s06 TIMEBOOST_cell_2029 ( .a(n_41978), .b(n_41774), .o(TIMEBOOST_net_629) );
no02m08 TIMEBOOST_cell_2991 ( .a(n_19329), .b(TIMEBOOST_net_786), .o(n_19414) );
no02m08 TIMEBOOST_cell_8495 ( .a(TIMEBOOST_net_2734), .b(n_32999), .o(n_33022) );
no02f06 TIMEBOOST_cell_2971 ( .a(TIMEBOOST_net_776), .b(n_24873), .o(n_24932) );
na02m06 g755690 ( .a(n_24461), .b(FE_OFN743_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24497) );
na02s02 g755691 ( .a(n_25311), .b(n_25368), .o(n_25369) );
no02s01 g755692 ( .a(n_25343), .b(n_25220), .o(n_25344) );
na02f08 TIMEBOOST_cell_2030 ( .a(TIMEBOOST_net_629), .b(n_41973), .o(n_42005) );
in01s01 g755695 ( .a(n_24553), .o(n_24554) );
na02f04 g755696 ( .a(n_24484), .b(n_23282), .o(n_24553) );
in01s01 g755697 ( .a(n_24592), .o(n_24593) );
na02m06 g755698 ( .a(n_24485), .b(n_23283), .o(n_24592) );
na02m08 TIMEBOOST_cell_6204 ( .a(TIMEBOOST_net_1953), .b(FE_OCP_RBN1822_n_24473), .o(n_24578) );
na02s01 g755700 ( .a(n_24549), .b(n_24550), .o(n_24551) );
no02s01 g755701 ( .a(n_24503), .b(n_24502), .o(n_24449) );
na02s01 g755702 ( .a(n_24446), .b(n_24447), .o(n_24448) );
na02s06 g755703 ( .a(n_24520), .b(n_24429), .o(n_24522) );
in01m04 g755704 ( .a(n_24547), .o(n_24548) );
no02s06 g755705 ( .a(n_24520), .b(n_24519), .o(n_24521) );
no02m06 g755706 ( .a(n_24520), .b(n_24519), .o(n_24547) );
no02s01 TIMEBOOST_cell_8501 ( .a(TIMEBOOST_net_2737), .b(n_23740), .o(FE_RN_218_0) );
na02m08 g755709 ( .a(n_24326), .b(n_23886), .o(n_24408) );
na02s06 TIMEBOOST_cell_4167 ( .a(n_40248), .b(n_40437), .o(TIMEBOOST_net_1174) );
in01s01 g755713 ( .a(n_24590), .o(n_24591) );
oa12s01 g755714 ( .a(n_24493), .b(n_24492), .c(n_24491), .o(n_24590) );
in01s03 g755715 ( .a(n_24465), .o(n_24466) );
in01s01 g755720 ( .a(n_24518), .o(n_24546) );
no02s06 g755722 ( .a(n_24346), .b(n_24014), .o(n_24375) );
na02s10 g755723 ( .a(n_24402), .b(n_24052), .o(n_24407) );
no02s02 g755724 ( .a(n_24325), .b(n_23885), .o(n_24327) );
na02s04 g755725 ( .a(n_24297), .b(n_23972), .o(n_24348) );
na02s06 g755726 ( .a(n_24325), .b(n_23820), .o(n_24326) );
in01s01 g755727 ( .a(n_25063), .o(n_25438) );
no02f02 g755728 ( .a(n_25006), .b(n_24954), .o(n_25063) );
no02m02 g755729 ( .a(n_25007), .b(n_25092), .o(n_25062) );
no02s06 g755730 ( .a(n_24462), .b(n_24305), .o(n_24464) );
na02f06 TIMEBOOST_cell_4166 ( .a(TIMEBOOST_net_1173), .b(n_40538), .o(n_40563) );
no02s01 TIMEBOOST_cell_3821 ( .a(n_46217), .b(n_46218), .o(TIMEBOOST_net_1001) );
in01s01 g755733 ( .a(n_25311), .o(n_25312) );
no02s01 g755734 ( .a(n_25222), .b(n_25771), .o(n_25311) );
na02s01 g755735 ( .a(n_25112), .b(n_25089), .o(n_25113) );
oa12m04 g755737 ( .a(n_23883), .b(n_24274), .c(FE_OCPN1721_n_23818), .o(n_24323) );
in01s02 g755738 ( .a(n_24405), .o(n_24406) );
no02f06 TIMEBOOST_cell_6701 ( .a(FE_OCP_RBN1595_n_14823), .b(FE_OCP_RBN4226_n_13962), .o(TIMEBOOST_net_2108) );
no02s01 g755741 ( .a(n_24444), .b(n_24494), .o(n_24550) );
na02s01 g755742 ( .a(n_24492), .b(n_24491), .o(n_24493) );
in01s01 g755744 ( .a(n_25309), .o(n_25310) );
oa12s01 g755745 ( .a(n_25290), .b(n_25192), .c(n_25160), .o(n_25309) );
na02s04 g755747 ( .a(n_25112), .b(n_25058), .o(n_25111) );
ao12s02 g755748 ( .a(n_25119), .b(n_25032), .c(n_25082), .o(n_25143) );
na02s02 g755749 ( .a(n_25219), .b(n_25161), .o(n_25343) );
na02s01 g755750 ( .a(n_24404), .b(n_24373), .o(n_24447) );
no02s06 TIMEBOOST_cell_8682 ( .a(n_21264), .b(FE_OCPN1382_n_45026), .o(TIMEBOOST_net_2828) );
in01m06 g755752 ( .a(n_24489), .o(n_24490) );
in01m06 g755753 ( .a(n_24463), .o(n_24489) );
no02m06 g755754 ( .a(n_24445), .b(n_23999), .o(n_24463) );
in01m04 g755756 ( .a(n_24520), .o(n_24488) );
na02m10 g755757 ( .a(n_24462), .b(n_24339), .o(n_24520) );
oa12s01 g755758 ( .a(n_25221), .b(n_25259), .c(n_25160), .o(n_26234) );
in01s01 g755759 ( .a(n_25286), .o(n_25287) );
ao12s01 g755760 ( .a(n_25160), .b(n_25259), .c(n_25258), .o(n_25286) );
in01s01 g755764 ( .a(n_24486), .o(n_24633) );
in01s02 g755765 ( .a(n_24461), .o(n_24486) );
oa22m06 g755766 ( .a(n_24364), .b(n_23846), .c(n_24363), .d(n_23847), .o(n_24461) );
in01m02 g755767 ( .a(n_24484), .o(n_24485) );
na03s06 TIMEBOOST_cell_5877 ( .a(n_22149), .b(FE_OCPN7089_n_20979), .c(n_22187), .o(n_22268) );
ao12f04 g755769 ( .a(n_24442), .b(n_24393), .c(n_24336), .o(n_24549) );
in01s01 g755770 ( .a(n_24432), .o(n_24433) );
oa12s01 g755771 ( .a(n_24343), .b(n_24342), .c(n_24341), .o(n_24432) );
in01s01 g755775 ( .a(FE_OCP_RBN2665_n_24372), .o(n_24529) );
no04m04 TIMEBOOST_cell_5809 ( .a(n_9658), .b(n_9404), .c(n_9657), .d(n_9405), .o(n_9907) );
in01s01 g755779 ( .a(n_25371), .o(n_25342) );
ao12s02 g755780 ( .a(n_25257), .b(n_25256), .c(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_25371) );
in01s01 g755781 ( .a(n_26162), .o(n_26192) );
oa12s01 g755782 ( .a(n_25061), .b(n_25060), .c(n_25059), .o(n_26162) );
in01s02 g755783 ( .a(n_24398), .o(n_24399) );
in01s01 TIMEBOOST_cell_7383 ( .a(TIMEBOOST_net_2318), .o(TIMEBOOST_net_2319) );
in01s02 g755785 ( .a(n_24369), .o(n_24370) );
no03f10 TIMEBOOST_cell_2216 ( .a(n_28068), .b(n_28067), .c(n_28120), .o(n_28192) );
in01s06 g755787 ( .a(n_24346), .o(n_24402) );
no02s10 g755788 ( .a(FE_OCP_RBN6640_n_24268), .b(n_24040), .o(n_24346) );
in01s02 g755789 ( .a(n_24325), .o(n_24297) );
no02m08 g755791 ( .a(n_24396), .b(n_23878), .o(n_24445) );
in01f01 g755792 ( .a(n_25006), .o(n_25007) );
no02f02 g755793 ( .a(n_24929), .b(n_24958), .o(n_25006) );
na02s01 g755794 ( .a(n_25060), .b(n_25059), .o(n_25061) );
no02s01 g755795 ( .a(n_25256), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_25257) );
in01s04 g755796 ( .a(n_24344), .o(n_24345) );
no02m06 g755797 ( .a(n_24322), .b(n_21975), .o(n_24344) );
no02m04 g755798 ( .a(n_24320), .b(n_24319), .o(n_24321) );
na02m01 TIMEBOOST_cell_5959 ( .a(FE_RN_1397_0), .b(FE_RN_1396_0), .o(TIMEBOOST_net_1831) );
no02f06 TIMEBOOST_cell_5325 ( .a(TIMEBOOST_net_1610), .b(n_10543), .o(n_10629) );
no02s03 g755801 ( .a(n_24293), .b(n_22111), .o(n_24318) );
in01s01 g755802 ( .a(n_24367), .o(n_24368) );
na02s04 g755803 ( .a(n_24310), .b(n_22111), .o(n_24367) );
no02m08 g755804 ( .a(n_24429), .b(n_22089), .o(n_24519) );
in01s01 g755805 ( .a(n_25221), .o(n_25222) );
na02s01 g755806 ( .a(n_25259), .b(n_25160), .o(n_25221) );
no02s03 g755807 ( .a(n_24274), .b(n_23926), .o(n_24272) );
na02f02 g755808 ( .a(n_24291), .b(n_23278), .o(n_24373) );
na02f06 g755809 ( .a(n_24292), .b(n_23279), .o(n_24404) );
na02s01 TIMEBOOST_cell_2003 ( .a(n_496), .b(n_484), .o(TIMEBOOST_net_616) );
no02s01 TIMEBOOST_cell_8858 ( .a(n_31716), .b(FE_RN_372_0), .o(TIMEBOOST_net_2916) );
in01s01 g755812 ( .a(n_24443), .o(n_24444) );
na02f04 g755813 ( .a(n_24426), .b(FE_OCPN5284_n_24425), .o(n_24443) );
no02s01 g755815 ( .a(n_24442), .b(n_24394), .o(n_24492) );
na02s01 g755816 ( .a(n_25316), .b(FE_OCPN1096_n_25318), .o(n_24316) );
na02s01 g755817 ( .a(n_24342), .b(n_24341), .o(n_24343) );
na03s02 TIMEBOOST_cell_6556 ( .a(FE_OCP_RBN4482_n_11439), .b(FE_OCPN3592_n_45301), .c(n_11451), .o(n_11600) );
na02f06 TIMEBOOST_cell_2020 ( .a(TIMEBOOST_net_624), .b(n_18876), .o(n_18981) );
in01m02 g755820 ( .a(n_24423), .o(n_24424) );
na02s04 g755821 ( .a(n_24396), .b(n_24017), .o(n_24423) );
in01f04 g755822 ( .a(n_24462), .o(n_24441) );
no02f10 g755823 ( .a(n_24360), .b(n_24289), .o(n_24462) );
oa12s01 g755824 ( .a(n_25368), .b(n_25160), .c(n_25304), .o(n_26237) );
no03m02 TIMEBOOST_cell_7892 ( .a(n_4407), .b(FE_RN_1939_0), .c(FE_RN_1940_0), .o(TIMEBOOST_net_2577) );
in01s01 g755828 ( .a(n_25142), .o(n_25169) );
no02s04 g755829 ( .a(n_25087), .b(n_25032), .o(n_25142) );
oa12s02 g755830 ( .a(n_25188), .b(n_25220), .c(n_25124), .o(n_25288) );
na02s02 g755831 ( .a(n_25005), .b(n_24998), .o(n_25058) );
na02s02 g755832 ( .a(n_25004), .b(n_24994), .o(n_25112) );
oa12s01 g755833 ( .a(n_25188), .b(n_25216), .c(n_24813), .o(n_25219) );
in01s01 g755838 ( .a(n_24395), .o(n_24422) );
in01s06 g755839 ( .a(n_24366), .o(n_24395) );
in01s01 g755842 ( .a(FE_OCPN5290_n_26125), .o(n_26214) );
ao12s01 g755843 ( .a(n_24391), .b(n_24390), .c(n_24389), .o(n_26125) );
no02m08 TIMEBOOST_cell_4940 ( .a(n_23462), .b(FE_RN_1317_0), .o(TIMEBOOST_net_1418) );
in01m04 g755849 ( .a(n_24438), .o(n_24458) );
in01m04 g755850 ( .a(n_24421), .o(n_24438) );
na02m08 g755854 ( .a(n_24340), .b(n_23822), .o(n_24396) );
in01s04 g755855 ( .a(n_24363), .o(n_24364) );
no02s04 g755856 ( .a(n_24340), .b(n_24016), .o(n_24363) );
in01s01 g755857 ( .a(n_24958), .o(n_25059) );
ao12m02 g755858 ( .a(n_24106), .b(n_24906), .c(n_24154), .o(n_24958) );
na02m08 g755859 ( .a(n_24305), .b(FE_OFN741_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24339) );
no02s02 g755860 ( .a(n_25167), .b(n_25134), .o(n_25168) );
na02s01 g755861 ( .a(n_25741), .b(n_25307), .o(n_25308) );
in01s01 g755862 ( .a(n_25199), .o(n_25200) );
no02s01 g755863 ( .a(n_25193), .b(n_25140), .o(n_25199) );
no02s01 TIMEBOOST_cell_3156 ( .a(n_34365), .b(n_34364), .o(TIMEBOOST_net_869) );
no02s02 g755865 ( .a(n_25056), .b(n_25029), .o(n_25057) );
no02s01 g755867 ( .a(n_25164), .b(n_25604), .o(n_25218) );
na02s02 g755868 ( .a(n_25197), .b(n_25162), .o(n_25198) );
no02s01 g755869 ( .a(n_25284), .b(n_25340), .o(n_25341) );
no02s01 g755870 ( .a(n_25195), .b(n_25216), .o(n_25196) );
na02s01 g755871 ( .a(n_25194), .b(n_25081), .o(n_25641) );
na02s01 g755872 ( .a(n_25306), .b(n_25166), .o(n_26072) );
no02s01 g755873 ( .a(n_25193), .b(n_25220), .o(n_25839) );
na02s01 g755874 ( .a(n_24955), .b(n_24930), .o(n_25060) );
na02s01 g755875 ( .a(n_25089), .b(n_25088), .o(n_25346) );
no02s01 g755876 ( .a(n_25217), .b(n_25216), .o(n_25799) );
no02s01 g755877 ( .a(n_25771), .b(n_25735), .o(n_26134) );
no02s01 g755878 ( .a(n_25055), .b(n_25033), .o(n_25471) );
no02s01 g755879 ( .a(n_25191), .b(n_25285), .o(n_25192) );
no02s02 g755881 ( .a(n_25086), .b(n_25085), .o(n_25087) );
na02s02 g755882 ( .a(n_25089), .b(n_24299), .o(n_25005) );
na02s02 g755883 ( .a(n_25003), .b(n_25002), .o(n_25004) );
no02s01 g755884 ( .a(n_25055), .b(n_25083), .o(n_25084) );
na02s01 g755885 ( .a(n_25081), .b(n_24605), .o(n_25082) );
na02s01 g755886 ( .a(n_25160), .b(n_25304), .o(n_25368) );
no02s01 g755887 ( .a(n_25436), .b(n_25086), .o(n_25493) );
na02s01 g755888 ( .a(n_25407), .b(n_25003), .o(n_25467) );
na02s01 g755889 ( .a(n_25522), .b(n_25548), .o(n_25637) );
no02s01 g755890 ( .a(n_25570), .b(n_25604), .o(n_25689) );
na02s01 g755891 ( .a(n_25254), .b(FE_RN_697_0), .o(n_25905) );
na02s01 g755892 ( .a(n_25741), .b(n_25680), .o(n_25950) );
no02f04 g755893 ( .a(n_24362), .b(FE_OCP_DRV_N1884_n_24361), .o(n_24442) );
in01s01 g755894 ( .a(n_24393), .o(n_24394) );
na02f04 g755895 ( .a(n_24362), .b(FE_OCP_DRV_N1884_n_24361), .o(n_24393) );
na02s01 g755896 ( .a(n_24305), .b(FE_OCP_RBN5671_n_24288), .o(n_24392) );
na02s01 g755897 ( .a(n_24419), .b(n_25386), .o(n_24420) );
no02s01 g755898 ( .a(n_24390), .b(n_24389), .o(n_24391) );
no02s03 TIMEBOOST_cell_4163 ( .a(n_32149), .b(FE_RN_369_0), .o(TIMEBOOST_net_1172) );
in01f02 g755900 ( .a(n_24311), .o(n_24312) );
in01f01 g755901 ( .a(n_24320), .o(n_24311) );
na02s02 TIMEBOOST_cell_7505 ( .a(TIMEBOOST_net_2383), .b(n_420), .o(n_446) );
in01m08 g755903 ( .a(n_24359), .o(n_24360) );
oa12s01 g755906 ( .a(n_25030), .b(n_25160), .c(n_25090), .o(n_25579) );
in01s01 g755907 ( .a(n_25710), .o(n_25711) );
oa12s01 g755908 ( .a(n_25307), .b(n_25160), .c(n_25251), .o(n_25710) );
ao12s01 g755909 ( .a(n_25056), .b(n_25160), .c(n_25001), .o(n_25572) );
ao12s01 g755910 ( .a(n_25053), .b(n_25188), .c(n_25028), .o(n_25606) );
ao12s01 g755911 ( .a(n_25167), .b(n_25188), .c(n_25122), .o(n_25716) );
oa12s01 g755912 ( .a(n_25163), .b(n_25160), .c(n_25133), .o(n_25772) );
oa12s01 g755913 ( .a(n_25197), .b(n_25160), .c(n_25132), .o(n_25802) );
oa12s01 g755914 ( .a(n_25141), .b(n_25160), .c(n_24844), .o(n_25883) );
in01s01 g755915 ( .a(n_25708), .o(n_25709) );
oa12s01 g755916 ( .a(n_25253), .b(n_25160), .c(n_25135), .o(n_25708) );
in01s01 g755917 ( .a(n_25739), .o(n_25740) );
ao12s01 g755918 ( .a(n_25340), .b(n_25188), .c(n_25285), .o(n_25739) );
in01s02 g755921 ( .a(n_24310), .o(n_24386) );
in01s06 g755925 ( .a(n_24293), .o(n_24310) );
oa12m04 g755927 ( .a(n_24143), .b(n_24270), .c(n_24144), .o(n_24446) );
in01f02 g755928 ( .a(n_24291), .o(n_24292) );
in01s01 g755930 ( .a(n_24457), .o(n_25390) );
in01s02 g755931 ( .a(n_24429), .o(n_24457) );
no02m08 g755934 ( .a(n_24309), .b(n_24290), .o(n_24429) );
oa12s01 g755936 ( .a(n_24250), .b(n_24270), .c(n_24249), .o(n_24342) );
oa22s01 g755937 ( .a(n_25188), .b(n_24153), .c(n_25139), .d(n_24131), .o(n_25256) );
ao12s01 g755938 ( .a(n_24909), .b(n_24908), .c(n_24907), .o(n_25259) );
oa22s01 g755939 ( .a(n_25160), .b(n_25085), .c(n_25188), .d(n_24382), .o(n_25576) );
oa22s01 g755940 ( .a(n_25160), .b(n_24236), .c(n_25188), .d(n_25092), .o(n_25437) );
ao22s01 g755941 ( .a(n_25160), .b(n_24258), .c(n_25188), .d(n_25002), .o(n_25525) );
in01s06 g755943 ( .a(n_24274), .o(n_24268) );
na02f06 TIMEBOOST_cell_8038 ( .a(n_31477), .b(n_31504), .o(TIMEBOOST_net_2650) );
no02f06 g755945 ( .a(n_24210), .b(n_24185), .o(n_24319) );
in01s01 g755946 ( .a(n_24267), .o(n_25316) );
in01s02 g755948 ( .a(n_24254), .o(n_24267) );
in01s03 g755963 ( .a(n_29630), .o(n_25859) );
in01s40 g755967 ( .a(n_29561), .o(n_29630) );
in01s40 g755972 ( .a(FE_OFN774_n_25834), .o(n_29561) );
in01s06 g755973 ( .a(FE_OFN774_n_25834), .o(n_25738) );
in01s02 g755979 ( .a(FE_OFN774_n_25834), .o(n_29379) );
na02s02 TIMEBOOST_cell_8717 ( .a(TIMEBOOST_net_2845), .b(n_1843), .o(n_1905) );
no02s04 g755983 ( .a(n_24264), .b(n_23789), .o(n_24290) );
no02m06 g755984 ( .a(n_24265), .b(n_23788), .o(n_24309) );
no02s01 g755987 ( .a(n_24908), .b(n_24907), .o(n_24909) );
no02s04 g755988 ( .a(n_24165), .b(FE_OFN743_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24185) );
no02f04 g755989 ( .a(FE_OCP_RBN1018_n_24165), .b(n_21852), .o(n_24210) );
no03m02 TIMEBOOST_cell_7746 ( .a(n_4743), .b(n_4609), .c(FE_RN_1915_0), .o(TIMEBOOST_net_2504) );
in01s01 g755991 ( .a(n_24229), .o(n_24230) );
na02s06 g755992 ( .a(n_24178), .b(n_21852), .o(n_24229) );
no02s06 TIMEBOOST_cell_4162 ( .a(TIMEBOOST_net_1171), .b(n_32087), .o(n_32219) );
no02s06 g755994 ( .a(n_24288), .b(n_21975), .o(n_24289) );
na02s02 TIMEBOOST_cell_7923 ( .a(TIMEBOOST_net_2592), .b(n_5064), .o(n_5243) );
in01s01 g755996 ( .a(n_25570), .o(n_25571) );
no02s01 g755997 ( .a(n_25160), .b(n_25129), .o(n_25570) );
in01s01 g755998 ( .a(n_25521), .o(n_25522) );
no02s01 g755999 ( .a(n_25160), .b(n_25109), .o(n_25521) );
na02s01 g756000 ( .a(n_25188), .b(n_24275), .o(n_25407) );
no02s02 g756001 ( .a(n_24994), .b(n_25001), .o(n_25056) );
na02s02 g756002 ( .a(n_24956), .b(n_24957), .o(n_25089) );
no02s01 g756003 ( .a(n_25160), .b(n_25000), .o(n_25436) );
na02s01 g756004 ( .a(n_25160), .b(n_25251), .o(n_25307) );
in01s01 g756005 ( .a(n_25003), .o(n_24982) );
na02s03 g756006 ( .a(n_24956), .b(n_24257), .o(n_25003) );
no02s01 g756007 ( .a(n_25188), .b(n_25285), .o(n_25340) );
in01s01 g756008 ( .a(n_25679), .o(n_25680) );
no02s01 g756009 ( .a(n_25160), .b(n_25250), .o(n_25679) );
in01s01 g756010 ( .a(n_25140), .o(n_25141) );
no02s01 g756011 ( .a(n_25032), .b(n_25124), .o(n_25140) );
in01s01 g756012 ( .a(n_25735), .o(n_25736) );
no02s01 g756013 ( .a(n_25160), .b(n_25258), .o(n_25735) );
in01s01 g756014 ( .a(n_25191), .o(n_25166) );
no02s01 g756015 ( .a(n_25139), .b(n_25138), .o(n_25191) );
na02s01 g756016 ( .a(n_25160), .b(n_25250), .o(n_25741) );
no02s01 g756017 ( .a(n_25026), .b(n_24768), .o(n_25220) );
no02s01 g756019 ( .a(n_25026), .b(n_25136), .o(n_25189) );
no02s01 g756020 ( .a(n_25032), .b(n_24767), .o(n_25193) );
na02s01 g756021 ( .a(n_25139), .b(n_25136), .o(n_25254) );
na02s01 g756022 ( .a(n_25139), .b(n_25135), .o(n_25253) );
no02s01 g756023 ( .a(n_25032), .b(n_25122), .o(n_25167) );
in01s01 g756024 ( .a(n_25134), .o(n_25194) );
no02s01 g756025 ( .a(n_25188), .b(n_25027), .o(n_25134) );
in01s01 g756026 ( .a(n_25031), .o(n_25086) );
na02s02 g756027 ( .a(n_24953), .b(n_25000), .o(n_25031) );
in01s01 g756028 ( .a(n_25033), .o(n_24999) );
no02s01 g756029 ( .a(n_24981), .b(n_24980), .o(n_25033) );
in01s02 g756030 ( .a(n_25030), .o(n_25083) );
na02s01 g756031 ( .a(n_24998), .b(n_25090), .o(n_25030) );
in01s01 g756032 ( .a(n_25029), .o(n_25088) );
no02s01 g756033 ( .a(n_24956), .b(n_24957), .o(n_25029) );
in01s01 g756034 ( .a(n_24929), .o(n_24930) );
no02s02 g756035 ( .a(n_24906), .b(n_23836), .o(n_24929) );
in01s01 g756036 ( .a(n_24954), .o(n_24955) );
no02s02 g756037 ( .a(n_24902), .b(n_23837), .o(n_24954) );
in01s01 g756038 ( .a(n_24997), .o(n_25055) );
na02s01 g756039 ( .a(n_24981), .b(n_24980), .o(n_24997) );
na02s01 g756040 ( .a(n_25026), .b(n_25109), .o(n_25548) );
no02s01 g756042 ( .a(n_25032), .b(n_25028), .o(n_25053) );
in01s01 g756043 ( .a(n_25081), .o(n_25052) );
na02s01 g756044 ( .a(n_25032), .b(n_25027), .o(n_25081) );
in01s01 g756045 ( .a(n_25163), .o(n_25164) );
na02s01 g756046 ( .a(n_25026), .b(n_25133), .o(n_25163) );
no02s01 g756047 ( .a(n_25032), .b(n_24627), .o(n_25604) );
na02s01 g756048 ( .a(n_25139), .b(n_25132), .o(n_25197) );
in01s01 g756049 ( .a(n_25162), .o(n_25217) );
na02s01 g756050 ( .a(n_25026), .b(n_25130), .o(n_25162) );
no02s01 g756051 ( .a(n_25026), .b(n_25130), .o(n_25216) );
in01s01 g756052 ( .a(n_25306), .o(n_25284) );
na02s01 g756053 ( .a(n_25160), .b(n_25138), .o(n_25306) );
no02s01 g756054 ( .a(n_25188), .b(n_24901), .o(n_25771) );
na02s01 g756055 ( .a(n_24270), .b(n_24249), .o(n_24250) );
in01s02 g756056 ( .a(n_24307), .o(n_24308) );
na02s06 g756057 ( .a(n_24285), .b(n_23947), .o(n_24307) );
in01s01 g756058 ( .a(n_25195), .o(n_25161) );
ao12s01 g756059 ( .a(n_25139), .b(n_25133), .c(n_25129), .o(n_25195) );
na02s01 g756060 ( .a(n_25188), .b(n_24793), .o(n_25290) );
ao12s01 g756061 ( .a(n_24998), .b(n_25085), .c(n_25000), .o(n_24996) );
no02s02 g756062 ( .a(n_24994), .b(n_24276), .o(n_24995) );
in01s01 g756063 ( .a(n_25119), .o(n_25120) );
ao12s01 g756064 ( .a(n_25026), .b(n_24541), .c(n_25109), .o(n_25119) );
na02m04 TIMEBOOST_cell_5148 ( .a(TIMEBOOST_net_1078), .b(n_38592), .o(TIMEBOOST_net_1522) );
in01s01 g756066 ( .a(n_24336), .o(n_24491) );
oa12m04 g756067 ( .a(n_24159), .b(n_24306), .c(n_24160), .o(n_24336) );
oa12s01 g756068 ( .a(n_24284), .b(n_24306), .c(n_24283), .o(n_24390) );
in01s01 g756069 ( .a(n_24979), .o(n_25304) );
oa12s01 g756070 ( .a(n_24905), .b(n_24904), .c(n_24903), .o(n_24979) );
in01s02 g756073 ( .a(n_24305), .o(n_24419) );
na02s06 g756078 ( .a(n_24183), .b(n_23734), .o(n_24208) );
in01m02 g756079 ( .a(n_24264), .o(n_24265) );
no02s04 g756080 ( .a(n_24248), .b(n_23946), .o(n_24264) );
no03s04 TIMEBOOST_cell_8391 ( .a(n_10770), .b(n_10390), .c(TIMEBOOST_net_1329), .o(n_10852) );
na02m08 g756082 ( .a(n_24248), .b(n_23762), .o(n_24285) );
na02s01 g756083 ( .a(n_24904), .b(n_24903), .o(n_24905) );
ao12s06 g756084 ( .a(n_23713), .b(n_24145), .c(n_23768), .o(n_24166) );
oa12s02 g756085 ( .a(n_23767), .b(n_24147), .c(n_23736), .o(n_24148) );
no02s06 TIMEBOOST_cell_8482 ( .a(n_11771), .b(n_11909), .o(TIMEBOOST_net_2728) );
no02f04 g756087 ( .a(FE_OCP_RBN1011_n_24246), .b(FE_OCP_RBN1007_n_24175), .o(n_24263) );
na02s01 g756088 ( .a(n_24306), .b(n_24283), .o(n_24284) );
oa12s02 g756089 ( .a(n_24352), .b(n_24864), .c(n_24045), .o(n_24908) );
oa12m02 g756091 ( .a(n_24100), .b(FE_OCP_RBN1020_n_24181), .c(n_21852), .o(n_24207) );
no02s02 TIMEBOOST_cell_1924 ( .a(TIMEBOOST_net_576), .b(n_11582), .o(n_11702) );
in01s02 g756095 ( .a(n_24981), .o(n_24953) );
in01s01 g756098 ( .a(n_24981), .o(n_24994) );
in01s04 g756129 ( .a(n_25188), .o(n_25160) );
in01s06 g756130 ( .a(n_25026), .o(n_25188) );
in01s02 g756132 ( .a(n_25032), .o(n_25139) );
in01s06 g756136 ( .a(n_25032), .o(n_25026) );
in01s06 g756137 ( .a(n_24998), .o(n_25032) );
in01s06 g756138 ( .a(n_24981), .o(n_24998) );
in01m08 g756139 ( .a(n_24956), .o(n_24981) );
in01m06 g756140 ( .a(n_24902), .o(n_24956) );
in01m04 g756141 ( .a(n_24906), .o(n_24902) );
no02f08 TIMEBOOST_cell_2014 ( .a(TIMEBOOST_net_621), .b(n_24646), .o(n_24723) );
in01s03 g756145 ( .a(FE_OCP_RBN1019_n_24165), .o(n_25265) );
in01s01 g756150 ( .a(n_24204), .o(n_25318) );
in01s03 g756151 ( .a(n_24178), .o(n_24204) );
oa22s06 g756152 ( .a(n_24145), .b(n_23790), .c(n_24147), .d(n_23791), .o(n_24178) );
oa22s02 g756153 ( .a(n_24181), .b(n_24100), .c(FE_OCP_RBN1020_n_24181), .d(n_24099), .o(n_24270) );
in01s01 g756154 ( .a(FE_OCP_RBN5671_n_24288), .o(n_25386) );
no02s01 TIMEBOOST_cell_1993 ( .a(n_38209), .b(n_37889), .o(TIMEBOOST_net_611) );
in01s01 g756160 ( .a(n_25258), .o(n_24901) );
ao12s01 g756161 ( .a(n_24846), .b(n_24864), .c(n_24845), .o(n_25258) );
no02s02 TIMEBOOST_cell_5613 ( .a(TIMEBOOST_net_1754), .b(n_27378), .o(n_27488) );
na02s02 TIMEBOOST_cell_1987 ( .a(n_29036), .b(n_28703), .o(TIMEBOOST_net_608) );
no02s06 TIMEBOOST_cell_8876 ( .a(FE_OCP_RBN3078_n_25816), .b(n_27086), .o(TIMEBOOST_net_2925) );
no02s01 g756167 ( .a(n_24864), .b(n_24845), .o(n_24846) );
no02m08 g756168 ( .a(n_24101), .b(n_21852), .o(n_24146) );
na02f04 TIMEBOOST_cell_5583 ( .a(TIMEBOOST_net_1739), .b(n_11139), .o(n_11297) );
no03f04 TIMEBOOST_cell_6525 ( .a(n_26198), .b(n_23447), .c(n_26219), .o(TIMEBOOST_net_1990) );
no02s02 g756171 ( .a(FE_OCP_RBN1021_n_24181), .b(FE_OCPN871_n_24098), .o(n_24201) );
na02s01 g756172 ( .a(n_25251), .b(n_25250), .o(n_24793) );
na02s06 g756173 ( .a(n_24145), .b(FE_OCPN1302_n_23771), .o(n_24183) );
in01s04 g756174 ( .a(n_24224), .o(n_24225) );
no02s06 TIMEBOOST_cell_1868 ( .a(TIMEBOOST_net_548), .b(n_40116), .o(n_40120) );
ao12f08 g756178 ( .a(n_22089), .b(n_24121), .c(n_24157), .o(n_24246) );
oa12s01 g756180 ( .a(n_24817), .b(n_24816), .c(n_24815), .o(n_25285) );
in01s01 g756181 ( .a(FE_OCP_RBN4157_n_24222), .o(n_24332) );
in01s02 g756189 ( .a(n_24145), .o(n_24127) );
in01s06 g756190 ( .a(n_24147), .o(n_24145) );
no02s06 TIMEBOOST_cell_5368 ( .a(FE_OCPN1705_n_14730), .b(FE_OCPN1733_n_14524), .o(TIMEBOOST_net_1632) );
na02m08 g756193 ( .a(n_24164), .b(n_23733), .o(n_24200) );
no02s02 g756194 ( .a(n_24164), .b(n_24162), .o(n_24163) );
na02s01 g756195 ( .a(n_24816), .b(n_24815), .o(n_24817) );
in01s01 g756196 ( .a(n_24791), .o(n_24792) );
na02f06 g756197 ( .a(n_24742), .b(n_24090), .o(n_24791) );
na02s02 g756198 ( .a(n_24743), .b(n_24192), .o(n_24864) );
in01f03 g756199 ( .a(n_24084), .o(n_24085) );
oa12f06 g756200 ( .a(n_23634), .b(n_24072), .c(n_23638), .o(n_24084) );
no02s04 g756201 ( .a(n_24341), .b(n_24142), .o(n_24144) );
na02s02 g756202 ( .a(n_24341), .b(FE_OCPN1346_n_24142), .o(n_24143) );
no02s01 g756203 ( .a(FE_OCP_RBN4149_n_24173), .b(FE_OCP_RBN1001_n_24079), .o(n_24221) );
in01s01 g756206 ( .a(n_24102), .o(n_24125) );
in01s04 g756207 ( .a(n_24102), .o(n_24101) );
in01s01 g756219 ( .a(n_24218), .o(n_24219) );
ao22s01 g756220 ( .a(n_24093), .b(n_24097), .c(FE_OCPN871_n_24098), .d(n_22752), .o(n_24218) );
ao12s01 g756221 ( .a(n_24677), .b(n_24676), .c(n_24675), .o(n_25251) );
ao12s01 g756222 ( .a(n_24741), .b(n_24740), .c(n_24739), .o(n_25138) );
in01s01 g756223 ( .a(n_25124), .o(n_24844) );
oa12s01 g756224 ( .a(n_24771), .b(n_24770), .c(n_24769), .o(n_25124) );
ao12s01 g756225 ( .a(n_24708), .b(n_24707), .c(n_24706), .o(n_25136) );
ao12s01 g756227 ( .a(n_24738), .b(n_24737), .c(n_24736), .o(n_25135) );
in01s01 g756228 ( .a(n_24813), .o(n_25132) );
oa12s01 g756229 ( .a(n_24735), .b(n_24734), .c(n_24733), .o(n_24813) );
na02m02 g756230 ( .a(n_24056), .b(n_23662), .o(n_24071) );
na03s02 TIMEBOOST_cell_8405 ( .a(FE_OCP_RBN4483_n_11439), .b(FE_OCP_RBN3330_n_11087), .c(n_11579), .o(n_11743) );
no02m08 g756232 ( .a(n_24122), .b(n_23679), .o(n_24164) );
in01s01 g756233 ( .a(n_24742), .o(n_24743) );
no02f06 g756234 ( .a(n_24355), .b(n_24670), .o(n_24742) );
no02s01 g756235 ( .a(n_24740), .b(n_24739), .o(n_24741) );
no02s01 g756236 ( .a(n_24707), .b(n_24706), .o(n_24708) );
in01m01 g756237 ( .a(n_24099), .o(n_24100) );
no02f04 g756240 ( .a(n_24070), .b(n_22089), .o(n_24099) );
no02s01 g756241 ( .a(n_24676), .b(n_24675), .o(n_24677) );
na02s01 g756242 ( .a(n_24770), .b(n_24769), .o(n_24771) );
no02s01 g756243 ( .a(n_24737), .b(n_24736), .o(n_24738) );
na02s01 g756244 ( .a(n_24734), .b(n_24733), .o(n_24735) );
na02s02 g756245 ( .a(FE_OCP_RBN5615_n_24070), .b(n_24097), .o(n_24341) );
no02s03 g756246 ( .a(n_24389), .b(FE_OCP_DRV_N1426_n_24158), .o(n_24160) );
na02s02 g756247 ( .a(n_24389), .b(FE_OCP_DRV_N1426_n_24158), .o(n_24159) );
no02s04 TIMEBOOST_cell_6695 ( .a(n_7895), .b(n_7957), .o(TIMEBOOST_net_2105) );
no02s02 TIMEBOOST_cell_1865 ( .a(n_40007), .b(FE_OCP_RBN6154_n_39816), .o(TIMEBOOST_net_547) );
oa22s01 g756252 ( .a(FE_OCP_RBN1003_n_24079), .b(n_22767), .c(FE_OCP_RBN1002_n_24079), .d(n_24119), .o(n_26090) );
ao12s01 g756253 ( .a(n_24666), .b(n_24665), .c(n_24664), .o(n_25250) );
in01s01 g756254 ( .a(n_24767), .o(n_24768) );
oa12s01 g756255 ( .a(n_24669), .b(n_24668), .c(n_24667), .o(n_24767) );
ao12s01 g756256 ( .a(n_24630), .b(n_24629), .c(n_24628), .o(n_25133) );
ao12s01 g756257 ( .a(n_24674), .b(n_24673), .c(n_24672), .o(n_25130) );
in01s01 g756261 ( .a(FE_OCP_RBN4149_n_24173), .o(n_24217) );
in01s04 g756263 ( .a(n_24157), .o(n_24173) );
na03f06 TIMEBOOST_cell_2652 ( .a(n_21092), .b(n_21164), .c(n_21016), .o(FE_RN_35_0) );
no02s02 TIMEBOOST_cell_1917 ( .a(n_17451), .b(n_17132), .o(TIMEBOOST_net_573) );
no02m06 g756268 ( .a(n_24080), .b(n_23775), .o(n_24094) );
na02m08 g756269 ( .a(n_24080), .b(n_23682), .o(n_24122) );
no02s01 g756270 ( .a(n_24673), .b(n_24672), .o(n_24674) );
in01s01 g756271 ( .a(n_24670), .o(n_24671) );
na02f06 g756272 ( .a(n_24606), .b(n_24091), .o(n_24670) );
na02s01 g756273 ( .a(n_24607), .b(n_24107), .o(n_24740) );
na02s01 g756274 ( .a(n_24668), .b(n_24667), .o(n_24669) );
no02s01 g756275 ( .a(n_24629), .b(n_24628), .o(n_24630) );
no02s01 g756276 ( .a(n_24665), .b(n_24664), .o(n_24666) );
in01s02 g756278 ( .a(n_24121), .o(n_24137) );
na02f08 g756279 ( .a(n_24079), .b(FE_OFN741_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24121) );
in01s04 g756280 ( .a(n_24072), .o(n_24043) );
no02s03 g756282 ( .a(FE_OCP_RBN1001_n_24079), .b(n_24119), .o(n_24389) );
in01m02 g756283 ( .a(n_24056), .o(n_24057) );
oa12m02 g756284 ( .a(n_23663), .b(n_23949), .c(n_23609), .o(n_24056) );
ao12s01 g756285 ( .a(n_23991), .b(n_24609), .c(n_24006), .o(n_24707) );
na02s01 g756286 ( .a(n_24608), .b(n_23992), .o(n_24737) );
oa12s01 g756287 ( .a(n_23705), .b(n_24586), .c(n_23908), .o(n_24734) );
oa12s01 g756288 ( .a(n_24008), .b(n_24588), .c(n_24074), .o(n_24676) );
no02s02 TIMEBOOST_cell_1862 ( .a(TIMEBOOST_net_545), .b(n_40118), .o(n_40083) );
in01s01 g756293 ( .a(FE_OCPN871_n_24098), .o(n_24093) );
ao22f02 g756295 ( .a(n_23949), .b(n_23688), .c(n_24005), .d(n_23687), .o(n_24070) );
no02s01 TIMEBOOST_cell_8818 ( .a(FE_OCP_RBN6715_n_3604), .b(FE_OCP_RBN4255_n_3705), .o(TIMEBOOST_net_2896) );
no02m08 g756297 ( .a(n_24042), .b(n_23582), .o(n_24080) );
no02s01 g756298 ( .a(n_24585), .b(n_23811), .o(n_24673) );
na02s01 g756299 ( .a(n_24609), .b(n_23862), .o(n_24610) );
na02s01 g756300 ( .a(n_24609), .b(n_24033), .o(n_24608) );
no02s01 g756301 ( .a(n_24609), .b(n_23911), .o(n_24668) );
no02s01 g756302 ( .a(n_24542), .b(n_24036), .o(n_24665) );
in01s01 g756304 ( .a(n_24606), .o(n_24607) );
no02f06 g756305 ( .a(n_24588), .b(n_24062), .o(n_24606) );
oa12s01 g756306 ( .a(n_24235), .b(n_24587), .c(n_24256), .o(n_24629) );
in01s01 g756314 ( .a(n_24605), .o(n_25122) );
ao12s01 g756315 ( .a(n_24515), .b(n_24514), .c(n_24513), .o(n_24605) );
in01s01 g756316 ( .a(n_25129), .o(n_24627) );
ao12s01 g756317 ( .a(n_24544), .b(n_24587), .c(n_24543), .o(n_25129) );
in01m02 g756318 ( .a(n_24042), .o(n_24068) );
na02m08 g756319 ( .a(n_24000), .b(FE_OCPN1362_n_23684), .o(n_24042) );
in01s01 g756320 ( .a(n_24585), .o(n_24586) );
no02s01 g756321 ( .a(n_24587), .b(n_23936), .o(n_24585) );
no02s02 g756322 ( .a(n_24587), .b(n_23957), .o(n_24609) );
no02s01 g756323 ( .a(n_24587), .b(n_24543), .o(n_24544) );
no02s01 g756324 ( .a(n_24514), .b(n_24513), .o(n_24515) );
in01s02 g756326 ( .a(n_23949), .o(n_24005) );
in01s01 g756330 ( .a(n_24588), .o(n_24542) );
na02m06 g756331 ( .a(n_24478), .b(n_24065), .o(n_24588) );
ao12s01 g756332 ( .a(n_23895), .b(n_23930), .c(n_23894), .o(n_25179) );
in01s01 g756333 ( .a(n_24054), .o(n_24055) );
oa12s01 g756334 ( .a(n_24003), .b(n_24002), .c(n_24001), .o(n_24054) );
oa12s01 g756335 ( .a(n_24481), .b(n_24480), .c(n_24479), .o(n_25027) );
in01s01 g756336 ( .a(n_24541), .o(n_25028) );
ao12s01 g756337 ( .a(n_24456), .b(n_24455), .c(n_24454), .o(n_24541) );
na02s01 g756338 ( .a(n_24002), .b(n_24001), .o(n_24003) );
no02s01 g756339 ( .a(n_23930), .b(n_23894), .o(n_23895) );
no02s01 g756340 ( .a(n_24455), .b(n_24454), .o(n_24456) );
in01f02 g756341 ( .a(n_24018), .o(n_24019) );
in01f02 g756342 ( .a(n_24000), .o(n_24018) );
na02s01 g756344 ( .a(n_24480), .b(n_24479), .o(n_24481) );
in01s01 g756345 ( .a(n_24478), .o(n_24587) );
oa12f04 g756346 ( .a(n_24030), .b(n_24453), .c(n_24026), .o(n_24478) );
oa12s01 g756347 ( .a(n_24031), .b(n_24453), .c(n_23981), .o(n_24514) );
na02s01 g756348 ( .a(n_24453), .b(n_23988), .o(n_24480) );
na02s03 g756349 ( .a(n_24066), .b(n_23966), .o(n_24092) );
ao12s01 g756351 ( .a(n_23594), .b(n_23948), .c(n_23635), .o(n_24002) );
ao12s01 g756352 ( .a(n_23955), .b(n_24417), .c(n_24215), .o(n_24455) );
ao12s01 g756354 ( .a(n_23798), .b(n_23827), .c(n_23797), .o(n_23892) );
oa22s01 g756355 ( .a(n_23948), .b(n_23652), .c(n_23889), .d(n_23651), .o(n_25126) );
ao12s01 g756356 ( .a(n_24384), .b(n_24417), .c(n_24383), .o(n_25109) );
ao12s01 g756357 ( .a(n_24416), .b(n_24415), .c(n_24414), .o(n_25090) );
na02f06 g756359 ( .a(n_24417), .b(n_23980), .o(n_24453) );
no02s01 g756360 ( .a(n_24417), .b(n_24383), .o(n_24384) );
na02s03 g756361 ( .a(n_24498), .b(n_23817), .o(n_24560) );
no02s01 g756362 ( .a(n_24415), .b(n_24414), .o(n_24416) );
in01s02 g756363 ( .a(n_24645), .o(n_24066) );
na02m02 g756364 ( .a(n_24498), .b(n_23927), .o(n_24645) );
no02s01 g756365 ( .a(n_23827), .b(n_23797), .o(n_23798) );
in01s01 g756366 ( .a(n_23890), .o(n_23891) );
oa12s01 g756367 ( .a(n_23796), .b(n_23795), .c(n_23794), .o(n_23890) );
in01s01 g756368 ( .a(n_25085), .o(n_24382) );
oa12s01 g756369 ( .a(n_24302), .b(n_24301), .c(n_24300), .o(n_25085) );
ao12s01 g756370 ( .a(n_24381), .b(n_24380), .c(n_24379), .o(n_24980) );
na02s01 g756371 ( .a(n_23795), .b(n_23794), .o(n_23796) );
no02s01 g756372 ( .a(n_24380), .b(n_24379), .o(n_24381) );
na02s01 g756373 ( .a(n_24301), .b(n_24300), .o(n_24302) );
no02s02 g756375 ( .a(n_24016), .b(n_23738), .o(n_24017) );
na02s01 g756376 ( .a(n_23973), .b(n_23856), .o(n_23999) );
in01s01 g756377 ( .a(n_23948), .o(n_23889) );
in01s01 g756378 ( .a(n_23859), .o(n_23948) );
oa12m06 g756380 ( .a(n_23959), .b(n_24277), .c(n_23953), .o(n_24417) );
no02m08 g756381 ( .a(n_24016), .b(n_23857), .o(n_24498) );
in01s01 g756382 ( .a(FE_OCP_DRV_N1476_n_23887), .o(n_23888) );
ao22s01 g756383 ( .a(n_23826), .b(n_23596), .c(n_23777), .d(n_23595), .o(n_23887) );
ao12s01 g756384 ( .a(n_23937), .b(n_24330), .c(n_23952), .o(n_24415) );
na02s01 g756385 ( .a(n_24052), .b(n_24012), .o(n_24053) );
na02s01 g756386 ( .a(n_23692), .b(n_23479), .o(n_23795) );
no02s01 g756387 ( .a(n_24330), .b(n_23958), .o(n_24380) );
no02s02 g756388 ( .a(n_23946), .b(n_23709), .o(n_23947) );
in01s06 g756389 ( .a(n_23973), .o(n_24016) );
no02s06 g756390 ( .a(n_23946), .b(n_23774), .o(n_23973) );
oa12s01 g756391 ( .a(n_23834), .b(FE_OCP_RBN5688_n_24259), .c(n_24169), .o(n_24301) );
oa12s02 g756392 ( .a(n_23695), .b(n_23694), .c(n_23693), .o(n_25064) );
oa12s01 g756393 ( .a(n_24241), .b(FE_OCP_RBN5688_n_24259), .c(n_24240), .o(n_25000) );
no02s02 g756394 ( .a(n_24014), .b(n_23945), .o(n_24015) );
no02s01 g756395 ( .a(n_24014), .b(n_24011), .o(n_24013) );
na02s01 g756396 ( .a(n_23694), .b(n_23693), .o(n_23695) );
in01s01 g756397 ( .a(n_24277), .o(n_24330) );
na02f04 g756398 ( .a(FE_OCP_RBN5687_n_24259), .b(n_23898), .o(n_24277) );
na02s01 g756399 ( .a(FE_OCP_RBN5688_n_24259), .b(n_24240), .o(n_24241) );
in01s01 g756400 ( .a(n_23691), .o(n_23692) );
na02s06 g756403 ( .a(n_23825), .b(n_23741), .o(n_23946) );
oa12s01 g756404 ( .a(FE_OCP_RBN6560_n_23572), .b(n_24011), .c(delay_add_ln22_unr14_stage6_stallmux_q_30_), .o(n_24012) );
in01s01 g756405 ( .a(n_23826), .o(n_23777) );
ao12f08 g756406 ( .a(n_23496), .b(n_23742), .c(n_23541), .o(n_23826) );
in01s01 g756407 ( .a(FE_OCP_DRV_N1474_n_23792), .o(n_23793) );
ao12s01 g756408 ( .a(n_23720), .b(n_23742), .c(n_23719), .o(n_23792) );
no02s01 g756409 ( .a(n_24040), .b(n_23998), .o(n_24041) );
in01s02 g756410 ( .a(n_24014), .o(n_24052) );
na02s06 g756411 ( .a(n_23928), .b(n_23972), .o(n_24014) );
no02s02 g756412 ( .a(n_24040), .b(n_23970), .o(n_23971) );
no02s01 g756413 ( .a(n_23742), .b(n_23719), .o(n_23720) );
in01s01 g756415 ( .a(n_24162), .o(n_23825) );
na02m06 g756416 ( .a(n_23737), .b(n_23739), .o(n_24162) );
oa12m01 g756417 ( .a(n_23856), .b(n_23766), .c(n_23821), .o(n_23857) );
no02s06 TIMEBOOST_cell_7402 ( .a(FE_OCP_RBN5181_n_44061), .b(delay_xor_ln22_unr15_stage6_stallmux_q_0_), .o(TIMEBOOST_net_2332) );
no02s01 g756420 ( .a(n_25002), .b(n_24275), .o(n_24276) );
in01s01 g756421 ( .a(n_23640), .o(n_23694) );
oa12f06 g756422 ( .a(n_23427), .b(n_23615), .c(n_23394), .o(n_23640) );
in01s01 g756423 ( .a(FE_OCP_DRV_N1900_n_23668), .o(n_23669) );
oa12s01 g756424 ( .a(n_23588), .b(n_23615), .c(n_23587), .o(n_23668) );
in01s01 g756425 ( .a(n_24299), .o(n_25001) );
ao12s01 g756426 ( .a(n_24239), .b(n_24238), .c(n_24237), .o(n_24299) );
oa12s01 g756427 ( .a(n_24115), .b(n_24114), .c(n_24113), .o(n_24957) );
na02s01 g756428 ( .a(n_23615), .b(n_23587), .o(n_23588) );
na02s01 g756429 ( .a(n_23997), .b(n_23994), .o(n_24039) );
no02s01 g756430 ( .a(n_24238), .b(n_24237), .o(n_24239) );
na02s03 g756431 ( .a(n_23770), .b(n_23757), .o(n_23824) );
na02s01 g756432 ( .a(n_24114), .b(n_24113), .o(n_24115) );
no03s04 TIMEBOOST_cell_8221 ( .a(n_12666), .b(n_12616), .c(FE_RN_1416_0), .o(FE_RN_1417_0) );
na02s06 g756435 ( .a(n_23855), .b(FE_OCPN1253_n_23815), .o(n_24040) );
ao12f08 g756436 ( .a(n_23471), .b(n_23666), .c(n_23512), .o(n_23742) );
na02f02 g756437 ( .a(n_24112), .b(n_24110), .o(n_24155) );
oa12s02 g756438 ( .a(FE_OCP_RBN6560_n_23572), .b(n_23884), .c(delay_add_ln22_unr14_stage6_stallmux_q_27_), .o(n_23928) );
ao12s01 g756439 ( .a(FE_OCP_RBN6559_n_23572), .b(n_23876), .c(n_22936), .o(n_24011) );
ao12s01 g756440 ( .a(n_23606), .b(n_23761), .c(n_23773), .o(n_23774) );
in01m02 g756442 ( .a(n_23775), .o(n_23739) );
no02s01 TIMEBOOST_cell_8577 ( .a(TIMEBOOST_net_2775), .b(n_21749), .o(n_21780) );
oa12m01 g756444 ( .a(n_23599), .b(n_23738), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_25_), .o(n_23856) );
oa12s01 g756445 ( .a(n_23783), .b(n_23922), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_29_), .o(n_23927) );
oa22s01 g756447 ( .a(n_23602), .b(n_23537), .c(n_23666), .d(n_23538), .o(n_25044) );
in01s01 g756448 ( .a(n_25002), .o(n_24258) );
ao12s01 g756449 ( .a(n_24196), .b(n_24195), .c(n_24194), .o(n_25002) );
in01s02 g756450 ( .a(n_23771), .o(n_23772) );
no02s04 g756451 ( .a(n_23736), .b(n_23735), .o(n_23771) );
no02m01 g756452 ( .a(n_23854), .b(n_23853), .o(n_23855) );
no02s01 g756453 ( .a(n_23885), .b(n_23884), .o(n_23886) );
in01s01 g756454 ( .a(n_23997), .o(n_23998) );
no02s01 g756455 ( .a(n_23969), .b(n_23970), .o(n_23997) );
no02s06 g756457 ( .a(n_23632), .b(n_23664), .o(n_23665) );
no02s01 g756460 ( .a(n_24195), .b(n_24194), .o(n_24196) );
in01s01 g756461 ( .a(n_23769), .o(n_23770) );
na02s02 g756462 ( .a(n_23711), .b(n_23734), .o(n_23769) );
in01s01 g756463 ( .a(n_23925), .o(n_23926) );
na02s01 g756464 ( .a(n_23883), .b(n_23819), .o(n_23925) );
no02s01 g756466 ( .a(n_23758), .b(n_23823), .o(n_23848) );
in01s02 g756467 ( .a(n_23689), .o(n_23690) );
na02s01 TIMEBOOST_cell_6849 ( .a(FE_OCP_RBN3247_n_26169), .b(n_27204), .o(TIMEBOOST_net_2182) );
in01m02 g756469 ( .a(n_23687), .o(n_23688) );
na02m02 g756470 ( .a(n_23663), .b(n_23584), .o(n_23687) );
in01s01 g756471 ( .a(n_23661), .o(n_23662) );
no02s02 g756472 ( .a(n_23639), .b(n_23613), .o(n_23661) );
in01s02 g756473 ( .a(n_23790), .o(n_23791) );
na02s06 g756474 ( .a(n_23768), .b(n_23767), .o(n_23790) );
no02s01 g756476 ( .a(n_23712), .b(n_24182), .o(n_23881) );
na03f08 TIMEBOOST_cell_8356 ( .a(n_45502), .b(n_14420), .c(n_45501), .o(n_15734) );
na02s06 TIMEBOOST_cell_5366 ( .a(n_27131), .b(FE_OCP_RBN6039_n_30733), .o(TIMEBOOST_net_1631) );
no02s02 g756479 ( .a(n_23765), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_27_), .o(n_23766) );
in01s01 g756480 ( .a(n_23923), .o(n_23924) );
no02s01 g756481 ( .a(n_23853), .b(n_23884), .o(n_23923) );
na02m02 g756482 ( .a(FE_OCPN1362_n_23684), .b(n_23656), .o(n_23685) );
no02s02 g756483 ( .a(n_23629), .b(n_23630), .o(n_23718) );
in01s01 g756484 ( .a(n_23967), .o(n_23968) );
no02s02 g756485 ( .a(n_23945), .b(n_23970), .o(n_23967) );
na02f02 g756486 ( .a(FE_OCP_RBN4130_n_24077), .b(n_24111), .o(n_24112) );
in01s01 g756487 ( .a(n_23879), .o(n_23880) );
no02s02 g756488 ( .a(n_23850), .b(n_23765), .o(n_23879) );
in01s02 g756489 ( .a(n_23763), .o(n_23764) );
na02s06 g756490 ( .a(n_23676), .b(n_23733), .o(n_23763) );
in01s01 g756491 ( .a(n_23716), .o(n_23717) );
na02s02 g756492 ( .a(n_23683), .b(n_23682), .o(n_23716) );
in01s01 g756493 ( .a(n_23788), .o(n_23789) );
na02s01 g756494 ( .a(n_23762), .b(n_23761), .o(n_23788) );
in01s01 g756495 ( .a(n_23846), .o(n_23847) );
na02s02 g756496 ( .a(n_23822), .b(n_23675), .o(n_23846) );
in01s01 g756497 ( .a(n_23943), .o(n_23944) );
no02s02 g756498 ( .a(n_23921), .b(n_23922), .o(n_23943) );
in01s01 g756499 ( .a(n_23995), .o(n_23996) );
na02s01 g756500 ( .a(n_23873), .b(n_23966), .o(n_23995) );
in01s02 g756501 ( .a(n_23731), .o(n_23732) );
na02s02 g756502 ( .a(n_23633), .b(n_23659), .o(n_23731) );
in01s01 g756503 ( .a(n_23786), .o(n_23787) );
ao12s02 g756504 ( .a(n_23735), .b(FE_OCP_RBN6557_n_23572), .c(delay_add_ln22_unr14_stage6_stallmux_q_21_), .o(n_23786) );
in01s01 g756505 ( .a(n_23919), .o(n_23920) );
ao12s01 g756506 ( .a(n_23854), .b(FE_OCP_RBN6560_n_23572), .c(delay_add_ln22_unr14_stage6_stallmux_q_27_), .o(n_23919) );
in01s01 g756507 ( .a(n_23680), .o(n_23681) );
no02f04 TIMEBOOST_cell_6058 ( .a(TIMEBOOST_net_1880), .b(n_29643), .o(n_29658) );
in01s01 g756509 ( .a(n_23917), .o(n_23918) );
ao12s01 g756510 ( .a(n_23878), .b(n_23783), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_25_), .o(n_23917) );
in01s01 g756511 ( .a(n_23759), .o(n_23760) );
ao22s01 g756512 ( .a(n_23606), .b(n_22717), .c(n_23599), .d(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_), .o(n_23759) );
no02s06 TIMEBOOST_cell_1812 ( .a(TIMEBOOST_net_520), .b(FE_RN_1968_0), .o(n_46957) );
in01s01 g756515 ( .a(n_23844), .o(n_23845) );
ao22s01 g756516 ( .a(n_23821), .b(n_23773), .c(n_23783), .d(delay_sub_ln21_0_unr14_stage6_stallmux_q_23_), .o(n_23844) );
in01s01 g756517 ( .a(n_24050), .o(n_24051) );
ao12s01 g756518 ( .a(n_23993), .b(FE_OCP_RBN6560_n_23572), .c(delay_add_ln22_unr14_stage6_stallmux_q_30_), .o(n_24050) );
in01s01 g756519 ( .a(n_23964), .o(n_23965) );
ao12m01 g756520 ( .a(n_23851), .b(n_23783), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_27_), .o(n_23964) );
ao12s02 g756522 ( .a(n_23874), .b(n_23783), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_29_), .o(n_23941) );
in01s01 g756523 ( .a(n_24009), .o(n_24010) );
ao12s01 g756524 ( .a(n_23969), .b(FE_OCP_RBN6560_n_23572), .c(delay_add_ln22_unr14_stage6_stallmux_q_29_), .o(n_24009) );
oa12f06 g756525 ( .a(n_23369), .b(n_23545), .c(n_23407), .o(n_23615) );
no02m06 TIMEBOOST_cell_1846 ( .a(TIMEBOOST_net_537), .b(n_5943), .o(n_5968) );
no02m08 TIMEBOOST_cell_1962 ( .a(TIMEBOOST_net_595), .b(n_37395), .o(n_37467) );
ao12s01 g756528 ( .a(n_23830), .b(n_24078), .c(n_23721), .o(n_24114) );
ao22s01 g756530 ( .a(FE_OCP_RBN6559_n_23572), .b(n_22858), .c(FE_OCP_RBN6557_n_23572), .d(delay_add_ln22_unr14_stage6_stallmux_q_25_), .o(n_23914) );
oa12s01 g756531 ( .a(n_23520), .b(n_23545), .c(n_23519), .o(n_24962) );
in01s01 g756532 ( .a(n_24048), .o(n_24049) );
oa22s01 g756533 ( .a(FE_OCP_RBN6560_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_31_), .c(FE_OCP_RBN6559_n_23572), .d(n_22929), .o(n_24048) );
in01s01 g756534 ( .a(n_23962), .o(n_23963) );
ao22s01 g756535 ( .a(n_23821), .b(n_22873), .c(n_23783), .d(delay_sub_ln21_0_unr14_stage6_stallmux_q_31_), .o(n_23962) );
in01s06 g756536 ( .a(n_23586), .o(n_23639) );
na02s10 g756537 ( .a(n_23563), .b(n_23562), .o(n_23586) );
no02s06 g756538 ( .a(n_23563), .b(n_23562), .o(n_23613) );
no02s02 g756539 ( .a(n_23551), .b(delay_add_ln22_unr14_stage6_stallmux_q_21_), .o(n_23735) );
no02s02 g756540 ( .a(FE_OCP_RBN6560_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_27_), .o(n_23854) );
no02s01 g756541 ( .a(FE_OCP_RBN6560_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_28_), .o(n_23970) );
na02s01 g756542 ( .a(FE_OCP_RBN6557_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_24_), .o(n_23883) );
na02s02 g756543 ( .a(n_23572), .b(n_23611), .o(n_23659) );
no02f08 TIMEBOOST_cell_5111 ( .a(TIMEBOOST_net_1503), .b(n_38205), .o(n_38288) );
no02s02 g756545 ( .a(n_23551), .b(delay_add_ln22_unr14_stage6_stallmux_q_18_), .o(n_23638) );
in01s01 g756546 ( .a(n_23767), .o(n_23713) );
na02s06 g756547 ( .a(FE_OCP_RBN6557_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_20_), .o(n_23767) );
in01s01 g756548 ( .a(n_23993), .o(n_23994) );
no02s01 g756549 ( .a(FE_OCP_RBN6560_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_30_), .o(n_23993) );
no02s02 g756550 ( .a(FE_OCP_RBN6559_n_23572), .b(n_22859), .o(n_23884) );
in01s01 g756551 ( .a(n_23853), .o(n_23820) );
no02s06 g756552 ( .a(FE_OCP_RBN6560_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_26_), .o(n_23853) );
in01s01 g756553 ( .a(n_23818), .o(n_23819) );
no02s01 g756554 ( .a(FE_OCP_RBN6557_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_24_), .o(n_23818) );
in01s02 g756555 ( .a(n_23736), .o(n_23768) );
no02s04 g756556 ( .a(n_23551), .b(delay_add_ln22_unr14_stage6_stallmux_q_20_), .o(n_23736) );
in01s01 g756557 ( .a(n_23876), .o(n_23945) );
na02s01 g756558 ( .a(FE_OCP_RBN6560_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_28_), .o(n_23876) );
in01s01 g756559 ( .a(n_23757), .o(n_23758) );
na02s01 g756560 ( .a(FE_OCP_RBN6557_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_23_), .o(n_23757) );
no02s06 g756561 ( .a(FE_OCP_RBN6557_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_22_), .o(n_24182) );
na02f06 g756562 ( .a(n_23636), .b(n_23635), .o(n_23637) );
no02s01 g756563 ( .a(FE_OCP_RBN6560_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_29_), .o(n_23969) );
no02s02 g756564 ( .a(FE_OCP_RBN6557_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_23_), .o(n_23823) );
in01s01 g756565 ( .a(n_23664), .o(n_23634) );
no02s03 g756566 ( .a(n_23563), .b(n_22669), .o(n_23664) );
in01s01 g756567 ( .a(n_23711), .o(n_23712) );
na02s03 g756568 ( .a(FE_OCP_RBN6557_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_22_), .o(n_23711) );
in01s01 g756569 ( .a(n_23632), .o(n_23633) );
no02s10 g756570 ( .a(n_23572), .b(n_23611), .o(n_23632) );
in01s01 g756572 ( .a(n_23584), .o(n_23609) );
na02f08 g756573 ( .a(n_23561), .b(n_23560), .o(n_23584) );
no02f02 TIMEBOOST_cell_6057 ( .a(FE_RN_2412_0), .b(FE_OFN774_n_25834), .o(TIMEBOOST_net_1880) );
no02m04 TIMEBOOST_cell_7519 ( .a(TIMEBOOST_net_2390), .b(n_23814), .o(n_23939) );
no02s02 g756576 ( .a(FE_OCPN1049_n_23581), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_), .o(n_23582) );
no02m01 g756577 ( .a(n_23783), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_25_), .o(n_23878) );
na02m01 g756579 ( .a(n_23606), .b(n_22754), .o(n_23762) );
no02s01 g756580 ( .a(n_23599), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_), .o(n_23677) );
na02m03 g756581 ( .a(n_23658), .b(n_23821), .o(n_23733) );
na02s03 g756582 ( .a(n_23574), .b(n_22630), .o(n_23682) );
no02s02 g756583 ( .a(n_23599), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_19_), .o(n_23679) );
na02f01 g756584 ( .a(n_23606), .b(n_23653), .o(n_23822) );
no02s02 g756585 ( .a(n_23599), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_26_), .o(n_23850) );
na02s01 g756586 ( .a(n_23636), .b(n_23601), .o(n_24001) );
no02f02 TIMEBOOST_cell_1813 ( .a(n_16080), .b(n_16123), .o(TIMEBOOST_net_521) );
no02s01 g756588 ( .a(n_23783), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_27_), .o(n_23851) );
in01s01 g756589 ( .a(n_23817), .o(n_23922) );
na02s01 g756590 ( .a(n_23599), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_28_), .o(n_23817) );
no02s02 g756591 ( .a(n_23783), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_28_), .o(n_23921) );
no02s02 g756593 ( .a(n_23783), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_29_), .o(n_23874) );
na02s01 g756594 ( .a(n_23783), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_30_), .o(n_23966) );
in01s01 g756595 ( .a(n_23872), .o(n_23873) );
no02s01 g756596 ( .a(n_23783), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_30_), .o(n_23872) );
in01s02 g756597 ( .a(n_23740), .o(n_23676) );
no02s06 g756598 ( .a(n_23606), .b(n_23658), .o(n_23740) );
na02s01 g756599 ( .a(n_23631), .b(n_23578), .o(n_23894) );
in01s01 g756600 ( .a(n_23761), .o(n_23709) );
na02s01 g756601 ( .a(n_23599), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_22_), .o(n_23761) );
in01m01 g756602 ( .a(n_23580), .o(n_23663) );
no02f06 g756603 ( .a(n_23561), .b(n_23560), .o(n_23580) );
in01s01 g756604 ( .a(n_23684), .o(n_23630) );
na02m02 g756605 ( .a(n_23604), .b(n_23603), .o(n_23684) );
na02s02 g756607 ( .a(FE_OCPN1050_n_23581), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_18_), .o(n_23683) );
in01m02 g756608 ( .a(n_23656), .o(n_24067) );
in01m02 g756610 ( .a(n_23629), .o(n_23656) );
no02m04 g756611 ( .a(n_23604), .b(n_23603), .o(n_23629) );
in01s02 g756612 ( .a(n_23708), .o(n_23765) );
na02f01 g756613 ( .a(n_23599), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_26_), .o(n_23708) );
in01s01 g756614 ( .a(n_23738), .o(n_23675) );
no02s01 g756615 ( .a(n_23606), .b(n_23653), .o(n_23738) );
no02s01 g756616 ( .a(n_24078), .b(n_24149), .o(n_24195) );
na02s01 g756617 ( .a(n_23545), .b(n_23519), .o(n_23520) );
in01s01 g756618 ( .a(n_23972), .o(n_23885) );
oa12s02 g756619 ( .a(FE_OCP_RBN6557_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_25_), .c(delay_add_ln22_unr14_stage6_stallmux_q_24_), .o(n_23972) );
ao12m01 g756621 ( .a(FE_OCP_RBN6560_n_23572), .b(delay_add_ln22_unr14_stage6_stallmux_q_25_), .c(delay_add_ln22_unr14_stage6_stallmux_q_24_), .o(n_23815) );
in01s01 g756622 ( .a(n_23666), .o(n_23602) );
ao12f08 g756623 ( .a(n_23418), .b(n_23579), .c(n_23455), .o(n_23666) );
na02s02 g756624 ( .a(n_24192), .b(n_24152), .o(n_24193) );
oa12s02 g756625 ( .a(n_23551), .b(delay_add_ln22_unr14_stage6_stallmux_q_20_), .c(delay_add_ln22_unr14_stage6_stallmux_q_21_), .o(n_23734) );
na02s06 g756626 ( .a(n_23572), .b(n_22773), .o(n_23707) );
na02m06 g756628 ( .a(n_24078), .b(n_23749), .o(n_24077) );
ao22s01 g756629 ( .a(n_23474), .b(n_23544), .c(n_23473), .d(n_23579), .o(n_25022) );
in01s01 g756630 ( .a(n_23627), .o(n_23628) );
ao12s01 g756631 ( .a(n_23559), .b(n_23558), .c(n_23557), .o(n_23627) );
ao12s02 g756632 ( .a(n_23508), .b(n_23507), .c(n_23506), .o(n_24893) );
in01s01 g756633 ( .a(n_24275), .o(n_24257) );
ao12s01 g756634 ( .a(n_24191), .b(n_24190), .c(n_24189), .o(n_24275) );
no02m06 g756635 ( .a(n_24190), .b(n_24037), .o(n_24078) );
na02f04 g756636 ( .a(n_23555), .b(n_23554), .o(n_23631) );
no02s01 g756637 ( .a(n_24190), .b(n_24189), .o(n_24191) );
in01s01 g756638 ( .a(n_23651), .o(n_23652) );
na02s01 g756639 ( .a(n_23635), .b(n_23626), .o(n_23651) );
no02s01 g756640 ( .a(n_23558), .b(n_23557), .o(n_23559) );
no02s01 g756641 ( .a(n_23518), .b(n_23556), .o(n_23797) );
in01s01 g756642 ( .a(FE_OCPN939_n_23577), .o(n_23578) );
no02m02 g756643 ( .a(n_23555), .b(n_23554), .o(n_23577) );
na02f06 g756644 ( .a(n_23576), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_15_), .o(n_23636) );
in01s01 g756645 ( .a(n_23600), .o(n_23601) );
no02s06 g756646 ( .a(n_23576), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_15_), .o(n_23600) );
na02f06 g756647 ( .a(n_23445), .b(n_23330), .o(n_23545) );
in01s06 g756650 ( .a(FE_OCPN1049_n_23581), .o(n_23574) );
in01s02 g756657 ( .a(n_23821), .o(n_23783) );
in01m03 g756660 ( .a(n_23599), .o(n_23821) );
in01m10 g756668 ( .a(n_23606), .o(n_23599) );
in01m10 g756669 ( .a(FE_OCPN1050_n_23581), .o(n_23606) );
no02s02 TIMEBOOST_cell_6900 ( .a(TIMEBOOST_net_2208), .b(n_18625), .o(n_18738) );
no02s01 g756671 ( .a(n_23507), .b(n_23506), .o(n_23508) );
in01s02 g756672 ( .a(n_24132), .o(n_24192) );
oa12s02 g756673 ( .a(n_24107), .b(n_24064), .c(FE_OFN780_n_23803), .o(n_24132) );
in01m10 g756701 ( .a(n_23551), .o(n_23572) );
in01m06 g756702 ( .a(n_23563), .o(n_23551) );
no02m04 TIMEBOOST_cell_6082 ( .a(TIMEBOOST_net_1892), .b(FE_OCP_RBN2747_n_8474), .o(n_8619) );
ao22f08 g756704 ( .a(n_23463), .b(n_23141), .c(n_23482), .d(n_23140), .o(n_23561) );
oa12m02 g756705 ( .a(n_23516), .b(n_23504), .c(n_23515), .o(n_23604) );
no02s01 TIMEBOOST_cell_1801 ( .a(FE_OCPN1238_n_30470), .b(FE_OCP_RBN6748_n_30170), .o(TIMEBOOST_net_515) );
in01s01 g756707 ( .a(n_23579), .o(n_23544) );
no02f04 TIMEBOOST_cell_7093 ( .a(FE_OCP_RBN7042_n_20336), .b(n_45060), .o(TIMEBOOST_net_2305) );
na02f08 g756710 ( .a(n_23480), .b(n_23479), .o(n_23481) );
in01s01 g756711 ( .a(n_23517), .o(n_23518) );
na02f10 g756712 ( .a(n_23502), .b(delay_add_ln22_unr14_stage6_stallmux_q_14_), .o(n_23517) );
in01s01 g756713 ( .a(n_23595), .o(n_23596) );
na02s01 g756714 ( .a(n_23571), .b(n_23543), .o(n_23595) );
no02s01 g756715 ( .a(n_23432), .b(n_23329), .o(n_23507) );
na02s01 g756716 ( .a(n_23480), .b(FE_OCPN1610_n_23503), .o(n_23794) );
no02s04 g756717 ( .a(n_23502), .b(delay_add_ln22_unr14_stage6_stallmux_q_14_), .o(n_23556) );
in01s01 g756718 ( .a(n_23626), .o(n_23594) );
na02f08 g756719 ( .a(n_23540), .b(n_22354), .o(n_23626) );
na02s01 TIMEBOOST_cell_3160 ( .a(FE_OCPN1628_n_34452), .b(n_34429), .o(TIMEBOOST_net_871) );
na02f04 g756721 ( .a(n_23539), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_14_), .o(n_23635) );
no02s01 g756722 ( .a(n_24036), .b(n_24007), .o(n_24008) );
oa12s01 g756723 ( .a(n_23373), .b(n_23514), .c(n_23371), .o(n_23558) );
in01s01 g756724 ( .a(n_24107), .o(n_24047) );
no02s02 g756725 ( .a(n_24036), .b(n_23984), .o(n_24107) );
na02f04 g756726 ( .a(n_23431), .b(n_23315), .o(n_23445) );
no02m06 g756727 ( .a(n_23939), .b(n_23813), .o(n_24190) );
ao12s01 g756728 ( .a(n_23499), .b(n_23514), .c(n_23498), .o(n_24943) );
oa12s01 g756729 ( .a(n_23430), .b(n_23429), .c(n_23428), .o(n_24825) );
no02s06 TIMEBOOST_cell_4930 ( .a(n_23313), .b(n_23096), .o(TIMEBOOST_net_1413) );
na02s06 TIMEBOOST_cell_4887 ( .a(TIMEBOOST_net_1391), .b(n_17537), .o(n_17734) );
in01s01 g756733 ( .a(n_23431), .o(n_23432) );
na02f04 g756734 ( .a(n_23397), .b(n_23287), .o(n_23431) );
na02s04 TIMEBOOST_cell_8165 ( .a(TIMEBOOST_net_2713), .b(n_11102), .o(n_11191) );
no02s01 TIMEBOOST_cell_6247 ( .a(n_4875), .b(n_4759), .o(TIMEBOOST_net_1975) );
na02m06 g756738 ( .a(n_23423), .b(n_22203), .o(n_23503) );
in01s01 g756739 ( .a(n_23542), .o(n_23543) );
no02f08 g756740 ( .a(n_23513), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_13_), .o(n_23542) );
na02s01 g756741 ( .a(n_23541), .b(n_23497), .o(n_23719) );
na02s01 g756742 ( .a(n_23479), .b(n_23444), .o(n_23693) );
in01m08 g756743 ( .a(n_23482), .o(n_23463) );
no02m20 g756744 ( .a(n_23426), .b(n_23114), .o(n_23482) );
na02f08 g756745 ( .a(n_23422), .b(delay_add_ln22_unr14_stage6_stallmux_q_13_), .o(n_23480) );
na02f04 g756747 ( .a(n_23513), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_13_), .o(n_23571) );
no02s01 g756748 ( .a(n_23991), .b(n_23990), .o(n_23992) );
na02s01 g756749 ( .a(n_23429), .b(n_23428), .o(n_23430) );
no02s01 g756750 ( .a(n_23514), .b(n_23498), .o(n_23499) );
oa12s02 g756752 ( .a(n_23938), .b(n_23866), .c(FE_OFN780_n_23803), .o(n_24036) );
na02s04 TIMEBOOST_cell_8782 ( .a(FE_OCP_RBN2803_n_3220), .b(FE_OCP_RBN2705_n_47023), .o(TIMEBOOST_net_2878) );
no02s02 g756754 ( .a(n_24035), .b(n_24032), .o(n_24065) );
ao12s01 g756755 ( .a(n_23459), .b(n_23458), .c(n_23457), .o(n_24919) );
ao12s01 g756756 ( .a(n_23410), .b(n_23409), .c(n_23408), .o(n_24747) );
in01s01 g756757 ( .a(n_25092), .o(n_24236) );
ao12s01 g756758 ( .a(n_24172), .b(n_24171), .c(n_24170), .o(n_25092) );
in01f04 g756759 ( .a(n_23539), .o(n_23540) );
no03s04 TIMEBOOST_cell_8310 ( .a(n_3273), .b(FE_OCP_RBN5724_n_47022), .c(n_3302), .o(n_3391) );
in01s01 g756762 ( .a(n_23443), .o(n_23444) );
no02s06 g756763 ( .a(n_23424), .b(delay_add_ln22_unr14_stage6_stallmux_q_12_), .o(n_23443) );
in01s01 g756764 ( .a(n_23537), .o(n_23538) );
na02s01 g756765 ( .a(n_23472), .b(n_23512), .o(n_23537) );
no02s01 g756766 ( .a(n_23458), .b(n_23457), .o(n_23459) );
na02s01 g756767 ( .a(n_23395), .b(n_23427), .o(n_23587) );
in01s01 g756768 ( .a(n_23496), .o(n_23497) );
no02s06 g756769 ( .a(n_23476), .b(n_23475), .o(n_23496) );
no02m08 g756770 ( .a(n_23439), .b(n_23462), .o(n_23500) );
na02s06 g756771 ( .a(n_23476), .b(n_23475), .o(n_23541) );
in01f04 g756773 ( .a(n_23426), .o(n_23441) );
na02m20 g756774 ( .a(n_23411), .b(FE_OCP_RBN2446_n_23079), .o(n_23426) );
na02f10 g756775 ( .a(n_23411), .b(n_23145), .o(n_23412) );
na02f08 g756777 ( .a(n_23424), .b(delay_add_ln22_unr14_stage6_stallmux_q_12_), .o(n_23479) );
no03f08 TIMEBOOST_cell_8443 ( .a(FE_OCP_RBN1040_n_26158), .b(n_26207), .c(n_26262), .o(n_26429) );
no02s01 g756779 ( .a(n_24171), .b(n_24170), .o(n_24172) );
na02s01 g756780 ( .a(n_24153), .b(n_24105), .o(n_24154) );
na02s02 g756781 ( .a(n_23956), .b(n_24034), .o(n_24035) );
in01s01 g756782 ( .a(n_23397), .o(n_23429) );
ao12f04 g756783 ( .a(n_23251), .b(n_23348), .c(n_23252), .o(n_23397) );
no02s01 g756784 ( .a(n_23409), .b(n_23408), .o(n_23410) );
in01s01 g756785 ( .a(n_23456), .o(n_23514) );
no02f06 g756786 ( .a(n_23405), .b(n_23264), .o(n_23456) );
in01s01 g756787 ( .a(n_23938), .o(n_23991) );
ao12s02 g756788 ( .a(n_23911), .b(n_23723), .c(n_23743), .o(n_23938) );
ao12s01 g756789 ( .a(n_24355), .b(n_24076), .c(n_24059), .o(n_24815) );
oa12s01 g756790 ( .a(n_24059), .b(n_24151), .c(n_24150), .o(n_24152) );
no02f02 TIMEBOOST_cell_1785 ( .a(n_15429), .b(n_14419), .o(TIMEBOOST_net_507) );
in01s02 g756792 ( .a(n_23422), .o(n_23423) );
na02f08 g756793 ( .a(n_23380), .b(n_23253), .o(n_23422) );
na02s01 TIMEBOOST_cell_4984 ( .a(TIMEBOOST_net_211), .b(n_37898), .o(TIMEBOOST_net_1440) );
no02s02 TIMEBOOST_cell_5164 ( .a(n_44100), .b(n_34127), .o(TIMEBOOST_net_1530) );
oa12f08 g756797 ( .a(n_23045), .b(FE_OCP_RBN5552_n_23328), .c(n_23378), .o(n_23380) );
in01m06 g756798 ( .a(n_23411), .o(n_23396) );
in01s01 g756800 ( .a(n_23473), .o(n_23474) );
na02s01 g756801 ( .a(n_23455), .b(n_23419), .o(n_23473) );
no02s01 g756802 ( .a(n_23370), .b(n_23407), .o(n_23519) );
no02s01 g756803 ( .a(n_23349), .b(n_23215), .o(n_23409) );
na02m04 g756804 ( .a(n_23377), .b(n_23376), .o(n_23427) );
in01s01 g756805 ( .a(n_23471), .o(n_23472) );
no02s08 g756806 ( .a(n_23452), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_11_), .o(n_23471) );
in01m04 g756808 ( .a(n_23439), .o(n_23453) );
na02m10 g756809 ( .a(n_47245), .b(n_23032), .o(n_23439) );
na02s06 g756810 ( .a(n_23452), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_11_), .o(n_23512) );
in01s01 g756811 ( .a(n_23394), .o(n_23395) );
no02s04 g756812 ( .a(n_23377), .b(n_23376), .o(n_23394) );
in01m02 g756813 ( .a(n_24171), .o(n_23814) );
no02m04 g756814 ( .a(n_23753), .b(n_23703), .o(n_24171) );
no02s04 g756815 ( .a(n_23754), .b(n_23812), .o(n_23813) );
in01s01 g756816 ( .a(n_24032), .o(n_24033) );
na02s01 g756817 ( .a(n_24006), .b(n_23950), .o(n_24032) );
no02s01 g756818 ( .a(n_24029), .b(n_23934), .o(n_24031) );
na02s01 g756819 ( .a(n_23865), .b(n_23909), .o(n_23937) );
na02s01 g756820 ( .a(n_24046), .b(n_24091), .o(n_24739) );
no02s01 g756821 ( .a(n_24059), .b(n_24076), .o(n_24355) );
no02s01 g756822 ( .a(n_24063), .b(n_24076), .o(n_24064) );
ao12s01 g756823 ( .a(n_23245), .b(n_23420), .c(n_23289), .o(n_23458) );
no02s02 g756824 ( .a(n_24029), .b(n_23987), .o(n_24030) );
no02s02 g756825 ( .a(n_23910), .b(n_23958), .o(n_23959) );
in01s02 g756826 ( .a(n_23838), .o(n_23911) );
ao12s02 g756827 ( .a(n_23811), .b(n_23724), .c(n_23671), .o(n_23838) );
ao12f04 g756829 ( .a(n_23291), .b(n_23365), .c(n_23281), .o(n_23405) );
in01s01 g756830 ( .a(n_24153), .o(n_24131) );
ao12s01 g756831 ( .a(n_24106), .b(n_24075), .c(n_24105), .o(n_24153) );
in01s01 g756832 ( .a(n_23956), .o(n_23957) );
no02s01 g756833 ( .a(n_23936), .b(n_23868), .o(n_23956) );
ao12s01 g756834 ( .a(n_24354), .b(n_24150), .c(n_24059), .o(n_24903) );
oa12s01 g756835 ( .a(n_24034), .b(n_23989), .c(n_24188), .o(n_24736) );
oa22s02 g756836 ( .a(n_23420), .b(n_23304), .c(n_23386), .d(n_23303), .o(n_24838) );
oa12s01 g756837 ( .a(n_23333), .b(n_23334), .c(n_23332), .o(n_24682) );
in01s01 g756838 ( .a(n_23836), .o(n_23837) );
oa12s01 g756839 ( .a(n_23752), .b(n_23751), .c(n_23750), .o(n_23836) );
oa12s06 g756840 ( .a(n_23336), .b(n_23385), .c(FE_OCPN1356_n_23335), .o(n_23476) );
no02f02 TIMEBOOST_cell_8554 ( .a(TIMEBOOST_net_2236), .b(n_8284), .o(TIMEBOOST_net_2764) );
na02s01 g756846 ( .a(n_23374), .b(n_23393), .o(n_23557) );
ao12s01 g756847 ( .a(n_23331), .b(n_23266), .c(delay_add_ln22_unr14_stage6_stallmux_q_9_), .o(n_23506) );
na02m06 g756848 ( .a(n_23328), .b(n_23179), .o(n_23350) );
in01s01 g756849 ( .a(n_23369), .o(n_23370) );
na02s04 g756850 ( .a(n_23363), .b(delay_add_ln22_unr14_stage6_stallmux_q_10_), .o(n_23369) );
in01s01 g756851 ( .a(n_23418), .o(n_23419) );
no02m08 g756852 ( .a(n_23404), .b(n_23403), .o(n_23418) );
na02m08 g756853 ( .a(n_23404), .b(n_23403), .o(n_23455) );
no02f04 g756858 ( .a(n_23363), .b(delay_add_ln22_unr14_stage6_stallmux_q_10_), .o(n_23407) );
no02s01 TIMEBOOST_cell_8503 ( .a(TIMEBOOST_net_2738), .b(n_7671), .o(n_7732) );
in01s01 g756860 ( .a(n_23348), .o(n_23349) );
in01s01 g756862 ( .a(n_23753), .o(n_23754) );
no02m04 g756863 ( .a(n_23750), .b(n_23702), .o(n_23753) );
na02s01 g756864 ( .a(n_23751), .b(n_23750), .o(n_23752) );
no02s01 g756865 ( .a(n_24075), .b(n_24105), .o(n_24106) );
no02s01 g756866 ( .a(n_23811), .b(n_23704), .o(n_23705) );
na02s01 g756867 ( .a(n_24061), .b(n_24044), .o(n_24062) );
no02s01 g756868 ( .a(n_23907), .b(n_23905), .o(n_24006) );
na02s01 g756869 ( .a(n_23867), .b(n_23832), .o(n_23868) );
no02s01 g756870 ( .a(n_23990), .b(n_23951), .o(n_24706) );
no02s01 g756871 ( .a(n_23990), .b(n_23701), .o(n_23866) );
na02s01 g756872 ( .a(FE_OFN780_n_23803), .b(n_24028), .o(n_24091) );
na02s01 g756873 ( .a(n_23989), .b(FE_OFN780_n_23803), .o(n_24034) );
no02s01 g756874 ( .a(n_24059), .b(n_24150), .o(n_24354) );
in01s01 g756875 ( .a(n_24063), .o(n_24046) );
no02s01 g756876 ( .a(n_24028), .b(FE_OFN780_n_23803), .o(n_24063) );
na02s01 g756877 ( .a(n_23334), .b(n_23332), .o(n_23333) );
oa12s01 g756878 ( .a(n_24061), .b(n_24188), .c(n_24023), .o(n_24675) );
oa12s01 g756879 ( .a(n_23906), .b(n_24188), .c(n_23863), .o(n_24769) );
oa12s01 g756880 ( .a(n_23867), .b(n_24188), .c(n_23810), .o(n_24733) );
in01s01 g756881 ( .a(n_23958), .o(n_23865) );
ao12s01 g756882 ( .a(n_23743), .b(n_23834), .c(n_23897), .o(n_23958) );
oa12s01 g756883 ( .a(FE_OFN780_n_23803), .b(n_24088), .c(n_24087), .o(n_24090) );
in01s01 g756884 ( .a(n_23988), .o(n_24029) );
oa12s01 g756885 ( .a(n_23743), .b(n_23955), .c(n_23954), .o(n_23988) );
ao12s01 g756886 ( .a(FE_OFN780_n_23803), .b(n_23986), .c(n_23985), .o(n_23987) );
ao12s01 g756887 ( .a(n_23743), .b(n_23909), .c(n_23901), .o(n_23910) );
ao12s01 g756888 ( .a(FE_OFN780_n_23803), .b(n_24086), .c(n_24088), .o(n_24151) );
ao12s01 g756889 ( .a(FE_OFN780_n_23803), .b(n_23899), .c(n_24023), .o(n_23984) );
ao12s01 g756890 ( .a(n_23368), .b(n_23367), .c(n_23366), .o(n_24764) );
ao12s02 g756891 ( .a(n_23311), .b(n_23310), .c(n_23309), .o(n_24613) );
oa12s01 g756892 ( .a(n_23649), .b(n_23648), .c(n_23647), .o(n_24076) );
no03m04 TIMEBOOST_cell_3562 ( .a(FE_OCP_RBN7030_n_44259), .b(n_33663), .c(n_33691), .o(n_33809) );
ao22s01 g756894 ( .a(n_24188), .b(n_24088), .c(n_24059), .d(n_23641), .o(n_24907) );
na02s02 TIMEBOOST_cell_7877 ( .a(TIMEBOOST_net_2569), .b(n_4247), .o(n_4434) );
no02s04 g756896 ( .a(n_23384), .b(n_23095), .o(n_23387) );
na03s03 TIMEBOOST_cell_8225 ( .a(n_28606), .b(FE_RN_1546_0), .c(n_28543), .o(FE_RN_1548_0) );
no02s01 TIMEBOOST_cell_1655 ( .a(n_3639), .b(n_3118), .o(TIMEBOOST_net_442) );
na02s01 TIMEBOOST_cell_4904 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_7_), .b(n_23087), .o(TIMEBOOST_net_1400) );
in01s01 g756900 ( .a(n_23330), .o(n_23331) );
na02s06 g756901 ( .a(n_23284), .b(n_21912), .o(n_23330) );
no02s01 g756902 ( .a(n_23371), .b(n_23325), .o(n_23498) );
no02s01 g756903 ( .a(n_23367), .b(n_23366), .o(n_23368) );
no02s01 g756904 ( .a(n_23329), .b(n_23288), .o(n_23428) );
no02s01 g756905 ( .a(n_23310), .b(n_23309), .o(n_23311) );
na02m02 g756906 ( .a(n_23347), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_9_), .o(n_23374) );
in01s01 g756907 ( .a(n_23420), .o(n_23386) );
in01s01 g756908 ( .a(n_23365), .o(n_23420) );
na02s01 g756910 ( .a(n_23648), .b(n_23647), .o(n_23649) );
no02s02 g756913 ( .a(n_23384), .b(n_23391), .o(n_23385) );
in01f02 g756914 ( .a(n_23361), .o(n_23393) );
no02f04 g756915 ( .a(n_23347), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_9_), .o(n_23361) );
na02m08 TIMEBOOST_cell_8615 ( .a(TIMEBOOST_net_2794), .b(n_21398), .o(n_21587) );
na02s01 g756918 ( .a(n_23833), .b(n_23864), .o(n_23936) );
na02s01 g756919 ( .a(n_24025), .b(n_24024), .o(n_24026) );
na02s02 g756920 ( .a(n_23952), .b(n_23932), .o(n_23953) );
no02s02 g756921 ( .a(n_23748), .b(n_23747), .o(n_23749) );
no02s01 g756922 ( .a(n_23704), .b(n_23908), .o(n_24672) );
no02s01 g756923 ( .a(n_23703), .b(n_23702), .o(n_23751) );
na02s01 g756924 ( .a(n_24024), .b(n_23986), .o(n_24479) );
no02s01 g756925 ( .a(n_23778), .b(n_23748), .o(n_24113) );
no02s01 g756926 ( .a(n_24234), .b(n_24256), .o(n_24543) );
na02s01 g756927 ( .a(n_24352), .b(n_24086), .o(n_24845) );
no02s01 g756928 ( .a(n_23900), .b(n_23831), .o(n_24379) );
na02s01 g756929 ( .a(FE_OFN780_n_23803), .b(n_24023), .o(n_24061) );
in01s01 g756930 ( .a(n_23950), .o(n_23951) );
na02s01 g756931 ( .a(n_23806), .b(FE_OFN780_n_23803), .o(n_23950) );
in01s01 g756932 ( .a(n_23906), .o(n_23907) );
na02s01 g756933 ( .a(FE_OFN780_n_23803), .b(n_23863), .o(n_23906) );
na02s01 g756934 ( .a(n_23700), .b(n_23810), .o(n_23867) );
na02s01 g756935 ( .a(n_23808), .b(n_23807), .o(n_23809) );
no02s01 g756936 ( .a(n_23806), .b(n_23700), .o(n_23990) );
na02s02 g756937 ( .a(n_23672), .b(n_23810), .o(n_23724) );
na02s01 g756938 ( .a(n_23722), .b(n_23863), .o(n_23723) );
no02s01 g756939 ( .a(n_24007), .b(n_24074), .o(n_24664) );
no02s01 g756940 ( .a(n_23697), .b(n_23905), .o(n_24667) );
no02s01 g756941 ( .a(n_24169), .b(n_23779), .o(n_24240) );
no02s01 g756942 ( .a(n_24149), .b(n_24037), .o(n_24189) );
na02s01 g756943 ( .a(n_24215), .b(n_23904), .o(n_24383) );
oa12s01 g756944 ( .a(n_23864), .b(n_24188), .c(n_23802), .o(n_24628) );
oa12s01 g756945 ( .a(n_24025), .b(n_24188), .c(n_23985), .o(n_24513) );
ao12s01 g756946 ( .a(n_23933), .b(n_24188), .c(n_23399), .o(n_24414) );
ao12s01 g756947 ( .a(n_23747), .b(FE_OFN779_n_23803), .c(n_23800), .o(n_24194) );
ao12s01 g756948 ( .a(n_23646), .b(n_23802), .c(n_23804), .o(n_23811) );
ao22s01 g756949 ( .a(FE_OFN779_n_23803), .b(n_23869), .c(n_24059), .d(n_23812), .o(n_24170) );
ao22s01 g756950 ( .a(n_24188), .b(n_23979), .c(n_24059), .d(n_23954), .o(n_24454) );
oa22s01 g756951 ( .a(n_24059), .b(n_23897), .c(n_24188), .d(n_23341), .o(n_24300) );
ao12s01 g756952 ( .a(n_23644), .b(n_23643), .c(n_23642), .o(n_24028) );
in01s01 g756953 ( .a(n_23701), .o(n_23989) );
oa12s01 g756954 ( .a(n_23620), .b(n_23619), .c(n_23618), .o(n_23701) );
oa12s01 g756955 ( .a(n_23593), .b(n_23592), .c(n_23591), .o(n_24150) );
oa22s01 g756956 ( .a(FE_OFN779_n_23803), .b(n_24111), .c(n_24059), .d(n_23807), .o(n_24237) );
oa22s01 g756957 ( .a(n_23743), .b(n_22811), .c(FE_OFN779_n_23803), .d(n_22885), .o(n_24075) );
na02m04 g756959 ( .a(n_23269), .b(n_23286), .o(n_23363) );
no02f06 g756993 ( .a(n_23215), .b(n_23250), .o(n_23252) );
na02m04 g756994 ( .a(n_23290), .b(n_23289), .o(n_23291) );
in01s01 g756995 ( .a(n_23287), .o(n_23288) );
na02s03 g756996 ( .a(n_47337), .b(n_23267), .o(n_23287) );
na02s01 g756997 ( .a(n_23346), .b(n_23213), .o(n_23367) );
na02s01 g756998 ( .a(n_23290), .b(n_23265), .o(n_23457) );
na02s01 g756999 ( .a(n_23197), .b(n_23270), .o(n_23310) );
na02s04 g757001 ( .a(n_23345), .b(n_23094), .o(n_23384) );
na02s01 g757002 ( .a(n_23619), .b(n_23618), .o(n_23620) );
na02s01 g757004 ( .a(n_23592), .b(n_23591), .o(n_23593) );
no02m06 g757006 ( .a(n_23305), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_8_), .o(n_23371) );
no02s01 g757007 ( .a(n_23251), .b(n_23250), .o(n_23408) );
oa12s02 g757008 ( .a(n_23074), .b(n_23195), .c(n_23307), .o(n_23269) );
no02f04 g757009 ( .a(n_47337), .b(n_23267), .o(n_23329) );
in01s01 g757010 ( .a(n_23373), .o(n_23325) );
na02s04 g757011 ( .a(n_23305), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_8_), .o(n_23373) );
no02f02 TIMEBOOST_cell_1648 ( .a(TIMEBOOST_net_438), .b(n_47262), .o(n_15045) );
in01s01 g757013 ( .a(n_24045), .o(n_24086) );
no02s01 g757014 ( .a(FE_OFN780_n_23803), .b(n_24087), .o(n_24045) );
na02s01 g757015 ( .a(n_24188), .b(n_23978), .o(n_24215) );
in01s01 g757016 ( .a(n_24234), .o(n_24235) );
no02s01 g757017 ( .a(n_24188), .b(n_23804), .o(n_24234) );
no02s01 g757018 ( .a(FE_OFN779_n_23803), .b(n_23746), .o(n_24169) );
no02s01 g757019 ( .a(n_24059), .b(n_23061), .o(n_24149) );
in01s01 g757020 ( .a(n_23747), .o(n_23721) );
no02s01 g757021 ( .a(n_23700), .b(n_23800), .o(n_23747) );
in01s01 g757022 ( .a(n_24044), .o(n_24074) );
na02s01 g757023 ( .a(FE_OFN780_n_23803), .b(n_23860), .o(n_24044) );
in01s01 g757024 ( .a(n_23905), .o(n_23862) );
no02s01 g757025 ( .a(n_23743), .b(n_23670), .o(n_23905) );
in01s01 g757026 ( .a(n_23833), .o(n_24256) );
na02s01 g757027 ( .a(FE_OFN780_n_23803), .b(n_23804), .o(n_23833) );
na02s01 g757028 ( .a(FE_OFN780_n_23803), .b(n_23802), .o(n_23864) );
in01s01 g757029 ( .a(n_23832), .o(n_23908) );
na02s01 g757030 ( .a(n_23700), .b(n_23645), .o(n_23832) );
in01s01 g757031 ( .a(n_23955), .o(n_23904) );
no02s01 g757032 ( .a(FE_OFN780_n_23803), .b(n_23978), .o(n_23955) );
in01s01 g757033 ( .a(n_23986), .o(n_23934) );
na02s01 g757034 ( .a(n_23743), .b(n_23903), .o(n_23986) );
na02s01 g757035 ( .a(FE_OFN780_n_23803), .b(n_23985), .o(n_24025) );
in01s01 g757036 ( .a(n_23981), .o(n_24024) );
no02s01 g757037 ( .a(n_23743), .b(n_23903), .o(n_23981) );
in01s01 g757038 ( .a(n_23834), .o(n_23779) );
na02s01 g757039 ( .a(n_23700), .b(n_23746), .o(n_23834) );
in01s01 g757040 ( .a(n_23909), .o(n_23831) );
na02s02 g757041 ( .a(FE_OFN779_n_23803), .b(n_23801), .o(n_23909) );
in01s01 g757042 ( .a(n_23932), .o(n_23933) );
na02s01 g757043 ( .a(n_23743), .b(n_23901), .o(n_23932) );
in01s01 g757044 ( .a(n_23900), .o(n_23952) );
no02s01 g757045 ( .a(FE_OFN779_n_23803), .b(n_23801), .o(n_23900) );
no02s01 g757046 ( .a(n_23700), .b(n_23699), .o(n_23748) );
no02s02 g757047 ( .a(n_23616), .b(n_22882), .o(n_23703) );
no02m04 g757048 ( .a(n_23646), .b(n_22883), .o(n_23702) );
no02s02 g757049 ( .a(n_23700), .b(n_23698), .o(n_24037) );
in01s01 g757050 ( .a(n_23808), .o(n_23778) );
na02s01 g757051 ( .a(n_23700), .b(n_23699), .o(n_23808) );
in01s01 g757052 ( .a(n_24007), .o(n_23899) );
no02s01 g757053 ( .a(n_23700), .b(n_23860), .o(n_24007) );
in01s01 g757054 ( .a(n_23704), .o(n_23672) );
no02s01 g757055 ( .a(n_23646), .b(n_23645), .o(n_23704) );
in01s01 g757056 ( .a(n_23722), .o(n_23697) );
na02s01 g757057 ( .a(n_23671), .b(n_23670), .o(n_23722) );
na02s01 g757058 ( .a(n_24188), .b(n_24087), .o(n_24352) );
no02s01 g757059 ( .a(n_23643), .b(n_23642), .o(n_23644) );
ao12s01 g757060 ( .a(n_23086), .b(n_23546), .c(n_23051), .o(n_23648) );
no02s06 TIMEBOOST_cell_8838 ( .a(FE_RN_2666_0), .b(FE_OCP_RBN4904_n_44256), .o(TIMEBOOST_net_2906) );
oa12s01 g757062 ( .a(FE_OFN780_n_23803), .b(n_23979), .c(n_23978), .o(n_23980) );
oa12s01 g757063 ( .a(n_23743), .b(n_23897), .c(n_23294), .o(n_23898) );
in01s01 g757064 ( .a(n_24110), .o(n_23830) );
oa12s01 g757065 ( .a(n_23700), .b(n_23800), .c(n_23698), .o(n_24110) );
in01s02 g757067 ( .a(n_23266), .o(n_23284) );
in01s01 g757069 ( .a(n_23359), .o(n_23360) );
ao12s01 g757070 ( .a(n_23302), .b(n_23301), .c(n_23300), .o(n_23359) );
in01s01 g757071 ( .a(n_23282), .o(n_23283) );
ao12s01 g757072 ( .a(n_23236), .b(n_23235), .c(n_23234), .o(n_23282) );
in01s01 g757073 ( .a(n_24088), .o(n_23641) );
ao12s01 g757074 ( .a(n_23570), .b(n_23569), .c(n_23568), .o(n_24088) );
ao12s01 g757075 ( .a(n_23567), .b(n_23566), .c(n_23565), .o(n_23806) );
ao12s01 g757077 ( .a(n_23550), .b(n_23549), .c(n_23548), .o(n_24023) );
ao22s01 g757078 ( .a(n_23521), .b(n_23150), .c(n_23522), .d(n_23151), .o(n_23863) );
ao22s01 g757079 ( .a(n_23523), .b(n_23148), .c(n_23524), .d(n_23149), .o(n_23810) );
no02s01 g757080 ( .a(n_23549), .b(n_23548), .o(n_23550) );
no02s01 g757081 ( .a(n_23569), .b(n_23568), .o(n_23570) );
no02f10 TIMEBOOST_cell_4891 ( .a(n_12108), .b(TIMEBOOST_net_1393), .o(n_12234) );
in01s01 g757083 ( .a(n_23303), .o(n_23304) );
na02s01 g757084 ( .a(n_23289), .b(n_23281), .o(n_23303) );
no02s01 g757085 ( .a(n_23301), .b(n_23300), .o(n_23302) );
no02s01 g757086 ( .a(n_23235), .b(n_23234), .o(n_23236) );
na02s01 g757087 ( .a(n_23249), .b(n_23232), .o(n_23332) );
na02m04 g757088 ( .a(n_23248), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_7_), .o(n_23290) );
no02f04 TIMEBOOST_cell_3970 ( .a(TIMEBOOST_net_1075), .b(n_19438), .o(n_19530) );
no02m10 g757091 ( .a(FE_OCP_RBN2449_n_23246), .b(FE_OCPN1906_n_23322), .o(n_23345) );
in01s01 g757092 ( .a(n_23264), .o(n_23265) );
no02s02 g757093 ( .a(n_23248), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_7_), .o(n_23264) );
na02f06 g757094 ( .a(n_23301), .b(n_23214), .o(n_23346) );
no02s01 g757097 ( .a(n_23566), .b(n_23565), .o(n_23567) );
in01m08 g757098 ( .a(n_23144), .o(n_23145) );
ao12f20 g757099 ( .a(n_23079), .b(FE_OCP_RBN6540_n_44083), .c(delay_xor_ln22_unr15_stage6_stallmux_q_14_), .o(n_23144) );
na02s01 g757100 ( .a(n_23547), .b(n_23085), .o(n_23643) );
in01s06 g757101 ( .a(n_23142), .o(n_23143) );
ao12m10 g757102 ( .a(n_23114), .b(FE_OCP_RBN6540_n_44083), .c(delay_xor_ln22_unr15_stage6_stallmux_q_15_), .o(n_23142) );
in01s06 g757103 ( .a(n_23178), .o(n_23179) );
no02s02 TIMEBOOST_cell_6762 ( .a(TIMEBOOST_net_2138), .b(FE_OCP_RBN3102_n_15768), .o(n_15907) );
in01s02 g757112 ( .a(FE_OFN1183_n_24059), .o(n_27845) );
in01s02 g757125 ( .a(n_24188), .o(n_24350) );
in01s03 g757128 ( .a(FE_OFN1183_n_24059), .o(n_27796) );
in01s02 g757135 ( .a(n_24059), .o(n_24188) );
in01s02 g757147 ( .a(FE_OFN780_n_23803), .o(n_24059) );
in01s02 g757159 ( .a(n_23743), .o(n_23803) );
in01s06 g757165 ( .a(n_23700), .o(n_23743) );
in01s08 g757168 ( .a(n_23671), .o(n_23700) );
in01s06 g757169 ( .a(n_23646), .o(n_23671) );
in01m06 g757170 ( .a(n_23616), .o(n_23646) );
oa12m08 g757171 ( .a(n_23185), .b(n_44996), .c(n_23118), .o(n_23616) );
ao12s01 g757172 ( .a(n_23182), .b(n_44995), .c(n_23117), .o(n_23592) );
ao12s01 g757173 ( .a(n_23531), .b(n_23530), .c(n_23529), .o(n_23860) );
ao12s01 g757174 ( .a(n_23534), .b(n_23533), .c(n_23532), .o(n_24087) );
oa12s01 g757175 ( .a(n_23528), .b(n_23527), .c(n_23526), .o(n_23670) );
ao22s01 g757176 ( .a(n_23493), .b(n_22880), .c(n_23492), .d(n_22881), .o(n_23645) );
ao22s02 g757178 ( .a(n_23489), .b(n_23152), .c(n_23488), .d(n_23153), .o(n_23802) );
no03s02 TIMEBOOST_cell_7978 ( .a(n_4368), .b(n_4846), .c(n_4369), .o(TIMEBOOST_net_2620) );
no02m02 TIMEBOOST_cell_1805 ( .a(n_21711), .b(n_21502), .o(TIMEBOOST_net_517) );
ao12f04 g757181 ( .a(n_23169), .b(n_23189), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_5_), .o(n_23216) );
in01s01 g757184 ( .a(n_23215), .o(n_23232) );
no02s04 g757185 ( .a(n_23193), .b(n_23192), .o(n_23215) );
na02s01 g757187 ( .a(FE_RN_72_0), .b(n_23190), .o(n_23366) );
na02s01 g757188 ( .a(n_23213), .b(n_23214), .o(n_23300) );
na02s01 g757189 ( .a(FE_RN_1657_0), .b(n_23133), .o(n_23309) );
na02s01 g757190 ( .a(n_23196), .b(n_23197), .o(n_23234) );
in01m04 g757195 ( .a(n_23195), .o(n_23212) );
na02m04 g757201 ( .a(n_23225), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_6_), .o(n_23289) );
in01m02 g757203 ( .a(n_23245), .o(n_23281) );
no02s04 g757204 ( .a(n_23225), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_6_), .o(n_23245) );
in01s06 g757205 ( .a(n_23378), .o(n_23113) );
no02s80 g757206 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_12_), .b(FE_OCP_RBN6540_n_44083), .o(n_23378) );
no02m80 g757209 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_14_), .b(FE_OCP_RBN6540_n_44083), .o(n_23079) );
no02s40 g757210 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_15_), .b(FE_OCP_RBN6540_n_44083), .o(n_23114) );
na02f06 g757211 ( .a(n_23193), .b(n_23192), .o(n_23249) );
na02s01 g757212 ( .a(n_23535), .b(n_22979), .o(n_23566) );
no02s01 g757213 ( .a(n_23533), .b(n_23532), .o(n_23534) );
in01s01 g757214 ( .a(n_23546), .o(n_23547) );
no02s01 g757215 ( .a(n_23491), .b(n_23181), .o(n_23546) );
in01m04 g757216 ( .a(n_23140), .o(n_23141) );
na02s08 g757217 ( .a(n_23112), .b(n_23111), .o(n_23140) );
no02s01 g757218 ( .a(n_23530), .b(n_23529), .o(n_23531) );
na02s01 g757219 ( .a(n_23527), .b(n_23526), .o(n_23528) );
no02s01 g757221 ( .a(n_44995), .b(n_23184), .o(n_23569) );
ao12f06 g757222 ( .a(n_23127), .b(n_44219), .c(n_23188), .o(n_23301) );
no02s01 g757223 ( .a(n_23490), .b(n_23060), .o(n_23549) );
in01s01 g757224 ( .a(n_23523), .o(n_23524) );
na02m04 TIMEBOOST_cell_3335 ( .a(TIMEBOOST_net_958), .b(n_11075), .o(n_11177) );
in01s01 g757226 ( .a(n_23521), .o(n_23522) );
ao12s01 g757227 ( .a(n_22954), .b(n_23495), .c(n_22809), .o(n_23521) );
na03m04 TIMEBOOST_cell_81 ( .a(n_12654), .b(n_12447), .c(n_12628), .o(n_12799) );
oa22s01 g757229 ( .a(n_44218), .b(n_23206), .c(n_44219), .d(n_23207), .o(n_24502) );
oa22s01 g757230 ( .a(n_23042), .b(n_23204), .c(n_23191), .d(n_23205), .o(n_24425) );
ao12m04 g757231 ( .a(n_23174), .b(n_23173), .c(n_23172), .o(n_23248) );
no02s08 TIMEBOOST_cell_2132 ( .a(TIMEBOOST_net_680), .b(n_10236), .o(n_10379) );
no02m06 g757236 ( .a(n_23173), .b(n_23172), .o(n_23174) );
na04s02 TIMEBOOST_cell_6557 ( .a(n_26884), .b(n_27033), .c(n_26885), .d(n_27034), .o(n_27093) );
na02s01 g757241 ( .a(n_23495), .b(n_22924), .o(n_23535) );
na02m08 g757243 ( .a(n_23110), .b(FE_OCP_RBN3979_n_22972), .o(n_23138) );
na02s01 g757244 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_5_), .b(n_23189), .o(n_23190) );
in01s01 g757245 ( .a(n_23210), .o(n_23211) );
no02s06 g757246 ( .a(n_23132), .b(n_23226), .o(n_23210) );
na02s01 g757247 ( .a(n_23494), .b(n_23183), .o(n_23533) );
in01s01 g757248 ( .a(n_23492), .o(n_23493) );
na02s01 g757249 ( .a(n_23469), .b(n_22852), .o(n_23492) );
no02m08 g757251 ( .a(n_23189), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_5_), .o(n_23208) );
no02m04 g757253 ( .a(n_23137), .b(delay_add_ln22_unr14_stage6_stallmux_q_5_), .o(n_23170) );
na02s02 g757254 ( .a(n_23136), .b(n_23135), .o(n_23214) );
na02s40 g757255 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_16_), .b(FE_OCP_RBN6540_n_44083), .o(n_23112) );
na02s20 g757256 ( .a(n_23004), .b(FE_OCP_RBN6539_n_44083), .o(n_23111) );
in01s01 g757257 ( .a(n_23169), .o(n_23213) );
no02m06 g757258 ( .a(n_23136), .b(n_23135), .o(n_23169) );
na02f06 g757260 ( .a(n_23069), .b(delay_add_ln22_unr14_stage6_stallmux_q_4_), .o(n_23197) );
na02s01 g757261 ( .a(n_23137), .b(delay_add_ln22_unr14_stage6_stallmux_q_5_), .o(n_23133) );
in01s01 g757263 ( .a(n_23490), .o(n_23491) );
no02s01 g757264 ( .a(n_23450), .b(n_23058), .o(n_23490) );
no02s01 g757265 ( .a(n_23451), .b(n_23026), .o(n_23530) );
no02s01 g757266 ( .a(n_23495), .b(n_22926), .o(n_23527) );
in01s01 g757267 ( .a(n_23488), .o(n_23489) );
oa12s02 g757268 ( .a(n_22732), .b(n_23468), .c(n_22843), .o(n_23488) );
ao12m08 g757270 ( .a(n_23023), .b(FE_OCP_RBN5533_n_44083), .c(delay_xor_ln22_unr15_stage6_stallmux_q_8_), .o(n_23047) );
in01m08 g757271 ( .a(n_23045), .o(n_23046) );
in01s01 g757273 ( .a(n_23107), .o(n_23108) );
in01m02 g757275 ( .a(n_23074), .o(n_23075) );
ao12m04 g757276 ( .a(n_23308), .b(FE_OCP_RBN5533_n_44083), .c(delay_xor_ln22_unr15_stage6_stallmux_q_10_), .o(n_23074) );
in01s01 g757277 ( .a(n_23278), .o(n_23279) );
ao12s01 g757278 ( .a(n_23224), .b(n_23223), .c(n_23222), .o(n_23278) );
ao12s01 g757279 ( .a(n_23073), .b(n_23072), .c(n_23071), .o(n_24361) );
ao12s01 g757280 ( .a(n_23449), .b(n_23468), .c(n_23448), .o(n_23804) );
ao22s01 g757283 ( .a(n_23417), .b(n_23201), .c(n_23416), .d(n_23202), .o(n_23985) );
in01s20 g757284 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_16_), .o(n_23004) );
in01s01 g757286 ( .a(n_23206), .o(n_23207) );
na02s01 g757287 ( .a(n_23188), .b(n_23128), .o(n_23206) );
no02s01 g757288 ( .a(n_23223), .b(n_23222), .o(n_23224) );
in01s01 g757289 ( .a(n_23204), .o(n_23205) );
na02s01 g757290 ( .a(FE_RN_1019_0), .b(n_23187), .o(n_23204) );
no02s01 g757291 ( .a(n_23072), .b(n_23071), .o(n_23073) );
na02s01 g757292 ( .a(n_23438), .b(n_22923), .o(n_23469) );
no02m80 g757294 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_8_), .b(FE_OCP_RBN3968_n_44061), .o(n_23023) );
no02s06 g757295 ( .a(FE_OCPN1653_n_23078), .b(n_23044), .o(n_23110) );
in01s03 g757296 ( .a(n_23173), .o(n_23132) );
no02s10 g757297 ( .a(n_23064), .b(FE_OCP_RBN2388_n_23227), .o(n_23173) );
in01s02 g757298 ( .a(n_23077), .o(n_23043) );
no02s40 g757299 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_11_), .b(FE_OCP_RBN5533_n_44083), .o(n_23077) );
no02m80 g757300 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_10_), .b(FE_OCP_RBN5533_n_44083), .o(n_23308) );
no02m40 g757301 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_13_), .b(FE_OCP_RBN5532_n_44083), .o(n_23022) );
no02s02 g757302 ( .a(n_23468), .b(n_22978), .o(n_23495) );
oa12s02 g757303 ( .a(n_23129), .b(n_23106), .c(FE_OCP_RBN6539_n_44083), .o(n_23335) );
ao12s10 g757305 ( .a(n_23462), .b(FE_OCP_RBN6541_n_44083), .c(delay_xor_ln21_unr15_stage6_stallmux_q_14_), .o(n_23167) );
in01s01 g757306 ( .a(n_23450), .o(n_23451) );
na02s01 g757307 ( .a(n_23438), .b(n_23437), .o(n_23450) );
no02s01 g757308 ( .a(n_23468), .b(n_23448), .o(n_23449) );
in01m01 g757309 ( .a(n_23165), .o(n_23166) );
ao12s20 g757310 ( .a(n_23131), .b(FE_OCP_RBN6541_n_44083), .c(delay_xor_ln21_unr15_stage6_stallmux_q_15_), .o(n_23165) );
in01s01 g757314 ( .a(n_23191), .o(n_23042) );
ao12m06 g757315 ( .a(n_22967), .b(n_23071), .c(n_23019), .o(n_23191) );
na02s04 TIMEBOOST_cell_7627 ( .a(TIMEBOOST_net_2444), .b(n_14363), .o(TIMEBOOST_net_850) );
no02s02 TIMEBOOST_cell_5071 ( .a(TIMEBOOST_net_1483), .b(n_13813), .o(n_13840) );
na02m06 g757333 ( .a(n_22970), .b(n_22937), .o(n_23002) );
na02s01 g757334 ( .a(n_23186), .b(n_23123), .o(n_23223) );
na02s01 g757335 ( .a(n_22968), .b(n_23019), .o(n_23072) );
na02m08 g757336 ( .a(n_23105), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_3_), .o(n_23188) );
in01s06 g757337 ( .a(n_23129), .o(n_23388) );
na02s40 g757338 ( .a(FE_OCP_RBN6539_n_44083), .b(n_23106), .o(n_23129) );
in01s01 g757339 ( .a(n_23127), .o(n_23128) );
no02f06 g757340 ( .a(n_23105), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_3_), .o(n_23127) );
no02s40 g757342 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_15_), .b(FE_OCP_RBN6541_n_44083), .o(n_23131) );
no02s40 g757343 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_14_), .b(FE_OCP_RBN6541_n_44083), .o(n_23462) );
in01m10 g757352 ( .a(n_23101), .o(n_23126) );
in01m10 g757353 ( .a(n_23064), .o(n_23101) );
no02f06 g757356 ( .a(n_23100), .b(delay_add_ln22_unr14_stage6_stallmux_q_3_), .o(n_23124) );
na02s06 g757357 ( .a(n_23100), .b(delay_add_ln22_unr14_stage6_stallmux_q_3_), .o(n_23187) );
na02s06 g757358 ( .a(n_23161), .b(n_23160), .o(n_23515) );
no02m10 g757360 ( .a(n_22912), .b(n_23078), .o(n_23000) );
in01s02 g757363 ( .a(n_23017), .o(n_23018) );
ao12s06 g757364 ( .a(n_23307), .b(FE_OCP_RBN5533_n_44083), .c(delay_xor_ln22_unr15_stage6_stallmux_q_9_), .o(n_23017) );
in01s01 g757365 ( .a(n_23416), .o(n_23417) );
ao12s01 g757366 ( .a(n_22918), .b(n_23400), .c(n_22808), .o(n_23416) );
in01m01 g757367 ( .a(n_23038), .o(n_23039) );
ao12m10 g757368 ( .a(n_23229), .b(FE_OCP_RBN2418_n_44083), .c(delay_xor_ln21_unr15_stage6_stallmux_q_8_), .o(n_23038) );
in01s01 g757369 ( .a(n_23438), .o(n_23468) );
ao12m06 g757370 ( .a(n_22953), .b(n_23400), .c(n_22922), .o(n_23438) );
in01s01 g757371 ( .a(FE_OCPN1346_n_24142), .o(n_24249) );
oa12s01 g757372 ( .a(n_23037), .b(n_23036), .c(n_23035), .o(n_24142) );
in01s01 g757374 ( .a(FE_OCP_DRV_N1426_n_24158), .o(n_24283) );
oa12s01 g757375 ( .a(n_22996), .b(n_22995), .c(n_22994), .o(n_24158) );
oa12s01 g757376 ( .a(n_23383), .b(n_23400), .c(n_23382), .o(n_23903) );
in01s01 g757377 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_31_), .o(n_22873) );
in01s40 g757381 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_12_), .o(n_23106) );
no02m10 g757383 ( .a(n_22828), .b(FE_OCP_RBN2369_n_44061), .o(n_22912) );
na02s01 g757384 ( .a(n_23036), .b(n_23035), .o(n_23037) );
na02s01 g757385 ( .a(n_22995), .b(n_22994), .o(n_22996) );
na02m06 g757386 ( .a(n_22942), .b(n_22941), .o(n_23019) );
in01m02 g757387 ( .a(n_22970), .o(n_22971) );
na02m08 g757388 ( .a(n_22945), .b(n_22944), .o(n_22970) );
no02s80 g757390 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_9_), .b(FE_OCP_RBN5528_n_44061), .o(n_23307) );
na02m06 g757391 ( .a(n_46964), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_2_), .o(n_23186) );
na02s10 g757392 ( .a(n_23034), .b(FE_OCP_RBN6539_n_44083), .o(n_23160) );
no02m40 g757393 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_8_), .b(FE_OCP_RBN3968_n_44061), .o(n_23229) );
na02m20 g757394 ( .a(n_23040), .b(n_23015), .o(n_23067) );
na02s10 g757395 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_16_), .b(FE_OCP_RBN6541_n_44083), .o(n_23161) );
in01s01 g757396 ( .a(n_23122), .o(n_23123) );
no02s06 g757397 ( .a(n_46964), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_2_), .o(n_23122) );
no02s80 g757399 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_6_), .b(FE_OCP_RBN3871_n_44061), .o(n_23078) );
no02s80 g757401 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_7_), .b(FE_OCP_RBN5529_n_44061), .o(n_22972) );
in01s01 g757402 ( .a(n_22967), .o(n_22968) );
no02m06 g757403 ( .a(n_22942), .b(n_22941), .o(n_22967) );
na02s01 g757404 ( .a(n_23400), .b(n_23382), .o(n_23383) );
ao12s03 g757406 ( .a(n_23461), .b(FE_OCP_RBN6541_n_44083), .c(delay_xor_ln21_unr15_stage6_stallmux_q_13_), .o(n_23097) );
in01m06 g757407 ( .a(n_22992), .o(n_22993) );
in01s02 g757409 ( .a(n_23095), .o(n_23096) );
ao12m01 g757410 ( .a(n_23391), .b(FE_OCP_RBN6541_n_44083), .c(delay_xor_ln21_unr15_stage6_stallmux_q_11_), .o(n_23095) );
in01s01 g757411 ( .a(n_23014), .o(n_23222) );
ao12m06 g757412 ( .a(n_22987), .b(n_22933), .c(n_22674), .o(n_23014) );
in01s04 g757413 ( .a(n_22965), .o(n_22966) );
na02f08 TIMEBOOST_cell_5099 ( .a(TIMEBOOST_net_1497), .b(n_29406), .o(n_29500) );
oa12s06 g757415 ( .a(n_23094), .b(n_23033), .c(n_44083), .o(n_23326) );
oa12m06 g757416 ( .a(n_22867), .b(n_22940), .c(n_22994), .o(n_23071) );
in01m02 g757421 ( .a(n_22914), .o(n_22871) );
na02m04 TIMEBOOST_cell_8744 ( .a(FE_OCP_RBN5630_n_33957), .b(n_33897), .o(TIMEBOOST_net_2859) );
ao12f08 g757428 ( .a(n_22991), .b(n_22990), .c(n_22989), .o(n_23105) );
in01s01 g757430 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_23_), .o(n_23773) );
in01m06 g757437 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_16_), .o(n_23034) );
in01m10 g757439 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_6_), .o(n_22828) );
no02m08 g757441 ( .a(n_22989), .b(n_22990), .o(n_22991) );
no02s02 TIMEBOOST_cell_6193 ( .a(n_35132), .b(n_47233), .o(TIMEBOOST_net_1948) );
na02s06 g757443 ( .a(n_22930), .b(n_22822), .o(n_22964) );
no02s01 g757444 ( .a(n_22934), .b(n_22987), .o(n_23036) );
no02s01 g757445 ( .a(n_22868), .b(n_22940), .o(n_22995) );
in01s20 g757446 ( .a(n_23094), .o(n_23390) );
na02s40 g757447 ( .a(n_23033), .b(n_44083), .o(n_23094) );
in01s06 g757448 ( .a(n_23461), .o(n_23032) );
no02s40 g757449 ( .a(FE_OCP_RBN5535_n_44083), .b(delay_xor_ln21_unr15_stage6_stallmux_q_13_), .o(n_23461) );
in01s01 g757450 ( .a(n_23391), .o(n_23031) );
no02s40 g757451 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_11_), .b(FE_OCP_RBN5534_n_44083), .o(n_23391) );
na02m40 g757452 ( .a(n_22939), .b(FE_OCP_RBN5175_n_44061), .o(n_23015) );
na02f02 TIMEBOOST_cell_7772 ( .a(FE_OCP_RBN5938_n_44563), .b(FE_OCP_RBN3136_n_10274), .o(TIMEBOOST_net_2517) );
in01s20 g757454 ( .a(n_22869), .o(n_22944) );
no02s40 g757455 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_4_), .b(FE_OCP_RBN6466_n_44061), .o(n_22869) );
oa12m06 g757456 ( .a(n_22951), .b(n_23299), .c(n_22921), .o(n_23400) );
oa12s06 g757457 ( .a(n_22959), .b(n_44083), .c(n_22935), .o(n_23172) );
in01s06 g757458 ( .a(n_23011), .o(n_23012) );
ao12s10 g757459 ( .a(FE_OCP_RBN2388_n_23227), .b(FE_OCP_RBN3968_n_44061), .c(delay_xor_ln21_unr15_stage6_stallmux_q_6_), .o(n_23011) );
in01s06 g757460 ( .a(n_22937), .o(n_22938) );
in01s01 g757465 ( .a(n_22835), .o(n_22804) );
in01s01 g757467 ( .a(n_23954), .o(n_23979) );
oa12s01 g757468 ( .a(n_23344), .b(n_23343), .c(n_23342), .o(n_23954) );
in01s01 g757469 ( .a(n_23901), .o(n_23399) );
ao12s01 g757470 ( .a(n_23358), .b(n_23357), .c(n_23356), .o(n_23901) );
in01s01 g757474 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_29_), .o(n_22936) );
in01s40 g757477 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_10_), .o(n_23033) );
in01s10 g757481 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_4_), .o(n_22803) );
in01s40 g757483 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_4_), .o(n_22939) );
in01m04 g757485 ( .a(n_22945), .o(n_22900) );
no02f10 g757486 ( .a(n_22823), .b(n_22822), .o(n_22945) );
in01m10 g757487 ( .a(n_22959), .o(n_23226) );
na02m40 g757488 ( .a(n_22935), .b(FE_OCP_RBN2369_n_44061), .o(n_22959) );
na02s02 TIMEBOOST_cell_5640 ( .a(n_6082), .b(n_5845), .o(TIMEBOOST_net_1768) );
no02m40 g757491 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_6_), .b(FE_OCP_RBN2250_n_44061), .o(n_23227) );
in01s01 g757492 ( .a(n_22933), .o(n_22934) );
na02m06 g757493 ( .a(n_22899), .b(n_22898), .o(n_22933) );
in01m06 g757494 ( .a(n_23040), .o(n_22985) );
no02s01 g757496 ( .a(n_23357), .b(n_23356), .o(n_23358) );
no02s06 g757497 ( .a(n_22899), .b(n_22898), .o(n_22987) );
in01s01 g757498 ( .a(n_22867), .o(n_22868) );
na02m06 g757499 ( .a(n_22827), .b(delay_add_ln22_unr14_stage6_stallmux_q_1_), .o(n_22867) );
no02m08 TIMEBOOST_cell_3912 ( .a(TIMEBOOST_net_1046), .b(FE_OCP_RBN4171_n_19390), .o(n_19605) );
no02m06 g757501 ( .a(n_22827), .b(delay_add_ln22_unr14_stage6_stallmux_q_1_), .o(n_22940) );
no02m10 g757502 ( .a(n_22864), .b(FE_OCP_RBN2390_FE_RN_1364_0), .o(n_22989) );
in01m01 g757503 ( .a(n_23029), .o(n_23030) );
ao12s10 g757504 ( .a(n_23322), .b(FE_OCP_RBN5536_n_44083), .c(delay_xor_ln21_unr15_stage6_stallmux_q_9_), .o(n_23029) );
in01m04 g757505 ( .a(n_22930), .o(n_22931) );
na02s01 g757507 ( .a(n_23343), .b(n_23342), .o(n_23344) );
in01f02 g757513 ( .a(n_22778), .o(n_22757) );
in01m02 g757515 ( .a(n_22806), .o(n_22776) );
in01m02 g757517 ( .a(n_22829), .o(n_22800) );
oa12s04 g757519 ( .a(n_22153), .b(n_22639), .c(n_22128), .o(n_22722) );
ao12m06 g757520 ( .a(n_22196), .b(FE_OCP_RBN6232_n_22639), .c(n_22129), .o(n_22756) );
ao22m04 g757522 ( .a(n_22686), .b(n_22343), .c(n_22720), .d(n_22306), .o(n_22755) );
oa12s02 g757523 ( .a(n_22305), .b(n_22720), .c(n_22221), .o(n_22721) );
ao12s02 g757524 ( .a(n_22342), .b(n_22686), .c(n_22220), .o(n_22687) );
oa12s02 g757525 ( .a(n_22349), .b(n_22686), .c(n_22194), .o(n_22685) );
ao12s02 g757526 ( .a(n_22313), .b(n_22720), .c(n_22214), .o(n_22719) );
ao12s01 g757527 ( .a(n_23297), .b(n_23298), .c(n_23296), .o(n_23978) );
oa12s01 g757528 ( .a(n_23321), .b(n_23320), .c(n_23319), .o(n_23801) );
in01s01 g757529 ( .a(n_23897), .o(n_23341) );
ao22s01 g757530 ( .a(n_23261), .b(n_22726), .c(n_23260), .d(n_22727), .o(n_23897) );
in01s01 g757531 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_22_), .o(n_22754) );
in01s01 g757533 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_), .o(n_22717) );
in01s01 g757535 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_24_), .o(n_23653) );
in01s40 g757539 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_7_), .o(n_22935) );
in01s01 g757541 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_31_), .o(n_22929) );
na02s01 g757545 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_19_), .b(delay_add_ln22_unr14_stage6_stallmux_q_18_), .o(n_22773) );
no02m06 g757546 ( .a(n_23298), .b(n_23295), .o(n_23299) );
na02s01 g757547 ( .a(n_23320), .b(n_23319), .o(n_23321) );
in01s02 g757549 ( .a(FE_OCPN1906_n_23322), .o(n_22984) );
no02s40 g757550 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_9_), .b(FE_OCP_RBN3968_n_44061), .o(n_23322) );
no02s40 g757553 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_3_), .b(FE_OCP_RBN3871_n_44061), .o(n_22823) );
no02s10 g757555 ( .a(FE_OCP_RBN6471_delay_xor_ln21_unr15_stage6_stallmux_q_3_), .b(n_44061), .o(n_22864) );
no02s01 g757561 ( .a(n_23298), .b(n_23296), .o(n_23297) );
in01m04 g757562 ( .a(n_22771), .o(n_22772) );
no02m20 g757565 ( .a(n_22817), .b(n_22796), .o(n_22927) );
no03m40 TIMEBOOST_cell_3456 ( .a(n_32820), .b(n_32613), .c(FE_OCP_RBN6526_n_44962), .o(n_32678) );
na02s02 TIMEBOOST_cell_3918 ( .a(TIMEBOOST_net_1049), .b(n_7804), .o(n_9003) );
in01s02 g757575 ( .a(n_22902), .o(n_22862) );
in01s02 g757577 ( .a(n_22901), .o(n_22861) );
oa12s01 g757582 ( .a(n_22888), .b(n_23243), .c(n_23295), .o(n_23343) );
in01s02 g757584 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_19_), .o(n_23611) );
in01s03 g757588 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_19_), .o(n_23605) );
in01s01 g757593 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_26_), .o(n_22859) );
in01s01 g757595 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_25_), .o(n_22858) );
no02s06 TIMEBOOST_cell_8816 ( .a(n_15114), .b(FE_OCPN1077_n_13831), .o(TIMEBOOST_net_2895) );
na02s01 g757599 ( .a(n_23276), .b(n_22812), .o(n_23320) );
in01s10 g757600 ( .a(n_22816), .o(n_22817) );
na02m40 g757601 ( .a(n_22795), .b(n_44061), .o(n_22816) );
no02s20 g757602 ( .a(n_22795), .b(n_44061), .o(n_22796) );
no02m06 g757603 ( .a(n_23242), .b(n_22887), .o(n_23298) );
no02s80 g757605 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_5_), .b(FE_OCP_RBN2250_n_44061), .o(n_22889) );
no02s06 g757608 ( .a(n_22601), .b(n_22473), .o(n_22686) );
in01s01 g757609 ( .a(n_23260), .o(n_23261) );
oa12s01 g757610 ( .a(n_22643), .b(n_23221), .c(n_22729), .o(n_23260) );
in01s01 g757611 ( .a(n_24097), .o(n_22752) );
oa12s01 g757612 ( .a(n_22633), .b(n_22632), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_0_), .o(n_24097) );
in01s01 g757613 ( .a(n_24119), .o(n_22767) );
ao12s01 g757614 ( .a(n_22676), .b(n_22675), .c(delay_add_ln22_unr14_stage6_stallmux_q_0_), .o(n_24119) );
na02m08 g757621 ( .a(n_22584), .b(n_22314), .o(n_22639) );
in01m02 g757622 ( .a(n_22684), .o(n_22637) );
oa12s04 g757626 ( .a(n_22047), .b(n_22564), .c(n_22164), .o(n_22603) );
ao12f04 g757627 ( .a(n_22078), .b(FE_OCP_RBN3417_n_22564), .c(n_22079), .o(n_22619) );
oa12s06 g757630 ( .a(n_22271), .b(n_45497), .c(n_22130), .o(n_22636) );
ao12s06 g757631 ( .a(n_22308), .b(n_45496), .c(n_22131), .o(n_22618) );
na02s06 TIMEBOOST_cell_2835 ( .a(n_7389), .b(TIMEBOOST_net_708), .o(n_7456) );
in01s02 g757633 ( .a(n_22774), .o(n_22751) );
in01s02 g757635 ( .a(n_22897), .o(n_22856) );
in01s01 g757637 ( .a(n_23746), .o(n_23294) );
oa22s01 g757638 ( .a(n_23244), .b(n_22762), .c(n_23220), .d(n_22761), .o(n_23746) );
in01s02 g757639 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_20_), .o(n_23658) );
in01m40 g757646 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_2_), .o(n_22795) );
na02s08 g757649 ( .a(n_22769), .b(n_22634), .o(n_22677) );
na02s20 g757651 ( .a(n_22820), .b(n_22708), .o(n_22748) );
na02s01 g757652 ( .a(n_23244), .b(n_22763), .o(n_23276) );
na02s01 g757653 ( .a(n_22632), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_0_), .o(n_22633) );
no02s01 g757654 ( .a(n_22675), .b(delay_add_ln22_unr14_stage6_stallmux_q_0_), .o(n_22676) );
in01s01 g757655 ( .a(n_22674), .o(n_23035) );
na02s06 g757657 ( .a(n_22613), .b(delay_add_ln22_unr14_stage6_stallmux_q_0_), .o(n_22994) );
na02m06 g757658 ( .a(n_45499), .b(n_22231), .o(n_22584) );
in01m06 g757659 ( .a(n_22672), .o(n_22673) );
in01m08 g757661 ( .a(n_22746), .o(n_22747) );
in01s01 g757663 ( .a(n_23242), .o(n_23243) );
oa12s02 g757665 ( .a(n_22439), .b(n_22705), .c(FE_OCP_RBN4485_n_22667), .o(n_22707) );
no02s04 g757666 ( .a(n_22668), .b(n_22413), .o(n_22745) );
oa12s02 g757668 ( .a(n_22330), .b(n_22461), .c(n_22705), .o(n_22706) );
in01f02 g757672 ( .a(n_22640), .o(n_22617) );
no02s04 g757674 ( .a(n_22542), .b(n_22273), .o(n_22601) );
in01f02 g757676 ( .a(n_22819), .o(n_22792) );
oa12s04 g757678 ( .a(n_22417), .b(n_22625), .c(n_22415), .o(n_22703) );
ao12f04 g757679 ( .a(FE_OCPN1248_n_22291), .b(FE_OCP_RBN4649_n_22625), .c(FE_OCPN4832_n_22294), .o(n_22743) );
in01f02 g757680 ( .a(n_22715), .o(n_22670) );
in01s02 g757684 ( .a(n_22790), .o(n_22857) );
in01s01 g757686 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_18_), .o(n_22669) );
in01s01 g757688 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_18_), .o(n_22630) );
in01s01 g757695 ( .a(n_23244), .o(n_23220) );
in01s01 g757696 ( .a(n_23221), .o(n_23244) );
ao12m04 g757697 ( .a(n_23088), .b(n_23090), .c(FE_OCP_RBN3879_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n_23221) );
no02s04 g757698 ( .a(n_22705), .b(FE_OCP_RBN4485_n_22667), .o(n_22668) );
oa22m02 g757701 ( .a(n_22540), .b(FE_OCPN1394_n_22801), .c(n_22514), .d(n_22580), .o(n_22581) );
in01f02 g757702 ( .a(n_22635), .o(n_22614) );
oa22f02 g757703 ( .a(n_22513), .b(n_22312), .c(n_22543), .d(n_22346), .o(n_22635) );
oa12m02 g757704 ( .a(n_22311), .b(n_22543), .c(n_22344), .o(n_22544) );
ao12m04 g757705 ( .a(n_22345), .b(n_22513), .c(n_22046), .o(n_22566) );
oa12f08 g757709 ( .a(n_22170), .b(n_22543), .c(n_22138), .o(n_22564) );
ao12s06 g757716 ( .a(n_22171), .b(n_22450), .c(n_22139), .o(n_22542) );
in01s01 g757717 ( .a(n_22613), .o(n_22675) );
no02m02 TIMEBOOST_cell_6682 ( .a(TIMEBOOST_net_2098), .b(n_8474), .o(TIMEBOOST_net_1892) );
oa12s01 g757724 ( .a(n_23156), .b(n_23155), .c(n_23154), .o(n_23699) );
in01s01 g757725 ( .a(n_23807), .o(n_24111) );
ao12s01 g757726 ( .a(n_23159), .b(n_23158), .c(n_23157), .o(n_23807) );
oa22f04 g757728 ( .a(n_22556), .b(n_22299), .c(FE_OCP_RBN5347_n_22556), .d(n_22335), .o(n_22709) );
oa12s02 g757729 ( .a(FE_OCP_RBN5216_n_22212), .b(n_22556), .c(FE_OCP_RBN5387_n_22149), .o(n_22598) );
ao12s04 g757730 ( .a(FE_OCP_RBN5217_n_22212), .b(FE_OCP_RBN5346_n_22556), .c(FE_OCP_RBN5388_n_22149), .o(n_22612) );
in01s03 g757731 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_), .o(n_22562) );
in01s40 g757736 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_1_), .o(n_22597) );
in01s06 g757738 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_17_), .o(n_23562) );
no02s04 TIMEBOOST_cell_6845 ( .a(n_26407), .b(n_23353), .o(TIMEBOOST_net_2180) );
no02m04 g757741 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_0_), .b(n_44061), .o(n_22560) );
na02m04 TIMEBOOST_cell_5175 ( .a(TIMEBOOST_net_1535), .b(n_8952), .o(n_9271) );
na02m40 g757744 ( .a(n_22537), .b(n_44061), .o(n_22820) );
no02s01 g757745 ( .a(n_23158), .b(n_23157), .o(n_23159) );
in01s06 g757746 ( .a(n_22769), .o(n_22575) );
na02s01 g757748 ( .a(n_23155), .b(n_23154), .o(n_23156) );
na02s06 g757752 ( .a(n_22591), .b(n_22470), .o(n_22705) );
oa12m08 g757756 ( .a(n_22327), .b(FE_OCP_RBN4646_n_22553), .c(FE_OCPN5238_n_22383), .o(n_22625) );
in01s02 g757757 ( .a(n_22739), .o(n_22789) );
in01m02 g757759 ( .a(n_46965), .o(n_22594) );
oa12m04 g757761 ( .a(n_44288), .b(n_22482), .c(n_22481), .o(n_22518) );
no02f04 g757762 ( .a(n_22483), .b(n_44287), .o(n_22538) );
oa12f08 g757763 ( .a(n_22466), .b(n_22589), .c(n_22406), .o(n_22661) );
ao12m04 g757764 ( .a(n_22432), .b(FE_OCP_RBN4647_n_22553), .c(n_22465), .o(n_22624) );
in01m02 g757766 ( .a(n_22631), .o(n_22611) );
oa12s01 g757768 ( .a(n_23093), .b(n_23092), .c(n_23091), .o(n_23800) );
oa12f04 g757769 ( .a(FE_OCP_RBN5215_n_22150), .b(n_22531), .c(n_22468), .o(n_22574) );
ao12s04 g757770 ( .a(FE_OCP_RBN5214_n_22150), .b(n_22511), .c(n_22507), .o(n_22558) );
in01m40 g757771 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_0_), .o(n_22537) );
na02s01 g757776 ( .a(n_23092), .b(n_23091), .o(n_23093) );
na02s01 g757777 ( .a(n_23089), .b(n_23087), .o(n_23158) );
na02m04 g757778 ( .a(n_23089), .b(n_22657), .o(n_23090) );
na02f02 g757780 ( .a(n_22482), .b(n_22347), .o(n_22536) );
no02f06 g757781 ( .a(n_22482), .b(n_22481), .o(n_22483) );
no03s04 TIMEBOOST_cell_7109 ( .a(n_17289), .b(n_17485), .c(n_17410), .o(n_17517) );
oa12s01 g757783 ( .a(n_23087), .b(n_23010), .c(n_22697), .o(n_23155) );
oa22f02 g757784 ( .a(n_22479), .b(n_20231), .c(n_22443), .d(n_22580), .o(n_22535) );
oa22f02 g757785 ( .a(n_22425), .b(FE_OCPN1394_n_22801), .c(n_22390), .d(n_22580), .o(n_22480) );
in01m02 g757786 ( .a(n_22540), .o(n_22514) );
oa22m04 g757787 ( .a(n_22358), .b(n_22108), .c(n_22391), .d(n_22109), .o(n_22540) );
in01f04 g757790 ( .a(n_22543), .o(n_22513) );
in01f06 g757791 ( .a(n_22450), .o(n_22543) );
oa12f06 g757793 ( .a(n_22436), .b(n_22554), .c(FE_OCP_RBN5344_n_22476), .o(n_22573) );
no02f06 TIMEBOOST_cell_6758 ( .a(TIMEBOOST_net_2136), .b(n_4713), .o(n_4887) );
in01f02 g757801 ( .a(n_22596), .o(n_22570) );
in01s01 g757805 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_16_), .o(n_23603) );
in01s01 g757807 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_16_), .o(n_23560) );
na02s06 TIMEBOOST_cell_8007 ( .a(TIMEBOOST_net_2634), .b(n_39964), .o(n_40063) );
no02m04 g757810 ( .a(n_23027), .b(n_22655), .o(n_23089) );
no02m04 g757811 ( .a(n_23121), .b(n_23120), .o(n_23185) );
na02s01 g757812 ( .a(n_23183), .b(n_23116), .o(n_23184) );
no02s01 g757813 ( .a(n_23009), .b(n_22693), .o(n_23092) );
na02s01 g757814 ( .a(n_23183), .b(n_23119), .o(n_23182) );
no02f08 g757817 ( .a(n_22357), .b(n_22172), .o(n_22482) );
na02s10 TIMEBOOST_cell_2863 ( .a(n_37489), .b(TIMEBOOST_net_722), .o(n_37593) );
oa22s02 g757819 ( .a(n_22392), .b(n_20231), .c(n_22355), .d(n_22580), .o(n_22449) );
oa22f02 g757820 ( .a(n_22359), .b(FE_OCPN1394_n_22801), .c(n_22317), .d(n_22580), .o(n_22424) );
in01m04 g757823 ( .a(n_22511), .o(n_22531) );
na02m08 g757824 ( .a(n_22423), .b(n_22388), .o(n_22511) );
in01s01 g757825 ( .a(n_23698), .o(n_23061) );
oa12s01 g757826 ( .a(n_22982), .b(n_22983), .c(n_22981), .o(n_23698) );
in01m06 g757829 ( .a(FE_OCP_RBN4647_n_22553), .o(n_22589) );
na02m08 g757832 ( .a(n_22447), .b(n_22472), .o(n_22553) );
in01s01 g757833 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_15_), .o(n_23554) );
na02s01 g757836 ( .a(n_23085), .b(n_23052), .o(n_23086) );
in01s01 g757837 ( .a(n_23009), .o(n_23010) );
no02s01 g757838 ( .a(n_22983), .b(n_22694), .o(n_23009) );
na02s01 g757839 ( .a(n_22983), .b(n_22981), .o(n_22982) );
no02f06 g757845 ( .a(n_22446), .b(n_22448), .o(n_22476) );
no02m06 g757846 ( .a(n_22983), .b(n_22765), .o(n_23027) );
na02s02 g757847 ( .a(n_22318), .b(n_21970), .o(n_22358) );
no02s04 g757848 ( .a(n_22319), .b(n_22002), .o(n_22391) );
in01f03 g757849 ( .a(n_22356), .o(n_22357) );
na02f08 g757850 ( .a(n_22279), .b(n_22084), .o(n_22356) );
na02m04 g757851 ( .a(n_22389), .b(FE_OCP_RBN5049_FE_RN_606_0), .o(n_22423) );
na02s06 g757852 ( .a(n_22446), .b(n_22445), .o(n_22447) );
na02s04 g757853 ( .a(n_22421), .b(n_22064), .o(n_22444) );
no02f04 g757854 ( .a(FE_OCP_RBN6211_n_22421), .b(n_22145), .o(n_22475) );
in01s01 g757855 ( .a(n_23121), .o(n_23183) );
oa12s04 g757856 ( .a(n_23085), .b(n_23007), .c(FE_OFN745_n_22641), .o(n_23121) );
in01f02 g757857 ( .a(n_22425), .o(n_22390) );
oa22f04 g757858 ( .a(n_22239), .b(n_22018), .c(n_22238), .d(n_22019), .o(n_22425) );
in01m02 g757859 ( .a(n_22479), .o(n_22443) );
oa22f02 g757860 ( .a(n_22237), .b(n_22183), .c(n_22316), .d(n_22184), .o(n_22479) );
na02s01 g757861 ( .a(n_23008), .b(n_22840), .o(n_23060) );
in01s02 g757862 ( .a(n_22318), .o(n_22319) );
in01s02 g757863 ( .a(n_22279), .o(n_22318) );
no02f08 g757864 ( .a(n_22205), .b(n_22003), .o(n_22279) );
no02s02 g757865 ( .a(n_22473), .b(n_22420), .o(n_22474) );
oa12m06 g757866 ( .a(n_22445), .b(n_22448), .c(n_22352), .o(n_22472) );
in01f02 g757868 ( .a(n_22389), .o(n_22421) );
no02f06 g757869 ( .a(n_22237), .b(n_22063), .o(n_22389) );
ao12s04 g757870 ( .a(n_23026), .b(n_22841), .c(n_22725), .o(n_23085) );
ao12s02 g757871 ( .a(FE_OFN745_n_22641), .b(n_23119), .c(n_23056), .o(n_23120) );
in01m02 g757873 ( .a(n_22359), .o(n_22317) );
oa22f04 g757874 ( .a(n_22169), .b(n_21971), .c(n_22140), .d(n_21972), .o(n_22359) );
in01s02 g757876 ( .a(n_22392), .o(n_22355) );
oa22s04 g757877 ( .a(n_22095), .b(n_22168), .c(n_22094), .d(n_22204), .o(n_22392) );
in01s01 g757879 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_14_), .o(n_22354) );
na02s01 g757881 ( .a(n_22979), .b(n_22879), .o(n_22980) );
in01m02 g757882 ( .a(n_22238), .o(n_22239) );
in01m02 g757883 ( .a(n_22205), .o(n_22238) );
oa12f08 g757884 ( .a(n_21954), .b(n_22088), .c(n_21941), .o(n_22205) );
in01s01 g757885 ( .a(n_22237), .o(n_22316) );
oa12f08 g757889 ( .a(n_22065), .b(n_22113), .c(n_22035), .o(n_22237) );
in01s01 g757890 ( .a(n_23026), .o(n_23008) );
na02s04 g757891 ( .a(n_22979), .b(n_22848), .o(n_23026) );
ao12s04 g757892 ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(n_22854), .c(n_22658), .o(n_22855) );
in01s01 g757894 ( .a(n_23812), .o(n_23869) );
ao12s01 g757895 ( .a(n_22814), .b(n_22854), .c(n_22813), .o(n_23812) );
na02m06 TIMEBOOST_cell_1492 ( .a(TIMEBOOST_net_360), .b(n_29634), .o(n_29648) );
na02s02 g757898 ( .a(n_23083), .b(n_23117), .o(n_23118) );
no02s01 g757899 ( .a(n_22887), .b(n_22730), .o(n_22888) );
na02s01 g757900 ( .a(n_22884), .b(n_22783), .o(n_22954) );
no03s10 TIMEBOOST_cell_5710 ( .a(TIMEBOOST_net_1197), .b(n_32716), .c(n_32871), .o(n_32990) );
oa12s04 g757902 ( .a(n_22170), .b(n_22082), .c(n_44277), .o(n_22171) );
na02s06 g757903 ( .a(n_22314), .b(n_22234), .o(n_22473) );
no03m04 TIMEBOOST_cell_8330 ( .a(n_42277), .b(n_41955), .c(n_42283), .o(n_42330) );
ao12s01 g757906 ( .a(n_23055), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_29_), .o(n_23568) );
ao12s06 g757908 ( .a(n_22926), .b(n_22784), .c(n_22725), .o(n_22979) );
no02s01 g757909 ( .a(n_22854), .b(n_22813), .o(n_22814) );
ao12s01 g757910 ( .a(n_23084), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_30_), .o(n_23591) );
oa12s02 g757911 ( .a(n_22725), .b(n_22952), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_29_), .o(n_23119) );
no02s02 g757912 ( .a(n_22978), .b(n_22925), .o(n_23437) );
ao12f08 g757913 ( .a(n_22186), .b(n_22388), .c(n_22269), .o(n_22448) );
oa22s01 g757914 ( .a(n_22110), .b(n_21998), .c(n_22086), .d(n_21997), .o(n_22236) );
oa12s02 g757915 ( .a(n_21936), .b(n_22086), .c(n_21937), .o(n_22140) );
ao12s02 g757916 ( .a(n_21921), .b(n_22110), .c(n_21922), .o(n_22169) );
oa22s01 g757917 ( .a(n_22106), .b(n_22032), .c(FE_OCP_RBN6179_n_22106), .d(n_22033), .o(n_22275) );
oa12s02 g757918 ( .a(n_22012), .b(n_22106), .c(n_21982), .o(n_22168) );
ao12s02 g757919 ( .a(n_21960), .b(FE_OCP_RBN6178_n_22106), .c(n_21961), .o(n_22204) );
no04s02 g757920 ( .a(n_23181), .b(n_23057), .c(n_23006), .d(n_23058), .o(n_23059) );
in01s01 g757921 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_13_), .o(n_22203) );
in01s01 g757923 ( .a(n_23083), .o(n_23084) );
na02s01 g757924 ( .a(n_23056), .b(FE_OFN745_n_22641), .o(n_23083) );
in01s01 g757925 ( .a(n_23055), .o(n_23117) );
no02s01 g757926 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_29_), .o(n_23055) );
na02s01 g757927 ( .a(n_22852), .b(n_22652), .o(n_22853) );
oa12s02 g757928 ( .a(n_22812), .b(n_22731), .c(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n_22887) );
ao12s06 g757929 ( .a(FE_OCP_RBN2386_n_22650), .b(n_22785), .c(n_22728), .o(n_22854) );
no02f06 g757930 ( .a(n_22049), .b(n_21921), .o(n_22088) );
ao12s01 g757931 ( .a(n_23057), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_27_), .o(n_23647) );
ao12s02 g757933 ( .a(n_22326), .b(n_22332), .c(n_22288), .o(n_22470) );
no02f08 g757934 ( .a(n_22080), .b(n_21960), .o(n_22113) );
in01s01 g757935 ( .a(n_22926), .o(n_22884) );
na02s06 g757936 ( .a(n_22852), .b(n_22736), .o(n_22926) );
na02s02 g757937 ( .a(n_22924), .b(n_22851), .o(n_22925) );
na02m06 g757938 ( .a(n_22268), .b(n_22351), .o(n_22352) );
in01s01 g757939 ( .a(n_22811), .o(n_22885) );
ao12s01 g757940 ( .a(n_22788), .b(n_22737), .c(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_22811) );
oa22s01 g757941 ( .a(n_22021), .b(n_21938), .c(n_22020), .d(n_21939), .o(n_22112) );
ao12m06 g757942 ( .a(n_22027), .b(n_22085), .c(n_21970), .o(n_22172) );
no02s06 g757944 ( .a(n_22138), .b(n_22081), .o(n_22139) );
in01s06 g757945 ( .a(n_22235), .o(n_22314) );
na02s01 TIMEBOOST_cell_1434 ( .a(TIMEBOOST_net_331), .b(n_34174), .o(n_34231) );
in01s02 g757947 ( .a(n_22233), .o(n_22234) );
no02m06 TIMEBOOST_cell_7023 ( .a(TIMEBOOST_net_1300), .b(n_26045), .o(TIMEBOOST_net_2270) );
in01s01 g757952 ( .a(n_22313), .o(n_22349) );
no02s02 g757953 ( .a(FE_OCP_RBN4462_n_44267), .b(n_22201), .o(n_22313) );
in01s01 g757954 ( .a(n_22882), .o(n_22883) );
ao12s01 g757955 ( .a(n_22787), .b(n_22786), .c(n_22785), .o(n_22882) );
in01s01 g757956 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_12_), .o(n_23475) );
in01s01 g757959 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_30_), .o(n_23056) );
no02s01 g757961 ( .a(n_22849), .b(n_22850), .o(n_22851) );
no02s01 g757962 ( .a(n_22950), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_27_), .o(n_23007) );
no02s01 g757963 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_27_), .o(n_23057) );
na02s01 g757964 ( .a(n_23116), .b(n_23054), .o(n_23532) );
no02s04 g757965 ( .a(n_22660), .b(n_22649), .o(n_22738) );
no02s01 g757966 ( .a(n_22737), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_22788) );
ao12s01 g757967 ( .a(n_23181), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_25_), .o(n_23548) );
in01s02 g757970 ( .a(n_22086), .o(n_22110) );
in01s01 g757971 ( .a(n_22049), .o(n_22086) );
oa12f04 g757972 ( .a(n_21925), .b(n_21974), .c(n_21906), .o(n_22049) );
in01s02 g757973 ( .a(n_22108), .o(n_22109) );
na02m02 g757974 ( .a(n_22085), .b(n_22084), .o(n_22108) );
no02f06 g757976 ( .a(n_22481), .b(n_44287), .o(n_22347) );
na02s01 g757978 ( .a(n_22311), .b(n_22046), .o(n_22312) );
no02s02 g757979 ( .a(n_22345), .b(n_22344), .o(n_22346) );
na02s06 g757980 ( .a(n_22083), .b(n_22046), .o(n_22138) );
na02s01 g757981 ( .a(n_22079), .b(n_22047), .o(n_22167) );
no02s02 g757982 ( .a(n_22164), .b(n_22078), .o(n_22165) );
no02s02 g757983 ( .a(n_22048), .b(FE_OCP_RBN7049_n_20941), .o(n_22082) );
na02s02 g757984 ( .a(n_22271), .b(n_22131), .o(n_22272) );
no02s01 g757985 ( .a(n_22308), .b(n_22130), .o(n_22309) );
na02s01 g757986 ( .a(n_22153), .b(n_22129), .o(n_22270) );
no02s02 g757987 ( .a(n_22196), .b(n_22128), .o(n_22307) );
no02m04 TIMEBOOST_cell_8633 ( .a(TIMEBOOST_net_2803), .b(n_4179), .o(n_4436) );
na02s06 g757989 ( .a(n_22305), .b(n_22220), .o(n_22306) );
no02s01 g757990 ( .a(n_22221), .b(n_22342), .o(n_22343) );
no02s06 TIMEBOOST_cell_1264 ( .a(TIMEBOOST_net_246), .b(FE_OCP_RBN4114_n_33533), .o(n_33628) );
no02s01 g757992 ( .a(n_22194), .b(n_47278), .o(n_22230) );
na02s01 g757994 ( .a(n_22923), .b(n_22847), .o(n_22978) );
na02s02 g757995 ( .a(n_22698), .b(n_22621), .o(n_22765) );
ao12s01 g757997 ( .a(n_22849), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_23_), .o(n_23618) );
no02s01 g757998 ( .a(n_22786), .b(n_22785), .o(n_22787) );
na02s01 TIMEBOOST_cell_1433 ( .a(n_33672), .b(n_33653), .o(TIMEBOOST_net_331) );
na02s06 g758000 ( .a(n_22047), .b(n_22022), .o(n_22081) );
oa12s01 g758001 ( .a(n_22725), .b(n_22759), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_23_), .o(n_22848) );
oa12s06 g758002 ( .a(n_22725), .b(n_22734), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_19_), .o(n_22736) );
na02s06 g758003 ( .a(n_22733), .b(n_22725), .o(n_22852) );
oa12s02 g758004 ( .a(n_22725), .b(n_22917), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_15_), .o(n_22922) );
na02f08 g758006 ( .a(n_22200), .b(n_22121), .o(n_22269) );
na02s01 g758007 ( .a(n_22263), .b(n_22083), .o(n_22303) );
no02s02 g758008 ( .a(n_22264), .b(n_22045), .o(n_22341) );
na02s02 g758009 ( .a(n_22261), .b(n_22300), .o(n_22340) );
no02s03 g758010 ( .a(n_22262), .b(n_22301), .o(n_22387) );
in01s01 g758011 ( .a(n_22338), .o(n_22339) );
na02s06 TIMEBOOST_cell_4966 ( .a(n_32912), .b(FE_OCP_RBN2453_n_32860), .o(TIMEBOOST_net_1431) );
in01s01 g758013 ( .a(n_22336), .o(n_22337) );
na02s01 TIMEBOOST_cell_1260 ( .a(TIMEBOOST_net_244), .b(n_33533), .o(n_33863) );
in01s01 g758015 ( .a(n_22385), .o(n_22386) );
na02s02 g758016 ( .a(n_22216), .b(n_22258), .o(n_22385) );
na02m08 g758017 ( .a(n_22155), .b(FE_OCP_RBN5050_FE_RN_606_0), .o(n_22388) );
na03m10 TIMEBOOST_cell_4573 ( .a(n_11774), .b(n_45224), .c(FE_RN_2499_0), .o(n_11788) );
oa22s01 g758020 ( .a(n_22015), .b(n_21962), .c(n_22014), .d(n_21963), .o(n_22107) );
in01s02 g758025 ( .a(n_22080), .o(n_22106) );
ao12f08 g758026 ( .a(n_21910), .b(n_21999), .c(n_21947), .o(n_22080) );
in01s02 g758028 ( .a(n_22381), .o(n_22382) );
na02m02 TIMEBOOST_cell_5492 ( .a(n_10667), .b(n_10736), .o(TIMEBOOST_net_1694) );
in01s01 g758030 ( .a(n_22379), .o(n_22380) );
in01s01 g758032 ( .a(n_22377), .o(n_22378) );
no02f06 TIMEBOOST_cell_7655 ( .a(TIMEBOOST_net_2458), .b(n_13548), .o(n_13547) );
no02s01 g758036 ( .a(n_22846), .b(n_22845), .o(n_22847) );
na02s01 g758037 ( .a(n_22812), .b(n_22699), .o(n_22700) );
no02s01 g758038 ( .a(n_22844), .b(n_22843), .o(n_22923) );
no02s01 g758039 ( .a(n_22842), .b(n_22839), .o(n_22924) );
na02s01 g758040 ( .a(n_22878), .b(n_22876), .o(n_22953) );
no02s01 g758041 ( .a(n_22647), .b(n_22697), .o(n_22698) );
no02s01 g758042 ( .a(n_22729), .b(n_22690), .o(n_22763) );
na02s01 g758044 ( .a(n_22920), .b(n_22645), .o(n_22921) );
na02s01 g758045 ( .a(n_22840), .b(n_22656), .o(n_22841) );
in01s01 g758046 ( .a(n_23053), .o(n_23054) );
no02s01 g758047 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_28_), .o(n_23053) );
na02s02 g758048 ( .a(n_22732), .b(n_22456), .o(n_22733) );
in01s01 g758049 ( .a(n_23116), .o(n_22952) );
na02s01 g758050 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_28_), .o(n_23116) );
no02s01 g758051 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_23_), .o(n_22849) );
no02s01 g758052 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_25_), .o(n_23181) );
no02s01 g758053 ( .a(n_22653), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_11_), .o(n_22731) );
na02s03 g758054 ( .a(n_22783), .b(n_22620), .o(n_22784) );
no02s01 g758055 ( .a(n_23058), .b(n_22807), .o(n_23529) );
na02s01 g758056 ( .a(n_23052), .b(n_23051), .o(n_23642) );
no02s01 g758057 ( .a(n_22688), .b(n_22843), .o(n_23448) );
na02s01 g758058 ( .a(n_22920), .b(n_22951), .o(n_23342) );
no02s01 g758059 ( .a(n_22760), .b(n_22839), .o(n_23526) );
in01s01 g758060 ( .a(n_22880), .o(n_22881) );
no02s01 g758061 ( .a(n_22845), .b(n_22734), .o(n_22880) );
no02s01 g758062 ( .a(n_22918), .b(n_22917), .o(n_23382) );
na02s01 g758063 ( .a(n_22879), .b(n_22810), .o(n_23565) );
na02s01 g758064 ( .a(n_22646), .b(n_22699), .o(n_23319) );
na02s01 g758065 ( .a(n_22654), .b(n_22648), .o(n_23154) );
no02s01 g758066 ( .a(n_23295), .b(n_22730), .o(n_23296) );
in01s01 g758067 ( .a(n_22761), .o(n_22762) );
no02s01 g758068 ( .a(n_22729), .b(n_22644), .o(n_22761) );
no02s01 g758069 ( .a(n_22694), .b(n_22693), .o(n_22981) );
na02s01 g758070 ( .a(n_22650), .b(n_22728), .o(n_22786) );
na02f04 g758071 ( .a(n_22507), .b(FE_OCP_RBN5215_n_22150), .o(n_22508) );
no02m04 g758072 ( .a(n_22468), .b(FE_OCP_RBN5214_n_22150), .o(n_22469) );
in01s01 g758073 ( .a(n_22504), .o(n_22505) );
na02s06 g758074 ( .a(n_22466), .b(n_22465), .o(n_22504) );
na02f06 g758075 ( .a(n_22150), .b(FE_OCP_RBN3720_n_20621), .o(n_22200) );
na02s04 g758076 ( .a(FE_OCP_RBN6184_n_44267), .b(n_20717), .o(n_22267) );
na02s01 g758077 ( .a(FE_OCP_RBN6185_n_44267), .b(n_21096), .o(n_22266) );
na02s02 g758078 ( .a(FE_OCP_RBN3210_n_21203), .b(n_44277), .o(n_22232) );
na02m04 g758079 ( .a(FE_OCP_RBN5207_n_20504), .b(n_22005), .o(n_22085) );
in01f04 g758080 ( .a(n_22027), .o(n_22084) );
no02f10 g758085 ( .a(n_44160), .b(FE_OCP_RBN6878_n_44267), .o(n_22481) );
no02f02 TIMEBOOST_cell_7656 ( .a(n_13535), .b(n_13489), .o(TIMEBOOST_net_2459) );
na02s01 g758087 ( .a(n_44275), .b(FE_OCP_RBN1162_n_20763), .o(n_22311) );
no02s02 g758088 ( .a(FE_OCP_RBN6184_n_44267), .b(FE_OCP_RBN1161_n_20763), .o(n_22345) );
in01s01 g758089 ( .a(n_22263), .o(n_22264) );
na02s02 g758090 ( .a(n_22043), .b(FE_OCP_RBN4467_n_44267), .o(n_22263) );
in01s01 g758091 ( .a(n_22079), .o(n_22164) );
in01s01 g758095 ( .a(n_22048), .o(n_22079) );
no02s02 g758096 ( .a(n_21973), .b(FE_OCPN6929_FE_OCP_RBN1152_n_20910), .o(n_22048) );
in01s01 g758101 ( .a(n_22047), .o(n_22078) );
na02s06 g758102 ( .a(FE_OCPN6929_FE_OCP_RBN1152_n_20910), .b(FE_OCP_RBN7056_FE_OCPN1068_n_21973), .o(n_22047) );
in01s01 g758103 ( .a(n_22261), .o(n_22262) );
na02s02 g758104 ( .a(FE_OCP_RBN4466_n_44267), .b(FE_OCP_RBN7049_n_20941), .o(n_22261) );
in01s01 g758105 ( .a(n_22300), .o(n_22301) );
na02s02 g758106 ( .a(FE_OCP_RBN7052_n_20941), .b(n_21973), .o(n_22022) );
na02s01 g758107 ( .a(FE_OCP_RBN6185_n_44267), .b(FE_OCP_RBN7051_n_20941), .o(n_22300) );
in01s02 g758110 ( .a(n_22131), .o(n_22130) );
in01s02 g758111 ( .a(n_22099), .o(n_22131) );
no02s03 g758112 ( .a(n_44277), .b(FE_OCP_RBN2115_n_20935), .o(n_22099) );
no02s01 TIMEBOOST_cell_8462 ( .a(n_32413), .b(n_32502), .o(TIMEBOOST_net_2718) );
in01s01 g758116 ( .a(n_22129), .o(n_22128) );
in01s01 g758117 ( .a(n_22098), .o(n_22129) );
no02s02 g758118 ( .a(n_44277), .b(FE_OCP_RBN6051_n_21118), .o(n_22098) );
na02m06 TIMEBOOST_cell_4974 ( .a(FE_RN_6_0), .b(FE_RN_7_0), .o(TIMEBOOST_net_1435) );
na02s06 g758120 ( .a(FE_OCPN1071_n_44267), .b(FE_OCP_RBN3222_n_21242), .o(n_22305) );
no02s01 g758121 ( .a(FE_OCP_RBN4468_n_44267), .b(n_21242), .o(n_22342) );
na02s01 g758122 ( .a(FE_OCP_RBN4462_n_44267), .b(n_21312), .o(n_22259) );
na02s01 TIMEBOOST_cell_1259 ( .a(n_33579), .b(n_33417), .o(TIMEBOOST_net_244) );
na02s01 g758126 ( .a(FE_OCP_RBN4462_n_44267), .b(n_21265), .o(n_22258) );
na02s02 g758127 ( .a(FE_OCP_RBN5216_n_22212), .b(FE_OCP_RBN5388_n_22149), .o(n_22299) );
no02s01 g758128 ( .a(n_22212), .b(FE_OCP_RBN5387_n_22149), .o(n_22335) );
in01s01 g758129 ( .a(n_23152), .o(n_23153) );
ao12s01 g758130 ( .a(n_22844), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_17_), .o(n_23152) );
in01s02 g758132 ( .a(n_22502), .o(n_22503) );
no02m06 g758133 ( .a(n_22411), .b(n_22554), .o(n_22502) );
ao12s01 g758134 ( .a(n_22692), .b(FE_OCP_RBN2266_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_11_), .o(n_23356) );
na02m06 g758135 ( .a(n_22154), .b(n_22064), .o(n_22155) );
in01s01 g758136 ( .a(n_23201), .o(n_23202) );
ao12s01 g758137 ( .a(n_22877), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_15_), .o(n_23201) );
na02s02 g758138 ( .a(FE_OCPN4832_n_22294), .b(n_22417), .o(n_22419) );
no02s01 g758139 ( .a(n_22415), .b(n_22291), .o(n_22416) );
na02s02 g758140 ( .a(n_22294), .b(FE_OCP_DRV_N1434_n_21283), .o(n_22332) );
na02s01 g758141 ( .a(n_22463), .b(n_22330), .o(n_22464) );
no02s01 g758142 ( .a(n_22461), .b(n_22370), .o(n_22462) );
in01s01 g758144 ( .a(n_22413), .o(n_22439) );
na02s02 g758145 ( .a(n_22330), .b(n_22293), .o(n_22413) );
in01s01 g758147 ( .a(n_22046), .o(n_22344) );
na02s04 g758148 ( .a(n_21973), .b(FE_OCP_RBN1161_n_20763), .o(n_22046) );
in01s02 g758149 ( .a(n_22295), .o(n_22296) );
na02m02 g758150 ( .a(FE_OCP_RBN5049_FE_RN_606_0), .b(n_22154), .o(n_22295) );
in01s01 g758152 ( .a(n_23150), .o(n_23151) );
ao12s01 g758153 ( .a(n_22842), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_21_), .o(n_23150) );
in01s01 g758154 ( .a(n_23148), .o(n_23149) );
ao12s01 g758155 ( .a(n_22846), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_19_), .o(n_23148) );
in01s01 g758156 ( .a(n_22726), .o(n_22727) );
ao12s01 g758157 ( .a(n_22690), .b(FE_OCP_RBN2264_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_9_), .o(n_22726) );
ao12s01 g758158 ( .a(n_22697), .b(FE_OCP_RBN3879_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_5_), .o(n_23091) );
no02s02 TIMEBOOST_cell_5590 ( .a(n_25650), .b(n_25651), .o(TIMEBOOST_net_1743) );
in01s02 g758162 ( .a(n_22221), .o(n_22220) );
no02s02 TIMEBOOST_cell_1263 ( .a(n_33416), .b(FE_OCP_RBN2532_n_33372), .o(TIMEBOOST_net_246) );
no02s06 g758164 ( .a(FE_OCP_RBN4462_n_44267), .b(FE_OCP_RBN3222_n_21242), .o(n_22221) );
no03f08 TIMEBOOST_cell_8436 ( .a(n_35553), .b(n_35533), .c(n_35575), .o(n_35576) );
in01s01 g758166 ( .a(n_22083), .o(n_22045) );
na02s02 g758167 ( .a(n_21973), .b(n_20882), .o(n_22083) );
na02s06 g758168 ( .a(FE_OCPN1071_n_44267), .b(FE_OCP_RBN2114_n_20935), .o(n_22271) );
no02s03 g758169 ( .a(FE_OCP_RBN2113_n_20935), .b(FE_OCP_RBN4466_n_44267), .o(n_22308) );
in01s01 g758173 ( .a(n_22153), .o(n_22196) );
na02s03 g758174 ( .a(n_44277), .b(FE_OCP_RBN6051_n_21118), .o(n_22153) );
na02s01 g758175 ( .a(FE_OCP_RBN4468_n_44267), .b(n_21264), .o(n_22216) );
in01s02 g758176 ( .a(n_22785), .o(n_22660) );
oa12m03 g758177 ( .a(n_21485), .b(n_21484), .c(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n_22785) );
na02s01 g758178 ( .a(n_22405), .b(n_22328), .o(n_22460) );
na02s04 TIMEBOOST_cell_8130 ( .a(FE_OCPN5114_n_22249), .b(FE_OCP_RBN3720_n_20621), .o(TIMEBOOST_net_2696) );
oa22s01 g758180 ( .a(FE_OCP_RBN3362_n_21951), .b(n_21916), .c(n_21990), .d(n_21917), .o(n_22044) );
in01s01 g758181 ( .a(n_22020), .o(n_22021) );
oa12s01 g758182 ( .a(FE_OCP_RBN3351_n_21812), .b(FE_OCP_RBN3362_n_21951), .c(n_21845), .o(n_22020) );
na02s03 g758184 ( .a(n_44277), .b(n_21076), .o(n_22231) );
in01s01 g758186 ( .a(n_22194), .o(n_22214) );
na02s02 g758188 ( .a(n_22404), .b(n_22253), .o(n_22459) );
no02s01 g758189 ( .a(n_22213), .b(n_22434), .o(n_22500) );
in01s01 g758190 ( .a(n_22498), .o(n_22499) );
na02s02 g758191 ( .a(n_22399), .b(n_22368), .o(n_22498) );
in01s01 g758192 ( .a(n_22457), .o(n_22458) );
no02f06 TIMEBOOST_cell_1254 ( .a(n_29192), .b(TIMEBOOST_net_241), .o(n_29233) );
in01s01 g758194 ( .a(n_22496), .o(n_22497) );
na03s20 TIMEBOOST_cell_4579 ( .a(n_16894), .b(n_16988), .c(n_16899), .o(n_17245) );
oa22s01 g758196 ( .a(n_22585), .b(n_21866), .c(n_22586), .d(n_21865), .o(n_22659) );
oa22s01 g758197 ( .a(n_22604), .b(n_21867), .c(FE_OCP_RBN3408_n_22604), .d(n_21868), .o(n_22689) );
na02s02 g758199 ( .a(n_21973), .b(n_20724), .o(n_22041) );
oa22s01 g758200 ( .a(n_21453), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .c(FE_OCP_RBN3881_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .d(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_), .o(n_22737) );
ao22s01 g758201 ( .a(FE_OCP_RBN3879_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_3_), .c(n_22658), .d(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n_22813) );
oa22s01 g758202 ( .a(n_22657), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .c(FE_OCP_RBN2258_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .d(delay_sub_ln23_0_unr16_stage6_stallmux_q_7_), .o(n_23157) );
in01s02 g758203 ( .a(n_22494), .o(n_22495) );
no02s01 TIMEBOOST_cell_8544 ( .a(n_38778), .b(FE_OFN5092_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(TIMEBOOST_net_2759) );
in01s02 g758205 ( .a(n_22492), .o(n_22493) );
no03s20 TIMEBOOST_cell_4581 ( .a(n_17197), .b(FE_RN_2175_0), .c(FE_OCP_RBN7102_n_44365), .o(n_17239) );
in01s02 g758207 ( .a(n_22490), .o(n_22491) );
na02s06 g758208 ( .a(n_22407), .b(n_22375), .o(n_22490) );
in01s01 g758211 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_25_), .o(n_22656) );
no02s02 g758214 ( .a(FE_OCP_RBN2266_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_12_), .o(n_23295) );
in01s01 g758215 ( .a(n_22877), .o(n_22878) );
no02s01 g758216 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_15_), .o(n_22877) );
in01s01 g758217 ( .a(n_22850), .o(n_22810) );
no02s01 g758218 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_22_), .o(n_22850) );
in01s01 g758219 ( .a(n_23006), .o(n_23051) );
no02s01 g758220 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_26_), .o(n_23006) );
in01s01 g758221 ( .a(n_22839), .o(n_22809) );
no02s01 g758222 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_20_), .o(n_22839) );
no02s01 g758223 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_18_), .o(n_22845) );
in01s01 g758224 ( .a(n_22732), .o(n_22688) );
na02s01 g758225 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_16_), .o(n_22732) );
in01s01 g758226 ( .a(n_22654), .o(n_22655) );
na02s01 g758227 ( .a(FE_OCP_RBN2259_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_6_), .o(n_22654) );
in01s01 g758228 ( .a(n_22699), .o(n_22653) );
na02s02 g758229 ( .a(FE_OCP_RBN2268_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_10_), .o(n_22699) );
no02s01 g758230 ( .a(FE_OCP_RBN2265_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_8_), .o(n_22729) );
in01s01 g758231 ( .a(n_22808), .o(n_22917) );
na02s01 g758232 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_14_), .o(n_22808) );
no02s01 g758233 ( .a(FE_OCP_RBN3879_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_5_), .o(n_22697) );
na02s01 g758234 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_13_), .o(n_22920) );
no02s01 g758235 ( .a(n_22608), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n_22693) );
in01s01 g758236 ( .a(n_23052), .o(n_22950) );
na02s01 g758237 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_26_), .o(n_23052) );
in01s01 g758238 ( .a(n_22840), .o(n_22807) );
na02s01 g758239 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_24_), .o(n_22840) );
in01s01 g758240 ( .a(n_22783), .o(n_22760) );
na02s01 g758241 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_20_), .o(n_22783) );
in01s01 g758242 ( .a(n_22734), .o(n_22652) );
no02s06 g758243 ( .a(n_22455), .b(FE_OFN745_n_22641), .o(n_22734) );
no02s01 g758244 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_19_), .o(n_22846) );
no02s01 g758245 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_17_), .o(n_22844) );
no02s01 g758246 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_16_), .o(n_22843) );
no02s01 g758247 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_21_), .o(n_22842) );
no02s01 g758248 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_24_), .o(n_23058) );
in01s01 g758249 ( .a(n_22918), .o(n_22876) );
no02s01 g758250 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_14_), .o(n_22918) );
na02s06 g758252 ( .a(FE_OCP_RBN5467_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_2_), .o(n_22650) );
in01m01 g758253 ( .a(n_22649), .o(n_22728) );
no02s03 g758254 ( .a(FE_OCP_RBN5466_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_2_), .o(n_22649) );
in01s01 g758255 ( .a(n_22647), .o(n_22648) );
no02s01 g758256 ( .a(FE_OCP_RBN2260_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_6_), .o(n_22647) );
in01s01 g758257 ( .a(n_22621), .o(n_22694) );
na02s01 g758258 ( .a(n_22608), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n_22621) );
no02s01 g758259 ( .a(FE_OCP_RBN2263_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_9_), .o(n_22690) );
in01s01 g758260 ( .a(n_22695), .o(n_22646) );
no02s01 g758261 ( .a(FE_OCP_RBN2267_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_10_), .o(n_22695) );
no02s01 g758262 ( .a(FE_OCP_RBN2266_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_11_), .o(n_22692) );
in01s01 g758263 ( .a(n_22645), .o(n_22730) );
na02s01 g758264 ( .a(FE_OCP_RBN2266_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_12_), .o(n_22645) );
na02s02 g758265 ( .a(FE_OFN745_n_22641), .b(n_22208), .o(n_22951) );
in01s01 g758266 ( .a(n_22643), .o(n_22644) );
na02s01 g758267 ( .a(FE_OCP_RBN3881_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_8_), .o(n_22643) );
in01s01 g758268 ( .a(n_22879), .o(n_22759) );
na02s03 g758269 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_22_), .o(n_22879) );
no03s20 TIMEBOOST_cell_4578 ( .a(n_11918), .b(FE_RN_2813_0), .c(FE_OCP_RBN6310_n_45224), .o(n_11770) );
na02s02 g758271 ( .a(FE_OCPN5113_n_22249), .b(FE_OCP_RBN6383_n_21087), .o(n_22375) );
in01s02 g758273 ( .a(n_22411), .o(n_22436) );
no02s08 g758274 ( .a(n_20867), .b(FE_OCPN5114_n_22249), .o(n_22411) );
no02f04 g758281 ( .a(n_21951), .b(n_21812), .o(n_21974) );
in01f02 g758282 ( .a(n_22018), .o(n_22019) );
no02f04 g758283 ( .a(n_22003), .b(n_22002), .o(n_22018) );
na02f06 g758286 ( .a(FE_OCP_RBN5341_n_22068), .b(n_20555), .o(n_22150) );
na02s01 g758287 ( .a(n_22249), .b(n_20862), .o(n_22374) );
in01s01 g758289 ( .a(n_22213), .o(n_22253) );
no02f08 TIMEBOOST_cell_7759 ( .a(n_19637), .b(TIMEBOOST_net_2510), .o(n_19700) );
na03m04 TIMEBOOST_cell_4580 ( .a(FE_RN_82_0), .b(delay_xor_ln21_unr15_stage6_stallmux_q_0_), .c(FE_OCP_RBN6464_n_44061), .o(FE_RN_83_0) );
na02m06 TIMEBOOST_cell_8810 ( .a(n_10879), .b(n_44511), .o(TIMEBOOST_net_2892) );
na02m08 g758294 ( .a(FE_OCPN5114_n_22249), .b(n_20614), .o(n_22507) );
no02m06 g758295 ( .a(n_22288), .b(FE_OCPN1388_n_20555), .o(n_22468) );
na02s01 g758296 ( .a(n_22288), .b(FE_OCP_RBN6384_n_21087), .o(n_22407) );
in01s02 g758297 ( .a(n_22465), .o(n_22406) );
na02s06 g758298 ( .a(n_21011), .b(FE_OCPN5113_n_22249), .o(n_22465) );
na02s01 g758299 ( .a(n_22288), .b(n_21324), .o(n_22405) );
no04m20 TIMEBOOST_cell_7332 ( .a(FE_RN_1034_0), .b(FE_OCP_RBN6463_n_44061), .c(delay_xor_ln22_unr15_stage6_stallmux_q_3_), .d(FE_OCP_RBN6467_n_44061), .o(n_22930) );
in01s01 g758302 ( .a(n_22294), .o(n_22415) );
na02s02 g758303 ( .a(n_22121), .b(FE_OCP_RBN1865_n_21163), .o(n_22294) );
na02s01 g758304 ( .a(n_22288), .b(n_20978), .o(n_22404) );
no02s01 g758305 ( .a(FE_OCPN5114_n_22249), .b(FE_OCPN7089_n_20979), .o(n_22434) );
no02s02 g758306 ( .a(n_22288), .b(FE_OCP_RBN3260_n_21360), .o(n_22438) );
na02s01 g758307 ( .a(n_22288), .b(FE_OCP_RBN6062_n_21194), .o(n_22463) );
no02s01 g758308 ( .a(FE_OCPN5113_n_22249), .b(n_21278), .o(n_22461) );
in01s01 g758312 ( .a(n_22330), .o(n_22370) );
na02m02 g758316 ( .a(FE_OCP_RBN5341_n_22068), .b(n_22126), .o(n_22149) );
na02s01 g758317 ( .a(n_22288), .b(n_21282), .o(n_22399) );
na02s01 g758318 ( .a(FE_OCPN5113_n_22249), .b(n_21281), .o(n_22368) );
na02s01 g758319 ( .a(n_22249), .b(n_21427), .o(n_22293) );
na02s01 g758320 ( .a(FE_OCPN5113_n_22249), .b(n_21427), .o(n_22367) );
no02f04 TIMEBOOST_cell_1253 ( .a(n_29091), .b(n_29379), .o(TIMEBOOST_net_241) );
na02m04 g758322 ( .a(n_22066), .b(FE_OCP_RBN4645_n_20420), .o(n_22154) );
oa12s01 g758323 ( .a(FE_OCP_RBN3879_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_4_), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_5_), .o(n_23087) );
oa12s01 g758324 ( .a(FE_OCP_RBN2262_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_8_), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_9_), .o(n_22812) );
in01s01 g758329 ( .a(n_22292), .o(n_22328) );
no02s02 g758330 ( .a(n_22187), .b(n_21324), .o(n_22292) );
in01s02 g758332 ( .a(FE_OCPN1248_n_22291), .o(n_22417) );
no02s02 g758333 ( .a(n_22187), .b(FE_OCP_RBN1865_n_21163), .o(n_22291) );
in01s01 g758334 ( .a(n_22466), .o(n_22432) );
na02s06 g758335 ( .a(n_22288), .b(n_21080), .o(n_22466) );
in01s02 g758337 ( .a(n_22326), .o(n_22327) );
no02s06 g758338 ( .a(n_22249), .b(FE_OCPN1386_n_21199), .o(n_22326) );
na02s06 g758370 ( .a(n_22187), .b(n_20868), .o(n_22351) );
no02s02 g758371 ( .a(n_22187), .b(FE_OCPN1214_n_21166), .o(n_22383) );
in01s04 g758372 ( .a(n_22185), .o(n_22186) );
na02f08 g758373 ( .a(FE_OCP_RBN5343_n_22068), .b(n_20691), .o(n_22185) );
oa22s01 g758374 ( .a(n_21966), .b(n_21894), .c(n_21965), .d(n_21893), .o(n_22016) );
no02s01 g758375 ( .a(n_22249), .b(n_21431), .o(n_22667) );
in01s01 g758376 ( .a(n_22014), .o(n_22015) );
in01s01 g758377 ( .a(n_21999), .o(n_22014) );
oa12f08 g758378 ( .a(n_21871), .b(n_21950), .c(n_21807), .o(n_21999) );
oa22s01 g758379 ( .a(n_22528), .b(n_21864), .c(n_22527), .d(n_21863), .o(n_22588) );
in01s01 g758380 ( .a(FE_OFN745_n_22641), .o(n_22782) );
in01s01 g758385 ( .a(n_23398), .o(n_23414) );
in01s02 g758391 ( .a(n_23509), .o(n_23486) );
in01s02 g758396 ( .a(FE_OCP_DRV_N6899_FE_OCPN5276_n_23590), .o(n_23564) );
in01s01 g758399 ( .a(n_23486), .o(n_23590) );
in01s02 g758401 ( .a(n_23447), .o(n_23509) );
in01s01 g758405 ( .a(FE_RN_1116_0), .o(n_26663) );
in01s03 g758411 ( .a(n_23398), .o(n_23447) );
in01s06 g758419 ( .a(FE_OFN747_n_22641), .o(n_23398) );
in01s06 g758429 ( .a(n_23259), .o(n_23317) );
in01s06 g758440 ( .a(n_23353), .o(n_23466) );
in01s06 g758441 ( .a(n_23339), .o(n_23353) );
in01s01 g758442 ( .a(n_23317), .o(n_23339) );
in01s06 g758452 ( .a(FE_OFN748_n_22641), .o(n_23259) );
in01s01 g758467 ( .a(FE_OFN748_n_22641), .o(n_23254) );
in01s01 g758469 ( .a(n_25824), .o(n_25831) );
in01s02 g758470 ( .a(FE_OFN748_n_22641), .o(n_25824) );
in01s01 g758471 ( .a(n_23271), .o(n_26054) );
in01s01 g758474 ( .a(n_25829), .o(n_23271) );
in01s02 g758475 ( .a(FE_OFN748_n_22641), .o(n_25829) );
in01s01 g758486 ( .a(FE_OFN745_n_22641), .o(n_23115) );
in01s04 g758495 ( .a(FE_OFN745_n_22641), .o(n_22725) );
in01s01 g758507 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_11_), .o(n_23376) );
in01s01 g758509 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_21_), .o(n_22620) );
na02f08 g758514 ( .a(n_21940), .b(n_21922), .o(n_21941) );
in01f02 g758515 ( .a(n_21971), .o(n_21972) );
na02f01 g758516 ( .a(n_21940), .b(n_21954), .o(n_21971) );
no02s06 g758517 ( .a(FE_OCP_RBN5211_n_20412), .b(n_21953), .o(n_22003) );
in01f02 g758519 ( .a(n_21970), .o(n_22002) );
na02f06 g758520 ( .a(FE_OCP_RBN5211_n_20412), .b(n_21953), .o(n_21970) );
in01m02 g758521 ( .a(n_22183), .o(n_22184) );
no02m04 g758522 ( .a(n_22145), .b(n_22063), .o(n_22183) );
oa22s01 g758523 ( .a(n_21919), .b(n_21813), .c(n_21918), .d(n_21814), .o(n_21969) );
in01s01 g758525 ( .a(FE_OCP_RBN3362_n_21951), .o(n_21990) );
ao12f04 g758527 ( .a(n_21738), .b(n_21900), .c(n_21792), .o(n_21951) );
in01s06 g758529 ( .a(FE_OCP_RBN5343_n_22068), .o(n_22121) );
in01m10 g758550 ( .a(n_22249), .o(n_22288) );
in01m10 g758551 ( .a(n_22187), .o(n_22249) );
in01m10 g758552 ( .a(FE_OCP_RBN5342_n_22068), .o(n_22187) );
oa22s01 g758560 ( .a(n_22488), .b(n_21827), .c(n_22487), .d(n_21828), .o(n_22568) );
oa22s01 g758561 ( .a(n_22523), .b(n_21853), .c(n_22524), .d(n_21854), .o(n_22587) );
oa22s01 g758562 ( .a(n_22526), .b(n_21859), .c(n_22525), .d(n_21860), .o(n_22606) );
in01s01 g758563 ( .a(n_22585), .o(n_22586) );
oa12s01 g758564 ( .a(n_21824), .b(n_22526), .c(n_21751), .o(n_22585) );
oa12s01 g758566 ( .a(n_21799), .b(n_22525), .c(n_21753), .o(n_22604) );
in01s01 g758569 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_10_), .o(n_23403) );
in01s01 g758573 ( .a(n_21938), .o(n_21939) );
na02s01 g758574 ( .a(n_21905), .b(n_21925), .o(n_21938) );
in01s01 g758575 ( .a(n_21997), .o(n_21998) );
na02s01 g758576 ( .a(n_21936), .b(n_21922), .o(n_21997) );
na02f04 g758577 ( .a(n_21815), .b(n_21905), .o(n_21906) );
na02m04 g758578 ( .a(n_21874), .b(FE_OCP_RBN7043_n_20336), .o(n_21940) );
na02f06 g758579 ( .a(n_21875), .b(FE_OCP_RBN1157_n_20336), .o(n_21954) );
in01s01 g758580 ( .a(n_22094), .o(n_22095) );
na02s02 g758581 ( .a(n_22034), .b(n_22065), .o(n_22094) );
in01m02 g758583 ( .a(n_22064), .o(n_22145) );
na02m06 g758584 ( .a(n_22037), .b(FE_OCP_RBN2094_n_47175), .o(n_22064) );
no02s06 g758588 ( .a(n_22037), .b(FE_OCP_RBN2094_n_47175), .o(n_22063) );
na02f08 g758589 ( .a(n_22034), .b(n_21961), .o(n_22035) );
in01m04 g758590 ( .a(n_21903), .o(n_21904) );
ao12m08 g758591 ( .a(n_21663), .b(n_21849), .c(n_21664), .o(n_21903) );
in01m02 g758592 ( .a(n_21923), .o(n_21924) );
in01s01 g758595 ( .a(n_22549), .o(n_22550) );
oa12f02 g758596 ( .a(n_21883), .b(n_22489), .c(n_21832), .o(n_22549) );
oa22s01 g758597 ( .a(n_21914), .b(n_21869), .c(n_21913), .d(n_21870), .o(n_21967) );
in01s01 g758598 ( .a(n_21965), .o(n_21966) );
in01s01 g758599 ( .a(n_21950), .o(n_21965) );
oa12f08 g758600 ( .a(n_21842), .b(n_21898), .c(n_21783), .o(n_21950) );
oa22s01 g758601 ( .a(n_22485), .b(n_21855), .c(n_22486), .d(n_21856), .o(n_22567) );
oa22s01 g758602 ( .a(n_22431), .b(n_21777), .c(n_22453), .d(n_21776), .o(n_22548) );
in01s01 g758603 ( .a(n_22527), .o(n_22528) );
oa12s01 g758604 ( .a(n_21692), .b(n_22431), .c(n_21748), .o(n_22527) );
na02f02 g758609 ( .a(n_21816), .b(n_20205), .o(n_21905) );
na02s06 g758610 ( .a(n_21817), .b(n_20206), .o(n_21925) );
in01s01 g758612 ( .a(n_21922), .o(n_21937) );
na02f06 g758613 ( .a(FE_OCP_RBN2098_n_20325), .b(n_21902), .o(n_21922) );
in01s01 g758616 ( .a(n_21921), .o(n_21936) );
no02f06 g758617 ( .a(FE_OCP_RBN2098_n_20325), .b(n_21902), .o(n_21921) );
in01s01 g758620 ( .a(n_22526), .o(n_22525) );
na02s01 g758621 ( .a(n_22489), .b(n_21796), .o(n_22526) );
na02f04 g758622 ( .a(n_21983), .b(n_20273), .o(n_22034) );
na02m08 g758623 ( .a(n_21984), .b(FE_OCP_RBN1838_n_20273), .o(n_22065) );
oa12m06 g758625 ( .a(n_21646), .b(n_21964), .c(n_21647), .o(n_21987) );
oa12m04 g758627 ( .a(n_21700), .b(n_21964), .c(n_21634), .o(n_21985) );
oa22s01 g758628 ( .a(n_21767), .b(n_21843), .c(n_21766), .d(n_21844), .o(n_21920) );
in01s01 g758629 ( .a(n_21918), .o(n_21919) );
in01s01 g758630 ( .a(n_21900), .o(n_21918) );
oa12f06 g758631 ( .a(n_21680), .b(n_21811), .c(n_21741), .o(n_21900) );
in01m02 g758632 ( .a(n_21874), .o(n_21875) );
in01s01 g758635 ( .a(n_22487), .o(n_22488) );
oa12s01 g758636 ( .a(n_21670), .b(n_22396), .c(n_21600), .o(n_22487) );
oa22s01 g758637 ( .a(n_22397), .b(n_21861), .c(n_22430), .d(n_21862), .o(n_22545) );
in01s01 g758638 ( .a(n_22523), .o(n_22524) );
oa12s01 g758639 ( .a(n_21825), .b(n_22430), .c(n_21772), .o(n_22523) );
oa22s01 g758640 ( .a(n_22396), .b(n_21695), .c(n_22428), .d(n_21696), .o(n_22522) );
in01s01 g758641 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_17_), .o(n_22456) );
in01s06 g758643 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_18_), .o(n_22455) );
in01f02 g758647 ( .a(n_21849), .o(n_21847) );
in01s01 g758649 ( .a(n_21916), .o(n_21917) );
na02s01 g758650 ( .a(n_21815), .b(FE_OCP_RBN3351_n_21812), .o(n_21916) );
in01s01 g758651 ( .a(n_22032), .o(n_22033) );
na02s01 g758652 ( .a(n_21961), .b(n_22012), .o(n_22032) );
in01s02 g758653 ( .a(n_21816), .o(n_21817) );
na02s01 TIMEBOOST_cell_1110 ( .a(TIMEBOOST_net_169), .b(n_37376), .o(n_37459) );
oa22s01 g758656 ( .a(n_21833), .b(n_21838), .c(n_21834), .d(n_21839), .o(n_21915) );
in01s01 g758657 ( .a(n_21913), .o(n_21914) );
in01s01 g758658 ( .a(n_21898), .o(n_21913) );
oa12f08 g758659 ( .a(n_21803), .b(n_21818), .c(n_21761), .o(n_21898) );
in01m02 g758660 ( .a(n_21983), .o(n_21984) );
oa22s01 g758662 ( .a(n_22286), .b(n_21821), .c(n_22287), .d(n_21822), .o(n_22398) );
oa22s01 g758663 ( .a(n_22426), .b(n_21627), .c(n_22395), .d(n_21628), .o(n_22521) );
in01s01 g758664 ( .a(n_22485), .o(n_22486) );
oa12s01 g758665 ( .a(n_21622), .b(n_22395), .c(n_21561), .o(n_22485) );
in01s01 g758667 ( .a(n_22431), .o(n_22453) );
oa12s01 g758668 ( .a(n_21782), .b(n_22363), .c(n_21779), .o(n_22431) );
na02f04 g758669 ( .a(n_21780), .b(n_22397), .o(n_22489) );
in01s01 g758670 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_9_), .o(n_21912) );
na02s01 TIMEBOOST_cell_1109 ( .a(n_37215), .b(n_36974), .o(TIMEBOOST_net_169) );
no02m04 g758673 ( .a(n_21743), .b(n_21553), .o(n_21793) );
in01s01 g758675 ( .a(n_21815), .o(n_21845) );
na02f02 g758676 ( .a(n_21791), .b(FE_OCPN5244_n_21790), .o(n_21815) );
in01s01 g758677 ( .a(n_21813), .o(n_21814) );
na02s01 g758678 ( .a(n_21792), .b(n_21687), .o(n_21813) );
no02m02 g758680 ( .a(n_21791), .b(FE_OCPN5292_n_21790), .o(n_21812) );
in01s01 g758681 ( .a(n_21962), .o(n_21963) );
na02s01 g758682 ( .a(n_21911), .b(n_21947), .o(n_21962) );
in01s01 g758684 ( .a(n_21961), .o(n_21982) );
na02f08 g758685 ( .a(FE_OCPN1216_n_21946), .b(FE_OCPN4931_n_20275), .o(n_21961) );
in01s01 g758687 ( .a(n_21960), .o(n_22012) );
no02f08 g758688 ( .a(FE_OCPN1216_n_21946), .b(FE_OCPN4931_n_20275), .o(n_21960) );
in01m02 g758689 ( .a(n_21944), .o(n_21945) );
in01m02 g758690 ( .a(n_21964), .o(n_21944) );
na02m08 g758691 ( .a(n_21644), .b(n_21873), .o(n_21964) );
in01s01 g758694 ( .a(n_22397), .o(n_22430) );
na02f06 g758695 ( .a(n_22363), .b(n_21725), .o(n_22397) );
oa12m02 g758696 ( .a(n_21501), .b(n_21713), .c(n_21711), .o(n_21745) );
no02s01 TIMEBOOST_cell_1098 ( .a(n_33003), .b(TIMEBOOST_net_163), .o(n_33125) );
in01s01 g758698 ( .a(n_21843), .o(n_21844) );
in01s01 g758699 ( .a(n_21811), .o(n_21843) );
oa22s01 g758702 ( .a(n_21683), .b(n_21734), .c(n_21682), .d(n_21735), .o(n_21810) );
oa22s01 g758703 ( .a(n_22242), .b(n_21857), .c(n_22243), .d(n_21858), .o(n_22362) );
oa22s01 g758704 ( .a(n_22247), .b(n_21716), .c(n_22248), .d(n_21715), .o(n_22361) );
in01s01 g758706 ( .a(n_22396), .o(n_22428) );
oa12s01 g758707 ( .a(n_21698), .b(n_22284), .c(n_21722), .o(n_22396) );
in01m02 g758711 ( .a(n_21742), .o(n_21743) );
no02m06 g758712 ( .a(n_21713), .b(n_21621), .o(n_21742) );
no02s01 TIMEBOOST_cell_6340 ( .a(TIMEBOOST_net_2021), .b(n_40154), .o(TIMEBOOST_net_984) );
in01s01 g758716 ( .a(n_21766), .o(n_21767) );
no02s01 g758717 ( .a(n_21741), .b(n_21620), .o(n_21766) );
in01s04 g758720 ( .a(n_21687), .o(n_21738) );
na02m04 g758721 ( .a(n_21656), .b(FE_OCP_DRV_N1494_n_20059), .o(n_21687) );
in01s01 g758723 ( .a(n_21910), .o(n_21911) );
no02s06 g758724 ( .a(n_21897), .b(FE_OCPN1384_n_21896), .o(n_21910) );
na02m06 g758725 ( .a(n_21897), .b(FE_OCPN1384_n_21896), .o(n_21947) );
in01s01 g758727 ( .a(n_22395), .o(n_22426) );
no02s01 g758728 ( .a(n_22285), .b(n_21629), .o(n_22395) );
oa12m02 g758729 ( .a(FE_OCP_RBN6385_n_21429), .b(n_21558), .c(n_21661), .o(n_21686) );
no02f02 g758730 ( .a(n_21662), .b(FE_OCP_RBN6386_n_21429), .o(n_21710) );
oa12m04 g758731 ( .a(n_21489), .b(FE_OCP_RBN6129_n_21804), .c(n_21490), .o(n_21895) );
no02s01 TIMEBOOST_cell_8066 ( .a(n_6244), .b(n_6223), .o(TIMEBOOST_net_2664) );
na02s01 TIMEBOOST_cell_1210 ( .a(TIMEBOOST_net_219), .b(n_38019), .o(n_38076) );
in01s01 g758735 ( .a(n_21833), .o(n_21834) );
in01s01 g758736 ( .a(n_21818), .o(n_21833) );
oa22s01 g758738 ( .a(n_21794), .b(n_21759), .c(n_21733), .d(n_21760), .o(n_21851) );
oa22m02 g758739 ( .a(FE_OCP_RBN6129_n_21804), .b(FE_OCP_RBN6123_n_21630), .c(n_21804), .d(n_21630), .o(n_21946) );
in01s01 g758740 ( .a(n_22286), .o(n_22287) );
oa12s01 g758741 ( .a(n_21451), .b(n_22210), .c(n_21697), .o(n_22286) );
na02f06 g758742 ( .a(n_22246), .b(n_21723), .o(n_22363) );
in01s01 g758743 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_8_), .o(n_23267) );
in01s02 g758746 ( .a(n_21665), .o(n_21711) );
no02f08 g758747 ( .a(n_21621), .b(n_21508), .o(n_21665) );
no02m04 g758748 ( .a(n_21615), .b(n_21505), .o(n_21664) );
na02s06 g758749 ( .a(n_21616), .b(n_21506), .o(n_21663) );
no02f02 g758750 ( .a(n_21558), .b(n_21661), .o(n_21662) );
na02f02 g758751 ( .a(n_21684), .b(n_21654), .o(n_21685) );
no02s02 g758752 ( .a(n_21618), .b(n_21617), .o(n_21709) );
na02m04 g758754 ( .a(FE_OCP_RBN3328_n_21616), .b(n_21708), .o(n_21736) );
na02f08 TIMEBOOST_cell_1217 ( .a(FE_RN_2380_0), .b(n_23517), .o(TIMEBOOST_net_223) );
na02s01 TIMEBOOST_cell_1209 ( .a(n_37878), .b(n_38021), .o(TIMEBOOST_net_219) );
in01s01 g758757 ( .a(n_21682), .o(n_21683) );
no02s01 g758758 ( .a(n_21660), .b(n_21659), .o(n_21682) );
in01f02 g758760 ( .a(n_21620), .o(n_21680) );
no02m02 g758761 ( .a(n_21581), .b(n_20018), .o(n_21620) );
in01s01 g758763 ( .a(n_21893), .o(n_21894) );
na02s01 g758764 ( .a(n_21871), .b(n_21808), .o(n_21893) );
in01s01 g758765 ( .a(n_22247), .o(n_22248) );
na02s01 g758766 ( .a(n_22210), .b(n_21566), .o(n_22247) );
in01m04 g758767 ( .a(n_21658), .o(n_21713) );
in01s01 g758769 ( .a(n_22284), .o(n_22285) );
in01s01 g758770 ( .a(n_22246), .o(n_22284) );
no02f06 g758771 ( .a(n_22210), .b(n_21669), .o(n_22246) );
in01s01 g758772 ( .a(n_21734), .o(n_21735) );
in01s01 g758773 ( .a(n_21707), .o(n_21734) );
ao12f06 g758774 ( .a(n_21473), .b(n_21679), .c(n_21544), .o(n_21707) );
oa22s01 g758777 ( .a(n_21580), .b(n_21612), .c(n_21579), .d(n_21679), .o(n_21706) );
no02m08 TIMEBOOST_cell_4552 ( .a(n_17147), .b(TIMEBOOST_net_1366), .o(n_17292) );
oa12s01 g758779 ( .a(n_22178), .b(n_22177), .c(n_22176), .o(n_22245) );
oa12s01 g758780 ( .a(n_22180), .b(n_22209), .c(n_22179), .o(n_22244) );
in01s01 g758781 ( .a(n_22242), .o(n_22243) );
oa12s01 g758782 ( .a(n_21379), .b(n_22209), .c(n_21795), .o(n_22242) );
in01s01 g758783 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_13_), .o(n_22208) );
na02f08 g758787 ( .a(n_21556), .b(n_21430), .o(n_21621) );
na02s02 g758788 ( .a(n_21556), .b(n_21554), .o(n_21588) );
no02s02 g758789 ( .a(n_21509), .b(n_21510), .o(n_21619) );
in01s01 g758790 ( .a(n_21684), .o(n_21618) );
na02m08 g758791 ( .a(n_21587), .b(FE_OCPN6925_n_45081), .o(n_21684) );
in01m01 g758793 ( .a(n_21617), .o(n_21654) );
no02m04 g758794 ( .a(n_21587), .b(FE_OCPN1638_n_45081), .o(n_21617) );
na02s04 g758798 ( .a(n_21586), .b(FE_OCPN1711_n_45073), .o(n_21616) );
in01m02 g758799 ( .a(n_21615), .o(n_21708) );
no02m02 g758800 ( .a(n_21586), .b(FE_OCPN1638_n_45081), .o(n_21615) );
na02s02 g758801 ( .a(n_21506), .b(n_21548), .o(n_21956) );
no02f04 g758803 ( .a(n_21503), .b(FE_OCPUNCON6887_n_19961), .o(n_21659) );
no02m06 g758804 ( .a(n_21504), .b(n_19962), .o(n_21660) );
na02s01 g758805 ( .a(n_22209), .b(n_22179), .o(n_22180) );
in01s01 g758806 ( .a(n_21869), .o(n_21870) );
na02s01 g758807 ( .a(n_21784), .b(n_21842), .o(n_21869) );
na02m06 g758808 ( .a(n_21789), .b(FE_OCPUNCON7071_n_21788), .o(n_21871) );
in01s01 g758809 ( .a(n_21807), .o(n_21808) );
no02m06 g758810 ( .a(n_21789), .b(FE_OCPUNCON7071_n_21788), .o(n_21807) );
na02s06 TIMEBOOST_cell_3351 ( .a(TIMEBOOST_net_966), .b(n_17140), .o(n_17282) );
na02s01 TIMEBOOST_cell_6356 ( .a(TIMEBOOST_net_2029), .b(n_17130), .o(n_17281) );
na02s01 g758813 ( .a(n_22177), .b(n_22176), .o(n_22178) );
na02f06 g758814 ( .a(n_22117), .b(n_21592), .o(n_22210) );
oa12f08 g758820 ( .a(n_21366), .b(n_21477), .c(n_21397), .o(n_21558) );
oa12s01 g758823 ( .a(n_21547), .b(n_21546), .c(n_21545), .o(n_21613) );
in01s01 g758824 ( .a(n_21794), .o(n_21733) );
oa22s01 g758826 ( .a(n_21648), .b(n_21632), .c(n_21705), .d(n_21633), .o(n_21732) );
in01m02 g758831 ( .a(n_21786), .o(n_21804) );
no02s01 TIMEBOOST_cell_1200 ( .a(n_41193), .b(TIMEBOOST_net_214), .o(n_41280) );
in01s01 g758835 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_7_), .o(n_21785) );
na02m06 g758838 ( .a(n_21477), .b(n_21331), .o(n_21511) );
in01s01 g758839 ( .a(n_21556), .o(n_21510) );
na02f06 g758840 ( .a(n_21476), .b(n_45026), .o(n_21556) );
in01s01 g758842 ( .a(n_21509), .o(n_21554) );
no02m06 g758843 ( .a(n_21476), .b(FE_OCPN1382_n_45026), .o(n_21509) );
in01s02 g758844 ( .a(n_21552), .o(n_21553) );
no02s02 g758845 ( .a(n_21508), .b(n_21507), .o(n_21552) );
na02s06 g758848 ( .a(n_21475), .b(FE_OCPN1638_n_45081), .o(n_21506) );
in01s02 g758850 ( .a(n_21505), .o(n_21548) );
no02m04 g758851 ( .a(n_21475), .b(FE_OCPN1638_n_45081), .o(n_21505) );
in01s02 g758852 ( .a(n_21730), .o(n_21731) );
no02s04 g758853 ( .a(n_21703), .b(n_21463), .o(n_21730) );
no02s01 TIMEBOOST_cell_1199 ( .a(n_41206), .b(n_40812), .o(TIMEBOOST_net_214) );
na02s01 g758855 ( .a(n_21546), .b(n_21545), .o(n_21547) );
in01s01 g758856 ( .a(n_21838), .o(n_21839) );
na02s01 g758857 ( .a(n_21803), .b(n_21762), .o(n_21838) );
in01s01 g758858 ( .a(n_21783), .o(n_21784) );
no02m06 g758859 ( .a(n_21764), .b(FE_OCP_DRV_N3538_n_21763), .o(n_21783) );
na02s06 g758860 ( .a(n_21764), .b(FE_OCP_DRV_N3538_n_21763), .o(n_21842) );
in01s01 g758861 ( .a(n_21579), .o(n_21580) );
na02s01 g758862 ( .a(n_21474), .b(n_21544), .o(n_21579) );
no02s10 TIMEBOOST_cell_8488 ( .a(FE_RN_27_0), .b(FE_RN_28_0), .o(TIMEBOOST_net_2731) );
in01s01 g758864 ( .a(n_21679), .o(n_21612) );
no02f08 g758865 ( .a(n_21500), .b(n_21432), .o(n_21679) );
in01m02 g758866 ( .a(n_21503), .o(n_21504) );
na03s10 TIMEBOOST_cell_7104 ( .a(FE_OCP_RBN6410_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(FE_RN_395_0), .c(n_1387), .o(n_1433) );
oa12s01 g758869 ( .a(n_21519), .b(n_22119), .c(n_21482), .o(n_22177) );
oa22s01 g758870 ( .a(n_22119), .b(n_21564), .c(n_22056), .d(n_21565), .o(n_22144) );
oa12s01 g758872 ( .a(n_22062), .b(n_22061), .c(n_22060), .o(n_22118) );
in01s01 g758873 ( .a(n_22117), .o(n_22209) );
ao12f04 g758874 ( .a(n_21518), .b(n_22030), .c(n_21483), .o(n_22117) );
na02m08 g758880 ( .a(n_21399), .b(n_21287), .o(n_21477) );
no02f04 g758881 ( .a(n_21330), .b(n_21365), .o(n_21366) );
na02s06 g758882 ( .a(n_21358), .b(n_45070), .o(n_21398) );
no02f04 TIMEBOOST_cell_8801 ( .a(TIMEBOOST_net_2887), .b(n_3640), .o(n_3828) );
no02m04 g758885 ( .a(n_21365), .b(n_21397), .o(n_21438) );
na02s02 g758886 ( .a(FE_OCP_RBN6385_n_21429), .b(n_21430), .o(n_21543) );
no02m02 g758887 ( .a(FE_OCP_RBN6386_n_21429), .b(n_21661), .o(n_21578) );
no02s06 g758888 ( .a(n_21361), .b(n_45072), .o(n_21508) );
in01s02 g758889 ( .a(n_21501), .o(n_21502) );
in01m02 g758890 ( .a(n_21507), .o(n_21501) );
no02f06 TIMEBOOST_cell_8485 ( .a(TIMEBOOST_net_2729), .b(FE_RN_2464_0), .o(FE_RN_2467_0) );
no02m08 g758893 ( .a(n_21609), .b(n_21462), .o(n_21703) );
na02s04 TIMEBOOST_cell_3263 ( .a(TIMEBOOST_net_922), .b(n_11123), .o(n_11169) );
no02f06 g758895 ( .a(n_21428), .b(n_21433), .o(n_21500) );
na02f04 g758896 ( .a(n_21435), .b(FE_OCPN5272_n_21434), .o(n_21544) );
in01s01 g758897 ( .a(n_21473), .o(n_21474) );
no02f04 g758898 ( .a(n_21435), .b(FE_OCPN5272_n_21434), .o(n_21473) );
no02s01 g758899 ( .a(n_21433), .b(n_21432), .o(n_21546) );
na02f04 g758900 ( .a(n_46966), .b(n_21728), .o(n_21803) );
in01s01 g758901 ( .a(n_21761), .o(n_21762) );
no02f04 g758902 ( .a(n_46966), .b(n_21728), .o(n_21761) );
no02s01 g758903 ( .a(FE_OCP_RBN1868_n_21358), .b(FE_OCP_RBN6061_n_21194), .o(n_21431) );
na02s01 g758904 ( .a(n_22061), .b(n_22060), .o(n_22062) );
in01s01 g758905 ( .a(n_21759), .o(n_21760) );
na02s01 g758906 ( .a(n_21677), .b(n_21727), .o(n_21759) );
na02f06 g758907 ( .a(n_21292), .b(n_21329), .o(n_21476) );
oa12s01 g758908 ( .a(n_21472), .b(n_21471), .c(n_21470), .o(n_21541) );
in01s01 g758909 ( .a(n_21705), .o(n_21648) );
oa12f06 g758910 ( .a(n_21569), .b(n_21642), .c(n_21487), .o(n_21705) );
no02s02 TIMEBOOST_cell_3348 ( .a(n_26794), .b(n_26868), .o(TIMEBOOST_net_965) );
oa12s01 g758912 ( .a(n_22059), .b(n_22058), .c(n_22057), .o(n_22116) );
oa12s01 g758913 ( .a(n_21643), .b(n_21642), .c(n_21641), .o(n_21702) );
no02m06 TIMEBOOST_cell_6290 ( .a(TIMEBOOST_net_1996), .b(n_10356), .o(n_10529) );
in01s01 g758915 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_6_), .o(n_23192) );
no02m08 g758918 ( .a(n_21572), .b(n_21490), .o(n_21611) );
no02m08 g758919 ( .a(n_21332), .b(FE_OCP_RBN6822_FE_RN_592_0), .o(n_21399) );
na02m04 g758921 ( .a(n_21332), .b(n_21192), .o(n_21363) );
in01s02 g758922 ( .a(n_21330), .o(n_21331) );
na02f04 g758923 ( .a(n_21288), .b(n_21240), .o(n_21330) );
na02m06 g758924 ( .a(n_21604), .b(n_21496), .o(n_21647) );
no02m06 g758925 ( .a(n_21605), .b(n_21495), .o(n_21646) );
na02s04 g758926 ( .a(n_21238), .b(n_45026), .o(n_21292) );
in01s02 g758929 ( .a(n_21430), .o(n_21661) );
na02m08 g758930 ( .a(n_21394), .b(n_45073), .o(n_21430) );
no02f02 g758931 ( .a(n_21233), .b(n_45024), .o(n_21365) );
no02m06 g758935 ( .a(n_21394), .b(n_45026), .o(n_21429) );
na02f04 g758936 ( .a(n_21237), .b(n_45070), .o(n_21329) );
na02m04 g758937 ( .a(n_21236), .b(n_45081), .o(n_21291) );
na02s02 g758938 ( .a(n_21700), .b(n_21604), .o(n_21701) );
no02s02 g758939 ( .a(n_21605), .b(n_21634), .o(n_21726) );
na02s01 g758940 ( .a(n_21606), .b(n_21644), .o(n_21645) );
no02m01 g758941 ( .a(n_21572), .b(n_21575), .o(n_21678) );
no02m04 TIMEBOOST_cell_6289 ( .a(n_10254), .b(n_10311), .o(TIMEBOOST_net_1996) );
no02m06 g758943 ( .a(n_21286), .b(n_19716), .o(n_21432) );
no02f04 g758944 ( .a(n_21285), .b(n_19715), .o(n_21433) );
na02s01 g758945 ( .a(n_21471), .b(n_21470), .o(n_21472) );
na02f02 g758946 ( .a(n_21640), .b(FE_OCP_DRV_N1486_n_21639), .o(n_21727) );
na02s01 g758947 ( .a(n_21641), .b(n_21642), .o(n_21643) );
in01s01 g758948 ( .a(n_21676), .o(n_21677) );
no02s02 g758949 ( .a(n_21640), .b(FE_OCP_DRV_N1486_n_21639), .o(n_21676) );
na02s02 TIMEBOOST_cell_3347 ( .a(TIMEBOOST_net_964), .b(n_36483), .o(n_36529) );
no02s06 TIMEBOOST_cell_7008 ( .a(TIMEBOOST_net_2262), .b(TIMEBOOST_net_1121), .o(n_10676) );
na02s01 g758952 ( .a(n_22058), .b(n_22057), .o(n_22059) );
oa12f06 g758955 ( .a(n_21391), .b(n_21280), .c(n_21470), .o(n_21428) );
ao12s01 g758957 ( .a(n_21448), .b(n_22011), .c(n_21516), .o(n_22061) );
in01s01 g758959 ( .a(FE_OCP_RBN3260_n_21360), .o(n_21393) );
in01s02 g758964 ( .a(n_21609), .o(n_21636) );
ao12m08 g758965 ( .a(n_21356), .b(n_21540), .c(n_21316), .o(n_21609) );
in01s01 g758968 ( .a(FE_OCP_RBN1869_n_21358), .o(n_21427) );
oa12s01 g758972 ( .a(n_22054), .b(n_22053), .c(n_22052), .o(n_22115) );
oa12s01 g758973 ( .a(n_21996), .b(n_22011), .c(n_21995), .o(n_22031) );
in01s01 g758974 ( .a(n_22119), .o(n_22056) );
in01s01 g758975 ( .a(n_22030), .o(n_22119) );
na03m04 TIMEBOOST_cell_2742 ( .a(n_11084), .b(n_11122), .c(n_11169), .o(n_11202) );
oa12s01 g758977 ( .a(n_22010), .b(n_22009), .c(n_22008), .o(n_22055) );
na02s01 g758978 ( .a(n_21392), .b(n_21322), .o(n_21545) );
na02m08 g758980 ( .a(n_21195), .b(FE_OCP_RBN6838_FE_RN_586_0), .o(n_21332) );
na02s02 g758984 ( .a(n_21535), .b(n_21269), .o(n_21576) );
no02s04 g758985 ( .a(n_21424), .b(n_21385), .o(n_21467) );
no02m04 g758987 ( .a(n_21202), .b(FE_OCP_RBN6823_FE_RN_592_0), .o(n_21289) );
in01m02 g758988 ( .a(n_21326), .o(n_21327) );
na02m02 g758989 ( .a(n_21288), .b(n_21287), .o(n_21326) );
in01s01 g758990 ( .a(n_21644), .o(n_21575) );
na02s03 g758991 ( .a(n_21537), .b(n_45072), .o(n_21644) );
in01s02 g758992 ( .a(n_21573), .o(n_21574) );
in01s01 g758994 ( .a(n_21538), .o(n_21539) );
na02s02 g758995 ( .a(n_21425), .b(n_21497), .o(n_21538) );
in01s01 g758997 ( .a(n_21572), .o(n_21606) );
no02m08 g758998 ( .a(n_21537), .b(n_45080), .o(n_21572) );
in01s02 g759000 ( .a(n_21605), .o(n_21700) );
no02s06 g759001 ( .a(n_21571), .b(n_45080), .o(n_21605) );
in01s02 g759004 ( .a(n_21604), .o(n_21634) );
na02s06 g759005 ( .a(n_21571), .b(n_45080), .o(n_21604) );
na02s04 g759006 ( .a(n_21531), .b(n_21496), .o(n_22039) );
no02s04 g759007 ( .a(n_21533), .b(n_21495), .o(n_22038) );
no02s01 g759008 ( .a(n_21279), .b(n_21323), .o(n_21471) );
na02s01 g759009 ( .a(n_21470), .b(n_21391), .o(n_21392) );
in01s01 g759010 ( .a(n_21632), .o(n_21633) );
na02s01 g759011 ( .a(n_21603), .b(n_21530), .o(n_21632) );
na02s01 g759012 ( .a(n_22053), .b(n_22052), .o(n_22054) );
na02s01 g759013 ( .a(n_22009), .b(n_22008), .o(n_22010) );
na02s01 g759014 ( .a(n_22011), .b(n_21995), .o(n_21996) );
in01m02 g759015 ( .a(n_21285), .o(n_21286) );
na02m08 g759017 ( .a(n_21232), .b(n_21200), .o(n_21394) );
oa12s01 g759018 ( .a(n_21355), .b(n_21354), .c(n_21353), .o(n_21426) );
in01s01 g759021 ( .a(n_21283), .o(n_21324) );
in01s01 g759022 ( .a(n_21238), .o(n_21283) );
in01f02 g759023 ( .a(n_21238), .o(n_21237) );
oa12f06 g759026 ( .a(n_21381), .b(n_21526), .c(n_21456), .o(n_21642) );
oa12s01 g759027 ( .a(n_21528), .b(n_21527), .c(n_21526), .o(n_21602) );
in01s01 g759028 ( .a(n_21281), .o(n_21282) );
in01m02 g759029 ( .a(n_21236), .o(n_21281) );
oa12s01 g759032 ( .a(n_21408), .b(n_21977), .c(n_21377), .o(n_22058) );
no02s10 TIMEBOOST_cell_5947 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_4_), .b(FE_OCP_RBN6517_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(TIMEBOOST_net_1825) );
in01s01 g759036 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_4_), .o(n_23135) );
no02m04 g759040 ( .a(n_21422), .b(n_21277), .o(n_21535) );
na02m08 g759041 ( .a(n_21318), .b(n_21317), .o(n_21356) );
na02m06 g759042 ( .a(FE_OCP_RBN1864_n_21163), .b(n_45026), .o(n_21232) );
no02f02 g759044 ( .a(n_21084), .b(n_45070), .o(n_21202) );
na02s02 g759045 ( .a(n_21127), .b(n_45091), .o(n_21288) );
na02s03 g759047 ( .a(n_21163), .b(n_45024), .o(n_21200) );
in01s01 g759049 ( .a(n_21496), .o(n_21533) );
na02s08 g759050 ( .a(n_21466), .b(n_45072), .o(n_21496) );
no02s08 g759051 ( .a(n_21421), .b(n_21219), .o(n_21540) );
in01s01 g759052 ( .a(n_21424), .o(n_21425) );
no02m02 g759053 ( .a(n_21390), .b(n_45072), .o(n_21424) );
na02s02 g759054 ( .a(n_21390), .b(n_45072), .o(n_21497) );
no02s02 g759056 ( .a(n_21521), .b(n_21490), .o(n_21630) );
in01s01 g759058 ( .a(n_21495), .o(n_21531) );
no02s08 g759059 ( .a(n_21466), .b(n_45080), .o(n_21495) );
no02s01 g759060 ( .a(FE_OCP_RBN6384_n_21087), .b(n_21080), .o(n_21199) );
in01s01 g759061 ( .a(n_21322), .o(n_21323) );
in01s01 g759062 ( .a(n_21280), .o(n_21322) );
no02m06 g759063 ( .a(n_21230), .b(FE_OCPN1707_n_21229), .o(n_21280) );
in01s01 g759064 ( .a(n_21391), .o(n_21279) );
na02f06 g759065 ( .a(n_21230), .b(FE_OCPN1707_n_21229), .o(n_21391) );
na02s01 g759066 ( .a(n_21354), .b(n_21353), .o(n_21355) );
in01s01 g759067 ( .a(n_21529), .o(n_21530) );
no02s06 g759068 ( .a(n_21494), .b(FE_OCPUNCON7069_n_21493), .o(n_21529) );
no02s01 g759069 ( .a(FE_OCP_RBN6383_n_21087), .b(n_21011), .o(n_21166) );
na02f04 g759070 ( .a(n_21494), .b(FE_OCPUNCON7069_n_21493), .o(n_21603) );
in01s03 g759071 ( .a(n_21197), .o(n_21198) );
ao12s08 g759072 ( .a(n_20661), .b(n_21143), .c(n_20786), .o(n_21197) );
na02s01 g759073 ( .a(n_21527), .b(n_21526), .o(n_21528) );
na02s01 g759074 ( .a(n_21488), .b(n_21569), .o(n_21641) );
no02s01 g759075 ( .a(n_21978), .b(n_21407), .o(n_22053) );
no02m08 g759076 ( .a(n_21131), .b(n_20667), .o(n_21196) );
na02s06 g759077 ( .a(n_21130), .b(FE_OCP_RBN6808_n_20667), .o(n_21165) );
in01f02 g759079 ( .a(n_21195), .o(n_21227) );
in01s01 g759082 ( .a(n_21959), .o(n_22011) );
ao12f04 g759083 ( .a(n_21452), .b(n_21909), .c(n_21410), .o(n_21959) );
no02m01 TIMEBOOST_cell_4201 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_30_), .b(FE_OFN736_n_17093), .o(TIMEBOOST_net_1191) );
oa12s01 g759085 ( .a(n_21958), .b(n_21909), .c(n_21957), .o(n_21994) );
ao12s01 g759086 ( .a(n_21774), .b(n_21909), .c(n_21826), .o(n_22009) );
in01s01 g759089 ( .a(FE_OCP_RBN6062_n_21194), .o(n_21278) );
ao22s06 g759092 ( .a(n_21093), .b(n_20749), .c(n_21143), .d(n_20751), .o(n_21194) );
na02s01 TIMEBOOST_cell_1140 ( .a(TIMEBOOST_net_184), .b(n_37472), .o(n_37474) );
in01s01 g759094 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_7_), .o(n_22657) );
in01m04 g759096 ( .a(n_21130), .o(n_21131) );
na02m08 g759097 ( .a(n_21093), .b(n_20750), .o(n_21130) );
no02m06 g759099 ( .a(n_21277), .b(n_21220), .o(n_21318) );
in01m02 g759100 ( .a(n_21132), .o(n_21133) );
na02f04 g759101 ( .a(n_21092), .b(n_21016), .o(n_21132) );
na02f04 g759103 ( .a(FE_OCP_RBN6837_FE_RN_586_0), .b(n_21192), .o(n_21224) );
na02s06 TIMEBOOST_cell_5407 ( .a(TIMEBOOST_net_1651), .b(n_30954), .o(n_31073) );
in01s02 g759105 ( .a(n_21421), .o(n_21422) );
na02m08 g759106 ( .a(n_21348), .b(FE_OCP_RBN5337_FE_RN_2064_0), .o(n_21421) );
na02s02 g759107 ( .a(n_21386), .b(n_21147), .o(n_21420) );
no02f04 g759108 ( .a(n_21387), .b(n_21175), .o(n_21464) );
na02m06 g759110 ( .a(n_21317), .b(n_21316), .o(n_21351) );
in01m02 g759111 ( .a(n_21491), .o(n_21492) );
no02m02 g759112 ( .a(n_21463), .b(n_21462), .o(n_21491) );
no02s08 g759117 ( .a(n_21461), .b(n_45080), .o(n_21490) );
in01s01 g759120 ( .a(n_21489), .o(n_21521) );
na02s08 g759121 ( .a(n_21461), .b(n_45080), .o(n_21489) );
no02m08 g759122 ( .a(n_21312), .b(n_45070), .o(n_21350) );
na02s01 TIMEBOOST_cell_1139 ( .a(n_37473), .b(n_37306), .o(TIMEBOOST_net_184) );
no02m04 TIMEBOOST_cell_1051 ( .a(FE_RN_2356_0), .b(FE_RN_2357_0), .o(TIMEBOOST_net_140) );
na02s01 g759126 ( .a(n_21909), .b(n_21957), .o(n_21958) );
in01s01 g759127 ( .a(n_21487), .o(n_21488) );
no02f06 g759128 ( .a(n_21459), .b(FE_OCPUNCON3488_n_21458), .o(n_21487) );
na02f06 g759129 ( .a(n_21459), .b(FE_OCPUNCON3488_n_21458), .o(n_21569) );
in01s01 g759130 ( .a(n_21977), .o(n_21978) );
na02s01 g759131 ( .a(n_21909), .b(n_21376), .o(n_21977) );
no02s01 g759132 ( .a(n_21160), .b(n_21187), .o(n_21354) );
no02s01 g759133 ( .a(n_21312), .b(FE_OCP_RBN3222_n_21242), .o(n_21419) );
in01m02 g759134 ( .a(n_21090), .o(n_21091) );
ao12m02 g759135 ( .a(n_20838), .b(n_21018), .c(n_20815), .o(n_21090) );
in01m03 g759136 ( .a(n_21088), .o(n_21089) );
oa12f06 g759137 ( .a(n_20674), .b(n_20983), .c(n_20575), .o(n_21088) );
no02s01 TIMEBOOST_cell_3238 ( .a(n_978), .b(n_1020), .o(TIMEBOOST_net_910) );
oa12s01 g759151 ( .a(n_21185), .b(n_21184), .c(n_21183), .o(n_21276) );
ao12f06 g759152 ( .a(n_21259), .b(n_21415), .c(n_21342), .o(n_21526) );
oa12s01 g759153 ( .a(n_21417), .b(n_21416), .c(n_21415), .o(n_21486) );
in01s06 g759162 ( .a(n_21093), .o(n_21143) );
no02m10 g759163 ( .a(n_21018), .b(n_20754), .o(n_21093) );
no02f04 TIMEBOOST_cell_6992 ( .a(TIMEBOOST_net_2254), .b(n_15149), .o(n_15338) );
na02s02 TIMEBOOST_cell_3237 ( .a(TIMEBOOST_net_909), .b(n_21069), .o(n_21177) );
na02m04 g759166 ( .a(n_21188), .b(n_21147), .o(n_21277) );
na02s04 g759169 ( .a(n_20951), .b(n_45013), .o(n_21016) );
na02m04 g759172 ( .a(n_21046), .b(n_45091), .o(n_21192) );
in01f02 g759175 ( .a(n_21386), .o(n_21387) );
in01f02 g759176 ( .a(n_21348), .o(n_21386) );
no02f08 g759177 ( .a(n_21266), .b(n_21214), .o(n_21348) );
in01s02 g759178 ( .a(n_21272), .o(n_21273) );
na02f02 g759179 ( .a(n_21188), .b(FE_OCP_RBN5338_FE_RN_2064_0), .o(n_21272) );
na02m04 g759180 ( .a(n_21157), .b(n_45023), .o(n_21317) );
no02s06 g759182 ( .a(n_21384), .b(n_45072), .o(n_21385) );
no02m02 g759183 ( .a(n_21384), .b(n_45072), .o(n_21463) );
no02s03 g759184 ( .a(n_21305), .b(FE_OCPN1711_n_45073), .o(n_21462) );
in01s01 g759185 ( .a(n_21186), .o(n_21187) );
na02m06 g759186 ( .a(n_21095), .b(n_19408), .o(n_21186) );
in01s01 g759187 ( .a(n_21159), .o(n_21160) );
na02f04 g759188 ( .a(n_21094), .b(n_19407), .o(n_21159) );
na02s01 g759189 ( .a(n_21184), .b(n_21183), .o(n_21185) );
na02s01 g759190 ( .a(n_21416), .b(n_21415), .o(n_21417) );
no02s01 g759191 ( .a(n_21382), .b(n_21456), .o(n_21527) );
no02f06 g759193 ( .a(n_20981), .b(n_20982), .o(n_21164) );
ao12f06 g759194 ( .a(n_21125), .b(n_21044), .c(n_21074), .o(n_21353) );
in01s01 g759196 ( .a(n_22156), .o(n_21413) );
in01s01 g759197 ( .a(n_21346), .o(n_22156) );
in01s02 g759198 ( .a(n_21346), .o(n_21345) );
na02f08 TIMEBOOST_cell_3332 ( .a(FE_RN_2670_0), .b(FE_RN_2669_0), .o(TIMEBOOST_net_957) );
na02s01 TIMEBOOST_cell_3218 ( .a(n_927), .b(n_963), .o(TIMEBOOST_net_900) );
no02f06 g759205 ( .a(n_21836), .b(n_21837), .o(n_21909) );
oa12s01 g759212 ( .a(n_21892), .b(n_21891), .c(n_21890), .o(n_21933) );
in01s04 g759215 ( .a(n_21014), .o(n_21015) );
in01s06 g759216 ( .a(n_20983), .o(n_21014) );
na02m10 g759217 ( .a(n_20947), .b(n_20712), .o(n_20983) );
no02m06 g759218 ( .a(n_20925), .b(n_20943), .o(n_20982) );
na02s04 g759219 ( .a(n_20980), .b(n_20944), .o(n_20981) );
na02s01 TIMEBOOST_cell_1086 ( .a(TIMEBOOST_net_157), .b(n_37289), .o(n_37348) );
in01s02 g759222 ( .a(n_21012), .o(n_21013) );
na02f02 g759223 ( .a(n_20980), .b(n_20924), .o(n_21012) );
na02m02 g759224 ( .a(n_21072), .b(n_45032), .o(n_21188) );
no02m02 g759227 ( .a(n_21220), .b(n_21219), .o(n_21269) );
no02m08 TIMEBOOST_cell_3217 ( .a(n_20684), .b(TIMEBOOST_net_899), .o(n_20821) );
no02s06 g759229 ( .a(n_21242), .b(FE_OCPN1382_n_45026), .o(n_21268) );
no02f04 g759230 ( .a(n_21344), .b(FE_OCP_DRV_N4510_n_21343), .o(n_21456) );
in01s01 g759231 ( .a(n_21381), .o(n_21382) );
na02f04 g759232 ( .a(n_21344), .b(FE_OCPN4515_n_21343), .o(n_21381) );
no02m04 g759233 ( .a(n_21801), .b(n_21835), .o(n_21837) );
na02s01 g759234 ( .a(n_21260), .b(n_21342), .o(n_21416) );
na02s01 g759235 ( .a(n_21891), .b(n_21890), .o(n_21892) );
no02s01 g759236 ( .a(n_21125), .b(n_21045), .o(n_21184) );
no02m10 g759237 ( .a(n_20947), .b(n_20607), .o(n_21018) );
ao12m06 g759239 ( .a(n_20531), .b(n_20926), .c(n_20535), .o(n_20945) );
in01s04 g759240 ( .a(n_21306), .o(n_21307) );
in01m04 g759241 ( .a(n_21266), .o(n_21306) );
na02f02 TIMEBOOST_cell_3328 ( .a(n_31232), .b(n_31099), .o(TIMEBOOST_net_955) );
in01m02 g759243 ( .a(n_21094), .o(n_21095) );
no02s01 TIMEBOOST_cell_6306 ( .a(TIMEBOOST_net_2004), .b(FE_OCP_RBN3308_n_43022), .o(n_43383) );
oa12s01 g759245 ( .a(n_21043), .b(n_21042), .c(n_21041), .o(n_21124) );
in01s01 g759246 ( .a(n_21264), .o(n_21265) );
in01s02 g759247 ( .a(n_21218), .o(n_21264) );
oa12f06 g759250 ( .a(n_21114), .b(n_21263), .c(n_21174), .o(n_21415) );
in01s04 g759251 ( .a(n_21305), .o(n_21384) );
oa12s01 g759253 ( .a(n_21258), .b(n_21263), .c(n_21257), .o(n_21341) );
in01s01 g759254 ( .a(FE_OCP_RBN3210_n_21203), .o(n_22134) );
ao12m04 g759258 ( .a(n_21374), .b(n_21755), .c(n_21835), .o(n_21836) );
oa12s01 g759259 ( .a(n_21758), .b(n_21757), .c(n_21756), .o(n_21802) );
in01s01 g759260 ( .a(n_21011), .o(n_21080) );
in01s01 g759263 ( .a(n_20984), .o(n_21011) );
in01m02 g759264 ( .a(n_20984), .o(n_20985) );
in01s01 g759268 ( .a(FE_OCPN7089_n_20979), .o(n_20978) );
in01s01 g759269 ( .a(n_20949), .o(n_20979) );
in01m02 g759270 ( .a(n_20949), .o(n_20950) );
na02m04 g759271 ( .a(n_20866), .b(n_20831), .o(n_20949) );
na02m04 g759273 ( .a(n_20948), .b(n_20922), .o(n_21046) );
no02m04 g759275 ( .a(n_20865), .b(n_20830), .o(n_20951) );
na02m02 g759279 ( .a(n_20802), .b(n_20578), .o(n_20831) );
na02s01 g759280 ( .a(n_21757), .b(n_21756), .o(n_21758) );
na02m04 g759281 ( .a(n_20803), .b(n_20579), .o(n_20866) );
in01m02 g759282 ( .a(n_20976), .o(n_20977) );
na02f04 g759283 ( .a(n_20944), .b(n_20943), .o(n_20976) );
no02f06 TIMEBOOST_cell_3239 ( .a(TIMEBOOST_net_910), .b(n_1255), .o(n_1266) );
no02f02 g759285 ( .a(n_20856), .b(n_20919), .o(n_20942) );
na02f04 g759286 ( .a(n_21077), .b(n_20995), .o(n_21078) );
no02m10 TIMEBOOST_cell_3327 ( .a(TIMEBOOST_net_954), .b(n_40398), .o(n_40409) );
na02s01 TIMEBOOST_cell_1085 ( .a(n_37230), .b(n_36973), .o(TIMEBOOST_net_157) );
na02m04 g759290 ( .a(FE_OCP_RBN6817_n_20889), .b(n_45091), .o(n_20948) );
no02s02 g759291 ( .a(n_20804), .b(n_45010), .o(n_20830) );
in01m02 g759292 ( .a(n_20924), .o(n_20925) );
na02f02 g759293 ( .a(n_20857), .b(n_45024), .o(n_20924) );
no02s04 g759295 ( .a(n_21064), .b(n_45024), .o(n_21220) );
no02m06 g759296 ( .a(n_21065), .b(n_45023), .o(n_21219) );
no02f08 g759298 ( .a(n_21214), .b(n_21175), .o(n_21261) );
in01f02 g759299 ( .a(n_21153), .o(n_21154) );
na02f02 g759300 ( .a(n_21040), .b(n_21077), .o(n_21153) );
no02m04 g759303 ( .a(n_20805), .b(n_45024), .o(n_20865) );
na02m02 g759304 ( .a(n_20889), .b(n_45069), .o(n_20922) );
in01s01 g759305 ( .a(n_21044), .o(n_21045) );
no02m04 g759307 ( .a(n_46969), .b(n_21007), .o(n_21125) );
na02s01 g759308 ( .a(n_21075), .b(FE_OCP_RBN2113_n_20935), .o(n_21076) );
na02s01 g759309 ( .a(n_21042), .b(n_21041), .o(n_21043) );
na02s01 g759310 ( .a(n_20862), .b(n_20867), .o(n_20868) );
in01s01 g759312 ( .a(n_21259), .o(n_21260) );
no02f04 g759313 ( .a(n_46968), .b(n_21212), .o(n_21259) );
na02f04 g759314 ( .a(n_46968), .b(n_21212), .o(n_21342) );
in01s01 g759315 ( .a(n_21801), .o(n_21891) );
na02m04 g759316 ( .a(n_21754), .b(n_21299), .o(n_21801) );
na02s01 g759317 ( .a(n_21257), .b(n_21263), .o(n_21258) );
in01s01 g759319 ( .a(n_21074), .o(n_21183) );
oa12f06 g759320 ( .a(n_20917), .b(n_20956), .c(n_21041), .o(n_21074) );
na02s02 TIMEBOOST_cell_5494 ( .a(n_16416), .b(n_16386), .o(TIMEBOOST_net_1695) );
na02s06 g759330 ( .a(n_21120), .b(n_21071), .o(n_21242) );
in01m04 g759331 ( .a(n_21149), .o(n_21150) );
in01s02 g759333 ( .a(n_21177), .o(n_21178) );
na03m08 TIMEBOOST_cell_6482 ( .a(n_24229), .b(FE_OFN743_delay_sub_ln23_0_unr15_stage6_stallmux_q), .c(n_24204), .o(n_24322) );
oa12s01 g759335 ( .a(n_21208), .b(n_21207), .c(n_21206), .o(n_21302) );
oa12s01 g759336 ( .a(n_21889), .b(n_21888), .c(n_21887), .o(n_21932) );
in01s01 g759337 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_4_), .o(n_22608) );
in01s01 g759339 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_2_), .o(n_22941) );
in01m01 g759341 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_1_), .o(n_22898) );
na02s01 g759343 ( .a(n_21888), .b(n_21887), .o(n_21889) );
na02f02 g759344 ( .a(n_21061), .b(n_21062), .o(n_21148) );
na02m06 g759345 ( .a(n_20829), .b(FE_OCP_RBN4362_FE_RN_1500_0), .o(n_20943) );
no02f04 TIMEBOOST_cell_6982 ( .a(TIMEBOOST_net_2249), .b(n_35008), .o(n_35097) );
in01s02 g759348 ( .a(n_20919), .o(n_20920) );
na02f02 g759349 ( .a(FE_OCP_RBN4361_FE_RN_1500_0), .b(n_20825), .o(n_20919) );
in01s06 g759352 ( .a(n_21147), .o(n_21175) );
na02m08 g759353 ( .a(n_21121), .b(n_45032), .o(n_21147) );
na02f02 g759354 ( .a(n_21006), .b(n_45091), .o(n_21077) );
in01f01 g759355 ( .a(n_21039), .o(n_21040) );
no02m02 g759356 ( .a(n_21006), .b(n_45091), .o(n_21039) );
no02s06 g759357 ( .a(n_21121), .b(n_45032), .o(n_21214) );
na02s06 g759358 ( .a(n_21069), .b(n_20665), .o(n_21071) );
na02s04 g759359 ( .a(n_20997), .b(n_20666), .o(n_21120) );
in01f02 g759360 ( .a(n_21754), .o(n_21755) );
no02m02 TIMEBOOST_cell_8673 ( .a(TIMEBOOST_net_2823), .b(n_26136), .o(n_26137) );
no03m04 TIMEBOOST_cell_3579 ( .a(FE_OCP_RBN5643_n_33977), .b(n_34003), .c(n_34011), .o(n_34086) );
na02s01 g759364 ( .a(n_21207), .b(n_21206), .o(n_21208) );
no02s01 g759365 ( .a(n_21115), .b(n_21174), .o(n_21257) );
no02s01 g759366 ( .a(n_20918), .b(n_20956), .o(n_21042) );
in01m02 g759367 ( .a(n_20926), .o(n_20861) );
na02m10 g759368 ( .a(n_20777), .b(n_20775), .o(n_20926) );
oa12s01 g759369 ( .a(n_21296), .b(n_21699), .c(n_21205), .o(n_21757) );
in01m02 g759370 ( .a(n_20802), .o(n_20803) );
ao12m02 g759371 ( .a(n_20539), .b(n_20693), .c(n_20492), .o(n_20802) );
ao12m08 g759374 ( .a(n_21035), .b(n_20967), .c(n_21036), .o(n_21119) );
in01s02 g759375 ( .a(n_21067), .o(n_21068) );
oa12s02 g759376 ( .a(n_20714), .b(n_20933), .c(n_20676), .o(n_21067) );
oa12s01 g759378 ( .a(n_21001), .b(n_21000), .c(n_20999), .o(n_21066) );
in01s01 g759379 ( .a(n_20889), .o(n_22126) );
na02f02 TIMEBOOST_cell_8026 ( .a(n_16827), .b(n_16825), .o(TIMEBOOST_net_2644) );
in01s01 g759383 ( .a(n_20862), .o(n_20859) );
in01s01 g759384 ( .a(n_20804), .o(n_20862) );
in01m02 g759385 ( .a(n_20804), .o(n_20805) );
in01s02 g759387 ( .a(n_21064), .o(n_21065) );
ao12f06 g759390 ( .a(n_21144), .b(n_21055), .c(n_21054), .o(n_21263) );
in01s01 g759392 ( .a(n_21075), .o(n_21096) );
in01s01 g759393 ( .a(n_21004), .o(n_21075) );
in01s02 g759394 ( .a(n_21004), .o(n_21003) );
oa12s04 g759399 ( .a(n_20459), .b(n_20973), .c(FE_OCP_RBN4353_FE_OCPN1263_n_20971), .o(n_21002) );
no02s01 TIMEBOOST_cell_1010 ( .a(TIMEBOOST_net_119), .b(n_37191), .o(n_37225) );
no03f10 TIMEBOOST_cell_6439 ( .a(FE_RN_426_0), .b(n_23639), .c(FE_RN_424_0), .o(TIMEBOOST_net_795) );
na02m03 TIMEBOOST_cell_8460 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n_6542), .o(TIMEBOOST_net_2717) );
in01f02 g759406 ( .a(n_20855), .o(n_20856) );
no02f04 g759407 ( .a(n_20829), .b(n_20828), .o(n_20855) );
na02f04 g759408 ( .a(n_20823), .b(n_20732), .o(n_20854) );
in01m02 g759410 ( .a(n_21062), .o(n_21063) );
no02m02 g759411 ( .a(n_21036), .b(n_21035), .o(n_21062) );
na02m02 g759414 ( .a(n_20771), .b(n_45066), .o(n_20825) );
na02s02 g759415 ( .a(n_20995), .b(n_20967), .o(n_21116) );
no02m02 g759416 ( .a(FE_OCP_RBN1603_n_20995), .b(n_20993), .o(n_21061) );
in01s01 g759417 ( .a(n_20917), .o(n_20918) );
na02f04 g759418 ( .a(n_20886), .b(n_20885), .o(n_20917) );
no02f04 g759419 ( .a(n_20886), .b(n_20885), .o(n_20956) );
na02s01 g759420 ( .a(n_21000), .b(n_20999), .o(n_21001) );
no02m06 TIMEBOOST_cell_3216 ( .a(n_20371), .b(n_20474), .o(TIMEBOOST_net_899) );
no02s04 g759423 ( .a(n_20991), .b(n_20963), .o(n_21034) );
in01s01 g759425 ( .a(n_21114), .o(n_21115) );
na02f04 g759426 ( .a(n_21059), .b(n_21058), .o(n_21114) );
no02s01 TIMEBOOST_cell_1009 ( .a(n_37224), .b(n_37167), .o(TIMEBOOST_net_119) );
no02s01 g759430 ( .a(n_21056), .b(n_21144), .o(n_21207) );
in01s04 g759432 ( .a(n_20997), .o(n_21069) );
no02m08 g759433 ( .a(n_20932), .b(n_20713), .o(n_20997) );
no02m08 g759434 ( .a(n_20696), .b(n_20654), .o(n_20775) );
oa12s01 g759435 ( .a(n_21699), .b(n_21714), .c(n_21819), .o(n_21888) );
na02m04 TIMEBOOST_cell_5623 ( .a(TIMEBOOST_net_1759), .b(n_16456), .o(n_16602) );
ao12f06 g759437 ( .a(n_20936), .b(n_20883), .c(n_20849), .o(n_21041) );
oa12s01 g759438 ( .a(n_20916), .b(n_20915), .c(n_20914), .o(n_20970) );
na02m08 g759445 ( .a(n_20939), .b(n_20968), .o(n_21121) );
oa12s01 g759447 ( .a(n_21111), .b(n_21110), .c(n_21109), .o(n_21173) );
oa12s01 g759448 ( .a(n_21886), .b(n_21885), .c(n_21884), .o(n_21931) );
na02s01 g759449 ( .a(n_21885), .b(n_21884), .o(n_21886) );
no02m08 g759450 ( .a(FE_OCP_RBN1140_n_19270), .b(n_20694), .o(n_20696) );
no02f06 g759451 ( .a(n_20732), .b(n_20774), .o(n_20829) );
no02f04 g759453 ( .a(n_20828), .b(n_20774), .o(n_20823) );
na02s06 g759454 ( .a(n_20910), .b(n_45032), .o(n_20939) );
na02m08 g759455 ( .a(FE_OCP_RBN1153_n_20910), .b(n_45069), .o(n_20968) );
na02f08 g759460 ( .a(n_20908), .b(n_45032), .o(n_20995) );
no02s08 g759461 ( .a(n_20966), .b(n_20879), .o(n_21036) );
in01s01 g759463 ( .a(n_20967), .o(n_20993) );
na02s08 g759464 ( .a(n_20907), .b(n_45069), .o(n_20967) );
na02m04 g759466 ( .a(n_20966), .b(FE_OCP_RBN5333_FE_RN_1490_0), .o(n_20991) );
na02s01 g759467 ( .a(n_20915), .b(n_20914), .o(n_20916) );
in01s01 g759468 ( .a(n_21055), .o(n_21056) );
na02f04 g759469 ( .a(n_21029), .b(n_21028), .o(n_21055) );
no02f04 g759470 ( .a(n_21029), .b(n_21028), .o(n_21144) );
na02s01 g759471 ( .a(n_21110), .b(n_21109), .o(n_21111) );
na02s08 g759473 ( .a(n_20913), .b(n_20608), .o(n_20973) );
no02s01 g759474 ( .a(n_20884), .b(n_20936), .o(n_21000) );
na02s02 TIMEBOOST_cell_3215 ( .a(n_20616), .b(TIMEBOOST_net_898), .o(FE_RN_572_0) );
in01s02 g759476 ( .a(n_20735), .o(n_20736) );
in01m02 g759477 ( .a(n_20693), .o(n_20735) );
ao12m04 g759478 ( .a(n_20654), .b(n_20652), .c(n_20442), .o(n_20693) );
na02f04 g759479 ( .a(n_21885), .b(n_21171), .o(n_21699) );
oa12m02 g759480 ( .a(n_20469), .b(n_20595), .c(FE_OCP_RBN2999_n_20374), .o(n_20620) );
ao12m04 g759481 ( .a(FE_OCP_RBN1842_FE_RN_442_0), .b(n_20374), .c(n_20652), .o(n_20653) );
oa12s01 g759483 ( .a(n_20962), .b(n_20961), .c(n_20960), .o(n_21027) );
in01s01 g759485 ( .a(n_20734), .o(n_20867) );
in01f02 g759486 ( .a(n_20734), .o(n_20733) );
na02f04 g759487 ( .a(n_20619), .b(n_20596), .o(n_20734) );
na02s01 TIMEBOOST_cell_1000 ( .a(TIMEBOOST_net_114), .b(n_1806), .o(n_1820) );
in01s01 g759494 ( .a(n_21054), .o(n_21206) );
oa12s04 g759498 ( .a(n_47258), .b(n_20821), .c(n_20396), .o(n_20891) );
in01s01 g759499 ( .a(n_20932), .o(n_20933) );
in01s01 g759503 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_3_), .o(n_22658) );
na02m04 g759505 ( .a(n_20552), .b(n_20470), .o(n_20619) );
na02m02 g759506 ( .a(n_20595), .b(n_20468), .o(n_20596) );
na02m08 g759507 ( .a(n_20912), .b(FE_OCP_RBN5333_FE_RN_1490_0), .o(n_21035) );
no02f06 g759508 ( .a(n_20651), .b(n_45067), .o(n_20828) );
no02m04 g759509 ( .a(n_20650), .b(n_45010), .o(n_20774) );
na02m06 g759510 ( .a(n_20878), .b(n_20842), .o(n_20966) );
na02f04 g759512 ( .a(n_20912), .b(FE_OCP_RBN1855_n_20879), .o(n_20963) );
na02s01 g759513 ( .a(FE_OCP_RBN3719_n_20621), .b(n_20555), .o(n_20691) );
in01s01 g759514 ( .a(n_20883), .o(n_20884) );
no02f04 g759516 ( .a(n_20853), .b(FE_OCPN5250_n_20852), .o(n_20936) );
na02s01 g759517 ( .a(n_20961), .b(n_20960), .o(n_20962) );
na02s01 TIMEBOOST_cell_999 ( .a(n_1550), .b(n_1527), .o(TIMEBOOST_net_114) );
na02s02 g759519 ( .a(n_20821), .b(FE_OCP_RBN5983_n_20495), .o(n_20822) );
no02s01 g759521 ( .a(n_20958), .b(n_20931), .o(n_21110) );
na02m10 g759522 ( .a(n_20850), .b(n_20426), .o(n_20913) );
na02m10 g759523 ( .a(n_20552), .b(n_20472), .o(n_20694) );
na02f04 g759524 ( .a(n_21455), .b(n_21380), .o(n_21885) );
in01s01 g759525 ( .a(n_20849), .o(n_20999) );
oa12m04 g759527 ( .a(FE_OCP_RBN4326_n_20333), .b(n_20767), .c(FE_OCPN4539_n_20332), .o(n_20799) );
na02m02 TIMEBOOST_cell_982 ( .a(n_23212), .b(TIMEBOOST_net_105), .o(n_23286) );
no02s01 TIMEBOOST_cell_984 ( .a(TIMEBOOST_net_106), .b(n_28298), .o(n_28339) );
in01s01 g759532 ( .a(n_22043), .o(n_20882) );
in01s01 g759533 ( .a(n_20848), .o(n_22043) );
in01f02 g759534 ( .a(n_20848), .o(n_20847) );
in01f04 g759536 ( .a(n_20907), .o(n_20908) );
no02s06 TIMEBOOST_cell_3182 ( .a(n_25731), .b(n_25824), .o(TIMEBOOST_net_882) );
no02s01 TIMEBOOST_cell_4391 ( .a(FE_OFN1196_n_27014), .b(n_30466), .o(TIMEBOOST_net_1286) );
oa12s01 g759539 ( .a(n_20798), .b(n_20820), .c(n_20797), .o(n_20915) );
na02f08 g759542 ( .a(FE_OCP_RBN1849_FE_RN_578_0), .b(n_20690), .o(n_20732) );
no02f04 TIMEBOOST_cell_5386 ( .a(n_16204), .b(n_16228), .o(TIMEBOOST_net_1641) );
no02f02 g759544 ( .a(n_20791), .b(n_20843), .o(n_20881) );
na02s02 TIMEBOOST_cell_4393 ( .a(n_4464), .b(n_4547), .o(TIMEBOOST_net_1287) );
no02s02 TIMEBOOST_cell_8529 ( .a(TIMEBOOST_net_2751), .b(n_2374), .o(n_2510) );
no02f08 g759548 ( .a(n_20846), .b(FE_OCPN1326_n_45050), .o(n_20879) );
na02m06 g759549 ( .a(n_20846), .b(FE_OCPN1326_n_45050), .o(n_20912) );
na02s01 g759550 ( .a(n_20820), .b(n_20797), .o(n_20798) );
na02m02 TIMEBOOST_cell_981 ( .a(n_23075), .b(FE_OCP_RBN5540_n_23307), .o(TIMEBOOST_net_105) );
no02s01 TIMEBOOST_cell_983 ( .a(n_28280), .b(n_27953), .o(TIMEBOOST_net_106) );
no02f02 TIMEBOOST_cell_5391 ( .a(TIMEBOOST_net_1643), .b(n_47013), .o(n_4283) );
in01s01 g759554 ( .a(n_20930), .o(n_20931) );
na02f04 g759555 ( .a(n_20872), .b(n_19098), .o(n_20930) );
in01s01 g759556 ( .a(n_20957), .o(n_20958) );
na02m06 g759557 ( .a(n_20873), .b(n_19099), .o(n_20957) );
no02s01 g759558 ( .a(n_21724), .b(n_21781), .o(n_21782) );
ao12s01 g759559 ( .a(n_21797), .b(n_21800), .c(n_21714), .o(n_21883) );
in01m04 g759560 ( .a(n_20595), .o(n_20652) );
in01m06 g759561 ( .a(n_20595), .o(n_20552) );
na02m08 g759563 ( .a(n_20447), .b(n_20341), .o(n_20595) );
oa12f02 g759564 ( .a(FE_OCP_RBN3131_n_21051), .b(n_21881), .c(n_21454), .o(n_21455) );
in01m02 g759565 ( .a(n_20730), .o(n_20731) );
na02f04 g759566 ( .a(n_20594), .b(FE_OCP_RBN1848_FE_RN_578_0), .o(n_20730) );
in01m02 g759567 ( .a(n_20904), .o(n_20905) );
in01s02 g759568 ( .a(n_20878), .o(n_20904) );
na02s01 TIMEBOOST_cell_5370 ( .a(n_27131), .b(FE_OCPN1340_n_27246), .o(TIMEBOOST_net_1633) );
in01f02 g759570 ( .a(n_20650), .o(n_20651) );
na02f06 TIMEBOOST_cell_4455 ( .a(n_39035), .b(n_39259), .o(TIMEBOOST_net_1318) );
na02s01 TIMEBOOST_cell_5076 ( .a(n_41300), .b(FE_OCP_RBN5676_n_41420), .o(TIMEBOOST_net_1486) );
ao12s01 g759579 ( .a(n_20841), .b(n_20877), .c(n_20876), .o(n_20961) );
in01m06 g759580 ( .a(n_20821), .o(n_20850) );
no02s01 TIMEBOOST_cell_978 ( .a(TIMEBOOST_net_103), .b(n_37333), .o(n_37442) );
in01s01 g759582 ( .a(n_20903), .o(n_21109) );
oa12s01 g759584 ( .a(n_21882), .b(n_21881), .c(n_21880), .o(n_21930) );
na02s06 g759586 ( .a(cordic_combinational_sub_ln23_0_unr20_z_0_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_), .o(n_21485) );
no02s03 g759587 ( .a(cordic_combinational_sub_ln23_0_unr20_z_0_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_), .o(n_21484) );
no02m02 g759588 ( .a(n_20445), .b(n_20439), .o(n_20481) );
na02m06 g759589 ( .a(n_20422), .b(n_20413), .o(n_20447) );
na02f06 TIMEBOOST_cell_8530 ( .a(FE_OCP_RBN2745_n_19747), .b(n_18230), .o(TIMEBOOST_net_2752) );
na02s01 g759591 ( .a(n_21881), .b(n_21880), .o(n_21882) );
na02s02 TIMEBOOST_cell_8705 ( .a(TIMEBOOST_net_2839), .b(FE_RN_67_0), .o(FE_RN_68_0) );
na02m02 g759593 ( .a(n_20641), .b(n_20548), .o(n_20687) );
no02m04 g759594 ( .a(n_20756), .b(n_20760), .o(n_20795) );
na03m06 TIMEBOOST_cell_8455 ( .a(n_27504), .b(n_27572), .c(n_27585), .o(n_27653) );
na02s02 g759596 ( .a(n_20549), .b(n_45066), .o(n_20594) );
na02f02 g759599 ( .a(n_20757), .b(n_20793), .o(n_20843) );
in01f02 g759600 ( .a(n_20874), .o(n_20875) );
na02f04 g759601 ( .a(FE_OCP_RBN5334_FE_RN_1490_0), .b(n_20842), .o(n_20874) );
no02s01 g759602 ( .a(n_20877), .b(n_20876), .o(n_20841) );
in01s06 g759604 ( .a(n_20767), .o(n_20764) );
na02m10 g759605 ( .a(n_20684), .b(n_20473), .o(n_20767) );
in01s01 g759606 ( .a(n_21724), .o(n_21725) );
oa12s02 g759607 ( .a(n_21698), .b(n_21601), .c(n_21374), .o(n_21724) );
na02f04 g759608 ( .a(n_20648), .b(n_20618), .o(n_20820) );
na02s02 TIMEBOOST_cell_6641 ( .a(n_41501), .b(n_41382), .o(TIMEBOOST_net_2078) );
no02s01 TIMEBOOST_cell_977 ( .a(n_37343), .b(n_37146), .o(TIMEBOOST_net_103) );
in01m02 g759618 ( .a(n_20872), .o(n_20873) );
na02m06 TIMEBOOST_cell_4457 ( .a(n_21497), .b(n_21467), .o(TIMEBOOST_net_1319) );
no02s03 TIMEBOOST_cell_5281 ( .a(TIMEBOOST_net_1588), .b(n_4385), .o(n_4604) );
in01s01 g759621 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_), .o(n_21453) );
na02s02 g759623 ( .a(n_21301), .b(n_21454), .o(n_21380) );
na02f04 g759624 ( .a(n_20598), .b(n_20317), .o(n_20648) );
na02m02 g759625 ( .a(n_20597), .b(n_20294), .o(n_20618) );
in01s02 g759626 ( .a(n_20690), .o(n_20647) );
no02f08 g759627 ( .a(n_20548), .b(n_20615), .o(n_20690) );
in01m02 g759628 ( .a(n_20790), .o(n_20791) );
no02f02 g759629 ( .a(n_20761), .b(n_20760), .o(n_20790) );
na02f08 TIMEBOOST_cell_4456 ( .a(TIMEBOOST_net_1318), .b(n_39356), .o(n_39446) );
na02s06 g759632 ( .a(n_20719), .b(n_45012), .o(n_20842) );
in01f01 g759633 ( .a(n_20756), .o(n_20757) );
no02f03 g759634 ( .a(n_20727), .b(n_45067), .o(n_20756) );
na02m02 g759635 ( .a(n_20727), .b(n_45067), .o(n_20793) );
na02f04 TIMEBOOST_cell_3103 ( .a(FE_OCP_RBN1164_n_24471), .b(TIMEBOOST_net_842), .o(n_24508) );
na02s04 g759637 ( .a(n_20640), .b(n_45012), .o(n_20683) );
na02s01 g759639 ( .a(n_20723), .b(n_44160), .o(n_20724) );
na02s01 g759640 ( .a(n_21752), .b(n_21831), .o(n_21832) );
na02m10 g759641 ( .a(n_20616), .b(n_20302), .o(n_20684) );
na02s02 TIMEBOOST_cell_5642 ( .a(n_6118), .b(n_5981), .o(TIMEBOOST_net_1769) );
no02s02 TIMEBOOST_cell_8612 ( .a(TIMEBOOST_net_2282), .b(n_5307), .o(TIMEBOOST_net_2793) );
in01f02 g759645 ( .a(n_20445), .o(n_20446) );
in01f01 g759646 ( .a(n_20422), .o(n_20445) );
ao12f06 g759647 ( .a(n_20264), .b(n_20321), .c(n_20240), .o(n_20422) );
no02s02 g759648 ( .a(n_21629), .b(n_21563), .o(n_21698) );
na02s01 g759649 ( .a(n_21799), .b(n_21798), .o(n_21800) );
na02m04 g759650 ( .a(n_21300), .b(n_21136), .o(n_21881) );
in01f02 g759651 ( .a(n_20641), .o(n_20642) );
in01s01 g759655 ( .a(n_20555), .o(n_20614) );
in01s01 g759659 ( .a(n_20510), .o(n_20555) );
na02m10 TIMEBOOST_cell_976 ( .a(n_32721), .b(TIMEBOOST_net_102), .o(FE_RN_770_0) );
oa12s01 g759663 ( .a(n_21879), .b(n_21878), .c(n_21877), .o(n_21929) );
na02s01 g759665 ( .a(n_21878), .b(n_21877), .o(n_21879) );
in01f04 g759666 ( .a(n_20553), .o(n_20548) );
no02f06 g759668 ( .a(n_20508), .b(n_20294), .o(n_20553) );
no02f04 g759669 ( .a(n_20682), .b(n_20638), .o(n_20761) );
no02f06 g759670 ( .a(n_20477), .b(n_45066), .o(n_20615) );
in01f02 g759672 ( .a(n_20721), .o(n_20722) );
no02f02 g759673 ( .a(n_20760), .b(n_20682), .o(n_20721) );
oa12s01 g759675 ( .a(n_21334), .b(n_21337), .c(n_21406), .o(n_21452) );
no02s02 g759676 ( .a(n_20349), .b(n_20281), .o(n_20383) );
no02s01 g759677 ( .a(n_21409), .b(n_21450), .o(n_21451) );
oa12s01 g759678 ( .a(n_21566), .b(n_21449), .c(n_21374), .o(n_21629) );
in01s01 g759679 ( .a(n_21796), .o(n_21797) );
no02s01 g759680 ( .a(n_21781), .b(n_21718), .o(n_21796) );
in01s01 g759681 ( .a(n_21300), .o(n_21301) );
na02m04 g759682 ( .a(n_21877), .b(n_21106), .o(n_21300) );
in01f02 g759683 ( .a(n_20597), .o(n_20598) );
no02s01 TIMEBOOST_cell_1012 ( .a(TIMEBOOST_net_120), .b(n_46253), .o(n_37284) );
no02s01 g759685 ( .a(n_21672), .b(n_21722), .o(n_21723) );
no02m03 TIMEBOOST_cell_6592 ( .a(TIMEBOOST_net_2053), .b(FE_RN_637_0), .o(FE_RN_639_0) );
in01s01 g759687 ( .a(n_21867), .o(n_21868) );
oa12s01 g759688 ( .a(n_21831), .b(n_21798), .c(n_21691), .o(n_21867) );
no02f06 g759692 ( .a(n_20611), .b(n_20591), .o(n_20719) );
in01s01 g759695 ( .a(FE_OCPN1942_n_20723), .o(n_20717) );
in01s01 g759696 ( .a(n_20640), .o(n_20723) );
oa12s01 g759699 ( .a(n_21256), .b(n_21255), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_21338) );
in01s01 g759700 ( .a(n_21865), .o(n_21866) );
oa22s01 g759701 ( .a(n_21750), .b(n_21714), .c(n_21721), .d(n_21691), .o(n_21865) );
in01s01 g759702 ( .a(n_21752), .o(n_21753) );
oa12s01 g759703 ( .a(n_21691), .b(n_21721), .c(n_21720), .o(n_21752) );
oa12s01 g759704 ( .a(n_21406), .b(n_21751), .c(n_21750), .o(n_21799) );
na02s01 g759705 ( .a(n_21255), .b(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_21256) );
na02f08 g759708 ( .a(n_20612), .b(n_20500), .o(n_20638) );
no02s01 TIMEBOOST_cell_1011 ( .a(n_46205), .b(n_46221), .o(TIMEBOOST_net_120) );
no02f04 g759710 ( .a(n_20417), .b(FE_OCPN869_n_45003), .o(n_20508) );
no02f02 g759711 ( .a(n_20545), .b(n_45008), .o(n_20591) );
no02f04 g759712 ( .a(n_44163), .b(n_45066), .o(n_20611) );
no02m02 g759716 ( .a(n_20542), .b(n_45066), .o(n_20682) );
no02f04 g759717 ( .a(n_20677), .b(FE_OCPN5246_n_18974), .o(n_20716) );
na02s02 g759718 ( .a(n_20755), .b(n_20787), .o(n_20838) );
na02s01 g759719 ( .a(n_21670), .b(n_21671), .o(n_21672) );
na02s01 g759720 ( .a(n_21798), .b(n_21691), .o(n_21831) );
oa12f02 g759721 ( .a(n_21107), .b(n_21172), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_21877) );
na02f02 g759723 ( .a(n_20587), .b(n_20612), .o(n_20678) );
in01s01 g759724 ( .a(n_21827), .o(n_21828) );
oa12s01 g759725 ( .a(n_21671), .b(n_21599), .c(n_21691), .o(n_21827) );
oa12s01 g759726 ( .a(n_20637), .b(n_20636), .c(n_20635), .o(n_20715) );
na02f04 g759728 ( .a(n_20348), .b(n_47174), .o(n_20477) );
no02s01 TIMEBOOST_cell_974 ( .a(TIMEBOOST_net_101), .b(n_17937), .o(n_18034) );
oa12s01 g759733 ( .a(FE_OCP_RBN3130_n_21051), .b(n_21482), .c(n_21481), .o(n_21483) );
no02s01 g759734 ( .a(n_21375), .b(n_21336), .o(n_21410) );
ao12f08 g759737 ( .a(n_20168), .b(n_20251), .c(n_20224), .o(n_20321) );
in01s01 g759738 ( .a(n_21409), .o(n_21566) );
ao12s01 g759739 ( .a(FE_OCP_RBN3126_n_21051), .b(n_21379), .c(n_21591), .o(n_21409) );
ao12s01 g759740 ( .a(n_21374), .b(n_21825), .c(n_21719), .o(n_21781) );
in01s01 g759741 ( .a(n_21863), .o(n_21864) );
ao12s01 g759742 ( .a(n_21778), .b(n_21694), .c(n_21714), .o(n_21863) );
no03s02 TIMEBOOST_cell_4715 ( .a(n_3887), .b(n_3871), .c(n_3864), .o(n_4015) );
na02f02 g759744 ( .a(n_47175), .b(n_45065), .o(n_20348) );
na02m06 g759746 ( .a(n_20501), .b(n_45060), .o(n_20612) );
na02f02 g759747 ( .a(n_20502), .b(n_45010), .o(n_20587) );
no02s01 g759748 ( .a(n_21600), .b(n_21104), .o(n_21601) );
no02s01 g759749 ( .a(n_21479), .b(n_21403), .o(n_22060) );
na02s01 g759750 ( .a(n_21775), .b(n_21826), .o(n_21957) );
na02m08 TIMEBOOST_cell_3998 ( .a(TIMEBOOST_net_1089), .b(FE_RN_474_0), .o(FE_RN_476_0) );
na02s01 g759752 ( .a(n_20635), .b(n_20636), .o(n_20637) );
no02s01 g759753 ( .a(n_21172), .b(n_21108), .o(n_21255) );
na02s01 g759754 ( .a(n_21404), .b(n_21516), .o(n_21480) );
no02s01 g759755 ( .a(n_21450), .b(n_20871), .o(n_21449) );
no02s01 TIMEBOOST_cell_973 ( .a(n_17359), .b(n_17431), .o(TIMEBOOST_net_101) );
no02s01 g759757 ( .a(n_21378), .b(n_21377), .o(n_22052) );
na02s01 g759758 ( .a(n_21299), .b(n_21253), .o(n_21756) );
no02f04 g759759 ( .a(n_20272), .b(FE_OCP_RBN5921_n_20236), .o(n_20320) );
na02s02 g759760 ( .a(n_21517), .b(n_21478), .o(n_21520) );
no02s01 g759761 ( .a(n_21407), .b(n_21378), .o(n_21408) );
in01s01 g759762 ( .a(n_21564), .o(n_21565) );
na02s01 g759763 ( .a(n_21519), .b(n_21402), .o(n_21564) );
no02s01 g759764 ( .a(n_21378), .b(n_20485), .o(n_21337) );
na02s01 g759765 ( .a(n_21519), .b(n_21447), .o(n_21518) );
na02s01 g759766 ( .a(n_21624), .b(n_21668), .o(n_21669) );
no02s06 TIMEBOOST_cell_4893 ( .a(TIMEBOOST_net_1394), .b(n_6790), .o(n_6907) );
in01s04 g759768 ( .a(n_20677), .o(n_20960) );
no02f06 g759769 ( .a(n_20636), .b(FE_OCPN5248_FE_OFN4715_n_18642), .o(n_20677) );
in01s01 g759770 ( .a(n_20754), .o(n_20755) );
na02s06 g759771 ( .a(n_20634), .b(n_20712), .o(n_20754) );
na02s01 g759772 ( .a(n_21252), .b(n_21253), .o(n_21254) );
in01s01 g759773 ( .a(n_21375), .o(n_21376) );
na02s01 g759774 ( .a(n_21248), .b(n_21826), .o(n_21375) );
na02s01 g759775 ( .a(n_21517), .b(n_21516), .o(n_21995) );
na02s01 g759776 ( .a(n_21335), .b(n_21297), .o(n_21336) );
no02s01 g759777 ( .a(n_21795), .b(n_21298), .o(n_22179) );
in01s01 g759778 ( .a(n_21715), .o(n_21716) );
no02s01 g759779 ( .a(n_21697), .b(n_21450), .o(n_21715) );
in01s01 g759780 ( .a(n_21627), .o(n_21628) );
na02s01 g759781 ( .a(n_21598), .b(n_21622), .o(n_21627) );
in01s01 g759782 ( .a(n_21695), .o(n_21696) );
na02s01 g759783 ( .a(n_21670), .b(n_21560), .o(n_21695) );
na02s01 g759784 ( .a(n_21599), .b(n_21374), .o(n_21671) );
in01s01 g759785 ( .a(n_21861), .o(n_21862) );
na02s01 g759786 ( .a(n_21773), .b(n_21825), .o(n_21861) );
in01s01 g759787 ( .a(n_21776), .o(n_21777) );
no02s01 g759788 ( .a(n_21749), .b(n_21748), .o(n_21776) );
no02s01 g759789 ( .a(n_21694), .b(FE_OCP_RBN3130_n_21051), .o(n_21778) );
in01s01 g759790 ( .a(n_21859), .o(n_21860) );
na02s01 g759791 ( .a(n_21824), .b(n_21693), .o(n_21859) );
oa12s01 g759792 ( .a(n_21622), .b(n_21374), .c(n_21562), .o(n_21563) );
ao12s01 g759793 ( .a(n_21142), .b(n_21141), .c(n_21140), .o(n_21798) );
in01f01 g759794 ( .a(n_20417), .o(n_20418) );
no02m06 TIMEBOOST_cell_6256 ( .a(TIMEBOOST_net_1979), .b(n_43441), .o(n_43626) );
ao12s01 g759796 ( .a(n_21446), .b(n_21714), .c(n_21481), .o(n_22176) );
in01s01 g759797 ( .a(n_21857), .o(n_21858) );
oa22s01 g759798 ( .a(n_21714), .b(n_20809), .c(n_21691), .d(n_21591), .o(n_21857) );
in01m02 g759799 ( .a(n_20505), .o(n_20506) );
in01m02 g759800 ( .a(n_20476), .o(n_20505) );
ao12f08 g759801 ( .a(n_20244), .b(n_20379), .c(n_20285), .o(n_20476) );
oa22s01 g759802 ( .a(n_21691), .b(n_21454), .c(n_21714), .d(n_20179), .o(n_21880) );
oa12s01 g759813 ( .a(n_21335), .b(n_21714), .c(n_21244), .o(n_22057) );
in01s01 g759814 ( .a(n_21821), .o(n_21822) );
oa12s01 g759815 ( .a(n_21668), .b(n_21691), .c(n_21595), .o(n_21821) );
in01s01 g759816 ( .a(n_21855), .o(n_21856) );
oa22s01 g759817 ( .a(n_21714), .b(n_21597), .c(n_21691), .d(n_21562), .o(n_21855) );
oa12s01 g759818 ( .a(n_21598), .b(FE_OCP_RBN3130_n_21051), .c(n_21597), .o(n_21722) );
in01s01 g759819 ( .a(n_21853), .o(n_21854) );
oa22s01 g759820 ( .a(n_21714), .b(n_21626), .c(n_21691), .d(n_21719), .o(n_21853) );
ao12s01 g759821 ( .a(FE_OCP_RBN3130_n_21051), .b(n_21626), .c(n_21625), .o(n_21779) );
in01s01 g759822 ( .a(n_21750), .o(n_21721) );
oa12s01 g759823 ( .a(n_21139), .b(n_21138), .c(n_21137), .o(n_21750) );
oa22s01 g759824 ( .a(n_21714), .b(n_21105), .c(n_21691), .d(n_21134), .o(n_21878) );
oa22s01 g759825 ( .a(n_21714), .b(n_21819), .c(n_21691), .d(n_20198), .o(n_21884) );
oa12s01 g759826 ( .a(n_21252), .b(n_21714), .c(n_21169), .o(n_21887) );
ao22s01 g759827 ( .a(n_21691), .b(n_21835), .c(n_21714), .d(n_20255), .o(n_21890) );
ao12s01 g759828 ( .a(n_21247), .b(n_21691), .c(n_21294), .o(n_22008) );
in01s02 g759837 ( .a(n_22280), .o(n_24620) );
in01s06 g759838 ( .a(n_22207), .o(n_22280) );
in01s01 g759845 ( .a(FE_OCPN1354_n_22484), .o(n_24691) );
in01s01 g759846 ( .a(n_22393), .o(n_22484) );
in01s02 g759849 ( .a(n_22207), .o(n_22393) );
in01s06 g759853 ( .a(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_22207) );
in01s03 g759858 ( .a(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_22089) );
in01s03 g759866 ( .a(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24624) );
in01s06 g759874 ( .a(FE_OFN5075_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_22111) );
in01s02 g759880 ( .a(FE_OFN741_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_21975) );
in01s02 g759888 ( .a(FE_OFN741_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_21852) );
na02f02 g759891 ( .a(n_20273), .b(FE_OCPN869_n_45003), .o(n_20297) );
no03m04 TIMEBOOST_cell_6255 ( .a(n_43329), .b(n_43370), .c(n_43364), .o(TIMEBOOST_net_1979) );
no02s01 g759893 ( .a(n_21141), .b(n_21140), .o(n_21142) );
na02s01 g759894 ( .a(n_21138), .b(n_21137), .o(n_21139) );
in01s01 g759895 ( .a(n_21379), .o(n_21298) );
na02s01 g759896 ( .a(FE_OCP_RBN3130_n_21051), .b(n_21251), .o(n_21379) );
na02s01 g759897 ( .a(n_21374), .b(n_21514), .o(n_21670) );
in01s01 g759898 ( .a(n_21598), .o(n_21561) );
na02s01 g759899 ( .a(n_21374), .b(n_20895), .o(n_21598) );
in01s01 g759900 ( .a(n_21478), .o(n_21479) );
na02s01 g759901 ( .a(n_21374), .b(n_21373), .o(n_21478) );
in01s01 g759902 ( .a(n_21774), .o(n_21775) );
no02s01 g759903 ( .a(n_21406), .b(n_21246), .o(n_21774) );
in01s01 g759904 ( .a(n_21751), .o(n_21693) );
no02s01 g759905 ( .a(n_21374), .b(n_21720), .o(n_21751) );
na02s01 g759906 ( .a(n_21406), .b(n_20894), .o(n_21622) );
na02s01 g759907 ( .a(n_21051), .b(n_21819), .o(n_21171) );
oa12m06 g759908 ( .a(n_20473), .b(n_20370), .c(FE_OCP_RBN4334_n_20242), .o(n_20474) );
no02m02 g759909 ( .a(n_21053), .b(n_21052), .o(n_21172) );
in01s01 g759910 ( .a(n_21107), .o(n_21108) );
na02m02 g759911 ( .a(n_21053), .b(n_21052), .o(n_21107) );
no02s10 TIMEBOOST_cell_908 ( .a(n_17442), .b(TIMEBOOST_net_68), .o(n_17579) );
na04m20 TIMEBOOST_cell_6401 ( .a(n_16988), .b(n_44721), .c(n_16900), .d(FE_OCP_RBN7105_n_44365), .o(FE_RN_1414_0) );
in01s01 g759914 ( .a(n_21297), .o(n_21377) );
na02s01 g759915 ( .a(n_21051), .b(n_21249), .o(n_21297) );
no02s01 g759916 ( .a(n_21051), .b(n_21249), .o(n_21378) );
na02s02 g759917 ( .a(n_21051), .b(n_21105), .o(n_21106) );
na02s02 g759918 ( .a(FE_OCP_RBN3127_n_21051), .b(n_21134), .o(n_21136) );
na02s01 g759919 ( .a(n_21051), .b(n_20156), .o(n_21253) );
in01s01 g759920 ( .a(n_21252), .o(n_21205) );
na02s01 g759921 ( .a(n_21051), .b(n_21169), .o(n_21252) );
na02s01 g759922 ( .a(FE_OCP_RBN3131_n_21051), .b(n_20157), .o(n_21299) );
in01s01 g759923 ( .a(n_21247), .o(n_21248) );
no02s01 g759924 ( .a(FE_OCP_RBN3131_n_21051), .b(n_21294), .o(n_21247) );
na02s01 g759925 ( .a(n_21051), .b(n_21246), .o(n_21826) );
na02s01 g759926 ( .a(n_21051), .b(n_21244), .o(n_21335) );
na02s01 g759927 ( .a(FE_OCP_RBN3130_n_21051), .b(n_21405), .o(n_21516) );
in01s01 g759928 ( .a(n_21448), .o(n_21517) );
no02s02 g759929 ( .a(n_21406), .b(n_21405), .o(n_21448) );
in01s01 g759930 ( .a(n_21403), .o(n_21404) );
no02s01 g759931 ( .a(n_21374), .b(n_21373), .o(n_21403) );
in01s01 g759932 ( .a(n_21482), .o(n_21402) );
no02s01 g759933 ( .a(FE_OCP_RBN3126_n_21051), .b(n_21371), .o(n_21482) );
na02s01 g759934 ( .a(n_21374), .b(n_21371), .o(n_21519) );
in01s01 g759935 ( .a(n_21446), .o(n_21447) );
no02s01 g759936 ( .a(n_21406), .b(n_21481), .o(n_21446) );
no02s01 g759937 ( .a(n_21406), .b(n_21251), .o(n_21795) );
no02s01 g759938 ( .a(FE_OCP_RBN3126_n_21051), .b(n_21370), .o(n_21450) );
in01s01 g759939 ( .a(n_21624), .o(n_21697) );
na02s01 g759940 ( .a(n_21374), .b(n_21370), .o(n_21624) );
na02s01 g759941 ( .a(n_21374), .b(n_21595), .o(n_21668) );
in01s01 g759942 ( .a(n_21600), .o(n_21560) );
no02s01 g759943 ( .a(n_21374), .b(n_21514), .o(n_21600) );
na02s01 g759944 ( .a(FE_OCP_RBN3130_n_21051), .b(n_21625), .o(n_21825) );
in01s01 g759945 ( .a(n_21772), .o(n_21773) );
no02s01 g759946 ( .a(n_21406), .b(n_21625), .o(n_21772) );
no02s01 g759947 ( .a(n_21374), .b(n_21593), .o(n_21748) );
in01s01 g759948 ( .a(n_21692), .o(n_21749) );
na02s01 g759949 ( .a(n_21374), .b(n_21593), .o(n_21692) );
na02s01 g759950 ( .a(n_21691), .b(n_21720), .o(n_21824) );
no02s02 g759951 ( .a(n_20753), .b(n_20667), .o(n_20815) );
in01s01 g759953 ( .a(n_21599), .o(n_21104) );
ao12s01 g759954 ( .a(n_20989), .b(n_20988), .c(n_20987), .o(n_21599) );
in01f02 g759955 ( .a(n_20271), .o(n_20272) );
in01m01 g759956 ( .a(n_20251), .o(n_20271) );
ao12f08 g759957 ( .a(n_20090), .b(n_20195), .c(n_20144), .o(n_20251) );
oa12s01 g759958 ( .a(n_21374), .b(n_21591), .c(n_20699), .o(n_21592) );
in01f02 g759959 ( .a(n_20501), .o(n_20502) );
na03m01 TIMEBOOST_cell_8445 ( .a(FE_OCPN945_n_27287), .b(n_26653), .c(n_27375), .o(n_27484) );
na02s01 g759961 ( .a(n_20709), .b(n_20456), .o(n_20787) );
in01s01 g759962 ( .a(n_21295), .o(n_21296) );
no02s01 g759963 ( .a(n_21051), .b(n_20199), .o(n_21295) );
in01s01 g759964 ( .a(n_21334), .o(n_21407) );
oa12s01 g759965 ( .a(FE_OCP_RBN3126_n_21051), .b(n_21294), .c(n_20327), .o(n_21334) );
oa12s01 g759969 ( .a(n_21103), .b(n_21102), .c(n_21101), .o(n_21694) );
no02f06 TIMEBOOST_cell_7654 ( .a(n_13480), .b(n_13507), .o(TIMEBOOST_net_2458) );
no02s01 g759971 ( .a(n_20988), .b(n_20987), .o(n_20989) );
in01s01 g759973 ( .a(n_20500), .o(n_20540) );
na02f06 g759974 ( .a(n_20435), .b(n_45101), .o(n_20500) );
no02s10 TIMEBOOST_cell_6864 ( .a(n_6734), .b(TIMEBOOST_net_2190), .o(n_6760) );
no02s01 TIMEBOOST_cell_6179 ( .a(FE_OCP_RBN5953_FE_OFN4772_n_44463), .b(n_44492), .o(TIMEBOOST_net_1941) );
na02s01 g759977 ( .a(n_21102), .b(n_21101), .o(n_21103) );
no02f02 g759978 ( .a(n_20163), .b(n_20215), .o(n_20229) );
na02s02 g759979 ( .a(n_20374), .b(n_20469), .o(n_20470) );
no02s02 g759980 ( .a(FE_OCP_RBN3000_n_20374), .b(FE_OCP_RBN1841_FE_RN_442_0), .o(n_20468) );
na02s01 g759981 ( .a(n_20675), .b(n_20657), .o(n_20676) );
no02s01 TIMEBOOST_cell_912 ( .a(TIMEBOOST_net_70), .b(n_32783), .o(n_32865) );
na02s06 g759983 ( .a(n_20529), .b(n_20606), .o(n_20607) );
in01s02 g759986 ( .a(n_20441), .o(n_20442) );
na02m06 g759987 ( .a(n_20375), .b(n_20374), .o(n_20441) );
in01s01 g759988 ( .a(n_20582), .o(n_20583) );
no02s06 g759989 ( .a(n_20491), .b(n_20539), .o(n_20582) );
no03f08 TIMEBOOST_cell_8433 ( .a(n_20026), .b(TIMEBOOST_net_2663), .c(n_20092), .o(n_20169) );
in01f02 g759991 ( .a(n_20414), .o(n_20415) );
in01s02 g759992 ( .a(n_20379), .o(n_20414) );
na02m08 g759993 ( .a(n_20291), .b(n_20267), .o(n_20379) );
no02s02 g759995 ( .a(n_20532), .b(n_20534), .o(n_20632) );
na02s01 g759997 ( .a(n_20674), .b(n_20533), .o(n_20710) );
na02s01 g759998 ( .a(FE_OCP_RBN1831_n_19663), .b(n_20660), .o(n_20709) );
na02s02 g759999 ( .a(n_20752), .b(n_20664), .o(n_20753) );
na02s02 g760000 ( .a(FE_OCP_RBN6808_n_20667), .b(n_20750), .o(n_20751) );
no02s02 g760001 ( .a(n_20667), .b(n_20669), .o(n_20749) );
no02s02 g760003 ( .a(n_20667), .b(n_20778), .o(n_20786) );
in01s02 g760013 ( .a(n_21406), .o(n_21691) );
in01s02 g760022 ( .a(n_21691), .o(n_21714) );
in01s02 g760024 ( .a(n_21374), .o(n_21406) );
in01s04 g760036 ( .a(FE_OCP_RBN3130_n_21051), .o(n_21374) );
in01m04 g760043 ( .a(n_21053), .o(n_21051) );
ao12f04 g760044 ( .a(n_20068), .b(n_20897), .c(n_21019), .o(n_21053) );
no02f04 g760045 ( .a(FE_OCP_RBN1837_n_20215), .b(n_20162), .o(n_20250) );
na02f02 g760047 ( .a(n_20413), .b(n_20342), .o(n_20439) );
ao12s01 g760048 ( .a(n_20037), .b(n_21050), .c(n_21019), .o(n_21141) );
oa12s01 g760049 ( .a(n_20254), .b(n_21050), .c(n_20218), .o(n_21138) );
oa12s01 g760051 ( .a(n_20914), .b(FE_OCPN4931_n_20275), .c(n_20293), .o(n_20378) );
in01s02 g760052 ( .a(n_20672), .o(n_20673) );
in01s01 g760054 ( .a(n_20836), .o(n_20837) );
na02m06 TIMEBOOST_cell_4917 ( .a(TIMEBOOST_net_1406), .b(n_1874), .o(n_1950) );
no02s02 g760056 ( .a(n_20409), .b(n_20406), .o(n_20465) );
no03s02 TIMEBOOST_cell_8222 ( .a(n_18912), .b(n_18913), .c(n_19416), .o(TIMEBOOST_net_2438) );
ao12s01 g760058 ( .a(n_21100), .b(n_21099), .c(n_21098), .o(n_21593) );
oa12f04 g760059 ( .a(n_20188), .b(n_20313), .c(n_20125), .o(n_20344) );
na02m06 TIMEBOOST_cell_888 ( .a(n_6889), .b(TIMEBOOST_net_58), .o(n_6980) );
no02m06 TIMEBOOST_cell_6806 ( .a(TIMEBOOST_net_2160), .b(n_10671), .o(n_10810) );
na02s02 g760065 ( .a(n_20752), .b(n_20705), .o(n_20812) );
in01s01 g760066 ( .a(n_20670), .o(n_20671) );
na02s02 g760067 ( .a(n_20606), .b(n_20573), .o(n_20670) );
in01s01 g760073 ( .a(n_21626), .o(n_21719) );
oa12s01 g760074 ( .a(n_21024), .b(n_21023), .c(n_21022), .o(n_21626) );
ao12s01 g760075 ( .a(n_21021), .b(n_21050), .c(n_21020), .o(n_21720) );
in01s02 g760076 ( .a(n_20784), .o(n_20785) );
na02s02 TIMEBOOST_cell_8709 ( .a(TIMEBOOST_net_2841), .b(FE_OCP_RBN2439_n_6937), .o(n_7002) );
in01s01 g760078 ( .a(n_20578), .o(n_20579) );
oa22s02 g760079 ( .a(n_20429), .b(FE_OCP_RBN1139_n_19270), .c(FE_OCP_RBN3018_n_20404), .d(FE_OCPN1665_FE_OCP_RBN1138_n_19270), .o(n_20578) );
in01s01 g760081 ( .a(n_20294), .o(n_20317) );
no02s03 g760082 ( .a(n_20245), .b(FE_OCPN869_n_45003), .o(n_20294) );
no02s01 g760083 ( .a(n_21099), .b(n_21098), .o(n_21100) );
na02s01 g760084 ( .a(n_21023), .b(n_21022), .o(n_21024) );
no02s01 g760085 ( .a(n_21050), .b(n_21020), .o(n_21021) );
in01s01 g760087 ( .a(n_20375), .o(n_20409) );
na02s04 g760088 ( .a(n_20340), .b(n_20343), .o(n_20375) );
na02f02 g760089 ( .a(n_20340), .b(FE_OCP_RBN5378_n_19055), .o(n_20342) );
na02s04 g760090 ( .a(FE_OCP_RBN5378_n_19055), .b(n_20340), .o(n_20341) );
na02s06 g760091 ( .a(FE_OCP_RBN4351_n_20456), .b(n_20536), .o(n_20606) );
in01s01 g760092 ( .a(n_20534), .o(n_20535) );
no02s02 g760094 ( .a(n_20429), .b(FE_OCP_RBN2064_n_19353), .o(n_20534) );
na03s08 TIMEBOOST_cell_8265 ( .a(n_8011), .b(n_7970), .c(n_7330), .o(n_8342) );
na02s02 g760098 ( .a(n_20275), .b(n_20293), .o(n_20914) );
in01s01 g760100 ( .a(n_20533), .o(n_20575) );
in01f01 g760103 ( .a(n_20195), .o(n_20215) );
ao12f08 g760104 ( .a(n_20029), .b(n_20107), .c(n_20006), .o(n_20195) );
na02m06 g760109 ( .a(n_20340), .b(FE_OCP_RBN1134_n_19077), .o(n_20374) );
na02f08 TIMEBOOST_cell_7912 ( .a(n_25998), .b(n_23466), .o(TIMEBOOST_net_2587) );
no02s02 g760111 ( .a(n_20404), .b(n_20343), .o(n_20406) );
in01s02 g760112 ( .a(n_20463), .o(n_20464) );
no02s06 g760113 ( .a(n_20332), .b(FE_OCP_RBN4325_n_20333), .o(n_20463) );
in01s02 g760114 ( .a(n_20337), .o(n_20338) );
no02s06 g760115 ( .a(n_20289), .b(n_47257), .o(n_20337) );
na02m02 TIMEBOOST_cell_5050 ( .a(n_13667), .b(FE_OCP_RBN4096_n_12880), .o(TIMEBOOST_net_1473) );
no02s06 g760117 ( .a(FE_OCP_RBN3017_n_20404), .b(n_19245), .o(n_20539) );
na02s06 TIMEBOOST_cell_887 ( .a(n_6634), .b(FE_RN_230_0), .o(TIMEBOOST_net_58) );
na02s40 TIMEBOOST_cell_7400 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_2_), .b(FE_OCP_RBN7005_n_44962), .o(TIMEBOOST_net_2331) );
no02f02 g760120 ( .a(n_20187), .b(n_20313), .o(n_20314) );
na02f01 g760121 ( .a(FE_RN_109_0), .b(n_20311), .o(n_20312) );
no02s02 g760122 ( .a(n_20309), .b(n_20269), .o(n_20310) );
na02s02 g760123 ( .a(n_20334), .b(n_20333), .o(n_20371) );
no02s06 g760124 ( .a(n_20332), .b(n_20369), .o(n_20370) );
na02s02 g760126 ( .a(n_20395), .b(n_47258), .o(n_20495) );
no02s02 g760127 ( .a(FE_OCP_RBN3018_n_20404), .b(FE_OCP_RBN1146_n_19353), .o(n_20532) );
no02s06 g760128 ( .a(FE_OCP_RBN4351_n_20456), .b(FE_OCP_RBN1146_n_19353), .o(n_20531) );
na02s02 TIMEBOOST_cell_6719 ( .a(n_2951), .b(n_3006), .o(TIMEBOOST_net_2117) );
na02s01 g760132 ( .a(n_20456), .b(FE_OCP_RBN1825_n_19513), .o(n_20573) );
na02s01 g760133 ( .a(n_20456), .b(FE_OCP_RBN4182_n_19599), .o(n_20708) );
in01s01 g760134 ( .a(n_20750), .o(n_20669) );
na02s02 g760135 ( .a(n_20456), .b(n_20630), .o(n_20750) );
in01s01 g760136 ( .a(n_20491), .o(n_20492) );
no02s01 TIMEBOOST_cell_911 ( .a(n_32796), .b(n_32486), .o(TIMEBOOST_net_70) );
no02s06 g760138 ( .a(n_20404), .b(n_19268), .o(n_20491) );
no02s02 g760144 ( .a(n_20456), .b(n_20630), .o(n_20667) );
no02s02 g760146 ( .a(FE_OCP_RBN5961_n_20459), .b(FE_OCP_RBN3003_n_20432), .o(n_20570) );
na02s01 g760147 ( .a(n_20456), .b(FE_OCP_RBN5705_n_19663), .o(n_20705) );
in01s02 g760148 ( .a(n_20665), .o(n_20666) );
na02s04 g760149 ( .a(n_20628), .b(FE_OCP_RBN6803_n_20565), .o(n_20665) );
na02s03 g760151 ( .a(n_20432), .b(n_20430), .o(n_20482) );
in01s01 g760152 ( .a(n_20778), .o(n_20664) );
no02s01 g760153 ( .a(n_20456), .b(n_19654), .o(n_20778) );
na02s01 g760154 ( .a(FE_OCP_RBN4351_n_20456), .b(FE_OCP_RBN1831_n_19663), .o(n_20752) );
na04s01 TIMEBOOST_cell_8358 ( .a(n_15964), .b(n_16615), .c(n_15965), .d(n_16630), .o(n_16721) );
no02s02 g760156 ( .a(n_20565), .b(n_20605), .o(n_20675) );
na02s06 g760158 ( .a(FE_OCP_RBN4351_n_20456), .b(n_20528), .o(n_20529) );
na02m01 g760159 ( .a(FE_OCP_RBN3018_n_20404), .b(n_20528), .o(n_20674) );
na02s04 g760160 ( .a(n_20299), .b(FE_OCP_RBN5379_n_19055), .o(n_20413) );
ao12s01 g760161 ( .a(n_20014), .b(n_20929), .c(n_19906), .o(n_20988) );
ao12s01 g760162 ( .a(n_20052), .b(n_20953), .c(n_19959), .o(n_21102) );
in01f02 g760163 ( .a(n_20461), .o(n_20462) );
in01f02 g760164 ( .a(n_20435), .o(n_20461) );
ao12s01 g760167 ( .a(n_20902), .b(n_20929), .c(n_20901), .o(n_21514) );
in01s01 g760168 ( .a(n_21562), .o(n_21597) );
ao12s01 g760169 ( .a(n_20900), .b(n_20899), .c(n_20898), .o(n_21562) );
no02s02 g760170 ( .a(n_20363), .b(n_20366), .o(n_20434) );
na02m01 g760171 ( .a(n_20334), .b(n_20399), .o(n_20460) );
na02m08 g760172 ( .a(n_20290), .b(n_20227), .o(n_20291) );
in01s01 g760177 ( .a(n_20660), .o(n_20661) );
na02s01 g760178 ( .a(n_19664), .b(n_20456), .o(n_20660) );
no02s01 TIMEBOOST_cell_8514 ( .a(n_38032), .b(n_37945), .o(TIMEBOOST_net_2744) );
in01s02 g760181 ( .a(n_20658), .o(n_20659) );
no02s02 g760182 ( .a(n_20605), .b(n_20567), .o(n_20658) );
in01s01 g760183 ( .a(n_20703), .o(n_20704) );
na02s02 TIMEBOOST_cell_2956 ( .a(FE_RN_773_0), .b(n_1979), .o(TIMEBOOST_net_769) );
na02s03 g760185 ( .a(n_20429), .b(n_19472), .o(n_20712) );
in01s01 g760186 ( .a(n_20744), .o(n_20745) );
na02s01 g760187 ( .a(n_20603), .b(n_20626), .o(n_20744) );
na02s04 g760189 ( .a(n_20288), .b(n_20304), .o(n_20400) );
na02s02 g760191 ( .a(n_20391), .b(n_20433), .o(n_20526) );
no02s01 g760192 ( .a(n_20929), .b(n_20901), .o(n_20902) );
na02s01 g760193 ( .a(n_20954), .b(n_20051), .o(n_21099) );
no02s01 g760194 ( .a(n_20899), .b(n_20898), .o(n_20900) );
oa12m04 g760195 ( .a(n_20896), .b(n_20834), .c(n_20055), .o(n_20897) );
na02s06 TIMEBOOST_cell_4073 ( .a(FE_RN_330_0), .b(FE_RN_331_0), .o(TIMEBOOST_net_1127) );
na02s01 g760197 ( .a(FE_OCP_RBN6791_n_20242), .b(n_20266), .o(n_20603) );
na02s01 g760198 ( .a(FE_OCP_RBN4337_n_20242), .b(FE_OCPN1316_n_20265), .o(n_20626) );
no02s01 g760199 ( .a(FE_OCP_RBN4337_n_20242), .b(n_19414), .o(n_20567) );
na02s02 g760200 ( .a(FE_OCP_RBN6790_n_20242), .b(n_20369), .o(n_20399) );
no02s01 g760201 ( .a(FE_OCP_RBN4335_n_20242), .b(n_19641), .o(n_20366) );
in01s01 g760203 ( .a(n_20334), .o(n_20363) );
na02s02 g760204 ( .a(n_20242), .b(n_19641), .o(n_20334) );
na02s03 g760208 ( .a(n_20242), .b(n_20307), .o(n_20333) );
no02m06 g760212 ( .a(n_20242), .b(n_20307), .o(n_20332) );
in01f02 g760213 ( .a(n_20290), .o(n_20313) );
in01m01 g760214 ( .a(n_20290), .o(n_20270) );
ao12f08 g760215 ( .a(n_20191), .b(n_20171), .c(n_20192), .o(n_20290) );
in01s01 g760216 ( .a(n_20311), .o(n_20269) );
in01m02 g760223 ( .a(n_20289), .o(n_20305) );
no02s06 g760224 ( .a(FE_OCP_RBN1150_n_18981), .b(n_20242), .o(n_20289) );
na02s04 g760225 ( .a(n_20242), .b(n_19134), .o(n_20304) );
na02s02 g760226 ( .a(n_19133), .b(n_20249), .o(n_20288) );
na02f02 g760227 ( .a(n_20285), .b(n_20262), .o(n_20286) );
no02f02 g760228 ( .a(n_20243), .b(n_20244), .o(n_20303) );
in01s01 g760229 ( .a(n_20395), .o(n_20396) );
na02s02 g760230 ( .a(FE_OCP_RBN4335_n_20242), .b(n_19345), .o(n_20395) );
na02s01 g760233 ( .a(FE_OCP_RBN4335_n_20242), .b(n_19346), .o(n_20433) );
na02s01 g760234 ( .a(FE_OCP_RBN6790_n_20242), .b(FE_OCP_RBN5682_n_19177), .o(n_20391) );
na02s03 g760238 ( .a(FE_OCP_RBN4337_n_20242), .b(FE_OCP_RBN3716_n_19241), .o(n_20459) );
na02s06 g760240 ( .a(FE_OCP_RBN6791_n_20242), .b(FE_OCP_RBN3714_n_19241), .o(n_20432) );
na02s02 g760241 ( .a(FE_OCP_RBN4337_n_20242), .b(FE_OCPN1924_n_20430), .o(n_20489) );
no02f06 TIMEBOOST_cell_8509 ( .a(TIMEBOOST_net_2741), .b(TIMEBOOST_net_1219), .o(n_29568) );
na02s02 g760243 ( .a(FE_OCP_RBN6791_n_20242), .b(n_20523), .o(n_20628) );
no02s02 g760245 ( .a(FE_OCP_RBN6791_n_20242), .b(n_20523), .o(n_20565) );
na02s01 g760246 ( .a(FE_OCP_RBN4337_n_20242), .b(n_19497), .o(n_20657) );
no02s01 g760247 ( .a(FE_OCP_RBN6791_n_20242), .b(n_19454), .o(n_20605) );
oa12s01 g760248 ( .a(n_20196), .b(n_20834), .c(n_20234), .o(n_21023) );
oa12s01 g760249 ( .a(n_20896), .b(n_20834), .c(n_20040), .o(n_21050) );
na02s03 g760250 ( .a(n_20242), .b(n_19236), .o(n_20302) );
oa12m06 g760251 ( .a(n_20222), .b(n_20261), .c(n_20186), .o(n_20267) );
na02s03 g760252 ( .a(n_20249), .b(n_19262), .o(n_20473) );
in01s10 g760257 ( .a(FE_OCP_RBN3018_n_20404), .o(n_20429) );
in01s06 g760269 ( .a(FE_OCP_RBN3018_n_20404), .o(n_20456) );
in01s10 g760279 ( .a(n_20372), .o(n_20404) );
in01m08 g760281 ( .a(n_20340), .o(n_20372) );
in01f08 g760282 ( .a(n_20299), .o(n_20340) );
na02s06 g760285 ( .a(FE_OCP_RBN6791_n_20242), .b(n_19347), .o(n_20608) );
na02s06 g760286 ( .a(FE_OCP_RBN4337_n_20242), .b(n_19317), .o(n_20426) );
in01s01 g760290 ( .a(n_20245), .o(n_20275) );
na02s04 TIMEBOOST_cell_5670 ( .a(n_11480), .b(n_11399), .o(TIMEBOOST_net_1783) );
oa12f01 g760292 ( .a(n_20106), .b(n_20081), .c(n_19967), .o(n_20174) );
no02f04 TIMEBOOST_cell_3166 ( .a(n_34795), .b(n_34363), .o(TIMEBOOST_net_874) );
in01s01 g760294 ( .a(n_20518), .o(n_20519) );
no02s01 g760295 ( .a(FE_OCP_RBN4337_n_20242), .b(n_19455), .o(n_20518) );
oa12s01 g760296 ( .a(n_20928), .b(n_20834), .c(n_20927), .o(n_21625) );
in01m02 g760297 ( .a(n_20281), .o(n_20282) );
no02m02 g760298 ( .a(n_20239), .b(n_20264), .o(n_20281) );
in01s01 g760299 ( .a(n_20953), .o(n_20954) );
no02s01 g760300 ( .a(n_20834), .b(n_19933), .o(n_20953) );
na02s01 g760301 ( .a(n_20834), .b(n_20927), .o(n_20928) );
na02f08 g760302 ( .a(n_20081), .b(n_20106), .o(n_20107) );
in01m01 g760304 ( .a(n_20244), .o(n_20262) );
no02f06 g760305 ( .a(FE_OCP_RBN5618_n_18899), .b(n_20228), .o(n_20244) );
in01m01 g760306 ( .a(n_20285), .o(n_20243) );
no02m06 g760308 ( .a(n_20214), .b(n_20125), .o(n_20227) );
no02s03 TIMEBOOST_cell_3915 ( .a(FE_RN_754_0), .b(FE_RN_753_0), .o(TIMEBOOST_net_1048) );
na02s06 TIMEBOOST_cell_7967 ( .a(TIMEBOOST_net_2614), .b(n_43142), .o(n_43369) );
no02m06 TIMEBOOST_cell_3165 ( .a(n_30603), .b(TIMEBOOST_net_873), .o(n_30670) );
ao12s01 g760314 ( .a(n_19989), .b(n_20835), .c(n_20053), .o(n_20929) );
ao12s01 g760315 ( .a(n_20176), .b(n_20835), .c(n_20220), .o(n_20899) );
in01m08 g760331 ( .a(n_20249), .o(n_20242) );
no02f10 g760340 ( .a(n_20153), .b(n_20172), .o(n_20249) );
ao12m02 g760341 ( .a(FE_OCP_RBN5381_n_20123), .b(n_20212), .c(n_20211), .o(n_20226) );
na02f02 g760342 ( .a(n_20213), .b(n_20123), .o(n_20241) );
ao12s01 g760343 ( .a(n_20105), .b(n_20104), .c(n_20103), .o(n_21896) );
in01s01 g760344 ( .a(n_20871), .o(n_21595) );
oa12s01 g760345 ( .a(n_20783), .b(n_20782), .c(n_20781), .o(n_20871) );
in01s01 g760346 ( .a(n_20894), .o(n_20895) );
oa12s01 g760347 ( .a(n_20811), .b(n_20835), .c(n_20810), .o(n_20894) );
no02s04 g760348 ( .a(n_20184), .b(FE_OCPN5101_n_18918), .o(n_20264) );
in01m04 g760349 ( .a(n_20239), .o(n_20240) );
no02f10 g760351 ( .a(FE_OCP_RBN2884_n_20127), .b(FE_OCP_RBN5764_n_19884), .o(n_20172) );
no02m08 g760352 ( .a(n_20127), .b(FE_OCP_RBN5763_n_19884), .o(n_20153) );
na02s01 g760353 ( .a(n_20835), .b(n_20810), .o(n_20811) );
na02s01 g760354 ( .a(n_20782), .b(n_20781), .o(n_20783) );
no02m04 g760355 ( .a(n_20204), .b(n_20161), .o(n_20238) );
no02f06 TIMEBOOST_cell_8821 ( .a(TIMEBOOST_net_2897), .b(n_15501), .o(n_15687) );
na02m02 g760358 ( .a(n_20224), .b(n_20190), .o(n_20236) );
in01m04 g760360 ( .a(n_20214), .o(n_20222) );
no02f06 g760361 ( .a(n_20164), .b(n_18949), .o(n_20214) );
no02f06 g760362 ( .a(n_20165), .b(n_18826), .o(n_20261) );
no02f06 g760363 ( .a(n_20170), .b(n_20160), .o(n_20171) );
na02f08 g760364 ( .a(n_20169), .b(n_20123), .o(n_20192) );
na02f02 g760365 ( .a(n_20212), .b(n_20211), .o(n_20213) );
no02f02 g760367 ( .a(n_20191), .b(n_20170), .o(n_20209) );
no02s01 g760368 ( .a(n_20104), .b(n_20103), .o(n_20105) );
in01s01 g760370 ( .a(n_20081), .o(n_20151) );
ao12f08 g760374 ( .a(n_20004), .b(n_20030), .c(n_19979), .o(n_20081) );
in01f04 g760375 ( .a(n_20207), .o(n_20208) );
na02s02 TIMEBOOST_cell_872 ( .a(TIMEBOOST_net_50), .b(n_17561), .o(n_17680) );
no02m06 g760380 ( .a(n_20740), .b(n_20042), .o(n_20834) );
in01s01 g760381 ( .a(n_20205), .o(n_20206) );
oa12s01 g760382 ( .a(n_20147), .b(FE_OCP_DRV_N3540_n_20146), .c(FE_OCP_DRV_N1761_n_20145), .o(n_20205) );
ao12s01 g760383 ( .a(n_20743), .b(n_20742), .c(n_20741), .o(n_21370) );
in01s01 g760384 ( .a(n_21591), .o(n_20809) );
ao12s01 g760385 ( .a(n_20702), .b(n_20701), .c(n_20700), .o(n_21591) );
na02f06 g760386 ( .a(n_20129), .b(n_20148), .o(n_20228) );
no02f08 g760387 ( .a(n_20149), .b(n_18140), .o(n_20150) );
na02f02 g760388 ( .a(n_20098), .b(FE_OCP_RBN5762_n_19884), .o(n_20129) );
na02m04 g760389 ( .a(FE_OCP_RBN5814_n_20098), .b(n_19884), .o(n_20148) );
no02s01 g760390 ( .a(n_20701), .b(n_20700), .o(n_20702) );
no02s01 g760391 ( .a(n_20742), .b(n_20741), .o(n_20743) );
na02s01 g760392 ( .a(n_20739), .b(n_20041), .o(n_20835) );
in01m02 g760393 ( .a(n_20203), .o(n_20204) );
in01m02 g760394 ( .a(n_20212), .o(n_20203) );
in01m02 g760395 ( .a(n_20169), .o(n_20212) );
na02s01 g760397 ( .a(n_20146), .b(n_20145), .o(n_20147) );
no02s06 g760398 ( .a(n_20167), .b(FE_OCP_RBN7027_n_18866), .o(n_20168) );
na02m02 g760399 ( .a(FE_OCP_RBN7040_n_20167), .b(FE_OCP_RBN7028_n_18866), .o(n_20190) );
na02s08 g760400 ( .a(n_20167), .b(FE_OCP_RBN7027_n_18866), .o(n_20224) );
no02f08 g760401 ( .a(n_20096), .b(FE_OCP_RBN4637_n_18600), .o(n_20191) );
no02m02 g760404 ( .a(n_20186), .b(n_20125), .o(n_20187) );
no02s01 g760405 ( .a(n_20031), .b(n_19919), .o(n_20104) );
na02m04 TIMEBOOST_cell_7077 ( .a(n_10932), .b(n_10931), .o(TIMEBOOST_net_2297) );
no02m06 g760410 ( .a(n_20739), .b(n_20054), .o(n_20740) );
in01f02 g760411 ( .a(n_20164), .o(n_20165) );
na02f04 TIMEBOOST_cell_5310 ( .a(n_39634), .b(FE_RN_1873_0), .o(TIMEBOOST_net_1603) );
oa12s01 g760413 ( .a(n_20034), .b(n_20033), .c(n_20032), .o(n_21788) );
ao12s01 g760414 ( .a(n_19958), .b(n_20655), .c(n_19926), .o(n_20782) );
na02f10 TIMEBOOST_cell_2847 ( .a(n_12623), .b(TIMEBOOST_net_714), .o(n_12753) );
no02f04 TIMEBOOST_cell_4196 ( .a(n_36569), .b(TIMEBOOST_net_1188), .o(TIMEBOOST_net_991) );
na02s06 TIMEBOOST_cell_3913 ( .a(n_33609), .b(n_33215), .o(TIMEBOOST_net_1047) );
no02f08 g760418 ( .a(n_20075), .b(n_20266), .o(n_20149) );
na02m02 g760420 ( .a(n_20079), .b(n_19973), .o(n_20098) );
no02s01 g760421 ( .a(n_20655), .b(n_19988), .o(n_20742) );
in01f02 g760422 ( .a(n_20162), .o(n_20163) );
na02f02 g760423 ( .a(n_20091), .b(n_20144), .o(n_20162) );
na02s02 g760424 ( .a(n_20211), .b(n_20123), .o(n_20183) );
no02m02 g760425 ( .a(FE_OCP_RBN5382_n_20123), .b(n_20160), .o(n_20161) );
na02s01 g760433 ( .a(n_20033), .b(n_20032), .o(n_20034) );
in01s01 g760434 ( .a(n_20030), .o(n_20031) );
na02f08 g760435 ( .a(n_20033), .b(n_19968), .o(n_20030) );
oa12s01 g760436 ( .a(n_20085), .b(n_20624), .c(n_20112), .o(n_20701) );
na02m06 g760437 ( .a(n_20655), .b(n_20013), .o(n_20739) );
in01s01 g760438 ( .a(n_21251), .o(n_20699) );
oa12s01 g760439 ( .a(n_20600), .b(n_20624), .c(n_20599), .o(n_21251) );
oa12s01 g760441 ( .a(n_20074), .b(n_20078), .c(n_20073), .o(n_21790) );
oa12s01 g760442 ( .a(n_20044), .b(n_20078), .c(FE_OCP_RBN5327_FE_RN_2034_0), .o(n_20145) );
oa12s01 g760443 ( .a(n_20560), .b(n_20559), .c(n_20558), .o(n_21481) );
in01m02 g760446 ( .a(n_20095), .o(n_20096) );
in01m02 g760448 ( .a(n_20075), .o(n_20076) );
na02m08 g760449 ( .a(n_20062), .b(n_19718), .o(n_20075) );
na02s06 g760450 ( .a(n_20049), .b(n_19866), .o(n_20079) );
in01m02 g760451 ( .a(n_20064), .o(n_20065) );
no02f06 g760452 ( .a(n_20049), .b(n_19888), .o(n_20064) );
na02s01 g760453 ( .a(n_20624), .b(n_20599), .o(n_20600) );
na02s01 g760454 ( .a(n_20559), .b(n_20558), .o(n_20560) );
na02f06 g760459 ( .a(n_20094), .b(FE_OCPN5270_n_18557), .o(n_20123) );
in01s02 g760460 ( .a(n_20160), .o(n_20211) );
no02f06 g760461 ( .a(n_20094), .b(FE_OCPN5270_n_18557), .o(n_20160) );
na02s01 g760462 ( .a(n_20078), .b(n_20073), .o(n_20074) );
no02s01 g760463 ( .a(n_20093), .b(n_20092), .o(n_20146) );
na02s06 g760464 ( .a(n_20072), .b(FE_OCPN5296_FE_OCP_RBN1105_n_18746), .o(n_20144) );
in01f01 g760465 ( .a(n_20090), .o(n_20091) );
no02f04 g760466 ( .a(n_20072), .b(FE_OCPN5296_FE_OCP_RBN1105_n_18746), .o(n_20090) );
in01f01 g760467 ( .a(n_20046), .o(n_20047) );
no02f01 g760468 ( .a(n_20029), .b(n_20005), .o(n_20046) );
no02s06 g760469 ( .a(n_20005), .b(n_19921), .o(n_20006) );
na02f04 TIMEBOOST_cell_7856 ( .a(n_35341), .b(n_35472), .o(TIMEBOOST_net_2559) );
no02m06 g760471 ( .a(n_20624), .b(n_19982), .o(n_20655) );
ao12s01 g760472 ( .a(n_20514), .b(n_20513), .c(n_20512), .o(n_21371) );
oa12s01 g760473 ( .a(n_20517), .b(n_20516), .c(n_20515), .o(n_21373) );
ao12s01 g760476 ( .a(n_19949), .b(n_19950), .c(n_19948), .o(n_21763) );
ao12f08 g760477 ( .a(n_19887), .b(n_19950), .c(n_19835), .o(n_20033) );
no02f08 g760480 ( .a(n_19972), .b(n_19816), .o(n_20049) );
na02s01 g760481 ( .a(n_20516), .b(n_20515), .o(n_20517) );
no02s06 g760482 ( .a(n_20021), .b(n_18409), .o(n_20092) );
no02f04 g760483 ( .a(n_20020), .b(n_18436), .o(n_20093) );
no02s01 g760484 ( .a(n_19950), .b(n_19948), .o(n_19949) );
no02s01 g760485 ( .a(n_20004), .b(n_19978), .o(n_20103) );
oa12m06 g760486 ( .a(n_19930), .b(n_20423), .c(n_19911), .o(n_20624) );
no02f06 g760487 ( .a(n_19978), .b(n_19919), .o(n_19979) );
no02s01 g760490 ( .a(n_20513), .b(n_20512), .o(n_20514) );
ao12f02 g760492 ( .a(n_19772), .b(n_19976), .c(n_19975), .o(n_20003) );
na02f04 g760493 ( .a(n_19977), .b(n_19773), .o(n_20028) );
na02s04 TIMEBOOST_cell_8082 ( .a(n_45024), .b(FE_OCP_RBN6050_n_21118), .o(TIMEBOOST_net_2672) );
oa12s01 g760495 ( .a(n_19910), .b(n_20451), .c(n_19872), .o(n_20559) );
no02m08 TIMEBOOST_cell_4189 ( .a(n_27308), .b(n_27513), .o(TIMEBOOST_net_1185) );
in01s01 g760498 ( .a(n_20026), .o(n_20078) );
oa12f06 g760499 ( .a(n_19941), .b(n_20007), .c(n_19880), .o(n_20026) );
oa12s01 g760501 ( .a(n_20000), .b(n_19999), .c(n_20007), .o(n_20059) );
in01s02 g760503 ( .a(n_20002), .o(n_20024) );
no02m08 g760504 ( .a(n_19944), .b(n_19685), .o(n_20002) );
na02m08 TIMEBOOST_cell_4188 ( .a(TIMEBOOST_net_1184), .b(FE_RN_1285_0), .o(n_27632) );
na02m04 g760506 ( .a(n_19970), .b(n_19803), .o(n_20001) );
na02f02 g760507 ( .a(n_19976), .b(n_19975), .o(n_19977) );
na02s01 g760508 ( .a(n_20451), .b(n_19821), .o(n_20513) );
na02s01 g760509 ( .a(n_20044), .b(n_19994), .o(n_20073) );
na02s01 g760510 ( .a(n_20007), .b(n_19999), .o(n_20000) );
no02f04 g760512 ( .a(n_19891), .b(n_18397), .o(n_19978) );
no02f06 g760513 ( .a(n_19892), .b(n_18553), .o(n_20004) );
na02s01 g760514 ( .a(n_19946), .b(n_19965), .o(n_20022) );
na02m04 TIMEBOOST_cell_3914 ( .a(n_33610), .b(TIMEBOOST_net_1047), .o(n_33657) );
in01m02 g760516 ( .a(n_19997), .o(n_19998) );
in01m02 g760517 ( .a(n_19972), .o(n_19997) );
ao12f06 g760518 ( .a(n_19842), .b(n_19924), .c(n_19786), .o(n_19972) );
oa12s01 g760519 ( .a(n_20133), .b(n_20450), .c(n_20178), .o(n_20516) );
in01s02 g760520 ( .a(n_20020), .o(n_20021) );
oa12s01 g760522 ( .a(n_19897), .b(n_19896), .c(n_19895), .o(n_21728) );
ao12f08 g760523 ( .a(n_19837), .b(n_19817), .c(n_19775), .o(n_19950) );
in01s01 g760526 ( .a(n_21244), .o(n_20485) );
ao12s01 g760527 ( .a(n_20386), .b(n_20385), .c(n_20384), .o(n_21244) );
ao12s01 g760528 ( .a(n_20425), .b(n_20450), .c(n_20424), .o(n_21405) );
in01m02 g760530 ( .a(n_19976), .o(n_19970) );
no02f06 g760531 ( .a(n_19924), .b(n_19784), .o(n_19976) );
no02s01 g760532 ( .a(n_20450), .b(n_20424), .o(n_20425) );
no02s01 g760533 ( .a(n_20385), .b(n_20384), .o(n_20386) );
in01s01 g760534 ( .a(n_19969), .o(n_20044) );
no02s03 g760535 ( .a(n_19915), .b(FE_OCP_DRV_N1898_n_18287), .o(n_19969) );
na02s01 g760536 ( .a(n_19896), .b(n_19895), .o(n_19897) );
na02s01 g760537 ( .a(n_19936), .b(n_19968), .o(n_20032) );
in01f02 g760540 ( .a(n_19946), .o(n_19967) );
in01f01 g760542 ( .a(n_19921), .o(n_19946) );
no02f04 g760543 ( .a(n_19894), .b(FE_OCP_RBN5028_n_18515), .o(n_19921) );
in01s01 g760545 ( .a(n_19945), .o(n_19965) );
in01m02 g760546 ( .a(n_20106), .o(n_19945) );
na02m04 g760547 ( .a(n_19894), .b(FE_OCP_RBN5028_n_18515), .o(n_20106) );
in01s01 g760548 ( .a(FE_OCP_RBN5327_FE_RN_2034_0), .o(n_19994) );
in01f02 g760550 ( .a(n_19963), .o(n_19964) );
in01f02 g760551 ( .a(n_19944), .o(n_19963) );
no02f08 g760552 ( .a(n_19868), .b(n_19861), .o(n_19944) );
in01m02 g760553 ( .a(n_19942), .o(n_19943) );
in01s01 TIMEBOOST_cell_6855 ( .a(TIMEBOOST_net_2185), .o(mux_while_ln12_psv_q_8_) );
na03f08 TIMEBOOST_cell_5832 ( .a(n_15037), .b(n_15010), .c(FE_OCP_RBN2928_n_14923), .o(n_15208) );
no02m06 g760556 ( .a(n_20450), .b(n_19935), .o(n_20423) );
ao12s01 g760557 ( .a(n_20353), .b(n_20354), .c(n_19934), .o(n_20451) );
ao12s01 g760559 ( .a(n_19940), .b(n_19939), .c(n_19938), .o(n_20018) );
oa12f08 g760560 ( .a(n_19882), .b(n_19854), .c(n_19833), .o(n_20007) );
oa12s01 g760561 ( .a(n_20330), .b(n_20329), .c(n_20328), .o(n_21294) );
ao12s01 g760562 ( .a(n_20357), .b(n_20356), .c(n_20355), .o(n_21249) );
in01m02 g760563 ( .a(n_19891), .o(n_19892) );
na02s04 g760565 ( .a(FE_RN_533_0), .b(n_19696), .o(n_19920) );
ao12f06 g760568 ( .a(n_19418), .b(n_19860), .c(n_19553), .o(n_19868) );
no02s01 TIMEBOOST_cell_6141 ( .a(FE_OCP_RBN5801_n_13962), .b(FE_OCP_RBN2834_n_13962), .o(TIMEBOOST_net_1922) );
na02s03 g760570 ( .a(FE_OCP_RBN5733_n_19806), .b(n_18140), .o(n_19866) );
na02s04 TIMEBOOST_cell_2062 ( .a(n_8885), .b(TIMEBOOST_net_645), .o(n_9010) );
no02s06 TIMEBOOST_cell_8467 ( .a(TIMEBOOST_net_2720), .b(TIMEBOOST_net_2332), .o(n_22613) );
na02f02 g760573 ( .a(n_19862), .b(n_19839), .o(n_19863) );
no02f02 g760574 ( .a(n_19816), .b(n_19888), .o(n_19889) );
na02s01 g760575 ( .a(n_20329), .b(n_20328), .o(n_20330) );
no02s01 g760576 ( .a(n_20356), .b(n_20355), .o(n_20357) );
no02m08 g760577 ( .a(n_20354), .b(n_20353), .o(n_20450) );
na02s01 g760578 ( .a(n_19881), .b(n_19941), .o(n_19999) );
no02s01 g760579 ( .a(n_19939), .b(n_19938), .o(n_19940) );
no02s01 g760580 ( .a(n_19836), .b(n_19887), .o(n_19948) );
in01s01 g760582 ( .a(n_19919), .o(n_19936) );
no02m04 g760583 ( .a(n_19886), .b(FE_OFN795_n_19885), .o(n_19919) );
na02m04 g760584 ( .a(n_19886), .b(FE_OFN795_n_19885), .o(n_19968) );
oa12f06 g760585 ( .a(n_19531), .b(n_19860), .c(n_19451), .o(n_19861) );
na02m06 g760586 ( .a(n_19812), .b(n_19785), .o(n_19842) );
in01m02 g760591 ( .a(n_19818), .o(n_19819) );
oa12f02 g760592 ( .a(n_19502), .b(n_19728), .c(n_19552), .o(n_19818) );
in01s01 g760595 ( .a(FE_OCPUNCON6887_n_19961), .o(n_19962) );
oa12s01 g760596 ( .a(n_19879), .b(n_19878), .c(n_19877), .o(n_19961) );
in01s01 g760597 ( .a(n_19817), .o(n_19895) );
ao12f06 g760598 ( .a(n_19750), .b(n_19701), .c(n_19809), .o(n_19817) );
ao12s01 g760599 ( .a(n_19811), .b(n_19810), .c(n_19809), .o(n_21639) );
oa12s01 g760601 ( .a(n_19852), .b(n_20301), .c(n_19824), .o(n_20385) );
no02m04 g760605 ( .a(n_19754), .b(n_19724), .o(n_19786) );
in01m01 g760607 ( .a(n_19816), .o(n_19839) );
no02f06 g760608 ( .a(n_19783), .b(n_18119), .o(n_19816) );
no02m04 g760609 ( .a(n_19784), .b(n_19703), .o(n_19785) );
no02m06 g760610 ( .a(n_19747), .b(n_18230), .o(n_19859) );
in01m04 g760611 ( .a(n_19862), .o(n_19888) );
na02m06 g760612 ( .a(n_19783), .b(n_18119), .o(n_19862) );
na02m03 g760614 ( .a(n_19778), .b(n_19812), .o(n_19813) );
no02s04 g760615 ( .a(n_19753), .b(n_19779), .o(n_19838) );
na02s01 g760616 ( .a(n_20301), .b(n_19876), .o(n_20356) );
na02s01 g760617 ( .a(n_19834), .b(n_19882), .o(n_19939) );
in01s01 g760618 ( .a(n_19880), .o(n_19881) );
no02m04 g760619 ( .a(n_19856), .b(FE_OCP_DRV_N1896_n_19855), .o(n_19880) );
na02s01 g760620 ( .a(n_19877), .b(n_19878), .o(n_19879) );
na02s04 g760621 ( .a(n_19856), .b(FE_OCP_DRV_N1896_n_19855), .o(n_19941) );
no02s01 g760622 ( .a(n_19776), .b(n_19837), .o(n_19896) );
no02s01 g760623 ( .a(n_19809), .b(n_19810), .o(n_19811) );
in01s01 g760624 ( .a(n_19835), .o(n_19836) );
na02f04 g760625 ( .a(n_19808), .b(FE_OCPUNCON1749_n_19807), .o(n_19835) );
no02s04 g760626 ( .a(n_19808), .b(FE_OCPUNCON1749_n_19807), .o(n_19887) );
no02m08 g760629 ( .a(n_20301), .b(n_19851), .o(n_20354) );
ao12s01 g760630 ( .a(n_20083), .b(n_20277), .c(n_20113), .o(n_20329) );
in01s01 g760631 ( .a(n_19854), .o(n_19938) );
no02m01 TIMEBOOST_cell_6591 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_15_), .o(TIMEBOOST_net_2053) );
no02f06 TIMEBOOST_cell_7791 ( .a(n_34828), .b(TIMEBOOST_net_2526), .o(TIMEBOOST_net_2263) );
in01s01 g760637 ( .a(n_21246), .o(n_20327) );
ao12s01 g760638 ( .a(n_20257), .b(n_20277), .c(n_20256), .o(n_21246) );
no02s02 g760639 ( .a(n_19726), .b(n_19346), .o(n_19755) );
no02s01 TIMEBOOST_cell_7790 ( .a(FE_OFN5086_delay_sub_ln23_0_unr22_stage8_stallmux_q), .b(n_30588), .o(TIMEBOOST_net_2526) );
in01s02 g760641 ( .a(n_19803), .o(n_19804) );
na02s06 g760642 ( .a(n_19975), .b(n_19744), .o(n_19803) );
in01s02 g760643 ( .a(n_19778), .o(n_19779) );
in01m02 g760644 ( .a(n_19754), .o(n_19778) );
no02m06 g760645 ( .a(n_19730), .b(n_18032), .o(n_19754) );
in01s01 g760646 ( .a(n_19812), .o(n_19753) );
na02s06 g760647 ( .a(n_19730), .b(FE_OCPN4528_n_18117), .o(n_19812) );
na02s03 g760648 ( .a(n_19663), .b(n_18119), .o(n_19708) );
no02s01 TIMEBOOST_cell_5192 ( .a(n_2913), .b(FE_OCP_RBN2629_n_2737), .o(TIMEBOOST_net_1544) );
no02s01 g760650 ( .a(n_20277), .b(n_20256), .o(n_20257) );
no02s01 g760651 ( .a(n_19771), .b(n_19740), .o(n_19878) );
in01s01 g760652 ( .a(n_19833), .o(n_19834) );
no02f06 g760653 ( .a(n_19802), .b(FE_OFN1185_n_19801), .o(n_19833) );
no02m06 g760655 ( .a(n_19752), .b(FE_OCP_DRV_N1464_n_19751), .o(n_19837) );
in01s01 g760656 ( .a(n_19775), .o(n_19776) );
na02m06 g760657 ( .a(n_19752), .b(FE_OCP_DRV_N1464_n_19751), .o(n_19775) );
no02s01 g760658 ( .a(FE_OCP_RBN6373_n_19701), .b(n_19750), .o(n_19810) );
na02s06 g760659 ( .a(n_19802), .b(FE_OFN1185_n_19801), .o(n_19882) );
in01s02 g760661 ( .a(n_19774), .o(n_19799) );
no02s01 TIMEBOOST_cell_4079 ( .a(n_4759), .b(n_4875), .o(TIMEBOOST_net_1130) );
no02f04 TIMEBOOST_cell_7056 ( .a(TIMEBOOST_net_2286), .b(n_20064), .o(TIMEBOOST_net_1243) );
in01m02 g760665 ( .a(n_19748), .o(n_19749) );
in01f02 g760666 ( .a(n_19728), .o(n_19748) );
oa12f02 g760667 ( .a(n_19570), .b(n_19673), .c(n_19556), .o(n_19728) );
na02m08 g760668 ( .a(n_20277), .b(n_19829), .o(n_20301) );
na02m04 g760669 ( .a(n_19745), .b(n_19746), .o(n_19856) );
ao12s01 g760670 ( .a(n_19743), .b(n_19742), .c(n_19741), .o(n_21434) );
ao12f06 g760671 ( .a(n_19594), .b(n_19656), .c(n_19719), .o(n_19809) );
na02f06 g760672 ( .a(n_19669), .b(n_19646), .o(n_19783) );
no02s01 TIMEBOOST_cell_5106 ( .a(n_7658), .b(n_7657), .o(TIMEBOOST_net_1501) );
oa12s01 g760675 ( .a(n_19721), .b(n_19720), .c(n_19719), .o(n_21493) );
no03m04 TIMEBOOST_cell_8434 ( .a(n_11283), .b(n_11158), .c(n_11215), .o(n_11285) );
na02s02 g760677 ( .a(n_19690), .b(FE_OCP_RBN2064_n_19353), .o(n_19746) );
na02s02 g760678 ( .a(n_19691), .b(FE_OCP_RBN2062_n_19353), .o(n_19745) );
in01s02 g760680 ( .a(n_19726), .o(n_19725) );
in01m06 g760681 ( .a(n_19707), .o(n_19726) );
na02f08 g760682 ( .a(n_19673), .b(n_19441), .o(n_19707) );
na02f02 g760684 ( .a(n_19635), .b(n_19101), .o(n_19672) );
no03f08 TIMEBOOST_cell_3598 ( .a(TIMEBOOST_net_642), .b(FE_RN_1099_0), .c(FE_RN_1101_0), .o(n_29645) );
no02s06 TIMEBOOST_cell_3883 ( .a(FE_RN_742_0), .b(TIMEBOOST_net_222), .o(TIMEBOOST_net_1032) );
in01s02 g760687 ( .a(n_19772), .o(n_19773) );
in01m02 g760688 ( .a(n_19744), .o(n_19772) );
in01s04 g760689 ( .a(n_19724), .o(n_19744) );
no02m06 g760690 ( .a(n_19634), .b(FE_OCPN1246_n_19645), .o(n_19724) );
na02m06 g760692 ( .a(n_19658), .b(n_19704), .o(n_19722) );
in01s02 g760693 ( .a(n_19703), .o(n_19975) );
no02m04 g760694 ( .a(n_19633), .b(n_19418), .o(n_19703) );
na02m02 g760695 ( .a(n_19601), .b(n_19645), .o(n_19646) );
na02f04 g760696 ( .a(FE_OCP_RBN2720_n_19601), .b(n_18140), .o(n_19669) );
no02s02 TIMEBOOST_cell_1994 ( .a(n_44869), .b(TIMEBOOST_net_611), .o(n_37909) );
na02s02 TIMEBOOST_cell_4549 ( .a(n_32190), .b(n_31840), .o(TIMEBOOST_net_1365) );
in01s01 g760699 ( .a(n_19770), .o(n_19771) );
na02m06 g760700 ( .a(n_19689), .b(n_18112), .o(n_19770) );
no02s01 g760701 ( .a(n_19742), .b(n_19741), .o(n_19743) );
in01s01 g760702 ( .a(n_19739), .o(n_19740) );
na02m04 g760703 ( .a(n_19688), .b(FE_OCP_DRV_N1460_n_18111), .o(n_19739) );
na02s01 g760704 ( .a(n_19719), .b(n_19720), .o(n_19721) );
na02f04 g760706 ( .a(n_19666), .b(FE_OCP_DRV_N1458_n_19665), .o(n_19701) );
no02m04 g760707 ( .a(n_19666), .b(FE_OCP_DRV_N1458_n_19665), .o(n_19750) );
na02s01 g760708 ( .a(FE_OCP_RBN2721_n_19601), .b(n_19587), .o(n_19664) );
no02s01 TIMEBOOST_cell_5210 ( .a(n_34562), .b(n_34563), .o(TIMEBOOST_net_1553) );
na02m04 g760710 ( .a(n_19693), .b(n_19661), .o(n_19738) );
no02s02 g760711 ( .a(n_19736), .b(n_19698), .o(n_19737) );
no02m08 g760712 ( .a(n_20182), .b(n_20181), .o(n_20277) );
no02s03 TIMEBOOST_cell_6620 ( .a(n_32920), .b(TIMEBOOST_net_2067), .o(FE_RN_648_0) );
ao12f04 g760714 ( .a(n_19692), .b(n_19623), .c(n_19555), .o(n_19877) );
no02s06 TIMEBOOST_cell_4164 ( .a(n_32150), .b(TIMEBOOST_net_1172), .o(FE_RN_371_0) );
na02s02 TIMEBOOST_cell_5152 ( .a(n_14125), .b(n_14062), .o(TIMEBOOST_net_1524) );
in01s01 g760721 ( .a(n_21835), .o(n_20255) );
oa12s02 g760722 ( .a(n_20202), .b(n_20201), .c(n_20200), .o(n_21835) );
no02s02 TIMEBOOST_cell_818 ( .a(TIMEBOOST_net_23), .b(n_6745), .o(n_6775) );
no02s01 TIMEBOOST_cell_6961 ( .a(n_47020), .b(n_3231), .o(TIMEBOOST_net_2239) );
no02s06 TIMEBOOST_cell_5209 ( .a(TIMEBOOST_net_1552), .b(FE_OCP_RBN2754_n_3016), .o(n_3128) );
no02s02 g760726 ( .a(n_19588), .b(FE_OCPN1727_n_18099), .o(n_19698) );
na02s02 g760727 ( .a(n_19589), .b(n_18119), .o(n_19661) );
no02s06 TIMEBOOST_cell_4980 ( .a(n_28271), .b(n_28031), .o(TIMEBOOST_net_1438) );
in01s01 g760729 ( .a(n_19695), .o(n_19696) );
in01s02 g760730 ( .a(n_19658), .o(n_19695) );
in01s04 g760731 ( .a(n_19639), .o(n_19658) );
no02m06 g760732 ( .a(n_19605), .b(n_18099), .o(n_19639) );
na02s06 g760733 ( .a(n_19605), .b(n_18099), .o(n_19704) );
na02s04 TIMEBOOST_cell_3036 ( .a(n_24015), .b(n_23971), .o(TIMEBOOST_net_809) );
na02s03 g760735 ( .a(n_19538), .b(FE_OFN738_n_17093), .o(n_19568) );
in01m02 g760737 ( .a(n_19736), .o(n_19693) );
no02m10 g760738 ( .a(n_19589), .b(FE_OCPN4528_n_18117), .o(n_19736) );
no02m06 g760739 ( .a(n_20155), .b(n_20136), .o(n_20182) );
na02s01 g760740 ( .a(n_20201), .b(n_20200), .o(n_20202) );
no02s01 g760741 ( .a(n_19692), .b(n_19624), .o(n_19742) );
no02s01 g760742 ( .a(n_20180), .b(n_20198), .o(n_20199) );
na02s01 g760743 ( .a(n_19595), .b(n_19656), .o(n_19720) );
no02s02 g760744 ( .a(n_19621), .b(n_19618), .o(n_19691) );
na03f08 TIMEBOOST_cell_6545 ( .a(n_39697), .b(n_39694), .c(n_39714), .o(n_39746) );
na02f08 g760747 ( .a(n_19603), .b(n_19322), .o(n_19673) );
in01s02 g760748 ( .a(n_19635), .o(n_19636) );
no02m02 g760749 ( .a(n_19603), .b(n_19362), .o(n_19635) );
oa12m06 g760750 ( .a(n_18119), .b(n_19653), .c(n_19581), .o(n_19718) );
no02s10 TIMEBOOST_cell_846 ( .a(TIMEBOOST_net_37), .b(n_11881), .o(n_11956) );
in01s02 g760752 ( .a(n_19688), .o(n_19689) );
na02m06 TIMEBOOST_cell_8625 ( .a(TIMEBOOST_net_2799), .b(n_10896), .o(n_10998) );
in01m02 g760754 ( .a(n_19633), .o(n_19634) );
in01s01 g760756 ( .a(n_20156), .o(n_20157) );
ao12s01 g760757 ( .a(n_20089), .b(n_20088), .c(n_20087), .o(n_20156) );
oa12f06 g760759 ( .a(n_19465), .b(n_19532), .c(n_19602), .o(n_19719) );
in01s01 g760761 ( .a(FE_OCP_RBN2721_n_19601), .o(n_19654) );
ao12s01 g760769 ( .a(n_19593), .b(n_19592), .c(n_19602), .o(n_21458) );
in01s01 g760770 ( .a(n_19715), .o(n_19716) );
ao12s01 g760771 ( .a(n_19627), .b(n_19626), .c(n_19625), .o(n_19715) );
no02s01 g760772 ( .a(n_20088), .b(n_20087), .o(n_20089) );
no02s01 TIMEBOOST_cell_817 ( .a(n_6716), .b(n_6715), .o(TIMEBOOST_net_23) );
no02f02 g760776 ( .a(n_19512), .b(n_19535), .o(n_19564) );
na02s06 TIMEBOOST_cell_1968 ( .a(TIMEBOOST_net_598), .b(n_37563), .o(n_37583) );
na02m02 g760779 ( .a(n_19615), .b(n_19616), .o(n_19687) );
no02m02 g760780 ( .a(n_19653), .b(n_19685), .o(n_19686) );
no02f04 g760781 ( .a(n_19530), .b(n_19442), .o(n_19570) );
in01s01 g760782 ( .a(n_20155), .o(n_20201) );
na02m06 g760783 ( .a(n_20137), .b(n_19762), .o(n_20155) );
no03s10 TIMEBOOST_cell_845 ( .a(n_11844), .b(n_11882), .c(n_11737), .o(TIMEBOOST_net_37) );
no02f02 g760785 ( .a(n_19591), .b(FE_OCP_DRV_N1454_n_19590), .o(n_19692) );
no02s01 g760786 ( .a(n_19626), .b(n_19625), .o(n_19627) );
in01s01 g760787 ( .a(n_19594), .o(n_19595) );
no02f04 g760788 ( .a(n_19563), .b(FE_OCP_DRV_N1456_n_19562), .o(n_19594) );
na02f04 g760789 ( .a(n_19563), .b(FE_OCP_DRV_N1456_n_19562), .o(n_19656) );
oa12s04 g760790 ( .a(n_18633), .b(FE_OCP_RBN2662_n_19393), .c(n_19478), .o(n_19519) );
na03s04 TIMEBOOST_cell_5798 ( .a(n_3370), .b(FE_OCP_RBN5731_n_4211), .c(n_3376), .o(n_3503) );
no02s01 g760792 ( .a(n_19592), .b(n_19602), .o(n_19593) );
in01s01 g760793 ( .a(n_19623), .o(n_19624) );
na02f02 g760794 ( .a(n_19591), .b(FE_OCP_DRV_N1454_n_19590), .o(n_19623) );
na02f10 g760798 ( .a(n_19537), .b(n_19468), .o(n_19637) );
na02s02 TIMEBOOST_cell_4491 ( .a(n_5805), .b(n_5606), .o(TIMEBOOST_net_1336) );
in01s06 g760802 ( .a(n_19588), .o(n_19589) );
in01m04 g760803 ( .a(n_19561), .o(n_19588) );
in01s01 g760805 ( .a(n_19587), .o(n_20630) );
in01s01 g760806 ( .a(FE_OCP_RBN1827_n_19538), .o(n_19587) );
in01s01 g760809 ( .a(n_20180), .o(n_21169) );
oa12s01 g760810 ( .a(n_20122), .b(n_20121), .c(n_20120), .o(n_20180) );
na03f06 TIMEBOOST_cell_6491 ( .a(n_24446), .b(n_24373), .c(n_24404), .o(n_24471) );
na02s01 g760812 ( .a(n_20121), .b(n_20120), .o(n_20122) );
in01m02 g760813 ( .a(n_19476), .o(n_19477) );
no03s20 TIMEBOOST_cell_6412 ( .a(n_28096), .b(FE_OCPN1400_n_28095), .c(n_28092), .o(n_28117) );
na02m04 g760815 ( .a(n_19435), .b(n_19201), .o(n_19518) );
no02m03 g760816 ( .a(n_19474), .b(n_19202), .o(n_19475) );
in01s02 g760817 ( .a(n_19617), .o(n_19618) );
no02f10 g760821 ( .a(n_19517), .b(n_19469), .o(n_19537) );
na02m02 g760823 ( .a(n_19517), .b(n_19430), .o(n_19535) );
no02f04 TIMEBOOST_cell_4058 ( .a(TIMEBOOST_net_1119), .b(n_20481), .o(n_20621) );
no02s01 TIMEBOOST_cell_8079 ( .a(TIMEBOOST_net_2670), .b(n_36100), .o(n_36246) );
no02m04 g760826 ( .a(n_19533), .b(n_19462), .o(n_19534) );
in01m01 g760827 ( .a(n_19685), .o(n_19616) );
no02m08 g760828 ( .a(n_19585), .b(n_18119), .o(n_19685) );
in01m06 g760831 ( .a(n_19615), .o(n_19653) );
na02s08 g760833 ( .a(n_19585), .b(n_18119), .o(n_19615) );
na02s02 g760835 ( .a(n_20265), .b(n_18140), .o(n_19583) );
na02s01 TIMEBOOST_cell_5034 ( .a(n_37551), .b(n_46416), .o(TIMEBOOST_net_1465) );
no02s01 g760837 ( .a(n_19532), .b(n_19466), .o(n_19592) );
na02s01 g760838 ( .a(FE_OCP_RBN1146_n_19353), .b(FE_OCP_RBN4170_n_19390), .o(n_19472) );
in01f02 g760839 ( .a(n_19441), .o(n_19442) );
ao12f06 g760840 ( .a(n_19565), .b(n_19287), .c(n_18032), .o(n_19441) );
ao12s01 g760841 ( .a(n_20058), .b(n_20057), .c(n_19731), .o(n_20088) );
in01s02 g760842 ( .a(n_19516), .o(n_19566) );
in01s01 g760844 ( .a(n_19530), .o(n_19531) );
na03m04 TIMEBOOST_cell_4734 ( .a(n_9268), .b(n_9330), .c(n_9241), .o(n_9485) );
oa12s01 g760847 ( .a(n_19510), .b(n_19509), .c(n_19508), .o(n_19626) );
in01s01 g760848 ( .a(n_19555), .o(n_19741) );
ao12f08 g760851 ( .a(n_19382), .b(n_19514), .c(n_19422), .o(n_19602) );
na02m04 g760853 ( .a(n_19363), .b(n_18675), .o(n_19470) );
oa12s01 g760854 ( .a(n_19507), .b(n_19506), .c(n_19514), .o(n_21343) );
in01m02 g760855 ( .a(n_19580), .o(n_19581) );
ao22m04 g760856 ( .a(n_19497), .b(FE_OCPN1727_n_18099), .c(n_19453), .d(FE_OCPN1246_n_19645), .o(n_19580) );
in01s01 g760858 ( .a(FE_OCP_RBN1825_n_19513), .o(n_20536) );
no02m06 g760860 ( .a(n_19364), .b(n_19391), .o(n_19513) );
no02m08 g760863 ( .a(n_19365), .b(n_18786), .o(n_19393) );
no02s03 g760864 ( .a(n_19333), .b(n_18540), .o(n_19364) );
no02s04 g760865 ( .a(n_19334), .b(n_18539), .o(n_19391) );
na02s02 g760866 ( .a(n_19365), .b(n_18455), .o(n_19363) );
no02s01 g760867 ( .a(n_20057), .b(n_20069), .o(n_20121) );
in01m01 g760868 ( .a(n_19511), .o(n_19512) );
no02m04 g760869 ( .a(n_19469), .b(n_19324), .o(n_19511) );
no02m06 g760870 ( .a(n_19450), .b(n_19552), .o(n_19553) );
no02m06 g760871 ( .a(n_19467), .b(n_18010), .o(n_19533) );
na02m01 TIMEBOOST_cell_8738 ( .a(FE_OCP_RBN4102_n_12880), .b(n_13916), .o(TIMEBOOST_net_2856) );
na02s06 g760873 ( .a(n_19467), .b(FE_OFN738_n_17093), .o(n_19468) );
na02s01 g760874 ( .a(n_19509), .b(n_19508), .o(n_19510) );
in01s01 g760875 ( .a(n_19465), .o(n_19466) );
na02f04 g760876 ( .a(n_19437), .b(n_19436), .o(n_19465) );
no02f04 g760877 ( .a(n_19437), .b(n_19436), .o(n_19532) );
na02s01 g760878 ( .a(n_19506), .b(n_19514), .o(n_19507) );
in01s01 TIMEBOOST_cell_8886 ( .a(n_1188), .o(TIMEBOOST_net_2930) );
no02m04 TIMEBOOST_cell_7391 ( .a(TIMEBOOST_net_2326), .b(delay_xor_ln22_unr18_stage7_stallmux_q_11_), .o(FE_RN_2015_0) );
in01m02 g760881 ( .a(n_19474), .o(n_19435) );
no03m08 TIMEBOOST_cell_342 ( .a(n_9627), .b(n_9582), .c(n_9507), .o(n_9855) );
na02f06 g760887 ( .a(n_19505), .b(n_19425), .o(n_19556) );
in01s01 g760888 ( .a(n_20198), .o(n_21819) );
oa12s01 g760889 ( .a(n_20119), .b(n_20118), .c(n_20117), .o(n_20198) );
oa12s01 g760890 ( .a(n_19500), .b(n_19499), .c(n_19498), .o(n_21229) );
in01s01 g760891 ( .a(FE_OCP_RBN1823_n_19434), .o(n_20528) );
na03f06 TIMEBOOST_cell_7230 ( .a(FE_OCP_RBN3148_n_15584), .b(n_15538), .c(n_15614), .o(n_15792) );
ao12s01 g760895 ( .a(n_19458), .b(n_19457), .c(n_19456), .o(n_21212) );
in01s02 g760897 ( .a(n_20265), .o(n_20266) );
na02m08 TIMEBOOST_cell_4928 ( .a(n_17865), .b(n_17864), .o(TIMEBOOST_net_1412) );
in01s02 g760899 ( .a(n_19462), .o(n_19463) );
in01s01 g760903 ( .a(FE_OCP_RBN4170_n_19390), .o(n_19461) );
no02m08 g760907 ( .a(n_19284), .b(n_18505), .o(n_19365) );
na02s01 g760908 ( .a(n_20118), .b(n_20117), .o(n_20119) );
in01m04 g760909 ( .a(n_20057), .o(n_20017) );
no02m06 g760910 ( .a(n_20118), .b(n_19993), .o(n_20057) );
no02m08 g760911 ( .a(n_19380), .b(n_17881), .o(n_19469) );
no02f06 TIMEBOOST_cell_6704 ( .a(TIMEBOOST_net_2109), .b(n_15053), .o(n_15108) );
in01f01 g760914 ( .a(n_19388), .o(n_19428) );
na02f06 g760915 ( .a(n_19330), .b(n_19279), .o(n_19388) );
na02m08 g760916 ( .a(n_19414), .b(n_18099), .o(n_19427) );
na02m08 TIMEBOOST_cell_4228 ( .a(n_37609), .b(TIMEBOOST_net_1204), .o(FE_RN_933_0) );
in01s01 g760918 ( .a(n_19501), .o(n_19502) );
no02f06 g760919 ( .a(n_19445), .b(n_17881), .o(n_19501) );
na02m02 g760920 ( .a(n_19313), .b(n_19286), .o(n_19362) );
na02f06 g760921 ( .a(n_19286), .b(n_19285), .o(n_19287) );
no02m04 g760922 ( .a(n_19360), .b(n_19218), .o(n_19438) );
na02s06 g760923 ( .a(n_19360), .b(n_18010), .o(n_19505) );
na02f04 g760924 ( .a(n_19378), .b(n_18010), .o(n_19425) );
no02s06 g760925 ( .a(n_19446), .b(FE_OFN738_n_17093), .o(n_19552) );
no02s02 TIMEBOOST_cell_1996 ( .a(n_44869), .b(TIMEBOOST_net_612), .o(n_37908) );
na02s01 g760927 ( .a(n_19499), .b(n_19498), .o(n_19500) );
no02m04 g760928 ( .a(n_19256), .b(n_18506), .o(n_19335) );
in01s02 g760929 ( .a(n_19333), .o(n_19334) );
no02f02 g760931 ( .a(n_19420), .b(n_19374), .o(n_19423) );
no02s10 TIMEBOOST_cell_1920 ( .a(TIMEBOOST_net_574), .b(FE_OCP_RBN6388_n_32238), .o(n_32324) );
no02s01 g760934 ( .a(n_19457), .b(n_19456), .o(n_19458) );
no02s01 g760935 ( .a(n_19454), .b(n_20523), .o(n_19455) );
na02s01 g760936 ( .a(n_19383), .b(n_19422), .o(n_19506) );
in01f02 g760937 ( .a(n_19386), .o(n_19387) );
in01f02 g760938 ( .a(n_19358), .o(n_19386) );
no02f04 TIMEBOOST_cell_5236 ( .a(FE_OCP_RBN3082_n_15314), .b(n_14452), .o(TIMEBOOST_net_1566) );
no02f02 g760940 ( .a(n_19420), .b(n_19385), .o(n_19421) );
no02s01 g760941 ( .a(n_19350), .b(n_19449), .o(n_19625) );
in01s01 g760944 ( .a(n_19497), .o(n_20124) );
in01m04 g760945 ( .a(n_19453), .o(n_19497) );
na02m06 g760947 ( .a(n_19357), .b(n_19332), .o(n_19453) );
in01s01 g760950 ( .a(n_19419), .o(n_19509) );
in01s03 g760952 ( .a(n_19450), .o(n_19451) );
na02f06 TIMEBOOST_cell_6927 ( .a(n_29030), .b(FE_OFN773_n_25834), .o(TIMEBOOST_net_2222) );
na02s02 g760955 ( .a(n_19327), .b(n_18937), .o(n_19332) );
na02m08 g760956 ( .a(n_19225), .b(n_18460), .o(n_19284) );
na02m04 g760957 ( .a(n_19328), .b(n_18936), .o(n_19357) );
in01m02 g760958 ( .a(n_19255), .o(n_19256) );
no02m04 g760959 ( .a(n_19225), .b(n_18462), .o(n_19255) );
na02s01 TIMEBOOST_cell_2061 ( .a(n_7573), .b(n_7548), .o(TIMEBOOST_net_645) );
no02m06 g760961 ( .a(FE_OCP_RBN1137_n_19270), .b(FE_RN_1458_0), .o(n_19331) );
na02s01 TIMEBOOST_cell_8670 ( .a(n_35684), .b(FE_OCP_RBN3171_n_44211), .o(TIMEBOOST_net_2822) );
na02f04 g760963 ( .a(n_19223), .b(n_19222), .o(n_19286) );
no02s01 g760965 ( .a(n_19374), .b(n_19498), .o(n_19449) );
na02f02 g760966 ( .a(n_19344), .b(FE_OCP_DRV_N1450_n_19384), .o(n_19385) );
in01s02 g760967 ( .a(n_19280), .o(n_19281) );
na03s08 TIMEBOOST_cell_8210 ( .a(FE_RN_2159_0), .b(FE_OCP_RBN2469_n_33034), .c(n_33099), .o(FE_RN_2161_0) );
no02f02 g760969 ( .a(n_19300), .b(n_19350), .o(n_19420) );
na02s01 g760970 ( .a(n_19344), .b(n_19375), .o(n_19499) );
in01s01 g760971 ( .a(n_19382), .o(n_19383) );
no02f06 g760972 ( .a(n_19355), .b(FE_OCPN1212_n_19354), .o(n_19382) );
na02f06 g760974 ( .a(n_19355), .b(FE_OCP_DRV_N1448_n_19354), .o(n_19422) );
no02s01 g760975 ( .a(n_19349), .b(n_19319), .o(n_19457) );
in01s01 g760976 ( .a(n_19416), .o(n_19417) );
no03f08 TIMEBOOST_cell_2217 ( .a(FE_OCP_RBN6542_n_23186), .b(n_23014), .c(n_23122), .o(n_44219) );
no02m04 g760978 ( .a(n_19914), .b(n_19853), .o(n_20118) );
ao12m04 g760979 ( .a(n_19272), .b(n_19278), .c(n_19169), .o(n_19279) );
in01s03 g760980 ( .a(n_19380), .o(n_19381) );
na02s01 TIMEBOOST_cell_2870 ( .a(n_28722), .b(n_28720), .o(TIMEBOOST_net_726) );
oa12f04 g760983 ( .a(n_17881), .b(n_19278), .c(n_19273), .o(n_19330) );
na02m08 g760990 ( .a(n_19250), .b(n_19215), .o(n_19353) );
in01s06 g760992 ( .a(n_19414), .o(n_19454) );
no02s01 TIMEBOOST_cell_5938 ( .a(TIMEBOOST_net_1820), .b(n_22885), .o(TIMEBOOST_net_231) );
in01m02 g760995 ( .a(n_19377), .o(n_19378) );
in01s02 g760997 ( .a(n_19445), .o(n_19446) );
na02s01 TIMEBOOST_cell_2886 ( .a(FE_OCP_RBN2562_n_13084), .b(n_13381), .o(TIMEBOOST_net_734) );
no02s01 TIMEBOOST_cell_6633 ( .a(FE_RN_201_0), .b(n_28460), .o(TIMEBOOST_net_2074) );
no02m04 TIMEBOOST_cell_8147 ( .a(n_18825), .b(TIMEBOOST_net_2704), .o(n_18938) );
no02s06 g761001 ( .a(n_19247), .b(n_18848), .o(n_19329) );
na03s08 TIMEBOOST_cell_2205 ( .a(FE_OCP_RBN2443_n_44798), .b(n_40761), .c(n_40873), .o(n_40853) );
na02f04 TIMEBOOST_cell_8571 ( .a(TIMEBOOST_net_2772), .b(n_29853), .o(n_29947) );
in01s02 g761004 ( .a(n_19327), .o(n_19328) );
no02s06 g761005 ( .a(n_19274), .b(n_18851), .o(n_19327) );
no02s01 g761007 ( .a(n_19273), .b(n_19272), .o(n_19325) );
na02m02 g761008 ( .a(n_19219), .b(n_19170), .o(n_19430) );
in01s01 g761009 ( .a(n_19323), .o(n_19324) );
na02s04 TIMEBOOST_cell_6720 ( .a(TIMEBOOST_net_2117), .b(n_2979), .o(n_3085) );
na02m06 TIMEBOOST_cell_3961 ( .a(FE_RN_1680_0), .b(FE_RN_1681_0), .o(TIMEBOOST_net_1071) );
na02s03 g761015 ( .a(n_19285), .b(n_19218), .o(n_19322) );
in01s01 TIMEBOOST_cell_5910 ( .a(TIMEBOOST_net_1798), .o(TIMEBOOST_net_1799) );
na02s01 TIMEBOOST_cell_6967 ( .a(n_8345), .b(n_8375), .o(TIMEBOOST_net_2242) );
na02m04 TIMEBOOST_cell_2885 ( .a(TIMEBOOST_net_733), .b(n_18110), .o(n_18161) );
na02s01 g761019 ( .a(n_20039), .b(n_19985), .o(n_20055) );
na02s06 g761020 ( .a(n_19178), .b(n_18459), .o(n_19215) );
na02m08 g761021 ( .a(FE_OCP_RBN1817_n_19178), .b(n_18458), .o(n_19250) );
no02s08 g761022 ( .a(n_19184), .b(n_18395), .o(n_19225) );
in01s01 g761024 ( .a(n_19350), .o(n_19375) );
no02f02 g761025 ( .a(n_19315), .b(FE_OCPN1252_n_19314), .o(n_19350) );
in01s01 g761026 ( .a(n_19348), .o(n_19349) );
in01s01 g761028 ( .a(n_19318), .o(n_19319) );
na02s01 g761030 ( .a(n_19346), .b(n_19345), .o(n_19347) );
na02s01 g761031 ( .a(FE_OCP_RBN5668_n_19101), .b(FE_OCP_RBN5679_n_19177), .o(n_19317) );
no02s01 g761032 ( .a(n_19992), .b(n_20010), .o(n_20896) );
in01s02 g761035 ( .a(n_19344), .o(n_19374) );
na02m02 g761036 ( .a(n_19315), .b(FE_OCPN1252_n_19314), .o(n_19344) );
ao12m02 g761037 ( .a(n_19609), .b(n_20115), .c(n_19913), .o(n_19914) );
na02f02 g761038 ( .a(n_19207), .b(n_19182), .o(n_19249) );
no02s06 TIMEBOOST_cell_4931 ( .a(TIMEBOOST_net_1413), .b(n_23387), .o(n_23452) );
in01s02 g761041 ( .a(n_19565), .o(n_19313) );
na02s01 TIMEBOOST_cell_8680 ( .a(n_22134), .b(n_22232), .o(TIMEBOOST_net_2827) );
in01s01 g761051 ( .a(n_19407), .o(n_19408) );
oa12s01 g761052 ( .a(n_19310), .b(n_19309), .c(n_19308), .o(n_19407) );
na02m02 TIMEBOOST_cell_6838 ( .a(TIMEBOOST_net_2176), .b(n_17048), .o(TIMEBOOST_net_1778) );
in01s01 g761054 ( .a(n_19372), .o(n_20523) );
in01m06 g761056 ( .a(n_19342), .o(n_19372) );
na02m08 g761058 ( .a(n_19248), .b(n_19212), .o(n_19342) );
in01s01 g761059 ( .a(n_21454), .o(n_20179) );
oa12s01 g761060 ( .a(n_20116), .b(n_20115), .c(n_20114), .o(n_21454) );
na02f08 g761061 ( .a(n_19089), .b(n_19119), .o(n_19223) );
no02s06 g761062 ( .a(n_19210), .b(n_18820), .o(n_19274) );
na02m06 TIMEBOOST_cell_8083 ( .a(TIMEBOOST_net_2672), .b(FE_RN_579_0), .o(n_21305) );
na02m06 g761064 ( .a(n_19116), .b(n_18428), .o(n_19154) );
na02m08 g761065 ( .a(n_19174), .b(n_18784), .o(n_19248) );
na02s03 g761066 ( .a(n_19173), .b(n_18785), .o(n_19212) );
na02s01 g761067 ( .a(n_20115), .b(n_20114), .o(n_20116) );
in01m02 g761068 ( .a(n_19181), .o(n_19182) );
na02f02 g761069 ( .a(n_19153), .b(n_19044), .o(n_19181) );
na02m04 g761072 ( .a(n_19064), .b(n_17881), .o(n_19089) );
na02f08 g761073 ( .a(n_19641), .b(n_17900), .o(n_19119) );
na02s01 g761074 ( .a(n_19309), .b(n_19308), .o(n_19310) );
in01s04 g761075 ( .a(n_19246), .o(n_19247) );
no02m04 g761077 ( .a(n_19140), .b(FE_OCP_RBN5620_n_18986), .o(n_19180) );
no02f04 TIMEBOOST_cell_5215 ( .a(TIMEBOOST_net_1555), .b(FE_OCP_RBN5967_n_14905), .o(n_15077) );
na02f04 g761079 ( .a(n_19168), .b(n_19056), .o(n_19273) );
ao12s01 g761083 ( .a(n_20016), .b(n_19912), .c(n_19980), .o(n_21101) );
ao12s01 g761084 ( .a(n_19787), .b(n_19766), .c(n_19991), .o(n_19992) );
na02s01 g761085 ( .a(n_19990), .b(n_20041), .o(n_20042) );
in01s01 g761086 ( .a(n_20039), .o(n_20040) );
no02s01 g761087 ( .a(n_19960), .b(n_20016), .o(n_20039) );
in01s06 g761090 ( .a(n_19184), .o(n_19178) );
ao12m10 g761091 ( .a(n_18396), .b(n_19088), .c(n_18394), .o(n_19184) );
in01s01 g761094 ( .a(n_19245), .o(n_19268) );
in01s01 g761095 ( .a(n_19206), .o(n_19245) );
no02m06 g761097 ( .a(n_19115), .b(n_19087), .o(n_19206) );
na02s01 TIMEBOOST_cell_3898 ( .a(TIMEBOOST_net_1039), .b(n_18916), .o(n_20345) );
in01s01 g761100 ( .a(n_19152), .o(n_19456) );
oa12f06 g761101 ( .a(n_19037), .b(n_19081), .c(n_19142), .o(n_19152) );
oa12s01 g761102 ( .a(n_19144), .b(n_19143), .c(n_19142), .o(n_21058) );
in01s01 g761104 ( .a(FE_OCP_RBN5680_n_19177), .o(n_19346) );
in01s01 g761118 ( .a(n_19301), .o(n_20430) );
in01s06 g761119 ( .a(n_19264), .o(n_19301) );
no02f08 TIMEBOOST_cell_8073 ( .a(TIMEBOOST_net_2667), .b(TIMEBOOST_net_663), .o(n_20763) );
in01s01 g761123 ( .a(n_19300), .o(n_19498) );
ao12f02 g761124 ( .a(n_19237), .b(n_19200), .c(n_19166), .o(n_19300) );
no02m08 g761126 ( .a(n_19146), .b(n_19171), .o(n_19285) );
in01s01 g761129 ( .a(n_19238), .o(n_20343) );
in01s01 g761130 ( .a(n_19203), .o(n_19238) );
in01s01 g761131 ( .a(n_19219), .o(n_19203) );
no02m08 g761135 ( .a(n_19106), .b(n_18707), .o(n_19175) );
no02m02 TIMEBOOST_cell_8559 ( .a(TIMEBOOST_net_2766), .b(n_3244), .o(n_3328) );
in01s03 g761137 ( .a(n_19173), .o(n_19174) );
no02s06 g761138 ( .a(n_19150), .b(n_18821), .o(n_19173) );
na02s08 g761139 ( .a(n_19150), .b(n_18742), .o(n_19210) );
no02m04 g761140 ( .a(FE_OCP_RBN5034_n_19062), .b(n_18391), .o(n_19115) );
no02s04 g761141 ( .a(n_19062), .b(n_18392), .o(n_19087) );
no02m04 g761142 ( .a(n_19797), .b(n_19714), .o(n_20115) );
no02s02 g761143 ( .a(n_19798), .b(n_19913), .o(n_19853) );
in01s02 g761144 ( .a(n_19201), .o(n_19202) );
in01s02 g761145 ( .a(n_19172), .o(n_19201) );
no02m04 g761146 ( .a(n_19148), .b(n_17900), .o(n_19172) );
na02m08 TIMEBOOST_cell_4986 ( .a(n_12293), .b(FE_RN_403_0), .o(TIMEBOOST_net_1441) );
no02m02 g761149 ( .a(n_19058), .b(FE_OCP_RBN4081_n_18899), .o(n_19147) );
no02s01 TIMEBOOST_cell_2803 ( .a(TIMEBOOST_net_692), .b(n_1512), .o(n_1597) );
no02m04 g761151 ( .a(n_19101), .b(n_17900), .o(n_19146) );
no02m08 g761152 ( .a(FE_OCP_RBN5665_n_19101), .b(n_19170), .o(n_19171) );
in01s01 TIMEBOOST_cell_8903 ( .a(TIMEBOOST_net_2946), .o(TIMEBOOST_net_2947) );
no02s01 g761154 ( .a(n_19912), .b(n_19845), .o(n_20016) );
no02s01 g761155 ( .a(n_19237), .b(n_19167), .o(n_19309) );
na02s01 g761156 ( .a(n_19133), .b(FE_OCP_RBN7033_n_18981), .o(n_19236) );
na02s01 g761157 ( .a(n_19134), .b(FE_OCP_RBN7035_n_18981), .o(n_19262) );
na02s01 g761158 ( .a(n_19143), .b(n_19142), .o(n_19144) );
ao12s01 g761159 ( .a(n_19989), .b(n_19907), .c(n_19845), .o(n_19990) );
in01m02 g761160 ( .a(n_19168), .o(n_19169) );
oa12m04 g761162 ( .a(n_17783), .b(n_18987), .c(n_19006), .o(n_19153) );
in01s02 g761163 ( .a(n_19140), .o(n_19141) );
in01m02 g761164 ( .a(n_19112), .o(n_19140) );
na02f08 g761165 ( .a(n_19046), .b(n_19058), .o(n_19112) );
na02s01 g761166 ( .a(n_20053), .b(n_20015), .o(n_20054) );
ao12s01 g761167 ( .a(n_19188), .b(n_19187), .c(n_19186), .o(n_21007) );
in01s01 g761168 ( .a(n_21105), .o(n_21134) );
ao12s01 g761169 ( .a(n_19768), .b(n_19769), .c(n_19767), .o(n_21105) );
ao12s01 g761170 ( .a(n_19084), .b(n_19083), .c(n_19082), .o(n_21028) );
in01s01 g761175 ( .a(n_19641), .o(n_20369) );
in01f06 g761176 ( .a(n_19064), .o(n_19641) );
oa12m04 g761181 ( .a(n_18310), .b(FE_OCP_RBN5033_n_18951), .c(n_18339), .o(n_19062) );
no02s08 g761182 ( .a(n_19080), .b(n_18674), .o(n_19150) );
in01s01 g761183 ( .a(n_19797), .o(n_19798) );
no02m04 g761184 ( .a(n_19769), .b(n_19713), .o(n_19797) );
no02s01 g761185 ( .a(n_19769), .b(n_19767), .o(n_19768) );
na02f04 g761186 ( .a(n_19005), .b(n_17815), .o(n_19046) );
no03f04 TIMEBOOST_cell_4794 ( .a(FE_RN_1104_0), .b(FE_OCP_RBN6036_n_10399), .c(FE_OCPN1066_n_44461), .o(n_10582) );
na02m02 g761189 ( .a(FE_OCP_RBN5621_n_18986), .b(n_17783), .o(n_19044) );
na02s01 g761190 ( .a(n_20051), .b(n_19991), .o(n_20052) );
no02s01 g761191 ( .a(n_20050), .b(n_20009), .o(n_21019) );
no02s01 g761192 ( .a(n_20014), .b(n_19957), .o(n_20015) );
na02s01 g761193 ( .a(n_19932), .b(n_19959), .o(n_19960) );
na02s01 g761194 ( .a(n_19991), .b(n_19959), .o(n_21098) );
no02s01 g761195 ( .a(n_19186), .b(n_19187), .o(n_19188) );
in01s01 g761196 ( .a(n_19166), .o(n_19167) );
na02s02 g761197 ( .a(n_19139), .b(FE_OCP_DRV_N1444_n_19138), .o(n_19166) );
no02s01 g761198 ( .a(n_19083), .b(n_19082), .o(n_19084) );
no02s01 g761199 ( .a(n_19038), .b(n_19081), .o(n_19143) );
na02m06 g761201 ( .a(n_18989), .b(n_18511), .o(n_19060) );
in01m04 g761202 ( .a(n_19107), .o(n_19108) );
na03m08 TIMEBOOST_cell_7286 ( .a(n_21291), .b(n_45072), .c(n_21281), .o(n_21475) );
in01m04 g761204 ( .a(n_19105), .o(n_19106) );
ao12s01 g761206 ( .a(n_19988), .b(n_19904), .c(n_19845), .o(n_20041) );
na02s02 g761207 ( .a(n_19832), .b(n_19876), .o(n_20353) );
no02m02 g761208 ( .a(n_19139), .b(FE_OCP_DRV_N1444_n_19138), .o(n_19237) );
oa12s02 g761209 ( .a(n_18298), .b(FE_OCP_RBN5032_n_18951), .c(n_19014), .o(n_19041) );
na02m06 TIMEBOOST_cell_8533 ( .a(TIMEBOOST_net_2753), .b(n_41812), .o(n_41858) );
na02m04 TIMEBOOST_cell_8809 ( .a(TIMEBOOST_net_2891), .b(n_10894), .o(n_10965) );
in01m01 g761213 ( .a(n_19104), .o(n_19135) );
ao12f04 g761214 ( .a(n_18945), .b(n_19025), .c(FE_OFN739_n_17093), .o(n_19104) );
in01m01 g761216 ( .a(n_19058), .o(n_19078) );
no02s01 TIMEBOOST_cell_1923 ( .a(n_11581), .b(n_11405), .o(TIMEBOOST_net_576) );
ao12s01 g761218 ( .a(n_20050), .b(n_20011), .c(n_19980), .o(n_21137) );
ao12s01 g761219 ( .a(n_19984), .b(n_20036), .c(n_19980), .o(n_21140) );
oa12s01 g761220 ( .a(n_19956), .b(n_19931), .c(n_20086), .o(n_20987) );
ao12s01 g761221 ( .a(n_19787), .b(n_19712), .c(n_19986), .o(n_20037) );
na02s02 TIMEBOOST_cell_4519 ( .a(n_11242), .b(n_11156), .o(TIMEBOOST_net_1350) );
in01s01 g761229 ( .a(n_19200), .o(n_19308) );
oa12f04 g761230 ( .a(n_19072), .b(n_19186), .c(n_19130), .o(n_19200) );
in01s03 g761231 ( .a(n_19133), .o(n_19134) );
in01s04 g761236 ( .a(n_19134), .o(n_19164) );
in01s02 g761238 ( .a(n_19148), .o(n_19133) );
ao12f06 g761240 ( .a(n_19035), .b(n_18980), .c(n_18984), .o(n_19142) );
in01s01 g761244 ( .a(FE_OCP_RBN5667_n_19101), .o(n_19345) );
no02s04 TIMEBOOST_cell_2050 ( .a(TIMEBOOST_net_639), .b(n_3377), .o(n_4905) );
in01s01 g761248 ( .a(n_19912), .o(n_19766) );
oa12s01 g761249 ( .a(n_19682), .b(n_19681), .c(n_19680), .o(n_19912) );
oa12s01 g761250 ( .a(n_19765), .b(n_19764), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_21052) );
in01s02 g761251 ( .a(n_19075), .o(n_19076) );
no02m06 TIMEBOOST_cell_1914 ( .a(TIMEBOOST_net_571), .b(n_11535), .o(n_11726) );
no02s02 g761254 ( .a(n_18951), .b(n_18324), .o(n_18990) );
na03s04 TIMEBOOST_cell_8178 ( .a(n_17560), .b(n_17458), .c(n_17593), .o(TIMEBOOST_net_50) );
no02m02 TIMEBOOST_cell_6625 ( .a(FE_RN_132_0), .b(n_12581), .o(TIMEBOOST_net_2070) );
na02s04 g761257 ( .a(n_18952), .b(n_18512), .o(n_18989) );
na02s01 g761258 ( .a(n_19764), .b(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_19765) );
na02m02 g761260 ( .a(n_19055), .b(n_17783), .o(n_19056) );
no02f06 TIMEBOOST_cell_8037 ( .a(TIMEBOOST_net_2649), .b(FE_RN_1380_0), .o(n_31207) );
na02s01 g761262 ( .a(n_19681), .b(n_19680), .o(n_19682) );
na02s01 g761263 ( .a(n_19910), .b(n_19909), .o(n_19911) );
na02s01 g761264 ( .a(n_19902), .b(n_19903), .o(n_19958) );
na02s01 g761265 ( .a(n_19934), .b(n_19905), .o(n_19935) );
no02s01 g761266 ( .a(n_19953), .b(n_20012), .o(n_20013) );
in01s01 g761267 ( .a(n_19932), .o(n_19933) );
no02s01 g761268 ( .a(n_19847), .b(n_20234), .o(n_19932) );
na02s01 g761269 ( .a(n_19679), .b(n_19845), .o(n_19991) );
na02s01 g761270 ( .a(n_19678), .b(n_19787), .o(n_19959) );
no02s01 g761271 ( .a(n_19875), .b(n_20014), .o(n_20901) );
in01s01 g761272 ( .a(n_19956), .o(n_19957) );
na02s01 g761273 ( .a(n_19931), .b(n_19787), .o(n_19956) );
in01s01 g761274 ( .a(n_19984), .o(n_19985) );
no02s01 g761275 ( .a(n_20036), .b(n_19845), .o(n_19984) );
no02s01 g761276 ( .a(n_20011), .b(n_19980), .o(n_20050) );
na02s01 g761277 ( .a(n_19906), .b(n_19931), .o(n_19907) );
no02f08 TIMEBOOST_cell_1894 ( .a(n_36015), .b(TIMEBOOST_net_561), .o(n_36208) );
no02s01 g761279 ( .a(n_19130), .b(n_19073), .o(n_19187) );
in01m04 g761280 ( .a(n_18955), .o(n_18956) );
ao12m08 g761281 ( .a(n_18473), .b(n_18832), .c(n_47246), .o(n_18955) );
no02f03 g761282 ( .a(n_19011), .b(FE_OCP_DRV_N1440_n_19010), .o(n_19081) );
in01s01 g761283 ( .a(n_19037), .o(n_19038) );
na02s03 g761284 ( .a(n_19011), .b(FE_OCP_DRV_N1440_n_19010), .o(n_19037) );
na02f02 TIMEBOOST_cell_6691 ( .a(n_14160), .b(n_14203), .o(TIMEBOOST_net_2103) );
no02s01 g761287 ( .a(n_19035), .b(n_18985), .o(n_19083) );
na02m10 g761288 ( .a(FE_OCP_RBN7037_n_18982), .b(n_18550), .o(n_19080) );
ao12f02 g761289 ( .a(n_19651), .b(n_19709), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_19769) );
ao12s01 g761290 ( .a(n_20012), .b(n_19952), .c(n_19980), .o(n_20781) );
oa12s01 g761291 ( .a(n_19846), .b(n_19983), .c(n_20086), .o(n_21022) );
in01s01 g761292 ( .a(n_20010), .o(n_20051) );
ao12s01 g761293 ( .a(n_19787), .b(n_19983), .c(n_19571), .o(n_20010) );
oa12s01 g761294 ( .a(n_19649), .b(n_19830), .c(n_19337), .o(n_19832) );
no02s01 TIMEBOOST_cell_4051 ( .a(n_25390), .b(n_25327), .o(TIMEBOOST_net_1116) );
oa12s01 g761296 ( .a(n_19129), .b(n_19128), .c(n_19127), .o(n_20885) );
in01s01 g761297 ( .a(n_19033), .o(n_20307) );
in01m04 g761298 ( .a(n_19008), .o(n_19033) );
no02m06 g761300 ( .a(n_18925), .b(n_18901), .o(n_19008) );
in01s01 g761303 ( .a(FE_OCP_RBN5621_n_18986), .o(n_19032) );
in01s01 g761306 ( .a(n_19098), .o(n_19099) );
ao12s01 g761307 ( .a(n_19029), .b(n_19028), .c(n_19027), .o(n_19098) );
in01m02 g761308 ( .a(n_19005), .o(n_19006) );
no03s04 TIMEBOOST_cell_5785 ( .a(TIMEBOOST_net_1554), .b(FE_OCP_RBN2753_n_3016), .c(n_3271), .o(n_3375) );
na02m01 g761312 ( .a(n_18945), .b(n_18918), .o(n_19030) );
no02f04 TIMEBOOST_cell_4050 ( .a(TIMEBOOST_net_1115), .b(n_25042), .o(n_25106) );
no02s01 g761314 ( .a(n_19828), .b(n_19792), .o(n_19829) );
no02s01 g761315 ( .a(n_19789), .b(n_19830), .o(n_19852) );
no02s01 g761316 ( .a(n_19899), .b(n_19954), .o(n_20053) );
na02s01 g761317 ( .a(n_19981), .b(n_19901), .o(n_19982) );
no02s01 g761318 ( .a(n_19827), .b(n_20178), .o(n_19934) );
na02s02 g761319 ( .a(n_19710), .b(n_19731), .o(n_19732) );
na02s01 g761320 ( .a(n_19849), .b(n_19850), .o(n_19851) );
no02s01 g761321 ( .a(n_19820), .b(n_19822), .o(n_19910) );
no02s01 g761322 ( .a(n_19848), .b(n_19845), .o(n_20014) );
na02s01 g761323 ( .a(n_20177), .b(n_20220), .o(n_20810) );
no02s01 g761324 ( .a(n_19714), .b(n_19713), .o(n_19767) );
na02s01 g761325 ( .a(n_19905), .b(n_19823), .o(n_20512) );
no02s01 g761326 ( .a(n_19953), .b(n_19871), .o(n_20741) );
no02s01 g761327 ( .a(n_20197), .b(n_20234), .o(n_20927) );
na02s01 g761328 ( .a(n_19849), .b(n_19763), .o(n_20355) );
no02s01 g761329 ( .a(n_19761), .b(n_19711), .o(n_20087) );
no02s01 g761330 ( .a(n_19952), .b(n_19845), .o(n_20012) );
na02s01 g761331 ( .a(n_19709), .b(n_19652), .o(n_19764) );
na02s01 g761332 ( .a(n_20082), .b(n_20113), .o(n_20256) );
in01s01 g761333 ( .a(n_19906), .o(n_19875) );
na02s01 g761334 ( .a(n_19848), .b(n_19845), .o(n_19906) );
na02s01 g761335 ( .a(n_19903), .b(n_19648), .o(n_19904) );
in01s01 g761336 ( .a(n_19846), .o(n_19847) );
na02s01 g761337 ( .a(n_19983), .b(n_19649), .o(n_19846) );
no02s01 g761338 ( .a(n_20069), .b(n_19993), .o(n_20117) );
no02s01 g761339 ( .a(n_20134), .b(n_20178), .o(n_20424) );
no02s01 g761340 ( .a(n_20084), .b(n_20112), .o(n_20599) );
na02s01 g761341 ( .a(n_20219), .b(n_20254), .o(n_21020) );
na02s01 g761342 ( .a(n_19909), .b(n_19930), .o(n_20558) );
in01s02 g761343 ( .a(n_19002), .o(n_19003) );
in01s01 g761345 ( .a(n_18984), .o(n_18985) );
na02f04 g761346 ( .a(n_18954), .b(n_18953), .o(n_18984) );
no02f04 g761347 ( .a(n_18954), .b(n_18953), .o(n_19035) );
in01m06 g761350 ( .a(n_18952), .o(n_18982) );
ao12m06 g761351 ( .a(n_18478), .b(FE_OCP_RBN4068_n_18829), .c(n_18516), .o(n_18952) );
no02s01 g761352 ( .a(n_19028), .b(n_19027), .o(n_19029) );
na02s01 g761353 ( .a(n_19128), .b(n_19127), .o(n_19129) );
in01s01 g761354 ( .a(n_19072), .o(n_19073) );
na02f02 g761355 ( .a(n_19054), .b(FE_OCP_DRV_N3536_n_19053), .o(n_19072) );
no02f02 g761356 ( .a(n_19054), .b(FE_OCP_DRV_N3536_n_19053), .o(n_19130) );
ao12s01 g761360 ( .a(n_18765), .b(n_19613), .c(n_18841), .o(n_19681) );
ao12s01 g761361 ( .a(n_19676), .b(n_20086), .c(n_19650), .o(n_20120) );
ao12s01 g761362 ( .a(n_19954), .b(n_19980), .c(n_19900), .o(n_20898) );
oa12s01 g761363 ( .a(n_19981), .b(n_20086), .c(n_19927), .o(n_20700) );
oa12s01 g761364 ( .a(n_19826), .b(n_19980), .c(n_19793), .o(n_20515) );
oa12s01 g761365 ( .a(n_19850), .b(n_19980), .c(n_19796), .o(n_20384) );
ao12s01 g761366 ( .a(n_19828), .b(n_20086), .c(n_19760), .o(n_20328) );
ao12s01 g761367 ( .a(n_19787), .b(n_19607), .c(n_19928), .o(n_19989) );
in01s01 g761368 ( .a(n_19988), .o(n_19902) );
ao12s01 g761369 ( .a(n_19787), .b(n_19927), .c(n_19873), .o(n_19988) );
no02f06 g761370 ( .a(n_19024), .b(n_19022), .o(n_19186) );
in01s01 g761375 ( .a(n_19712), .o(n_20011) );
ao12s01 g761376 ( .a(n_19612), .b(n_19611), .c(n_19610), .o(n_19712) );
no02s06 TIMEBOOST_cell_1961 ( .a(n_37040), .b(FE_RN_284_0), .o(TIMEBOOST_net_595) );
in01s01 g761384 ( .a(n_18980), .o(n_19082) );
oa12f06 g761385 ( .a(n_18863), .b(n_18862), .c(n_18948), .o(n_18980) );
ao22s01 g761386 ( .a(n_19787), .b(n_18886), .c(n_19980), .d(n_19913), .o(n_20114) );
oa12s01 g761387 ( .a(n_19579), .b(n_19578), .c(n_19577), .o(n_20036) );
in01s01 g761388 ( .a(n_19678), .o(n_19679) );
ao12s01 g761389 ( .a(n_19576), .b(n_19613), .c(n_19575), .o(n_19678) );
ao12s01 g761390 ( .a(n_19574), .b(n_19573), .c(n_19572), .o(n_19931) );
ao22s01 g761391 ( .a(n_20086), .b(n_20136), .c(n_19980), .d(n_20135), .o(n_20200) );
in01s01 g761392 ( .a(n_19025), .o(n_19026) );
na02f08 g761394 ( .a(n_18875), .b(n_18831), .o(n_18987) );
na03m06 TIMEBOOST_cell_6553 ( .a(n_10694), .b(n_10737), .c(TIMEBOOST_net_1694), .o(n_10902) );
na02f04 g761434 ( .a(n_18829), .b(n_18370), .o(n_18876) );
na03s01 TIMEBOOST_cell_7302 ( .a(n_39956), .b(n_39858), .c(n_40085), .o(n_40161) );
na02m06 g761436 ( .a(n_18799), .b(n_18710), .o(n_18832) );
na03s08 TIMEBOOST_cell_7140 ( .a(n_28458), .b(n_28525), .c(n_28632), .o(n_28651) );
na02m04 g761439 ( .a(n_18797), .b(FE_OFN737_n_17093), .o(n_18831) );
na02f06 g761440 ( .a(n_17661), .b(n_18761), .o(n_18875) );
na02s01 g761441 ( .a(n_19578), .b(n_19577), .o(n_19579) );
no02s01 g761442 ( .a(n_19611), .b(n_19610), .o(n_19612) );
in01s01 g761443 ( .a(n_20176), .o(n_20177) );
no02s01 g761444 ( .a(n_20086), .b(n_19928), .o(n_20176) );
na02s01 g761445 ( .a(n_19787), .b(n_19927), .o(n_19981) );
in01s01 g761446 ( .a(n_20218), .o(n_20219) );
no02s01 g761447 ( .a(n_20086), .b(n_19986), .o(n_20218) );
in01s01 g761448 ( .a(n_19901), .o(n_20112) );
na02s01 g761449 ( .a(n_19787), .b(n_19873), .o(n_19901) );
in01s01 g761450 ( .a(n_20084), .o(n_20085) );
no02s01 g761451 ( .a(n_20086), .b(n_19873), .o(n_20084) );
in01s01 g761452 ( .a(n_20133), .o(n_20134) );
na02s01 g761453 ( .a(n_20086), .b(n_19825), .o(n_20133) );
no02s02 g761454 ( .a(n_19609), .b(n_18778), .o(n_19714) );
in01s01 g761455 ( .a(n_19710), .o(n_19711) );
na02s01 g761456 ( .a(n_19647), .b(n_19677), .o(n_19710) );
na02s01 g761457 ( .a(n_19647), .b(n_19796), .o(n_19850) );
in01s01 g761458 ( .a(n_19651), .o(n_19652) );
no02s02 g761459 ( .a(n_19609), .b(n_19608), .o(n_19651) );
in01s01 g761460 ( .a(n_19830), .o(n_19763) );
no02s01 g761461 ( .a(n_19647), .b(n_19735), .o(n_19830) );
na02m04 g761462 ( .a(n_19609), .b(n_19608), .o(n_19709) );
no02s01 g761463 ( .a(n_19647), .b(n_19794), .o(n_20234) );
in01s01 g761464 ( .a(n_19905), .o(n_19872) );
na02s01 g761465 ( .a(n_19647), .b(n_19790), .o(n_19905) );
na02s01 g761466 ( .a(n_19845), .b(n_19398), .o(n_19909) );
in01s01 g761467 ( .a(n_20254), .o(n_20009) );
na02s01 g761468 ( .a(n_19986), .b(n_19787), .o(n_20254) );
in01s01 g761469 ( .a(n_20196), .o(n_20197) );
na02s01 g761470 ( .a(n_19980), .b(n_19794), .o(n_20196) );
in01s01 g761471 ( .a(n_19761), .o(n_19762) );
no02s01 g761472 ( .a(n_19647), .b(n_19677), .o(n_19761) );
in01s01 g761473 ( .a(n_19953), .o(n_19926) );
no02s01 g761474 ( .a(n_19845), .b(n_19844), .o(n_19953) );
in01s01 g761475 ( .a(n_19903), .o(n_19871) );
na02s01 g761476 ( .a(n_19845), .b(n_19844), .o(n_19903) );
no02s01 g761477 ( .a(n_19845), .b(n_19900), .o(n_19954) );
in01s01 g761478 ( .a(n_19826), .o(n_19827) );
na02s01 g761479 ( .a(n_19647), .b(n_19793), .o(n_19826) );
no02s01 g761480 ( .a(n_19649), .b(n_19825), .o(n_20178) );
no02s01 g761481 ( .a(n_19649), .b(n_19760), .o(n_19828) );
in01s01 g761482 ( .a(n_19792), .o(n_20113) );
no02s01 g761483 ( .a(n_19649), .b(n_19758), .o(n_19792) );
in01s01 g761484 ( .a(n_19676), .o(n_19731) );
no02s01 g761485 ( .a(n_19649), .b(n_19650), .o(n_19676) );
no02s01 g761486 ( .a(n_19649), .b(n_18935), .o(n_19993) );
no02s02 g761487 ( .a(n_19569), .b(n_18777), .o(n_19713) );
in01s01 g761488 ( .a(n_19849), .o(n_19824) );
na02s01 g761489 ( .a(n_19647), .b(n_19735), .o(n_19849) );
in01s01 g761490 ( .a(n_19822), .o(n_19823) );
no02s01 g761491 ( .a(n_19647), .b(n_19790), .o(n_19822) );
na02s02 g761492 ( .a(n_19787), .b(n_19399), .o(n_19930) );
no02s01 g761493 ( .a(n_19980), .b(n_19733), .o(n_20069) );
in01s01 g761494 ( .a(n_20082), .o(n_20083) );
na02s01 g761495 ( .a(n_20086), .b(n_19758), .o(n_20082) );
in01s01 g761496 ( .a(n_20220), .o(n_19899) );
na02s01 g761497 ( .a(n_19928), .b(n_19787), .o(n_20220) );
no02s01 g761498 ( .a(n_19613), .b(n_19575), .o(n_19576) );
no02f04 g761499 ( .a(n_18971), .b(n_18996), .o(n_19024) );
oa12m04 g761501 ( .a(n_18434), .b(FE_OCP_RBN6371_FE_RN_1425_0), .c(n_18346), .o(n_18873) );
no02s01 g761502 ( .a(n_19573), .b(n_19572), .o(n_19574) );
na02s01 g761503 ( .a(n_18997), .b(n_19023), .o(n_19128) );
no02s04 TIMEBOOST_cell_1953 ( .a(FE_OCPN1653_n_23078), .b(n_22972), .o(TIMEBOOST_net_591) );
in01s01 g761506 ( .a(n_18945), .o(n_18978) );
in01s01 g761508 ( .a(n_19820), .o(n_19821) );
ao12s01 g761509 ( .a(n_19647), .b(n_19793), .c(n_19291), .o(n_19820) );
in01s01 g761510 ( .a(n_19876), .o(n_19789) );
oa12s01 g761511 ( .a(n_19649), .b(n_19760), .c(n_19758), .o(n_19876) );
ao12s01 g761512 ( .a(n_19647), .b(n_19051), .c(n_19733), .o(n_20058) );
na03s02 TIMEBOOST_cell_4605 ( .a(FE_RN_1580_0), .b(FE_OCP_RBN2478_n_1862), .c(n_1851), .o(n_1915) );
ao12s01 g761514 ( .a(n_19000), .b(n_18999), .c(n_18998), .o(n_20852) );
no02f06 g761521 ( .a(n_18801), .b(n_18760), .o(n_18899) );
no02m04 g761522 ( .a(n_18828), .b(n_18798), .o(n_18954) );
ao12s01 g761523 ( .a(n_18920), .b(n_18948), .c(n_18919), .o(n_19028) );
in01s01 g761524 ( .a(n_18974), .o(n_20876) );
oa12s01 g761525 ( .a(n_18896), .b(n_18895), .c(n_18894), .o(n_18974) );
ao12s01 g761526 ( .a(n_19549), .b(n_19548), .c(n_19547), .o(n_19983) );
oa12s01 g761527 ( .a(n_19546), .b(n_19545), .c(n_19544), .o(n_19848) );
in01s01 g761528 ( .a(n_19648), .o(n_19952) );
ao12s01 g761529 ( .a(n_19543), .b(n_19542), .c(n_19541), .o(n_19648) );
in01s02 g761530 ( .a(FE_OCP_RBN4067_n_18829), .o(n_18869) );
na03s06 TIMEBOOST_cell_5753 ( .a(n_7852), .b(FE_OCP_RBN6604_n_7881), .c(n_7836), .o(n_8017) );
no02f04 g761534 ( .a(FE_OCP_RBN6372_FE_RN_1425_0), .b(n_18320), .o(n_18801) );
in01s02 g761536 ( .a(n_18799), .o(n_18871) );
no02m02 g761539 ( .a(n_18754), .b(n_18716), .o(n_18798) );
no02m02 g761540 ( .a(FE_OCP_RBN1809_n_18754), .b(n_18682), .o(n_18828) );
no02s01 g761541 ( .a(n_19548), .b(n_19547), .o(n_19549) );
na02s01 g761542 ( .a(n_19545), .b(n_19544), .o(n_19546) );
no02s01 g761546 ( .a(n_18999), .b(n_18998), .o(n_19000) );
no02s06 TIMEBOOST_cell_8692 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_4_), .b(FE_OCP_RBN6516_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(TIMEBOOST_net_2833) );
in01s01 g761548 ( .a(n_18996), .o(n_18997) );
no02m04 g761549 ( .a(n_18938), .b(FE_OCP_DRV_N1438_n_17643), .o(n_18996) );
no02s01 g761550 ( .a(n_19542), .b(n_19541), .o(n_19543) );
na02f04 g761551 ( .a(n_18861), .b(FE_OCPN1636_n_18860), .o(n_18863) );
no02s06 g761552 ( .a(n_18861), .b(FE_OCPN1646_n_18860), .o(n_18862) );
no02s01 g761553 ( .a(n_18948), .b(n_18919), .o(n_18920) );
na02s01 g761554 ( .a(n_18895), .b(n_18894), .o(n_18896) );
in01s01 g761555 ( .a(n_19022), .o(n_19023) );
no02m06 g761556 ( .a(n_18939), .b(n_17644), .o(n_19022) );
no02f01 g761557 ( .a(n_18858), .b(n_18866), .o(n_18942) );
in01f01 g761558 ( .a(n_18950), .o(n_18859) );
na02f08 g761559 ( .a(FE_OCP_RBN1810_n_18754), .b(n_18721), .o(n_18950) );
in01s03 g761569 ( .a(n_20231), .o(n_22580) );
in01s02 g761573 ( .a(n_20086), .o(n_20231) );
in01s02 g761576 ( .a(n_20231), .o(n_22833) );
in01s02 g761577 ( .a(n_20231), .o(n_22793) );
in01s02 g761580 ( .a(n_20252), .o(n_22961) );
in01s01 g761582 ( .a(n_22580), .o(n_22907) );
in01s01 g761586 ( .a(n_20252), .o(n_22801) );
in01s01 g761587 ( .a(n_20231), .o(n_20252) );
in01s02 g761599 ( .a(n_19980), .o(n_20086) );
in01s02 g761603 ( .a(n_19787), .o(n_19980) );
in01s01 g761611 ( .a(n_19787), .o(n_19845) );
in01s02 g761612 ( .a(n_19647), .o(n_19787) );
in01s03 g761618 ( .a(n_19649), .o(n_19647) );
in01s02 g761619 ( .a(n_19609), .o(n_19649) );
in01s01 g761620 ( .a(n_19609), .o(n_19569) );
oa12s01 g761622 ( .a(n_18843), .b(n_19526), .c(n_18932), .o(n_19578) );
ao12s01 g761623 ( .a(n_18818), .b(n_19540), .c(n_18816), .o(n_19611) );
ao12s01 g761624 ( .a(n_19096), .b(n_19496), .c(n_18623), .o(n_19613) );
ao12s01 g761625 ( .a(n_18934), .b(n_19494), .c(n_18664), .o(n_19573) );
oa12s01 g761626 ( .a(n_19522), .b(n_19521), .c(n_19520), .o(n_19844) );
in01s01 g761627 ( .a(n_19607), .o(n_19900) );
ao12s01 g761628 ( .a(n_19525), .b(n_19524), .c(n_19523), .o(n_19607) );
in01s01 g761632 ( .a(n_18893), .o(n_18918) );
in01f02 g761633 ( .a(n_18893), .o(n_18892) );
na02s02 TIMEBOOST_cell_6813 ( .a(n_11026), .b(n_11000), .o(TIMEBOOST_net_2164) );
in01s01 g761635 ( .a(n_18971), .o(n_19127) );
ao12f02 g761636 ( .a(n_18940), .b(n_18887), .c(n_18822), .o(n_18971) );
in01s04 g761638 ( .a(n_18949), .o(n_18826) );
in01m02 g761639 ( .a(n_18797), .o(n_18949) );
in01m02 g761640 ( .a(n_18797), .o(n_18761) );
no02f04 g761641 ( .a(n_18652), .b(n_18683), .o(n_18797) );
in01s01 g761642 ( .a(n_19794), .o(n_19571) );
oa12s01 g761643 ( .a(n_19493), .b(n_19492), .c(n_19491), .o(n_19794) );
ao12s01 g761644 ( .a(n_19490), .b(n_19489), .c(n_19488), .o(n_19928) );
ao12s01 g761645 ( .a(n_19487), .b(n_19486), .c(n_19485), .o(n_19927) );
ao22s01 g761646 ( .a(n_19540), .b(n_18838), .c(n_19526), .d(n_18837), .o(n_19986) );
no02m08 g761648 ( .a(n_18756), .b(n_18265), .o(n_18758) );
na03m04 TIMEBOOST_cell_5752 ( .a(FE_RN_1922_0), .b(FE_RN_1921_0), .c(FE_RN_541_0), .o(n_19419) );
na02m06 g761651 ( .a(n_18682), .b(FE_OFN737_n_17093), .o(n_18721) );
no02s01 g761652 ( .a(n_19496), .b(n_19049), .o(n_19548) );
no02s01 g761654 ( .a(n_19494), .b(n_18883), .o(n_19545) );
na02s01 g761655 ( .a(n_19492), .b(n_19491), .o(n_19493) );
no02s01 g761656 ( .a(n_19524), .b(n_19523), .o(n_19525) );
na02s01 g761657 ( .a(n_19521), .b(n_19520), .o(n_19522) );
no02s01 g761658 ( .a(n_19489), .b(n_19488), .o(n_19490) );
no02s01 g761659 ( .a(n_19486), .b(n_19485), .o(n_19487) );
no03s02 TIMEBOOST_cell_8364 ( .a(FE_OCP_RBN5870_n_3704), .b(FE_OCP_RBN6765_n_3704), .c(FE_OCP_RBN2938_n_47013), .o(TIMEBOOST_net_1643) );
no02s01 g761661 ( .a(n_18940), .b(n_18888), .o(n_18999) );
no02s04 TIMEBOOST_cell_1915 ( .a(n_11366), .b(n_11386), .o(TIMEBOOST_net_572) );
na02s02 g761663 ( .a(n_18756), .b(n_18276), .o(n_18757) );
in01s01 g761665 ( .a(n_18858), .o(n_18890) );
na02f06 g761669 ( .a(n_18681), .b(n_18649), .o(n_18754) );
ao12s01 g761670 ( .a(n_18776), .b(n_19370), .c(n_18581), .o(n_19542) );
in01s01 g761671 ( .a(FE_RN_2617_0), .o(n_20797) );
in01s01 TIMEBOOST_cell_5915 ( .a(FE_OFN1_n_43918), .o(TIMEBOOST_net_1804) );
in01s01 g761678 ( .a(n_18861), .o(n_19027) );
oa12f06 g761679 ( .a(n_18561), .b(n_18560), .c(n_18795), .o(n_18861) );
no02s04 g761680 ( .a(n_18794), .b(n_18750), .o(n_18948) );
oa12s01 g761681 ( .a(n_18749), .b(n_18795), .c(n_18748), .o(n_18895) );
in01s02 g761682 ( .a(n_18938), .o(n_18939) );
na03m08 TIMEBOOST_cell_4831 ( .a(FE_RN_2703_0), .b(FE_RN_2704_0), .c(FE_RN_614_0), .o(n_31677) );
in01f01 g761684 ( .a(n_18756), .o(n_18717) );
oa12f08 g761685 ( .a(n_18243), .b(n_18647), .c(n_18221), .o(n_18756) );
na02f08 g761688 ( .a(n_18602), .b(n_18271), .o(n_18650) );
na02m08 TIMEBOOST_cell_1969 ( .a(n_37337), .b(n_37156), .o(TIMEBOOST_net_599) );
no04m10 TIMEBOOST_cell_3649 ( .a(FE_OCP_RBN6763_FE_RN_2259_0), .b(FE_OCP_RBN4309_n_25178), .c(n_25265), .d(n_25295), .o(FE_RN_323_0) );
na02m04 g761692 ( .a(n_18600), .b(FE_OFN737_n_17093), .o(n_18649) );
no02f01 g761693 ( .a(n_18824), .b(n_18713), .o(n_18825) );
na02s01 g761694 ( .a(n_19405), .b(n_19406), .o(n_19492) );
no02s01 g761695 ( .a(n_19405), .b(n_18737), .o(n_19496) );
no02s01 g761696 ( .a(n_19404), .b(n_18571), .o(n_19494) );
na02s01 TIMEBOOST_cell_4441 ( .a(n_9173), .b(n_9111), .o(TIMEBOOST_net_1311) );
na02s01 g761698 ( .a(n_18853), .b(n_18432), .o(n_18916) );
no02s02 g761699 ( .a(n_18681), .b(n_18600), .o(n_18794) );
no02s02 g761700 ( .a(FE_OCP_RBN4639_n_18681), .b(FE_OCP_RBN4636_n_18600), .o(n_18750) );
na02s01 g761701 ( .a(n_18795), .b(n_18748), .o(n_18749) );
in01s01 g761702 ( .a(n_18887), .o(n_18888) );
na02f02 g761703 ( .a(n_18855), .b(FE_OCPN1258_n_18854), .o(n_18887) );
no02f02 g761704 ( .a(n_18855), .b(FE_OCPN1258_n_18854), .o(n_18940) );
na02m04 TIMEBOOST_cell_3266 ( .a(n_30297), .b(n_30280), .o(TIMEBOOST_net_924) );
no02s04 TIMEBOOST_cell_1845 ( .a(n_5818), .b(FE_OCPN3584_n_4556), .o(TIMEBOOST_net_537) );
oa12s01 g761708 ( .a(n_19402), .b(n_19401), .c(n_18739), .o(n_19489) );
oa12s01 g761709 ( .a(n_19400), .b(n_19401), .c(n_18694), .o(n_19486) );
in01s01 g761713 ( .a(n_18682), .o(n_18716) );
ao12s01 g761715 ( .a(n_19368), .b(n_19401), .c(n_19367), .o(n_19873) );
in01s01 g761716 ( .a(n_19398), .o(n_19399) );
oa12s01 g761717 ( .a(n_19297), .b(n_19296), .c(n_19295), .o(n_19398) );
in01s01 g761718 ( .a(n_19526), .o(n_19540) );
oa12s01 g761719 ( .a(n_18992), .b(n_19401), .c(n_18964), .o(n_19526) );
no02m02 g761721 ( .a(n_18647), .b(n_18214), .o(n_18653) );
no02f06 g761722 ( .a(n_18439), .b(n_18311), .o(n_18602) );
na02s01 g761723 ( .a(n_19339), .b(n_18910), .o(n_19405) );
in01s01 g761724 ( .a(n_19369), .o(n_19370) );
na02s01 g761725 ( .a(n_19339), .b(n_18663), .o(n_19369) );
na02s01 g761726 ( .a(n_19339), .b(n_18774), .o(n_19404) );
no02s01 g761727 ( .a(n_19401), .b(n_19367), .o(n_19368) );
na02s01 g761728 ( .a(n_19296), .b(n_19295), .o(n_19297) );
in01s01 g761729 ( .a(n_18824), .o(n_18791) );
no02s02 TIMEBOOST_cell_1928 ( .a(TIMEBOOST_net_578), .b(n_11823), .o(n_11982) );
in01s01 g761739 ( .a(n_18713), .o(n_18746) );
in01s01 g761741 ( .a(n_18852), .o(n_18853) );
oa12s01 g761742 ( .a(n_18745), .b(n_18789), .c(n_18744), .o(n_18852) );
na02f02 g761743 ( .a(n_18709), .b(n_18684), .o(n_18855) );
in01s01 g761744 ( .a(n_18822), .o(n_18998) );
oa12m02 g761745 ( .a(n_18480), .b(n_18789), .c(n_18482), .o(n_18822) );
no02f06 g761751 ( .a(n_18565), .b(n_18599), .o(n_18795) );
ao12s01 g761752 ( .a(n_19294), .b(n_19293), .c(n_19292), .o(n_19790) );
in01s01 g761753 ( .a(n_19337), .o(n_19796) );
oa12s01 g761754 ( .a(n_19230), .b(n_19229), .c(n_19228), .o(n_19337) );
ao12s01 g761755 ( .a(n_19233), .b(n_19232), .c(n_19231), .o(n_19793) );
no02f08 g761756 ( .a(n_18518), .b(n_18215), .o(n_18647) );
in01s02 g761757 ( .a(n_18519), .o(n_18520) );
in01m01 g761758 ( .a(n_18439), .o(n_18519) );
oa12f04 g761759 ( .a(n_18246), .b(n_18348), .c(n_18223), .o(n_18439) );
na02m06 g761760 ( .a(n_18710), .b(n_18472), .o(n_18870) );
na02m08 TIMEBOOST_cell_1970 ( .a(TIMEBOOST_net_599), .b(n_37488), .o(n_37536) );
no02m02 g761763 ( .a(n_18564), .b(n_18437), .o(n_18565) );
no02m06 g761764 ( .a(n_18517), .b(n_18484), .o(n_18599) );
no02s01 g761765 ( .a(n_19293), .b(n_19292), .o(n_19294) );
na02s01 g761766 ( .a(n_18789), .b(n_18744), .o(n_18745) );
na02s02 g761767 ( .a(FE_OCP_RBN5030_n_18678), .b(n_18645), .o(n_18709) );
no02s01 g761768 ( .a(n_19232), .b(n_19231), .o(n_19233) );
na02s01 g761769 ( .a(n_19229), .b(n_19228), .o(n_19230) );
na02f01 g761770 ( .a(n_18646), .b(n_18678), .o(n_18684) );
ao12s01 g761771 ( .a(n_18885), .b(n_19191), .c(n_18809), .o(n_19296) );
oa12s01 g761772 ( .a(n_19161), .b(n_19160), .c(n_19159), .o(n_19760) );
ao12s01 g761773 ( .a(n_19195), .b(n_19194), .c(n_19193), .o(n_19735) );
in01s01 g761774 ( .a(n_19339), .o(n_19401) );
in01s01 g761776 ( .a(n_19291), .o(n_19825) );
ao12s01 g761777 ( .a(n_19198), .b(n_19197), .c(n_19196), .o(n_19291) );
na02m06 g761778 ( .a(n_18555), .b(n_18477), .o(n_18710) );
in01s02 g761780 ( .a(n_18562), .o(n_18563) );
in01m01 g761781 ( .a(n_18518), .o(n_18562) );
ao12f06 g761782 ( .a(n_18185), .b(n_18376), .c(n_18213), .o(n_18518) );
in01s01 g761783 ( .a(n_18850), .o(n_18851) );
no02s01 g761784 ( .a(n_18821), .b(n_18743), .o(n_18850) );
na02s01 g761785 ( .a(n_19158), .b(n_18884), .o(n_19293) );
na02s01 g761786 ( .a(n_19160), .b(n_19159), .o(n_19161) );
na02m02 g761787 ( .a(n_18894), .b(n_18559), .o(n_18561) );
no02s03 g761788 ( .a(n_18894), .b(FE_OCP_DRV_N3534_n_18559), .o(n_18560) );
no02s01 g761789 ( .a(n_19197), .b(n_19196), .o(n_19198) );
no02s01 g761790 ( .a(n_19194), .b(n_19193), .o(n_19195) );
oa12m02 g761791 ( .a(n_18217), .b(n_18379), .c(n_18377), .o(n_18412) );
na02s01 TIMEBOOST_cell_1839 ( .a(n_15479), .b(FE_OCP_RBN3134_n_46982), .o(TIMEBOOST_net_534) );
in01f04 g761793 ( .a(n_18645), .o(n_18646) );
oa12s01 g761797 ( .a(n_18815), .b(n_19125), .c(n_18655), .o(n_19232) );
in01s01 g761803 ( .a(n_18517), .o(n_18557) );
in01m02 g761805 ( .a(n_18564), .o(n_18517) );
no02f04 g761806 ( .a(n_18411), .b(n_18380), .o(n_18564) );
in01s01 g761807 ( .a(FE_OCPN5248_FE_OFN4715_n_18642), .o(n_20635) );
ao22s01 g761808 ( .a(n_18436), .b(n_16968), .c(n_18409), .d(n_18483), .o(n_18642) );
oa12s01 g761809 ( .a(n_18700), .b(n_19126), .c(n_18610), .o(n_19229) );
no02s02 g761811 ( .a(n_18379), .b(n_18244), .o(n_18380) );
no02m02 g761812 ( .a(n_18347), .b(n_18245), .o(n_18411) );
no02f04 g761813 ( .a(n_18322), .b(n_18193), .o(n_18348) );
no02m04 TIMEBOOST_cell_1836 ( .a(TIMEBOOST_net_532), .b(n_31863), .o(n_31951) );
in01m02 g761815 ( .a(n_18554), .o(n_18555) );
na02m08 g761816 ( .a(n_18435), .b(n_18373), .o(n_18554) );
ao12s02 g761817 ( .a(n_18398), .b(n_18406), .c(n_18284), .o(n_18516) );
na02m01 g761818 ( .a(n_18641), .b(n_18431), .o(n_18821) );
in01s02 g761820 ( .a(n_18437), .o(n_18484) );
no02m06 g761821 ( .a(n_18375), .b(n_17423), .o(n_18437) );
na02s01 g761822 ( .a(n_19126), .b(n_18619), .o(n_19194) );
no02s02 g761823 ( .a(n_18375), .b(n_18483), .o(n_18894) );
na02s01 g761824 ( .a(n_19125), .b(n_18731), .o(n_19197) );
in01s01 g761825 ( .a(n_19191), .o(n_19158) );
no02m06 g761826 ( .a(n_19125), .b(n_18730), .o(n_19191) );
ao12s01 g761827 ( .a(n_18583), .b(n_19097), .c(n_18657), .o(n_19160) );
oa12s01 g761828 ( .a(n_19071), .b(n_19097), .c(n_19070), .o(n_19758) );
ao12s01 g761829 ( .a(n_18786), .b(n_18672), .c(n_18355), .o(n_18787) );
na02s01 g761830 ( .a(n_19097), .b(n_18697), .o(n_19126) );
no02s02 g761831 ( .a(n_18481), .b(n_18479), .o(n_18482) );
na02s01 g761832 ( .a(n_18481), .b(n_18479), .o(n_18480) );
na02s01 g761833 ( .a(n_19097), .b(n_19070), .o(n_19071) );
na03s08 TIMEBOOST_cell_6433 ( .a(n_18134), .b(FE_RN_355_0), .c(FE_RN_354_0), .o(n_18188) );
oa12f06 g761835 ( .a(n_18126), .b(n_18318), .c(n_18127), .o(n_18376) );
in01m01 g761836 ( .a(n_18379), .o(n_18347) );
in01m01 g761837 ( .a(n_18322), .o(n_18379) );
oa12f04 g761838 ( .a(n_18202), .b(n_18269), .c(n_18171), .o(n_18322) );
in01s02 g761839 ( .a(n_18475), .o(n_18476) );
ao12s02 g761840 ( .a(n_18127), .b(n_18318), .c(n_18126), .o(n_18475) );
oa12s01 g761841 ( .a(n_18284), .b(n_18595), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_27_), .o(n_18641) );
ao12s01 g761842 ( .a(n_18704), .b(n_18741), .c(n_17748), .o(n_18743) );
oa22s01 g761843 ( .a(n_18553), .b(n_16931), .c(n_18397), .d(n_18404), .o(n_20293) );
in01s01 g761851 ( .a(n_18409), .o(n_18436) );
in01s01 g761853 ( .a(n_18375), .o(n_18409) );
ao12s01 g761856 ( .a(n_18995), .b(n_18994), .c(n_18993), .o(n_19677) );
in01s01 g761857 ( .a(n_20135), .o(n_20136) );
ao12s01 g761858 ( .a(n_19021), .b(n_19020), .c(n_19019), .o(n_20135) );
no02m06 g761859 ( .a(n_18321), .b(n_18346), .o(n_18718) );
na02s02 g761860 ( .a(n_18472), .b(n_18470), .o(n_18473) );
no02s02 g761862 ( .a(n_18549), .b(n_18548), .o(n_18550) );
na02s04 TIMEBOOST_cell_6775 ( .a(n_9289), .b(n_9348), .o(TIMEBOOST_net_2145) );
in01m02 g761864 ( .a(n_18407), .o(n_18408) );
na02m01 g761865 ( .a(n_18373), .b(n_18372), .o(n_18407) );
no02s01 g761866 ( .a(n_18786), .b(n_18593), .o(n_18675) );
na02s01 g761867 ( .a(n_18368), .b(n_18367), .o(n_18406) );
in01s01 g761868 ( .a(n_18784), .o(n_18785) );
na02s02 g761869 ( .a(n_18742), .b(n_18741), .o(n_18784) );
in01s01 g761870 ( .a(n_18513), .o(n_18514) );
na02s06 g761871 ( .a(n_47246), .b(n_18470), .o(n_18513) );
in01s02 g761872 ( .a(n_18370), .o(n_18371) );
na02s06 g761873 ( .a(n_47247), .b(n_18345), .o(n_18370) );
in01s01 g761874 ( .a(n_18936), .o(n_18937) );
na02s01 g761875 ( .a(n_18915), .b(n_18914), .o(n_18936) );
in01s01 g761876 ( .a(n_18546), .o(n_18547) );
na02s06 g761877 ( .a(n_18511), .b(n_18512), .o(n_18546) );
in01s01 g761878 ( .a(n_18639), .o(n_18640) );
no02s01 g761879 ( .a(FE_RN_1842_0), .b(n_18549), .o(n_18639) );
no02s01 g761880 ( .a(n_18994), .b(n_18993), .o(n_18995) );
no02s01 g761881 ( .a(n_19020), .b(n_19019), .o(n_19021) );
in01s01 g761883 ( .a(n_18433), .o(n_18468) );
na02m04 g761884 ( .a(n_18405), .b(FE_OFN737_n_17093), .o(n_18433) );
in01s01 g761885 ( .a(n_18848), .o(n_18849) );
ao12s01 g761886 ( .a(n_18820), .b(n_18284), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_29_), .o(n_18848) );
in01s02 g761887 ( .a(n_18509), .o(n_18510) );
no02s06 TIMEBOOST_cell_8854 ( .a(FE_OCP_RBN4391_n_16230), .b(n_14618), .o(TIMEBOOST_net_2914) );
in01s01 g761889 ( .a(n_18707), .o(n_18708) );
ao12f01 g761890 ( .a(n_18674), .b(n_18284), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_27_), .o(n_18707) );
in01s01 g761891 ( .a(n_18481), .o(n_18432) );
na02m01 g761892 ( .a(n_18405), .b(n_18404), .o(n_18481) );
in01s01 g761894 ( .a(n_19650), .o(n_19051) );
oa12s01 g761895 ( .a(n_18970), .b(n_18969), .c(n_18968), .o(n_19650) );
in01s01 g761896 ( .a(n_18912), .o(n_18913) );
ao22s01 g761897 ( .a(n_18704), .b(n_17724), .c(n_18284), .d(delay_sub_ln21_0_unr11_stage5_stallmux_q_31_), .o(n_18912) );
in01s01 g761898 ( .a(n_18544), .o(n_18545) );
oa12s02 g761899 ( .a(n_18401), .b(n_18284), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n_18544) );
in01s01 g761900 ( .a(n_18637), .o(n_18638) );
oa12s01 g761901 ( .a(n_18467), .b(n_18284), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_), .o(n_18637) );
na02s01 g761903 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_28_), .o(n_18741) );
in01m04 g761904 ( .a(n_18321), .o(n_18373) );
no02m08 g761905 ( .a(n_18302), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_19_), .o(n_18321) );
na02s01 g761908 ( .a(n_18704), .b(n_17749), .o(n_18915) );
na02s06 g761909 ( .a(FE_OFN777_n_18268), .b(n_18291), .o(n_18345) );
na02s01 g761910 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_30_), .o(n_18914) );
no02s01 g761911 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_29_), .o(n_18820) );
na02f01 g761912 ( .a(FE_OFN777_n_18268), .b(n_17696), .o(n_18742) );
na02m08 g761913 ( .a(n_18302), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_19_), .o(n_18372) );
na02s06 g761915 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_22_), .o(n_18470) );
na02s01 g761918 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n_18401) );
in01s01 g761919 ( .a(n_18319), .o(n_18320) );
na02m02 g761920 ( .a(n_18434), .b(n_18301), .o(n_18319) );
na02s01 TIMEBOOST_cell_7597 ( .a(TIMEBOOST_net_2429), .b(n_34532), .o(n_34653) );
na02s02 g761922 ( .a(FE_OFN777_n_18268), .b(n_18367), .o(n_18440) );
na02s03 g761923 ( .a(n_18508), .b(n_18424), .o(n_18786) );
na02s01 g761924 ( .a(n_18634), .b(n_17856), .o(n_18672) );
na02s06 g761925 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_24_), .o(n_18511) );
na02s06 g761926 ( .a(FE_OFN777_n_18268), .b(n_17772), .o(n_18512) );
na02s01 g761927 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_), .o(n_18467) );
no02s01 g761928 ( .a(FE_OFN777_n_18268), .b(n_17722), .o(n_18595) );
no02s01 g761929 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_26_), .o(n_18549) );
no02m01 g761930 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_27_), .o(n_18674) );
na02s01 g761931 ( .a(n_18969), .b(n_18968), .o(n_18970) );
na02s01 g761933 ( .a(n_19050), .b(n_18839), .o(n_19096) );
oa12s04 g761934 ( .a(FE_OFN777_n_18268), .b(n_18291), .c(n_17508), .o(n_18477) );
na02s02 g761935 ( .a(FE_OFN777_n_18268), .b(n_17556), .o(n_18366) );
na02f08 TIMEBOOST_cell_4929 ( .a(n_17843), .b(TIMEBOOST_net_1412), .o(n_17997) );
in01s02 g761940 ( .a(n_18398), .o(n_18472) );
no02s03 g761941 ( .a(FE_OFN777_n_18268), .b(n_17555), .o(n_18398) );
no02s01 g761942 ( .a(n_18284), .b(n_17773), .o(n_18548) );
in01s01 g761943 ( .a(n_18431), .o(n_18594) );
oa12s02 g761944 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_24_), .o(n_18431) );
in01m01 g761946 ( .a(n_18318), .o(n_18360) );
oa12f08 g761949 ( .a(n_18109), .b(n_18267), .c(n_18071), .o(n_18318) );
oa12f06 g761952 ( .a(n_18136), .b(n_18248), .c(n_18091), .o(n_18269) );
oa12s01 g761953 ( .a(n_18735), .b(n_18911), .c(n_18533), .o(n_18994) );
no02s01 g761954 ( .a(n_18966), .b(n_18736), .o(n_19020) );
oa22s01 g761956 ( .a(FE_OCP_RBN7022_n_18248), .b(n_18149), .c(n_18248), .d(n_18150), .o(n_18287) );
in01s01 g761958 ( .a(n_18397), .o(n_18553) );
in01s01 g761959 ( .a(n_18405), .o(n_18397) );
no02m04 TIMEBOOST_cell_6297 ( .a(n_10966), .b(n_10917), .o(TIMEBOOST_net_2000) );
na02s04 g761962 ( .a(n_18357), .b(n_18393), .o(n_18396) );
in01s02 g761963 ( .a(n_18301), .o(n_18346) );
na02s06 g761964 ( .a(n_18224), .b(n_17186), .o(n_18301) );
na02m08 g761965 ( .a(n_18225), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_18_), .o(n_18434) );
in01m02 g761966 ( .a(n_18316), .o(n_18317) );
no02m02 g761967 ( .a(n_18300), .b(n_18285), .o(n_18316) );
no02s01 g761968 ( .a(n_18705), .b(n_18589), .o(n_18706) );
na02s01 g761969 ( .a(n_18911), .b(n_18622), .o(n_18969) );
no02s01 g761970 ( .a(n_18963), .b(n_18931), .o(n_18992) );
in01s01 g761972 ( .a(n_19049), .o(n_19050) );
na02s01 g761973 ( .a(n_19406), .b(n_18840), .o(n_19049) );
in01s01 g761983 ( .a(n_18284), .o(n_18704) );
in01m10 g761984 ( .a(FE_OFN777_n_18268), .o(n_18284) );
ao12m06 g762000 ( .a(n_18005), .b(n_18226), .c(n_18050), .o(n_18268) );
no02m04 g762001 ( .a(n_18911), .b(n_18587), .o(n_18966) );
oa12s02 g762002 ( .a(n_18355), .b(n_18461), .c(delay_add_ln22_unr11_stage5_stallmux_q_27_), .o(n_18508) );
in01s01 g762003 ( .a(n_18634), .o(n_19478) );
oa12s01 g762004 ( .a(n_18355), .b(n_18593), .c(delay_add_ln22_unr11_stage5_stallmux_q_29_), .o(n_18634) );
no02s02 TIMEBOOST_cell_7518 ( .a(n_23869), .b(n_23671), .o(TIMEBOOST_net_2390) );
in01s01 g762006 ( .a(n_18935), .o(n_19733) );
oa12s01 g762007 ( .a(n_18846), .b(n_18847), .c(n_18845), .o(n_18935) );
in01s01 g762008 ( .a(n_19913), .o(n_18886) );
ao12s01 g762009 ( .a(n_18781), .b(n_18780), .c(n_18779), .o(n_19913) );
na02s01 g762010 ( .a(n_18332), .b(n_18354), .o(n_18395) );
no02s02 g762015 ( .a(n_18309), .b(n_18337), .o(n_18357) );
in01s01 g762016 ( .a(n_18633), .o(n_18705) );
no02s01 g762017 ( .a(n_18541), .b(n_18590), .o(n_18633) );
in01s01 g762019 ( .a(n_18506), .o(n_18507) );
na02s01 g762020 ( .a(n_18390), .b(n_18460), .o(n_18506) );
in01s01 g762021 ( .a(n_18427), .o(n_18428) );
na02s06 g762022 ( .a(n_18393), .b(n_18394), .o(n_18427) );
no02s06 g762023 ( .a(n_18205), .b(n_16990), .o(n_18285) );
in01s01 g762024 ( .a(n_18391), .o(n_18392) );
no02s01 g762025 ( .a(n_18356), .b(n_18337), .o(n_18391) );
in01s01 g762026 ( .a(n_18458), .o(n_18459) );
no02s02 g762027 ( .a(n_18426), .b(n_18425), .o(n_18458) );
in01s01 g762028 ( .a(n_18335), .o(n_18336) );
na02m01 g762029 ( .a(n_18279), .b(n_18313), .o(n_18335) );
in01m02 g762030 ( .a(n_18300), .o(n_18271) );
no02m08 g762031 ( .a(n_18206), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_17_), .o(n_18300) );
in01s02 g762032 ( .a(n_18333), .o(n_18334) );
no02m02 g762033 ( .a(n_18263), .b(n_18311), .o(n_18333) );
in01s01 g762034 ( .a(n_18591), .o(n_18592) );
no02s01 g762035 ( .a(n_18541), .b(n_18593), .o(n_18591) );
in01s01 g762036 ( .a(n_18323), .o(n_18324) );
no02s06 g762037 ( .a(n_19014), .b(n_18280), .o(n_18323) );
no02s01 g762038 ( .a(n_18780), .b(n_18779), .o(n_18781) );
na02m04 g762039 ( .a(n_18847), .b(n_18614), .o(n_18911) );
na02s01 g762040 ( .a(n_18847), .b(n_18845), .o(n_18846) );
no02m08 g762041 ( .a(n_18195), .b(n_18076), .o(n_18204) );
na02s01 TIMEBOOST_cell_6038 ( .a(TIMEBOOST_net_1870), .b(n_37945), .o(TIMEBOOST_net_1051) );
na02s01 g762043 ( .a(n_18930), .b(n_18807), .o(n_18934) );
na02s04 g762044 ( .a(n_18738), .b(n_18910), .o(n_18964) );
in01s01 g762045 ( .a(n_18539), .o(n_18540) );
ao12s01 g762046 ( .a(n_18505), .b(n_18355), .c(delay_add_ln22_unr11_stage5_stallmux_q_27_), .o(n_18539) );
in01s01 g762047 ( .a(n_18537), .o(n_18538) );
ao22s01 g762048 ( .a(FE_OCP_RBN2496_n_18242), .b(n_18331), .c(n_18355), .d(delay_add_ln22_unr11_stage5_stallmux_q_25_), .o(n_18537) );
in01s01 g762049 ( .a(n_18456), .o(n_18457) );
ao12s01 g762050 ( .a(n_47248), .b(n_18355), .c(delay_add_ln22_unr11_stage5_stallmux_q_21_), .o(n_18456) );
ao12s01 g762052 ( .a(n_18590), .b(n_18355), .c(delay_add_ln22_unr11_stage5_stallmux_q_29_), .o(n_18631) );
in01s01 g762053 ( .a(n_18629), .o(n_18630) );
ao12s01 g762054 ( .a(n_18589), .b(n_18355), .c(delay_add_ln22_unr11_stage5_stallmux_q_30_), .o(n_18629) );
oa12f08 g762056 ( .a(n_18114), .b(n_18196), .c(n_18078), .o(n_18248) );
in01s01 g762057 ( .a(n_18282), .o(n_18283) );
in01s01 g762058 ( .a(n_18267), .o(n_18282) );
oa12f08 g762059 ( .a(n_18105), .b(n_18247), .c(n_18067), .o(n_18267) );
in01s02 g762061 ( .a(n_18963), .o(n_19406) );
na02s04 g762062 ( .a(n_18930), .b(n_18836), .o(n_18963) );
ao12s01 g762063 ( .a(n_18180), .b(n_18196), .c(n_18179), .o(n_19855) );
in01s01 g762064 ( .a(n_18669), .o(n_18670) );
oa22s01 g762065 ( .a(n_18355), .b(delay_add_ln22_unr11_stage5_stallmux_q_31_), .c(FE_OCP_RBN2496_n_18242), .d(n_17852), .o(n_18669) );
ao22s01 g762066 ( .a(n_18247), .b(n_18125), .c(n_18201), .d(n_18124), .o(n_19885) );
in01m04 g762067 ( .a(n_18224), .o(n_18225) );
no02s02 g762069 ( .a(n_18355), .b(delay_add_ln22_unr11_stage5_stallmux_q_27_), .o(n_18505) );
in01s01 g762070 ( .a(n_18390), .o(n_18461) );
na02s01 g762071 ( .a(n_18355), .b(delay_add_ln22_unr11_stage5_stallmux_q_26_), .o(n_18390) );
na02s01 g762072 ( .a(FE_OCP_RBN2496_n_18242), .b(n_18331), .o(n_18332) );
no02s01 g762073 ( .a(FE_OCP_RBN2496_n_18242), .b(n_18329), .o(n_18426) );
in01s01 g762074 ( .a(n_18354), .o(n_18425) );
na02s02 g762075 ( .a(FE_OCP_RBN2496_n_18242), .b(n_18329), .o(n_18354) );
no02s10 g762076 ( .a(FE_OCP_RBN2495_n_18242), .b(delay_add_ln22_unr11_stage5_stallmux_q_20_), .o(n_19014) );
no02s02 g762079 ( .a(FE_OCP_RBN2495_n_18242), .b(delay_add_ln22_unr11_stage5_stallmux_q_22_), .o(n_18356) );
na02s10 g762080 ( .a(FE_OCP_RBN2496_n_18242), .b(n_17692), .o(n_18394) );
na02s03 g762081 ( .a(FE_OCP_RBN2497_n_18242), .b(delay_add_ln22_unr11_stage5_stallmux_q_23_), .o(n_18393) );
no02s01 g762082 ( .a(n_18242), .b(n_17625), .o(n_18337) );
in01s01 g762084 ( .a(n_18280), .o(n_18298) );
no02s02 g762085 ( .a(n_18242), .b(n_17416), .o(n_18280) );
na02f04 g762086 ( .a(n_18216), .b(n_18222), .o(n_18223) );
in01s01 g762087 ( .a(n_18541), .o(n_18455) );
no02s01 g762088 ( .a(n_18355), .b(delay_add_ln22_unr11_stage5_stallmux_q_28_), .o(n_18541) );
no02s01 g762089 ( .a(FE_OCP_RBN2496_n_18242), .b(n_17805), .o(n_18593) );
no02s01 g762090 ( .a(n_18355), .b(delay_add_ln22_unr11_stage5_stallmux_q_29_), .o(n_18590) );
no02s01 g762091 ( .a(n_18355), .b(delay_add_ln22_unr11_stage5_stallmux_q_30_), .o(n_18589) );
na02m01 g762092 ( .a(FE_OCP_RBN2496_n_18242), .b(n_17806), .o(n_18460) );
no02s01 g762093 ( .a(n_18196), .b(n_18179), .o(n_18180) );
in01s01 g762094 ( .a(n_18278), .o(n_18279) );
no02s06 g762095 ( .a(n_18266), .b(delay_add_ln22_unr11_stage5_stallmux_q_19_), .o(n_18278) );
na02s04 g762096 ( .a(n_18266), .b(delay_add_ln22_unr11_stage5_stallmux_q_19_), .o(n_18313) );
in01s02 g762097 ( .a(n_18276), .o(n_18277) );
no02s06 g762098 ( .a(n_18265), .b(n_18264), .o(n_18276) );
no02m06 g762099 ( .a(n_18208), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_16_), .o(n_18311) );
na02m06 g762100 ( .a(n_18177), .b(n_18176), .o(n_18178) );
in01m08 g762101 ( .a(n_18195), .o(n_18226) );
na02m10 g762102 ( .a(n_18177), .b(n_18060), .o(n_18195) );
no02s06 g762106 ( .a(n_46972), .b(n_16830), .o(n_18263) );
in01s02 g762107 ( .a(n_18261), .o(n_18262) );
na02m02 g762108 ( .a(n_18246), .b(n_18222), .o(n_18261) );
na02s01 g762109 ( .a(n_18884), .b(n_18810), .o(n_18885) );
in01s01 g762110 ( .a(n_18462), .o(n_18424) );
no02s01 g762111 ( .a(FE_OCP_RBN2496_n_18242), .b(n_17813), .o(n_18462) );
in01s01 g762112 ( .a(n_18309), .o(n_18310) );
no02s01 g762113 ( .a(n_18242), .b(n_17568), .o(n_18309) );
na02m04 g762114 ( .a(n_18702), .b(n_18500), .o(n_18847) );
ao12s01 g762115 ( .a(n_18499), .b(n_18703), .c(n_18701), .o(n_18780) );
in01s02 g762116 ( .a(n_18883), .o(n_18930) );
na02s02 g762117 ( .a(n_19402), .b(n_18767), .o(n_18883) );
no02s04 g762118 ( .a(n_18775), .b(n_18666), .o(n_18910) );
in01s01 g762120 ( .a(n_18777), .o(n_18778) );
oa12s01 g762121 ( .a(n_18668), .b(n_18703), .c(n_18667), .o(n_18777) );
in01m04 g762122 ( .a(n_18205), .o(n_18206) );
oa12m08 g762123 ( .a(n_18175), .b(n_18174), .c(n_18173), .o(n_18205) );
na02m06 g762124 ( .a(n_18220), .b(n_18187), .o(n_18221) );
na02m08 g762125 ( .a(n_18174), .b(n_18173), .o(n_18175) );
in01m02 g762126 ( .a(n_18218), .o(n_18219) );
in01m02 g762128 ( .a(n_18244), .o(n_18245) );
na02m02 g762129 ( .a(n_18217), .b(n_18216), .o(n_18244) );
no02m06 g762130 ( .a(n_18189), .b(n_17050), .o(n_18264) );
no02s06 g762131 ( .a(n_18188), .b(delay_add_ln22_unr11_stage5_stallmux_q_18_), .o(n_18265) );
in01s02 g762132 ( .a(n_18259), .o(n_18260) );
na02m02 g762133 ( .a(n_18243), .b(n_18220), .o(n_18259) );
na02f04 g762134 ( .a(n_18164), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_15_), .o(n_18222) );
na02s06 g762136 ( .a(n_18165), .b(n_16779), .o(n_18246) );
na02s01 g762137 ( .a(n_18703), .b(n_18667), .o(n_18668) );
no02s02 g762138 ( .a(n_18776), .b(n_18766), .o(n_19402) );
no02s01 g762140 ( .a(n_18771), .b(n_18818), .o(n_18843) );
na02s01 g762141 ( .a(n_18817), .b(n_18816), .o(n_18932) );
no02s01 g762142 ( .a(n_18882), .b(n_18812), .o(n_19577) );
no02s01 g762143 ( .a(n_18814), .b(n_18577), .o(n_18815) );
na02s01 g762144 ( .a(n_18817), .b(n_18772), .o(n_19610) );
in01s02 g762145 ( .a(n_18774), .o(n_18775) );
no02s02 g762146 ( .a(n_18739), .b(n_18576), .o(n_18774) );
in01m02 g762155 ( .a(FE_OCP_RBN2496_n_18242), .o(n_18355) );
no02f06 TIMEBOOST_cell_5377 ( .a(TIMEBOOST_net_1636), .b(n_21793), .o(n_21902) );
oa12f08 g762168 ( .a(n_18088), .b(n_18138), .c(n_18045), .o(n_18196) );
in01s01 g762169 ( .a(n_18247), .o(n_18201) );
oa12f08 g762170 ( .a(n_18066), .b(n_18194), .c(n_18016), .o(n_18247) );
no02s01 TIMEBOOST_cell_1773 ( .a(n_21694), .b(n_21374), .o(TIMEBOOST_net_501) );
no02s04 g762173 ( .a(n_18814), .b(n_18618), .o(n_18884) );
oa22s01 g762174 ( .a(n_18138), .b(n_18108), .c(n_18095), .d(n_18107), .o(n_19801) );
na02m06 TIMEBOOST_cell_6034 ( .a(TIMEBOOST_net_1868), .b(n_19191), .o(n_19339) );
oa12s01 g762176 ( .a(n_18169), .b(n_18194), .c(n_18168), .o(n_19807) );
ao12s01 g762177 ( .a(n_18627), .b(n_18626), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_19608) );
na02m08 TIMEBOOST_cell_8623 ( .a(TIMEBOOST_net_2798), .b(n_11033), .o(n_11132) );
in01s02 g762180 ( .a(n_46972), .o(n_18208) );
na02s06 g762182 ( .a(n_18153), .b(n_18152), .o(n_18202) );
na02s06 g762183 ( .a(n_18162), .b(n_16921), .o(n_18243) );
in01s02 g762184 ( .a(n_18217), .o(n_18200) );
in01s02 g762185 ( .a(n_18193), .o(n_18217) );
no02s04 g762186 ( .a(n_18167), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_14_), .o(n_18193) );
na02m04 g762187 ( .a(n_18161), .b(delay_add_ln22_unr11_stage5_stallmux_q_17_), .o(n_18220) );
no02m06 g762189 ( .a(n_18153), .b(n_18152), .o(n_18171) );
in01m02 g762190 ( .a(n_18240), .o(n_18241) );
no02m02 g762191 ( .a(n_18215), .b(n_18214), .o(n_18240) );
na02s02 TIMEBOOST_cell_4231 ( .a(n_33396), .b(FE_OCP_RBN2505_n_33226), .o(TIMEBOOST_net_1206) );
no02s10 g762194 ( .a(n_18113), .b(n_18137), .o(n_18174) );
na02s01 g762195 ( .a(n_18194), .b(n_18168), .o(n_18169) );
in01s01 g762196 ( .a(n_18216), .o(n_18377) );
na02s04 g762197 ( .a(n_18167), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_14_), .o(n_18216) );
no02m06 TIMEBOOST_cell_6950 ( .a(TIMEBOOST_net_2233), .b(n_29473), .o(FE_RN_1101_0) );
no02s01 g762199 ( .a(n_18626), .b(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_18627) );
na02s06 TIMEBOOST_cell_8006 ( .a(FE_OCP_RBN4431_n_39942), .b(n_39992), .o(TIMEBOOST_net_2634) );
no03s02 TIMEBOOST_cell_8259 ( .a(FE_OCP_RBN2654_FE_OCPN914_n_8091), .b(FE_OCP_RBN2655_FE_OCPN914_n_8091), .c(n_7985), .o(TIMEBOOST_net_2106) );
na02s01 g762202 ( .a(n_18624), .b(n_18623), .o(n_18625) );
na02s01 g762203 ( .a(n_18735), .b(n_18620), .o(n_18736) );
no02s01 g762204 ( .a(n_18698), .b(n_18443), .o(n_18700) );
na02s01 g762205 ( .a(n_18813), .b(n_18624), .o(n_19680) );
no02s01 g762206 ( .a(n_18773), .b(n_45002), .o(n_18882) );
in01s01 g762207 ( .a(n_18837), .o(n_18838) );
na02s01 g762208 ( .a(n_18695), .b(n_18816), .o(n_18837) );
in01s01 g762209 ( .a(n_18811), .o(n_18812) );
na02s01 g762210 ( .a(n_18773), .b(n_45002), .o(n_18811) );
in01s01 g762211 ( .a(n_18771), .o(n_18772) );
no02s01 g762212 ( .a(n_18734), .b(n_45003), .o(n_18771) );
na02s01 g762213 ( .a(n_18734), .b(n_45003), .o(n_18817) );
na02m04 g762214 ( .a(n_18445), .b(n_18501), .o(n_18703) );
na02m04 TIMEBOOST_cell_7714 ( .a(n_29527), .b(FE_OFN775_n_25834), .o(TIMEBOOST_net_2488) );
na02s02 g762216 ( .a(n_18615), .b(n_19400), .o(n_18776) );
na02s02 g762218 ( .a(n_18663), .b(n_18586), .o(n_18739) );
in01m02 g762220 ( .a(n_18731), .o(n_18814) );
no02s04 g762221 ( .a(n_18698), .b(n_18536), .o(n_18731) );
in01s02 g762222 ( .a(n_18164), .o(n_18165) );
in01m02 g762224 ( .a(n_18188), .o(n_18189) );
no02m02 TIMEBOOST_cell_6055 ( .a(n_2359), .b(n_2273), .o(TIMEBOOST_net_1879) );
no02m01 TIMEBOOST_cell_5663 ( .a(TIMEBOOST_net_1779), .b(n_17120), .o(n_17190) );
na02s01 g762228 ( .a(n_18114), .b(n_18079), .o(n_18179) );
in01s01 g762229 ( .a(n_18149), .o(n_18150) );
na02s01 g762230 ( .a(n_18092), .b(n_18136), .o(n_18149) );
in01m02 g762231 ( .a(n_18148), .o(n_18190) );
na02m03 g762232 ( .a(n_18135), .b(n_17946), .o(n_18148) );
na02s06 g762233 ( .a(n_18135), .b(n_18133), .o(n_18134) );
in01m02 g762234 ( .a(n_18187), .o(n_18214) );
na02m04 g762235 ( .a(n_18163), .b(delay_add_ln22_unr11_stage5_stallmux_q_16_), .o(n_18187) );
no02m04 g762236 ( .a(n_18163), .b(delay_add_ln22_unr11_stage5_stallmux_q_16_), .o(n_18215) );
in01s02 g762237 ( .a(n_18238), .o(n_18239) );
na02m02 g762238 ( .a(n_18213), .b(n_18186), .o(n_18238) );
na02s10 g762241 ( .a(n_18096), .b(FE_RN_235_0), .o(n_18113) );
na02m01 g762242 ( .a(n_18451), .b(n_17427), .o(n_18501) );
no02s01 g762243 ( .a(n_18835), .b(n_18834), .o(n_18836) );
na02s01 g762245 ( .a(n_18578), .b(n_18580), .o(n_18587) );
no02s01 g762246 ( .a(n_18453), .b(n_18585), .o(n_18586) );
no02s01 g762247 ( .a(n_18496), .b(n_18694), .o(n_18663) );
in01s01 g762249 ( .a(n_18696), .o(n_18697) );
na02s01 g762250 ( .a(n_18608), .b(n_18657), .o(n_18696) );
in01s01 g762251 ( .a(n_18661), .o(n_18735) );
na02s02 g762252 ( .a(n_18579), .b(n_18622), .o(n_18661) );
na02s01 g762254 ( .a(n_18728), .b(n_18729), .o(n_18730) );
na02s01 g762256 ( .a(n_18535), .b(n_18534), .o(n_18536) );
in01m02 g762257 ( .a(n_18619), .o(n_18698) );
no02s02 g762258 ( .a(n_18584), .b(n_18583), .o(n_18619) );
na02s01 g762259 ( .a(n_18616), .b(n_18617), .o(n_18618) );
no02s01 g762260 ( .a(n_18523), .b(n_18497), .o(n_18615) );
no02s01 g762261 ( .a(n_18726), .b(n_18725), .o(n_18767) );
no02s01 g762262 ( .a(n_18499), .b(n_18498), .o(n_18500) );
na02s01 g762263 ( .a(n_18582), .b(n_18495), .o(n_19485) );
na02s01 g762264 ( .a(n_18522), .b(n_18581), .o(n_19520) );
no02s01 g762265 ( .a(n_18766), .b(n_18585), .o(n_19541) );
in01s01 g762266 ( .a(n_18818), .o(n_18695) );
no02s01 g762267 ( .a(n_18660), .b(n_45003), .o(n_18818) );
na02s01 g762268 ( .a(n_18840), .b(n_18611), .o(n_19491) );
na02s01 g762269 ( .a(n_18810), .b(n_18809), .o(n_19292) );
na02s01 g762270 ( .a(n_45003), .b(n_18660), .o(n_18816) );
na02s01 g762271 ( .a(n_18622), .b(n_18614), .o(n_18845) );
na02s01 g762272 ( .a(n_18727), .b(n_18665), .o(n_19523) );
no02s01 g762273 ( .a(n_18693), .b(n_18528), .o(n_19547) );
no02s01 g762274 ( .a(n_18723), .b(n_18769), .o(n_19295) );
no02s01 g762275 ( .a(n_18692), .b(n_18765), .o(n_19575) );
na02s01 g762276 ( .a(n_45002), .b(n_18414), .o(n_18624) );
na02s01 g762277 ( .a(n_18535), .b(n_18659), .o(n_19228) );
na02s01 g762278 ( .a(n_18620), .b(n_18580), .o(n_18993) );
na02s01 g762279 ( .a(n_18534), .b(n_18658), .o(n_19193) );
no02s01 g762280 ( .a(n_18584), .b(n_18609), .o(n_19159) );
na02s01 g762281 ( .a(n_45003), .b(n_18415), .o(n_18813) );
no02s01 g762282 ( .a(n_18835), .b(n_18569), .o(n_19572) );
na02s01 g762283 ( .a(n_18617), .b(n_18729), .o(n_19231) );
no02s01 g762284 ( .a(n_18613), .b(n_18524), .o(n_19019) );
na02s01 g762285 ( .a(n_18579), .b(n_18578), .o(n_18968) );
na02s01 g762286 ( .a(n_18446), .b(n_18701), .o(n_18667) );
no02s01 g762287 ( .a(n_18444), .b(n_18452), .o(n_18626) );
no02s01 g762288 ( .a(n_18834), .b(n_18490), .o(n_19544) );
na02s01 g762289 ( .a(n_18808), .b(n_18575), .o(n_19488) );
no02s01 g762290 ( .a(n_18607), .b(n_18694), .o(n_19367) );
na02s01 g762291 ( .a(n_18532), .b(n_18657), .o(n_19070) );
no02s01 g762292 ( .a(n_18498), .b(n_18450), .o(n_18779) );
na02s01 g762293 ( .a(n_18616), .b(n_18728), .o(n_19196) );
oa12s10 g762294 ( .a(n_18060), .b(n_18008), .c(FE_OCP_RBN2436_FE_OCPN833_n_45450), .o(n_18176) );
oa12m06 g762295 ( .a(n_18025), .b(n_18009), .c(FE_OCP_RBN2436_FE_OCPN833_n_45450), .o(n_18173) );
in01s01 g762296 ( .a(n_18138), .o(n_18095) );
oa12f08 g762297 ( .a(n_17999), .b(n_18080), .c(n_17952), .o(n_18138) );
oa12f08 g762298 ( .a(n_18015), .b(n_18130), .c(n_17964), .o(n_18194) );
in01s01 g762299 ( .a(FE_OCP_DRV_N1460_n_18111), .o(n_18112) );
oa12s01 g762300 ( .a(n_18058), .b(n_18080), .c(n_18057), .o(n_18111) );
in01s02 g762301 ( .a(n_18161), .o(n_18162) );
na02m08 TIMEBOOST_cell_6604 ( .a(TIMEBOOST_net_2059), .b(n_22964), .o(n_23100) );
na02m08 g762303 ( .a(n_18059), .b(n_18061), .o(n_18153) );
ao22s01 g762304 ( .a(n_18087), .b(n_18036), .c(n_18130), .d(n_18037), .o(n_19751) );
ao12s01 g762305 ( .a(n_18387), .b(n_18386), .c(n_18385), .o(n_18773) );
oa12s01 g762306 ( .a(n_18384), .b(n_18383), .c(n_18382), .o(n_18734) );
no02m04 g762307 ( .a(n_18093), .b(n_18054), .o(n_18167) );
no02s08 TIMEBOOST_cell_1716 ( .a(TIMEBOOST_net_472), .b(n_38901), .o(n_39053) );
na02s02 g762309 ( .a(n_18074), .b(n_17945), .o(n_18110) );
no02s02 TIMEBOOST_cell_6228 ( .a(TIMEBOOST_net_1965), .b(n_3777), .o(n_4008) );
oa12s02 g762311 ( .a(n_18001), .b(n_17971), .c(n_18052), .o(n_18059) );
in01s01 g762312 ( .a(n_18078), .o(n_18079) );
no02s06 g762313 ( .a(n_18056), .b(n_18055), .o(n_18078) );
na02m02 TIMEBOOST_cell_8655 ( .a(TIMEBOOST_net_2814), .b(n_36732), .o(n_36748) );
na02s01 g762315 ( .a(n_18080), .b(n_18057), .o(n_18058) );
na02s06 g762316 ( .a(n_18056), .b(n_18055), .o(n_18114) );
in01s01 g762317 ( .a(n_18091), .o(n_18092) );
no02m08 g762318 ( .a(n_18077), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_12_), .o(n_18091) );
na02m08 g762319 ( .a(n_18077), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_12_), .o(n_18136) );
no02m08 g762320 ( .a(n_18090), .b(n_17920), .o(n_18135) );
na02s06 g762321 ( .a(n_18160), .b(n_18159), .o(n_18213) );
in01m01 g762322 ( .a(n_18185), .o(n_18186) );
no02s06 g762323 ( .a(n_18160), .b(n_18159), .o(n_18185) );
in01s02 g762324 ( .a(n_18128), .o(n_18129) );
na02s02 g762325 ( .a(n_18072), .b(n_18109), .o(n_18128) );
in01m01 g762326 ( .a(n_18198), .o(n_18199) );
na02m02 g762327 ( .a(n_18126), .b(n_18146), .o(n_18198) );
no02s01 TIMEBOOST_cell_1651 ( .a(n_4307), .b(n_3297), .o(TIMEBOOST_net_440) );
in01s06 g762329 ( .a(n_18096), .o(n_18115) );
in01m10 g762331 ( .a(n_18025), .o(n_18026) );
na02m20 g762332 ( .a(n_18009), .b(FE_OCP_RBN2436_FE_OCPN833_n_45450), .o(n_18025) );
na02s40 g762333 ( .a(n_18008), .b(FE_OCP_RBN2436_FE_OCPN833_n_45450), .o(n_18060) );
no02s01 g762334 ( .a(n_18386), .b(n_18385), .o(n_18387) );
na02s01 g762335 ( .a(n_18383), .b(n_18382), .o(n_18384) );
in01s01 g762336 ( .a(n_18075), .o(n_18076) );
na02s10 g762337 ( .a(n_18006), .b(n_18050), .o(n_18075) );
in01s01 g762338 ( .a(n_18834), .o(n_18807) );
no02s01 g762339 ( .a(n_45002), .b(n_18441), .o(n_18834) );
in01s01 g762340 ( .a(n_18453), .o(n_18581) );
no02s01 g762341 ( .a(FE_OCP_RBN2517_n_45120), .b(n_18422), .o(n_18453) );
in01s01 g762342 ( .a(n_18451), .o(n_18452) );
na02m01 g762343 ( .a(n_18421), .b(n_18418), .o(n_18451) );
in01s01 g762344 ( .a(n_18726), .o(n_18727) );
no02s01 g762345 ( .a(n_18526), .b(n_45002), .o(n_18726) );
in01s01 g762346 ( .a(n_18725), .o(n_18808) );
no02s01 g762347 ( .a(n_45002), .b(n_18529), .o(n_18725) );
in01s01 g762348 ( .a(n_18497), .o(n_18582) );
no02s01 g762349 ( .a(n_45120), .b(n_18448), .o(n_18497) );
no02s01 g762350 ( .a(n_18521), .b(n_45002), .o(n_18835) );
no02s01 g762351 ( .a(n_18252), .b(n_45002), .o(n_18766) );
in01s01 g762352 ( .a(n_18449), .o(n_18450) );
na02s01 g762353 ( .a(n_18421), .b(n_18419), .o(n_18449) );
in01s01 g762354 ( .a(n_18495), .o(n_18496) );
na02s01 g762355 ( .a(n_45120), .b(n_18448), .o(n_18495) );
in01s01 g762356 ( .a(n_18578), .o(n_18533) );
na02s02 g762357 ( .a(FE_OCP_RBN2515_n_45120), .b(n_17860), .o(n_18578) );
in01s01 g762358 ( .a(n_18583), .o(n_18532) );
no02s02 g762359 ( .a(FE_OCP_RBN2515_n_45120), .b(n_18494), .o(n_18583) );
na02s02 g762360 ( .a(FE_OCP_RBN2515_n_45120), .b(n_17883), .o(n_18580) );
na02s01 g762361 ( .a(n_45118), .b(n_17859), .o(n_18579) );
in01s01 g762362 ( .a(n_18616), .o(n_18577) );
na02s01 g762363 ( .a(n_45002), .b(n_18531), .o(n_18616) );
na02s01 g762364 ( .a(n_45002), .b(n_18102), .o(n_18617) );
in01s01 g762365 ( .a(n_18839), .o(n_18693) );
na02s01 g762366 ( .a(n_18492), .b(n_45003), .o(n_18839) );
in01s01 g762367 ( .a(n_18612), .o(n_18613) );
na02s01 g762368 ( .a(FE_OCP_RBN2515_n_45120), .b(n_18488), .o(n_18612) );
no02s01 g762369 ( .a(n_45002), .b(n_18689), .o(n_18769) );
in01s01 g762370 ( .a(n_18841), .o(n_18692) );
na02s01 g762371 ( .a(n_18572), .b(n_45003), .o(n_18841) );
in01s01 g762372 ( .a(n_18575), .o(n_18576) );
na02s01 g762373 ( .a(n_45118), .b(n_18529), .o(n_18575) );
in01s01 g762374 ( .a(n_18737), .o(n_18611) );
no02s01 g762375 ( .a(n_45003), .b(n_18574), .o(n_18737) );
no02s01 g762376 ( .a(n_18572), .b(n_45003), .o(n_18765) );
in01s01 g762377 ( .a(n_18528), .o(n_18623) );
no02s01 g762378 ( .a(FE_OCP_RBN2517_n_45120), .b(n_18492), .o(n_18528) );
no02s01 g762379 ( .a(FE_OCP_RBN2517_n_45120), .b(n_18251), .o(n_18585) );
no02s01 g762380 ( .a(FE_OCP_RBN2517_n_45120), .b(n_18420), .o(n_18694) );
in01s01 g762381 ( .a(n_18665), .o(n_18571) );
na02s01 g762382 ( .a(n_18526), .b(n_45118), .o(n_18665) );
in01s01 g762383 ( .a(n_18664), .o(n_18490) );
na02s01 g762384 ( .a(n_45118), .b(n_18441), .o(n_18664) );
in01s01 g762385 ( .a(n_18724), .o(n_18809) );
no02s01 g762386 ( .a(n_45002), .b(n_18688), .o(n_18724) );
na02s01 g762387 ( .a(FE_OCP_RBN2515_n_45120), .b(n_18065), .o(n_18659) );
in01s01 g762388 ( .a(n_18658), .o(n_18610) );
na02s01 g762389 ( .a(FE_OCP_RBN2515_n_45120), .b(n_18416), .o(n_18658) );
in01s01 g762390 ( .a(n_18608), .o(n_18609) );
na02s01 g762391 ( .a(FE_OCP_RBN2515_n_45120), .b(n_18487), .o(n_18608) );
na02s01 g762392 ( .a(FE_OCP_RBN2515_n_45120), .b(n_18494), .o(n_18657) );
na02s01 g762393 ( .a(n_45118), .b(n_17785), .o(n_18622) );
no02s01 g762395 ( .a(FE_OCP_RBN2515_n_45120), .b(n_18488), .o(n_18524) );
na02s01 g762396 ( .a(n_45118), .b(n_17882), .o(n_18620) );
in01s01 g762397 ( .a(n_18499), .o(n_18446) );
no02s01 g762398 ( .a(n_18421), .b(n_18417), .o(n_18499) );
no02s01 g762399 ( .a(n_18421), .b(n_18419), .o(n_18498) );
in01s01 g762400 ( .a(n_18444), .o(n_18445) );
no02s01 g762401 ( .a(n_18421), .b(n_18418), .o(n_18444) );
na02s01 g762402 ( .a(n_18421), .b(n_18417), .o(n_18701) );
na02s02 g762403 ( .a(FE_OCP_RBN2515_n_45120), .b(n_17786), .o(n_18614) );
na02s01 g762404 ( .a(n_45003), .b(n_18103), .o(n_18729) );
in01s01 g762405 ( .a(n_18655), .o(n_18728) );
no02s01 g762406 ( .a(n_45002), .b(n_18531), .o(n_18655) );
in01s01 g762407 ( .a(n_18722), .o(n_18723) );
na02s01 g762408 ( .a(n_45002), .b(n_18689), .o(n_18722) );
no02s02 g762409 ( .a(FE_OCP_RBN2515_n_45120), .b(n_18487), .o(n_18584) );
na02s01 g762410 ( .a(n_45003), .b(n_18574), .o(n_18840) );
in01s01 g762411 ( .a(n_19400), .o(n_18607) );
na02s01 g762412 ( .a(FE_OCP_RBN2517_n_45120), .b(n_18420), .o(n_19400) );
in01s01 g762413 ( .a(n_18522), .o(n_18523) );
na02s01 g762414 ( .a(FE_OCP_RBN2517_n_45120), .b(n_18422), .o(n_18522) );
in01s01 g762415 ( .a(n_18443), .o(n_18534) );
no02s01 g762416 ( .a(n_18421), .b(n_18416), .o(n_18443) );
in01s01 g762417 ( .a(n_18568), .o(n_18569) );
na02s02 g762418 ( .a(n_45118), .b(n_18521), .o(n_18568) );
na02s01 g762419 ( .a(n_45120), .b(n_18064), .o(n_18535) );
na02s01 g762420 ( .a(n_45002), .b(n_18688), .o(n_18810) );
in01m02 g762421 ( .a(n_18023), .o(n_18024) );
ao12m08 g762422 ( .a(n_17977), .b(FE_OCP_RBN2435_FE_OCPN833_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_15_), .o(n_18023) );
in01s01 g762423 ( .a(n_18414), .o(n_18415) );
ao12s02 g762424 ( .a(n_18328), .b(n_18327), .c(n_18326), .o(n_18414) );
oa12s01 g762425 ( .a(n_18352), .b(n_18351), .c(n_18350), .o(n_18660) );
na03m04 TIMEBOOST_cell_8248 ( .a(n_7692), .b(n_7728), .c(n_7704), .o(n_7820) );
in01m20 g762427 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_17_), .o(n_18009) );
in01s40 g762429 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_18_), .o(n_18008) );
in01s01 g762431 ( .a(n_18090), .o(n_18074) );
na02m08 g762432 ( .a(n_18021), .b(n_17873), .o(n_18090) );
in01s03 g762433 ( .a(n_18005), .o(n_18006) );
no02s20 g762434 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_19_), .b(FE_OCP_RBN2438_FE_OCPN833_n_45450), .o(n_18005) );
na02m01 g762435 ( .a(n_18021), .b(n_17919), .o(n_18089) );
na03s02 TIMEBOOST_cell_7164 ( .a(n_7718), .b(n_8389), .c(n_7777), .o(n_7875) );
in01s01 g762438 ( .a(n_18127), .o(n_18146) );
no02m08 g762439 ( .a(n_18106), .b(delay_add_ln22_unr11_stage5_stallmux_q_14_), .o(n_18127) );
na02s03 g762440 ( .a(n_18049), .b(n_18048), .o(n_18109) );
in01s01 g762441 ( .a(n_18071), .o(n_18072) );
no02s04 g762442 ( .a(n_18049), .b(n_18048), .o(n_18071) );
in01s01 g762443 ( .a(n_18107), .o(n_18108) );
na02s01 g762444 ( .a(n_18046), .b(n_18088), .o(n_18107) );
na02s06 g762448 ( .a(n_18106), .b(delay_add_ln22_unr11_stage5_stallmux_q_14_), .o(n_18126) );
na02s01 g762449 ( .a(n_18351), .b(n_18350), .o(n_18352) );
no02m20 g762452 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_15_), .b(FE_OCP_RBN2435_FE_OCPN833_n_45450), .o(n_17977) );
na02s06 g762453 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_19_), .b(FE_OCP_RBN2438_FE_OCPN833_n_45450), .o(n_18050) );
in01s02 g762454 ( .a(n_18003), .o(n_18004) );
ao12s06 g762455 ( .a(n_17975), .b(FE_OCP_RBN2435_FE_OCPN833_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_14_), .o(n_18003) );
in01s06 g762456 ( .a(n_18001), .o(n_18002) );
ao12s10 g762457 ( .a(n_18051), .b(FE_OCPN6277_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_13_), .o(n_18001) );
ao12s06 g762459 ( .a(n_18137), .b(FE_OCP_RBN2435_FE_OCPN833_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_16_), .o(n_17973) );
no02s01 g762460 ( .a(n_18327), .b(n_18326), .o(n_18328) );
oa12f08 g762461 ( .a(n_17896), .b(n_18000), .c(n_17849), .o(n_18080) );
in01s01 g762462 ( .a(n_18130), .o(n_18087) );
oa12f08 g762463 ( .a(n_17966), .b(n_18070), .c(n_17912), .o(n_18130) );
ao12s01 g762464 ( .a(n_17710), .b(n_45524), .c(n_17611), .o(n_18386) );
no03f04 TIMEBOOST_cell_2430 ( .a(n_19078), .b(FE_OCP_RBN5617_n_18899), .c(n_19147), .o(n_19243) );
ao22s01 g762598 ( .a(n_18000), .b(n_17925), .c(n_17949), .d(n_17924), .o(n_19590) );
oa12s01 g762599 ( .a(n_18042), .b(n_18070), .c(n_18041), .o(n_19665) );
oa12s01 g762600 ( .a(n_18295), .b(n_18294), .c(n_18293), .o(n_18572) );
ao12s01 g762601 ( .a(n_17709), .b(n_45524), .c(n_17531), .o(n_18383) );
oa22s01 g762603 ( .a(n_18253), .b(n_17707), .c(n_18254), .d(n_17706), .o(n_18492) );
no02s02 g762608 ( .a(n_18039), .b(n_17950), .o(n_18069) );
no02f04 TIMEBOOST_cell_7968 ( .a(n_30598), .b(TIMEBOOST_net_1286), .o(TIMEBOOST_net_2615) );
no02s01 g762610 ( .a(n_45524), .b(n_17734), .o(n_18351) );
no02s40 g762611 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_14_), .b(FE_OCP_RBN2435_FE_OCPN833_n_45450), .o(n_17975) );
in01s01 g762612 ( .a(n_18045), .o(n_18046) );
no02s06 g762613 ( .a(n_18022), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_10_), .o(n_18045) );
na02s06 g762614 ( .a(n_18022), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_10_), .o(n_18088) );
no02s06 g762615 ( .a(n_17971), .b(n_17970), .o(n_17972) );
in01s01 g762617 ( .a(n_18021), .o(n_18043) );
na02s01 g762619 ( .a(n_17999), .b(n_17953), .o(n_18057) );
no02s20 g762620 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_16_), .b(FE_OCP_RBN2435_FE_OCPN833_n_45450), .o(n_18137) );
na02s01 g762621 ( .a(n_18070), .b(n_18041), .o(n_18042) );
in01s01 g762622 ( .a(n_18124), .o(n_18125) );
na02s01 g762623 ( .a(n_18105), .b(n_18068), .o(n_18124) );
no02s40 g762624 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_13_), .b(FE_OCP_RBN2435_FE_OCPN833_n_45450), .o(n_18051) );
na02s01 g762625 ( .a(n_18294), .b(n_18293), .o(n_18295) );
oa12s02 g762627 ( .a(n_17608), .b(n_45529), .c(n_17605), .o(n_18327) );
ao22s02 g762630 ( .a(n_17914), .b(n_17916), .c(FE_OCP_RBN5551_n_17914), .d(n_17915), .o(n_18049) );
ao12s01 g762631 ( .a(n_18257), .b(n_18256), .c(n_18255), .o(n_18521) );
ao22s02 g762632 ( .a(n_18232), .b(n_17704), .c(n_18231), .d(n_17705), .o(n_18526) );
in01s01 g762635 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_30_), .o(n_17856) );
na02s06 g762640 ( .a(n_17932), .b(n_17931), .o(n_17999) );
in01s01 g762641 ( .a(n_17952), .o(n_17953) );
no02s06 g762642 ( .a(n_17932), .b(n_17931), .o(n_17952) );
no02m02 TIMEBOOST_cell_1631 ( .a(FE_OCP_RBN4146_n_7743), .b(n_8870), .o(TIMEBOOST_net_430) );
in01s02 g762647 ( .a(n_18039), .o(n_18040) );
na02s02 g762648 ( .a(n_18020), .b(n_17917), .o(n_18039) );
na02s03 g762649 ( .a(n_18020), .b(n_18018), .o(n_18019) );
na02m06 g762650 ( .a(n_18038), .b(delay_add_ln22_unr11_stage5_stallmux_q_12_), .o(n_18105) );
in01s01 g762651 ( .a(n_18067), .o(n_18068) );
no02m06 g762652 ( .a(n_18038), .b(delay_add_ln22_unr11_stage5_stallmux_q_12_), .o(n_18067) );
na02s01 g762653 ( .a(n_18017), .b(n_18066), .o(n_18168) );
no02s01 g762654 ( .a(n_45528), .b(n_17607), .o(n_18294) );
no02s01 g762655 ( .a(n_18256), .b(n_18255), .o(n_18257) );
ao12s03 g762657 ( .a(n_17851), .b(FE_OCPN6277_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_11_), .o(n_17897) );
ao12s10 g762658 ( .a(n_18052), .b(FE_OCPN6277_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_12_), .o(n_17970) );
in01s01 g762659 ( .a(n_17950), .o(n_17951) );
ao12s01 g762660 ( .a(n_17929), .b(FE_OCPN836_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_15_), .o(n_17950) );
in01s01 g762661 ( .a(n_18253), .o(n_18254) );
oa12s01 g762662 ( .a(n_17353), .b(n_18237), .c(n_17572), .o(n_18253) );
in01s01 g762664 ( .a(n_18000), .o(n_17949) );
oa12f08 g762665 ( .a(n_17870), .b(n_17928), .c(n_17822), .o(n_18000) );
oa12f08 g762666 ( .a(n_17906), .b(n_17997), .c(n_17866), .o(n_18070) );
in01s01 g762669 ( .a(FE_OCPN1290_n_19384), .o(n_19508) );
ao12s01 g762670 ( .a(n_17927), .b(n_17928), .c(n_17926), .o(n_19384) );
ao22s01 g762671 ( .a(n_17997), .b(n_17941), .c(n_17943), .d(n_17940), .o(n_19562) );
oa12s01 g762672 ( .a(n_18212), .b(n_18237), .c(n_18211), .o(n_18574) );
ao12s01 g762673 ( .a(n_18236), .b(n_18235), .c(n_18234), .o(n_18441) );
in01s01 g762675 ( .a(n_18251), .o(n_18252) );
oa22s02 g762676 ( .a(n_18183), .b(n_17703), .c(n_18184), .d(n_17702), .o(n_18251) );
in01s01 g762678 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_31_), .o(n_17852) );
no02s01 g762680 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_24_), .b(delay_add_ln22_unr11_stage5_stallmux_q_25_), .o(n_17813) );
no02s01 g762681 ( .a(n_17928), .b(n_17926), .o(n_17927) );
in01s01 g762682 ( .a(n_17924), .o(n_17925) );
na02s01 g762683 ( .a(n_17850), .b(n_17896), .o(n_17924) );
in01s03 g762684 ( .a(n_17851), .o(n_17930) );
no02f03 g762685 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_11_), .b(FE_OCPN867_n_45450), .o(n_17851) );
in01s02 g762686 ( .a(n_17895), .o(n_17923) );
in01s02 g762688 ( .a(n_18052), .o(n_17893) );
no02s40 g762689 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_12_), .b(FE_OCPN867_n_45450), .o(n_18052) );
no02m04 g762690 ( .a(FE_OCP_RBN5550_n_17914), .b(n_17967), .o(n_18020) );
no02f03 g762691 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_15_), .b(FE_OCPN6277_n_45450), .o(n_17929) );
na02s06 g762692 ( .a(n_17996), .b(n_17995), .o(n_18066) );
in01s01 g762693 ( .a(n_18016), .o(n_18017) );
no02m06 g762694 ( .a(n_17996), .b(n_17995), .o(n_18016) );
in01s01 g762695 ( .a(n_17947), .o(n_17948) );
na02m03 g762696 ( .a(n_17921), .b(n_17922), .o(n_17947) );
na02s01 g762697 ( .a(n_18237), .b(n_18211), .o(n_18212) );
no02s01 g762698 ( .a(n_18235), .b(n_18234), .o(n_18236) );
oa12m03 g762699 ( .a(n_17946), .b(n_17892), .c(FE_OCP_RBN2436_FE_OCPN833_n_45450), .o(n_18133) );
in01s01 g762700 ( .a(n_17944), .o(n_17945) );
ao12s02 g762701 ( .a(n_17920), .b(FE_OCP_RBN2435_FE_OCPN833_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_17_), .o(n_17944) );
in01m01 g762702 ( .a(n_17918), .o(n_17919) );
ao12m02 g762703 ( .a(n_17872), .b(FE_OCPN836_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_16_), .o(n_17918) );
oa12s02 g762704 ( .a(n_17917), .b(n_17875), .c(FE_OCP_RBN2436_FE_OCPN833_n_45450), .o(n_18018) );
in01s02 g762705 ( .a(n_17915), .o(n_17916) );
ao12s03 g762706 ( .a(n_17967), .b(FE_OCPN6277_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_13_), .o(n_17915) );
in01s01 g762709 ( .a(n_18231), .o(n_18232) );
oa12s01 g762710 ( .a(n_17155), .b(n_18210), .c(n_17309), .o(n_18231) );
in01s01 g762715 ( .a(n_17812), .o(n_17809) );
ao22s01 g762718 ( .a(n_18210), .b(n_17356), .c(n_18157), .d(n_17357), .o(n_18529) );
oa22s01 g762720 ( .a(n_17632), .b(n_17539), .c(n_18197), .d(n_17358), .o(n_18256) );
in01s01 g762722 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_25_), .o(n_18331) );
in01s01 g762724 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_26_), .o(n_17806) );
in01s01 g762726 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_28_), .o(n_17805) );
na03f02 TIMEBOOST_cell_8294 ( .a(TIMEBOOST_net_2464), .b(n_14612), .c(n_45520), .o(n_14818) );
na02s06 g762732 ( .a(n_17827), .b(n_17779), .o(n_17828) );
na02s06 g762735 ( .a(n_17826), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_8_), .o(n_17896) );
in01s01 g762736 ( .a(n_17849), .o(n_17850) );
no02s06 g762737 ( .a(n_17826), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_8_), .o(n_17849) );
na02m03 g762738 ( .a(n_17824), .b(FE_OCP_RBN2436_FE_OCPN833_n_45450), .o(n_17921) );
na02s06 g762739 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_19_), .b(FE_OCP_RBN2437_FE_OCPN833_n_45450), .o(n_17922) );
na02s40 g762740 ( .a(n_17892), .b(FE_OCP_RBN2436_FE_OCPN833_n_45450), .o(n_17946) );
in01s06 g762741 ( .a(n_17917), .o(n_17891) );
na02s40 g762742 ( .a(n_17875), .b(FE_OCP_RBN2436_FE_OCPN833_n_45450), .o(n_17917) );
no02s40 g762743 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_13_), .b(FE_OCPN867_n_45450), .o(n_17967) );
in01m08 g762744 ( .a(n_17872), .o(n_17873) );
no02m20 g762745 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_16_), .b(FE_OCPN836_n_45450), .o(n_17872) );
no02m03 g762746 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_17_), .b(FE_OCP_RBN2435_FE_OCPN833_n_45450), .o(n_17920) );
in01s01 g762747 ( .a(n_18036), .o(n_18037) );
na02s01 g762748 ( .a(n_18015), .b(n_17965), .o(n_18036) );
na02s01 g762749 ( .a(n_17913), .b(n_17966), .o(n_18041) );
na02s01 g762750 ( .a(n_18197), .b(n_17615), .o(n_18235) );
in01s06 g762751 ( .a(n_17847), .o(n_17848) );
ao12s03 g762752 ( .a(n_17825), .b(FE_OCPN1202_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_10_), .o(n_17847) );
in01s01 g762753 ( .a(n_18183), .o(n_18184) );
oa12s01 g762754 ( .a(n_17261), .b(n_18158), .c(n_17260), .o(n_18183) );
oa12f08 g762755 ( .a(n_17766), .b(n_17846), .c(n_17718), .o(n_17928) );
in01s01 g762756 ( .a(n_17997), .o(n_17943) );
no02s01 TIMEBOOST_cell_3985 ( .a(n_42468), .b(n_42419), .o(TIMEBOOST_net_1083) );
oa12f08 g762758 ( .a(n_17540), .b(n_18156), .c(n_17633), .o(n_18237) );
in01s01 g762759 ( .a(n_17811), .o(n_17781) );
in01s02 g762761 ( .a(n_17834), .o(n_17803) );
oa12s01 g762764 ( .a(n_17911), .b(n_17910), .c(n_17909), .o(n_19436) );
oa12s01 g762765 ( .a(n_18142), .b(n_18158), .c(n_18141), .o(n_18422) );
oa22s01 g762766 ( .a(n_17799), .b(n_17794), .c(n_17846), .d(n_17795), .o(n_19314) );
in01s06 g762767 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_19_), .o(n_17824) );
in01s40 g762769 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_18_), .o(n_17892) );
in01s40 g762771 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_14_), .o(n_17875) );
no02s04 g762776 ( .a(n_17889), .b(n_17888), .o(n_17890) );
in01s01 g762777 ( .a(n_18157), .o(n_18210) );
na02s01 g762778 ( .a(n_18123), .b(n_17502), .o(n_18157) );
in01m01 g762779 ( .a(n_17825), .o(n_17802) );
no02s40 g762780 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_10_), .b(FE_OCPN1202_n_45450), .o(n_17825) );
na02s01 g762781 ( .a(n_17720), .b(n_17894), .o(n_17780) );
in01s01 g762784 ( .a(n_17964), .o(n_17965) );
no02m06 g762785 ( .a(n_17942), .b(delay_add_ln22_unr11_stage5_stallmux_q_10_), .o(n_17964) );
na02s06 g762786 ( .a(n_17887), .b(n_17886), .o(n_17966) );
in01s01 g762787 ( .a(n_17912), .o(n_17913) );
no02m06 g762788 ( .a(n_17887), .b(n_17886), .o(n_17912) );
na02s02 TIMEBOOST_cell_5264 ( .a(n_24574), .b(n_24395), .o(TIMEBOOST_net_1580) );
na02m06 g762790 ( .a(n_17942), .b(delay_add_ln22_unr11_stage5_stallmux_q_10_), .o(n_18015) );
na02s01 g762791 ( .a(n_17870), .b(n_17823), .o(n_17926) );
na02s01 g762792 ( .a(n_18156), .b(n_17614), .o(n_18197) );
na02s01 g762793 ( .a(n_17910), .b(n_17909), .o(n_17911) );
na02s01 g762794 ( .a(n_18158), .b(n_18141), .o(n_18142) );
in01s01 g762795 ( .a(n_17778), .o(n_17779) );
ao12m03 g762796 ( .a(n_17758), .b(FE_OCPN1202_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_9_), .o(n_17778) );
in01s02 g762797 ( .a(n_17868), .o(n_17869) );
ao12s03 g762798 ( .a(n_17845), .b(FE_OCPN6277_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_12_), .o(n_17868) );
in01s01 g762804 ( .a(n_17782), .o(n_17756) );
oa12s02 g762808 ( .a(n_17323), .b(n_17659), .c(n_16996), .o(n_17660) );
ao12s06 g762809 ( .a(n_17388), .b(n_17694), .c(n_17035), .o(n_17695) );
oa12s06 g762810 ( .a(n_17235), .b(n_17694), .c(n_17120), .o(n_17693) );
ao12s02 g762811 ( .a(n_17195), .b(n_17659), .c(n_17174), .o(n_17658) );
ao12s01 g762812 ( .a(n_18085), .b(n_18084), .c(n_18083), .o(n_18448) );
ao12s06 g762813 ( .a(n_17727), .b(n_17656), .c(n_17726), .o(n_17826) );
in01s01 g762814 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_23_), .o(n_17692) );
in01s01 g762816 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_24_), .o(n_18329) );
no02s01 g762820 ( .a(n_17700), .b(n_17772), .o(n_17773) );
in01m03 g762821 ( .a(n_17758), .o(n_17894) );
no02s40 g762822 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_9_), .b(FE_OCPN1296_n_45450), .o(n_17758) );
na02s06 g762824 ( .a(n_17801), .b(n_17800), .o(n_17870) );
in01s01 g762825 ( .a(n_17822), .o(n_17823) );
no02s06 g762826 ( .a(n_17801), .b(n_17800), .o(n_17822) );
in01s04 g762827 ( .a(n_17907), .o(n_17908) );
no02s06 g762828 ( .a(n_17889), .b(n_17885), .o(n_17907) );
no02s40 g762829 ( .a(FE_OCPN867_n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_12_), .o(n_17845) );
in01m06 g762830 ( .a(n_18123), .o(n_18156) );
na02f08 g762831 ( .a(n_18104), .b(n_17470), .o(n_18123) );
in01s01 g762832 ( .a(n_17940), .o(n_17941) );
na02s01 g762833 ( .a(n_17906), .b(n_17867), .o(n_17940) );
no02m01 g762834 ( .a(n_18104), .b(n_17469), .o(n_18158) );
no02s01 g762835 ( .a(n_18084), .b(n_18083), .o(n_18085) );
na02s02 g762836 ( .a(n_17597), .b(n_17135), .o(n_17629) );
no02s02 g762837 ( .a(n_17598), .b(n_17036), .o(n_17657) );
ao12s06 g762838 ( .a(n_17885), .b(FE_OCPN6277_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_11_), .o(n_17888) );
in01s01 g762839 ( .a(n_17846), .o(n_17799) );
oa12f08 g762840 ( .a(n_17672), .b(n_17622), .c(n_17771), .o(n_17846) );
in01s01 g762841 ( .a(n_17843), .o(n_17910) );
ao12f08 g762842 ( .a(n_17740), .b(n_17839), .c(n_17791), .o(n_17843) );
ao12m04 g762851 ( .a(n_17798), .b(n_17797), .c(n_17796), .o(n_17887) );
ao12s01 g762852 ( .a(n_17747), .b(n_17771), .c(n_17746), .o(n_19138) );
ao12s01 g762853 ( .a(n_17840), .b(n_17839), .c(n_17838), .o(n_19354) );
in01s01 g762855 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_30_), .o(n_17749) );
in01s01 g762857 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_28_), .o(n_17696) );
in01s01 g762859 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_31_), .o(n_17724) );
in01s01 g762863 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_29_), .o(n_17748) );
in01s01 g762865 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_), .o(n_17700) );
in01s01 g762867 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_26_), .o(n_17722) );
no02m04 g762869 ( .a(n_17797), .b(n_17796), .o(n_17798) );
in01s02 g762870 ( .a(n_17720), .o(n_17721) );
in01s06 g762872 ( .a(n_17827), .o(n_17698) );
no02s10 g762874 ( .a(n_17655), .b(n_17656), .o(n_17827) );
no02s40 g762875 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_11_), .b(FE_OCPN867_n_45450), .o(n_17885) );
na02s08 g762876 ( .a(n_17842), .b(n_17744), .o(n_17889) );
na02s06 g762877 ( .a(n_17841), .b(delay_add_ln22_unr11_stage5_stallmux_q_8_), .o(n_17906) );
in01s01 g762878 ( .a(n_17866), .o(n_17867) );
no02s06 g762879 ( .a(n_17841), .b(delay_add_ln22_unr11_stage5_stallmux_q_8_), .o(n_17866) );
na02s01 g762881 ( .a(n_17865), .b(n_17864), .o(n_17909) );
no02s01 g762882 ( .a(n_17839), .b(n_17838), .o(n_17840) );
no02s01 g762883 ( .a(n_18013), .b(n_17463), .o(n_18084) );
in01s01 g762884 ( .a(n_17794), .o(n_17795) );
na02s01 g762885 ( .a(n_17766), .b(n_17719), .o(n_17794) );
no02s01 g762886 ( .a(n_17746), .b(n_17771), .o(n_17747) );
na02s06 g762887 ( .a(n_17523), .b(n_17282), .o(n_17659) );
no02m03 g762888 ( .a(n_17595), .b(n_17444), .o(n_17694) );
ao12s10 g762889 ( .a(n_17655), .b(FE_OCPN1296_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_8_), .o(n_17726) );
in01m02 g762891 ( .a(n_17630), .o(n_17628) );
in01s01 g762893 ( .a(n_17728), .o(n_17682) );
oa12s02 g762895 ( .a(n_17329), .b(FE_OCP_RBN1025_n_17417), .c(n_17325), .o(n_17627) );
ao12s02 g762896 ( .a(n_17326), .b(FE_OCP_RBN1026_n_17417), .c(n_17328), .o(n_17601) );
ao12s02 g762898 ( .a(n_17070), .b(FE_OCP_RBN1025_n_17417), .c(n_16991), .o(n_17626) );
in01s01 g762899 ( .a(n_17597), .o(n_17598) );
oa12s02 g762900 ( .a(n_17140), .b(FE_OCP_RBN1025_n_17417), .c(n_17070), .o(n_17597) );
oa12s01 g762902 ( .a(n_17993), .b(n_17994), .c(n_17992), .o(n_18420) );
na02s06 g762903 ( .a(n_17680), .b(n_17624), .o(n_17801) );
in01s01 g762906 ( .a(n_18102), .o(n_18103) );
oa12s01 g762907 ( .a(n_18035), .b(n_18034), .c(n_18033), .o(n_18102) );
oa12s01 g762908 ( .a(n_17991), .b(n_17990), .c(n_17989), .o(n_18689) );
in01s01 g762909 ( .a(n_18064), .o(n_18065) );
oa12s01 g762910 ( .a(n_17988), .b(n_17987), .c(n_17986), .o(n_18064) );
in01s01 g762911 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_22_), .o(n_17625) );
no02s01 TIMEBOOST_cell_1593 ( .a(n_34993), .b(n_34704), .o(TIMEBOOST_net_411) );
na02s02 g762915 ( .a(n_17683), .b(n_17592), .o(n_17624) );
no02s01 g762916 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_20_), .b(delay_add_ln22_unr11_stage5_stallmux_q_21_), .o(n_17568) );
no02f08 g762918 ( .a(n_17994), .b(n_17464), .o(n_18013) );
na02s01 g762919 ( .a(n_17994), .b(n_17992), .o(n_17993) );
no02s20 g762920 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_8_), .b(FE_OCP_RBN5514_n_44365), .o(n_17655) );
in01s01 g762921 ( .a(n_17718), .o(n_17719) );
no02m08 g762922 ( .a(n_17679), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_6_), .o(n_17718) );
na02m08 g762923 ( .a(n_17679), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_6_), .o(n_17766) );
in01s10 g762924 ( .a(n_17842), .o(n_17884) );
no02s10 g762925 ( .a(n_17797), .b(n_17745), .o(n_17842) );
na02m08 g762926 ( .a(n_17763), .b(n_15892), .o(n_17864) );
na02s06 g762927 ( .a(n_17762), .b(delay_add_ln22_unr11_stage5_stallmux_q_7_), .o(n_17865) );
na02s01 g762928 ( .a(n_17990), .b(n_17989), .o(n_17991) );
na02s01 g762929 ( .a(n_17987), .b(n_17986), .o(n_17988) );
na02s01 g762930 ( .a(n_18034), .b(n_18033), .o(n_18035) );
in01s06 g762931 ( .a(n_17792), .o(n_17793) );
ao12m03 g762932 ( .a(n_17765), .b(FE_OCPN867_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_10_), .o(n_17792) );
ao12m10 g762933 ( .a(n_17745), .b(FE_OCPN867_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_9_), .o(n_17796) );
oa12m08 g762934 ( .a(n_17619), .b(n_17678), .c(n_17548), .o(n_17771) );
ao12f08 g762935 ( .a(n_17639), .b(n_17717), .c(n_17715), .o(n_17839) );
oa22m02 g762936 ( .a(n_17460), .b(n_17584), .c(n_17456), .d(n_16339), .o(n_17567) );
oa22s01 g762938 ( .a(n_17678), .b(n_17638), .c(n_17621), .d(n_17637), .o(n_19053) );
in01m01 g762939 ( .a(n_17523), .o(n_17595) );
in01s01 g762949 ( .a(n_17725), .o(n_17674) );
in01s01 g762951 ( .a(n_17687), .o(n_17649) );
ao12s01 g762953 ( .a(n_17963), .b(n_17962), .c(n_17961), .o(n_18416) );
oa12s01 g762954 ( .a(n_17960), .b(n_17959), .c(n_17958), .o(n_18688) );
ao22s01 g762956 ( .a(n_17717), .b(n_17738), .c(FE_OCP_RBN7020_n_17717), .d(n_17737), .o(n_17836) );
ao12s01 g762957 ( .a(n_17985), .b(n_17984), .c(n_17983), .o(n_18487) );
oa12s01 g762958 ( .a(n_17982), .b(n_17981), .c(n_17980), .o(n_18531) );
in01s01 g762962 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_24_), .o(n_17772) );
no02s20 g762965 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_9_), .b(FE_OCPN1202_n_45450), .o(n_17745) );
in01s01 g762966 ( .a(n_17765), .o(n_17744) );
no02s40 g762967 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_10_), .b(FE_OCPN867_n_45450), .o(n_17765) );
na02s02 g762968 ( .a(n_17742), .b(n_17741), .o(n_17743) );
na02s01 g762969 ( .a(n_17623), .b(n_17672), .o(n_17746) );
na02s01 g762970 ( .a(n_17739), .b(n_17791), .o(n_17838) );
no02s01 g762971 ( .a(n_17984), .b(n_17983), .o(n_17985) );
no02s01 g762972 ( .a(n_17962), .b(n_17961), .o(n_17963) );
na02s01 g762973 ( .a(n_17981), .b(n_17980), .o(n_17982) );
ao12f08 g762974 ( .a(n_17542), .b(n_17939), .c(n_17364), .o(n_17994) );
oa12m02 g762975 ( .a(n_16902), .b(n_17489), .c(FE_OCP_RBN6876_n_16920), .o(n_17522) );
no02m04 g762976 ( .a(n_17490), .b(n_16942), .o(n_17566) );
na02s01 g762977 ( .a(n_17959), .b(n_17958), .o(n_17960) );
in01s02 g762978 ( .a(n_17592), .o(n_17593) );
ao12s02 g762979 ( .a(n_17684), .b(FE_OCP_RBN5511_n_44365), .c(delay_xor_ln21_unr12_stage5_stallmux_q_7_), .o(n_17592) );
ao12s01 g762980 ( .a(n_17543), .b(n_17939), .c(n_17301), .o(n_17990) );
no02s08 TIMEBOOST_cell_1744 ( .a(TIMEBOOST_net_486), .b(n_26354), .o(n_26456) );
in01m02 g762983 ( .a(n_17594), .o(n_17565) );
oa12s02 g762985 ( .a(n_17332), .b(n_17349), .c(n_17390), .o(n_17457) );
ao12s06 g762994 ( .a(n_16993), .b(n_17292), .c(n_17090), .o(n_17417) );
in01m04 g762995 ( .a(n_17762), .o(n_17763) );
ao12s01 g762997 ( .a(n_17370), .b(n_17905), .c(n_17299), .o(n_17987) );
no02m08 g762998 ( .a(n_17517), .b(n_17562), .o(n_17679) );
in01s01 g763001 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_23_), .o(n_18367) );
no03f08 TIMEBOOST_cell_85 ( .a(n_379), .b(n_371), .c(FE_RN_69_0), .o(FE_RN_71_0) );
no02s06 g763007 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_7_), .b(FE_OCP_RBN7104_n_44365), .o(n_17684) );
na02s06 g763008 ( .a(n_17590), .b(n_17589), .o(n_17672) );
in01s01 g763009 ( .a(n_17622), .o(n_17623) );
no02s06 g763010 ( .a(n_17590), .b(n_17589), .o(n_17622) );
ao12m04 g763011 ( .a(n_17486), .b(n_17561), .c(n_17560), .o(n_17562) );
in01s04 g763014 ( .a(n_17739), .o(n_17740) );
na02s04 g763015 ( .a(n_17667), .b(delay_add_ln22_unr11_stage5_stallmux_q_6_), .o(n_17739) );
in01s01 g763017 ( .a(n_17737), .o(n_17738) );
na02s01 g763018 ( .a(n_17715), .b(n_17640), .o(n_17737) );
na02s01 g763019 ( .a(n_17937), .b(n_17430), .o(n_17981) );
no02s01 g763020 ( .a(n_17905), .b(n_17266), .o(n_17962) );
oa12s02 g763021 ( .a(n_16986), .b(n_17483), .c(n_17515), .o(n_17516) );
no02s02 g763022 ( .a(n_17484), .b(n_17023), .o(n_17559) );
in01s02 g763023 ( .a(n_17557), .o(n_17558) );
oa12s06 g763024 ( .a(n_17082), .b(n_17403), .c(n_17515), .o(n_17557) );
no02s01 g763025 ( .a(n_17939), .b(n_17471), .o(n_17959) );
ao12s06 g763026 ( .a(n_17641), .b(FE_OCPN1296_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_8_), .o(n_17741) );
oa12s01 g763027 ( .a(n_17056), .b(n_17863), .c(n_17530), .o(n_17984) );
in01s01 g763028 ( .a(n_17678), .o(n_17621) );
oa12m08 g763029 ( .a(n_17482), .b(n_17588), .c(n_17406), .o(n_17678) );
ao12f08 g763031 ( .a(n_17504), .b(n_17635), .c(n_17580), .o(n_17717) );
oa12m02 g763032 ( .a(n_16976), .b(n_17452), .c(n_17454), .o(n_17493) );
no02s04 g763033 ( .a(n_17455), .b(n_17022), .o(n_17514) );
oa12f04 g763034 ( .a(n_17121), .b(n_17452), .c(n_17451), .o(n_17492) );
no02m06 TIMEBOOST_cell_1516 ( .a(TIMEBOOST_net_372), .b(n_29899), .o(n_29967) );
no02s04 g763036 ( .a(n_17489), .b(FE_OCP_RBN6876_n_16920), .o(n_17490) );
oa12s01 g763037 ( .a(n_17233), .b(n_17452), .c(n_17449), .o(n_17487) );
no02s02 g763038 ( .a(n_17450), .b(FE_OCP_RBN3401_n_17233), .o(n_17512) );
no02s06 g763040 ( .a(n_17415), .b(n_17405), .o(n_17510) );
oa22m02 g763041 ( .a(n_17294), .b(n_17584), .c(n_17290), .d(n_17753), .o(n_17418) );
in01s02 g763042 ( .a(n_17460), .o(n_17456) );
no02f08 TIMEBOOST_cell_1530 ( .a(TIMEBOOST_net_379), .b(n_38604), .o(n_38655) );
oa12s01 g763046 ( .a(n_17636), .b(n_17635), .c(n_17634), .o(n_19010) );
ao12s01 g763047 ( .a(n_17904), .b(n_17903), .c(n_17902), .o(n_18494) );
in01s01 g763048 ( .a(FE_OCP_DRV_N1438_n_17643), .o(n_17644) );
oa12s01 g763049 ( .a(n_17554), .b(n_17588), .c(n_17553), .o(n_17643) );
in01s01 g763050 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_20_), .o(n_17416) );
na02s01 g763053 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n_17556) );
no02s01 g763054 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n_17555) );
in01s06 g763057 ( .a(n_17641), .o(n_17642) );
no02s10 g763058 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_8_), .b(FE_OCP_RBN5513_n_44365), .o(n_17641) );
na02s04 g763059 ( .a(n_17579), .b(n_17669), .o(n_17742) );
in01s01 g763060 ( .a(n_17639), .o(n_17640) );
no02s06 g763061 ( .a(n_17620), .b(delay_add_ln22_unr11_stage5_stallmux_q_5_), .o(n_17639) );
na02s06 g763062 ( .a(n_17620), .b(delay_add_ln22_unr11_stage5_stallmux_q_5_), .o(n_17715) );
in01s01 g763063 ( .a(n_17637), .o(n_17638) );
na02s01 g763064 ( .a(n_17549), .b(n_17619), .o(n_17637) );
na02s01 g763065 ( .a(n_17862), .b(n_17499), .o(n_17937) );
na02s01 g763066 ( .a(n_17634), .b(n_17635), .o(n_17636) );
na02s01 g763067 ( .a(n_17553), .b(n_17588), .o(n_17554) );
no02s01 g763068 ( .a(n_17863), .b(n_17426), .o(n_17905) );
no02s04 g763069 ( .a(n_17452), .b(n_17454), .o(n_17455) );
no02m04 TIMEBOOST_cell_1515 ( .a(n_29898), .b(n_29896), .o(TIMEBOOST_net_372) );
no02m04 g763071 ( .a(n_17414), .b(n_17132), .o(n_17489) );
no02s02 g763072 ( .a(n_17452), .b(n_17449), .o(n_17450) );
na02s02 g763073 ( .a(n_17200), .b(n_17044), .o(n_17252) );
no02m04 TIMEBOOST_cell_1529 ( .a(n_38583), .b(n_38778), .o(TIMEBOOST_net_379) );
in01s01 g763075 ( .a(n_17485), .o(n_17486) );
no02s01 g763079 ( .a(n_17903), .b(n_17902), .o(n_17904) );
no02s02 g763080 ( .a(n_17515), .b(n_17483), .o(n_17484) );
no02s02 g763081 ( .a(n_17414), .b(n_17234), .o(n_17415) );
in01s02 g763085 ( .a(n_17349), .o(n_17350) );
in01m02 g763088 ( .a(n_17292), .o(n_17349) );
na02s01 TIMEBOOST_cell_1180 ( .a(TIMEBOOST_net_204), .b(n_12761), .o(n_46985) );
no02m04 TIMEBOOST_cell_3965 ( .a(n_8159), .b(FE_RN_974_0), .o(TIMEBOOST_net_1073) );
ao12s01 g763093 ( .a(n_17546), .b(n_17545), .c(n_17544), .o(n_18953) );
ao22s01 g763094 ( .a(n_17816), .b(n_17602), .c(n_17817), .d(n_17603), .o(n_18488) );
in01s01 g763097 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n_17508) );
in01s01 g763100 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_22_), .o(n_18368) );
no02s01 TIMEBOOST_cell_3964 ( .a(TIMEBOOST_net_1072), .b(n_34283), .o(n_34394) );
no03s02 TIMEBOOST_cell_7936 ( .a(n_5277), .b(n_5230), .c(n_5276), .o(TIMEBOOST_net_2599) );
na02s03 g763104 ( .a(FE_OCP_RBN7103_n_44365), .b(n_17409), .o(n_17458) );
na02s06 g763105 ( .a(n_17507), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_4_), .o(n_17619) );
in01s01 g763106 ( .a(n_17548), .o(n_17549) );
no02s08 g763107 ( .a(n_17507), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_4_), .o(n_17548) );
in01s02 g763108 ( .a(n_17547), .o(n_17669) );
no02s40 g763109 ( .a(FE_OCP_RBN5513_n_44365), .b(delay_xor_ln22_unr12_stage5_stallmux_q_7_), .o(n_17547) );
no02m04 TIMEBOOST_cell_3916 ( .a(TIMEBOOST_net_1048), .b(FE_OCP_RBN2581_n_37913), .o(FE_RN_757_0) );
na02s01 g763111 ( .a(n_17482), .b(n_17407), .o(n_17553) );
na02s01 g763112 ( .a(n_17505), .b(n_17580), .o(n_17634) );
no02s01 g763113 ( .a(n_17545), .b(n_17544), .o(n_17546) );
in01s02 g763116 ( .a(n_17452), .o(n_17446) );
in01f08 g763117 ( .a(n_17414), .o(n_17452) );
no02f08 g763118 ( .a(n_17250), .b(n_17249), .o(n_17414) );
in01s02 g763119 ( .a(n_17200), .o(n_17201) );
na02s02 g763120 ( .a(n_17146), .b(n_16880), .o(n_17200) );
no02m06 g763121 ( .a(n_17045), .b(n_17146), .o(n_17147) );
no02s06 g763122 ( .a(n_17343), .b(n_17444), .o(n_17445) );
oa12m08 g763124 ( .a(n_17398), .b(n_17481), .c(n_17279), .o(n_17588) );
ao12f08 g763125 ( .a(n_17399), .b(n_17433), .c(n_17477), .o(n_17635) );
in01s01 g763126 ( .a(n_17862), .o(n_17903) );
in01s01 g763128 ( .a(n_17863), .o(n_17862) );
ao12f08 g763129 ( .a(n_17368), .b(n_17787), .c(n_17298), .o(n_17863) );
oa22m02 g763130 ( .a(n_17199), .b(n_17336), .c(n_17142), .d(n_17753), .o(n_17291) );
in01m02 g763131 ( .a(n_17294), .o(n_17290) );
na02s06 TIMEBOOST_cell_2824 ( .a(n_7016), .b(n_7017), .o(TIMEBOOST_net_703) );
na02s02 TIMEBOOST_cell_7566 ( .a(FE_RN_858_0), .b(n_18811), .o(TIMEBOOST_net_2414) );
ao22s01 g763134 ( .a(n_17481), .b(n_17435), .c(n_17397), .d(n_17434), .o(n_18854) );
in01s01 g763135 ( .a(n_17882), .o(n_17883) );
oa12s01 g763136 ( .a(n_17820), .b(n_17819), .c(n_17818), .o(n_17882) );
in01s01 g763137 ( .a(n_17859), .o(n_17860) );
oa12s01 g763138 ( .a(n_17790), .b(n_17789), .c(n_17788), .o(n_17859) );
in01m06 g763140 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_6_), .o(n_17409) );
na02s06 g763143 ( .a(n_17401), .b(n_17396), .o(n_17480) );
na02f08 TIMEBOOST_cell_7565 ( .a(TIMEBOOST_net_2413), .b(n_23640), .o(FE_RN_2382_0) );
in01s01 g763145 ( .a(n_17406), .o(n_17407) );
no02s06 g763146 ( .a(n_17348), .b(n_17347), .o(n_17406) );
na02s06 g763147 ( .a(n_17348), .b(n_17347), .o(n_17482) );
na02s06 g763151 ( .a(n_17479), .b(n_17478), .o(n_17580) );
in01s01 g763152 ( .a(n_17504), .o(n_17505) );
no02s06 g763153 ( .a(n_17479), .b(n_17478), .o(n_17504) );
na02s01 g763154 ( .a(n_17477), .b(n_17400), .o(n_17544) );
na02s01 g763155 ( .a(n_17789), .b(n_17788), .o(n_17790) );
na02s01 g763156 ( .a(n_17819), .b(n_17818), .o(n_17820) );
na02s02 TIMEBOOST_cell_5575 ( .a(TIMEBOOST_net_1735), .b(n_6360), .o(n_6476) );
na02m08 TIMEBOOST_cell_2823 ( .a(n_7127), .b(TIMEBOOST_net_702), .o(n_7209) );
na02m06 g763159 ( .a(n_17009), .b(n_16879), .o(n_17146) );
in01s03 g763160 ( .a(n_17345), .o(n_17346) );
ao12s06 g763161 ( .a(n_17289), .b(FE_OCP_RBN7110_n_44365), .c(delay_xor_ln21_unr12_stage5_stallmux_q_5_), .o(n_17345) );
na02s02 g763163 ( .a(n_17281), .b(n_17274), .o(n_17405) );
in01s01 g763164 ( .a(n_17816), .o(n_17817) );
no02s01 g763165 ( .a(n_17787), .b(n_17369), .o(n_17816) );
oa12s02 g763167 ( .a(n_17172), .b(n_17287), .c(n_16839), .o(n_17344) );
no02m04 g763168 ( .a(n_17118), .b(n_17288), .o(n_17404) );
na02s06 g763169 ( .a(n_17402), .b(n_17284), .o(n_17403) );
no02s01 TIMEBOOST_cell_1212 ( .a(n_28591), .b(TIMEBOOST_net_220), .o(n_28714) );
in01s02 g763172 ( .a(n_17459), .o(n_17441) );
oa22s04 g763173 ( .a(n_17237), .b(n_16950), .c(n_17238), .d(n_16995), .o(n_17459) );
in01m02 g763174 ( .a(n_17475), .o(n_17550) );
no02m04 TIMEBOOST_cell_1312 ( .a(TIMEBOOST_net_270), .b(FE_OCP_RBN2662_n_19393), .o(n_19539) );
in01s01 g763178 ( .a(FE_OCPN1636_n_18860), .o(n_18919) );
oa12s01 g763179 ( .a(n_17474), .b(n_17473), .c(n_17472), .o(n_18860) );
in01s01 g763180 ( .a(n_18479), .o(n_18744) );
oa12s01 g763181 ( .a(n_17439), .b(n_17438), .c(n_17437), .o(n_18479) );
no02f06 TIMEBOOST_cell_8055 ( .a(TIMEBOOST_net_2658), .b(n_6231), .o(n_6358) );
in01s01 g763183 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_), .o(n_18291) );
na02s01 g763185 ( .a(n_17438), .b(n_17437), .o(n_17439) );
in01s06 g763186 ( .a(n_17289), .o(n_17560) );
no02s03 g763187 ( .a(FE_OCP_RBN7110_n_44365), .b(delay_xor_ln21_unr12_stage5_stallmux_q_5_), .o(n_17289) );
ao12s06 g763189 ( .a(n_17240), .b(n_17247), .c(n_17040), .o(n_17341) );
no02s06 TIMEBOOST_cell_6116 ( .a(TIMEBOOST_net_1909), .b(n_3915), .o(n_4101) );
in01s01 g763192 ( .a(n_17399), .o(n_17400) );
no02m08 g763193 ( .a(n_17340), .b(delay_add_ln22_unr11_stage5_stallmux_q_3_), .o(n_17399) );
na02s08 g763194 ( .a(n_17340), .b(delay_add_ln22_unr11_stage5_stallmux_q_3_), .o(n_17477) );
na02s01 g763195 ( .a(n_17473), .b(n_17472), .o(n_17474) );
in01s01 g763196 ( .a(n_17434), .o(n_17435) );
na02s01 g763197 ( .a(n_17280), .b(n_17398), .o(n_17434) );
no02s04 TIMEBOOST_cell_1683 ( .a(n_9578), .b(n_9726), .o(TIMEBOOST_net_456) );
no02m02 g763200 ( .a(n_17287), .b(n_16839), .o(n_17288) );
na02s06 g763201 ( .a(n_17249), .b(n_17233), .o(n_17402) );
no02s01 TIMEBOOST_cell_1211 ( .a(n_28615), .b(n_28105), .o(TIMEBOOST_net_220) );
in01s01 g763203 ( .a(n_17481), .o(n_17397) );
ao12m08 g763204 ( .a(n_17335), .b(n_17231), .c(n_16857), .o(n_17481) );
in01s02 g763205 ( .a(n_17395), .o(n_17396) );
ao12s06 g763206 ( .a(n_17339), .b(FE_OCP_RBN5511_n_44365), .c(delay_xor_ln22_unr12_stage5_stallmux_q_5_), .o(n_17395) );
no02s02 g763208 ( .a(n_17283), .b(FE_OCP_RBN3387_n_17130), .o(n_17284) );
oa12s01 g763209 ( .a(n_17159), .b(n_17736), .c(n_17462), .o(n_17789) );
in01s01 g763210 ( .a(n_17433), .o(n_17545) );
ao12f08 g763211 ( .a(n_17272), .b(n_17472), .c(n_17393), .o(n_17433) );
oa22f02 g763212 ( .a(n_46974), .b(n_17336), .c(n_17003), .d(FE_OCP_RBN3196_n_15599), .o(n_17144) );
in01m02 g763214 ( .a(n_17199), .o(n_17142) );
na02s02 TIMEBOOST_cell_2888 ( .a(n_1953), .b(n_1952), .o(TIMEBOOST_net_735) );
in01s01 g763216 ( .a(n_17048), .o(n_17049) );
in01s01 g763217 ( .a(n_17009), .o(n_17048) );
oa12m06 g763218 ( .a(n_16809), .b(n_16884), .c(n_16760), .o(n_17009) );
in01s06 g763219 ( .a(n_17282), .o(n_17444) );
oa12f06 g763222 ( .a(n_16869), .b(n_17001), .c(n_16951), .o(n_17091) );
in01s01 g763223 ( .a(n_17785), .o(n_17786) );
oa12s01 g763224 ( .a(n_17712), .b(n_17736), .c(n_17711), .o(n_17785) );
na02m04 TIMEBOOST_cell_8643 ( .a(TIMEBOOST_net_2808), .b(n_5468), .o(n_47000) );
no02m04 TIMEBOOST_cell_1696 ( .a(TIMEBOOST_net_462), .b(n_20149), .o(n_20184) );
in01s01 g763227 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_18_), .o(n_17050) );
in01s03 g763230 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_6_), .o(n_17394) );
in01s08 g763233 ( .a(n_17561), .o(n_17410) );
in01s01 g763235 ( .a(n_17279), .o(n_17280) );
no02m08 g763236 ( .a(n_17243), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_2_), .o(n_17279) );
na02m08 g763237 ( .a(n_17243), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_2_), .o(n_17398) );
no02s10 g763239 ( .a(FE_OCP_RBN7111_n_44365), .b(delay_xor_ln22_unr12_stage5_stallmux_q_5_), .o(n_17339) );
no02s04 TIMEBOOST_cell_1684 ( .a(TIMEBOOST_net_456), .b(n_9672), .o(n_9727) );
no02s01 g763242 ( .a(n_17232), .b(n_17335), .o(n_17438) );
na02s01 g763243 ( .a(n_17273), .b(n_17393), .o(n_17473) );
no02s01 TIMEBOOST_cell_1681 ( .a(n_30356), .b(n_30076), .o(TIMEBOOST_net_455) );
na02s01 g763245 ( .a(n_17736), .b(n_17711), .o(n_17712) );
no02m06 g763246 ( .a(n_17006), .b(n_16998), .o(n_17249) );
na02m04 g763247 ( .a(n_16917), .b(n_16833), .o(n_16954) );
na02s02 TIMEBOOST_cell_2887 ( .a(n_13259), .b(TIMEBOOST_net_734), .o(n_13470) );
in01s06 g763250 ( .a(n_17239), .o(n_17240) );
no02s01 TIMEBOOST_cell_1311 ( .a(n_19478), .b(n_18705), .o(TIMEBOOST_net_270) );
in01s02 g763255 ( .a(n_17287), .o(n_17275) );
na02m06 g763256 ( .a(n_17088), .b(n_17002), .o(n_17287) );
in01s04 g763257 ( .a(n_17237), .o(n_17238) );
ao12s08 g763258 ( .a(n_16782), .b(n_17083), .c(n_16832), .o(n_17237) );
na02s01 TIMEBOOST_cell_1179 ( .a(n_12461), .b(n_12495), .o(TIMEBOOST_net_204) );
na02s06 g763260 ( .a(n_17007), .b(n_16923), .o(n_17090) );
in01s01 g763263 ( .a(n_17195), .o(n_17235) );
no02s06 g763264 ( .a(FE_OCP_RBN6172_n_16923), .b(n_17041), .o(n_17195) );
in01f02 g763266 ( .a(n_17334), .o(n_17440) );
in01s02 g763268 ( .a(n_17274), .o(n_17449) );
in01s02 g763269 ( .a(n_17283), .o(n_17274) );
no02m04 TIMEBOOST_cell_5672 ( .a(n_26694), .b(n_26615), .o(TIMEBOOST_net_1784) );
na02s02 g763271 ( .a(n_17233), .b(n_17134), .o(n_17234) );
in01s01 g763272 ( .a(FE_OCP_DRV_N3534_n_18559), .o(n_18748) );
oa12s01 g763273 ( .a(n_17228), .b(n_17227), .c(n_17226), .o(n_18559) );
no02s20 g763275 ( .a(FE_OCP_RBN7104_n_44365), .b(delay_xor_ln21_unr12_stage5_stallmux_q_4_), .o(n_17197) );
no02m08 g763277 ( .a(n_17194), .b(n_17193), .o(n_17335) );
in01s01 g763278 ( .a(n_17231), .o(n_17232) );
na02m08 g763279 ( .a(n_17194), .b(n_17193), .o(n_17231) );
na02m08 g763282 ( .a(n_17230), .b(n_17229), .o(n_17393) );
in01s01 g763283 ( .a(n_17272), .o(n_17273) );
no02m08 g763284 ( .a(n_17229), .b(n_17230), .o(n_17272) );
na02s01 g763285 ( .a(n_17227), .b(n_17226), .o(n_17228) );
na02m04 g763287 ( .a(n_16911), .b(n_17039), .o(n_17088) );
in01s01 g763288 ( .a(n_17043), .o(n_17044) );
no02m02 g763289 ( .a(n_17045), .b(n_16952), .o(n_17043) );
no02m06 g763290 ( .a(n_16952), .b(n_16808), .o(n_16953) );
na02s02 g763291 ( .a(n_17332), .b(n_17331), .o(n_17333) );
no02m02 g763292 ( .a(n_17391), .b(n_17390), .o(n_17392) );
no02s01 TIMEBOOST_cell_1176 ( .a(TIMEBOOST_net_202), .b(n_37785), .o(n_37825) );
na02s01 g763294 ( .a(n_17329), .b(n_17328), .o(n_17330) );
no02s01 g763295 ( .a(n_17326), .b(n_17325), .o(n_17327) );
na02s01 g763296 ( .a(n_17037), .b(n_17135), .o(n_17136) );
no02s01 g763297 ( .a(n_16957), .b(n_17036), .o(n_17191) );
no02s06 g763298 ( .a(n_17042), .b(n_16957), .o(n_17140) );
no02m08 TIMEBOOST_cell_1304 ( .a(TIMEBOOST_net_266), .b(n_24246), .o(n_24262) );
na02s01 g763300 ( .a(n_17323), .b(n_17035), .o(n_17324) );
no02s01 g763301 ( .a(n_16996), .b(n_17388), .o(n_17389) );
na02m04 TIMEBOOST_cell_8616 ( .a(TIMEBOOST_net_1126), .b(n_21360), .o(TIMEBOOST_net_2795) );
no02s06 g763303 ( .a(FE_OCP_RBN6078_n_16084), .b(n_16996), .o(n_17041) );
na02f08 TIMEBOOST_cell_1188 ( .a(FE_RN_1717_0), .b(TIMEBOOST_net_208), .o(n_33518) );
in01s06 g763305 ( .a(n_17085), .o(n_17086) );
na02s10 g763306 ( .a(n_16915), .b(n_17040), .o(n_17085) );
in01s06 g763307 ( .a(n_17188), .o(n_17189) );
ao12s10 g763308 ( .a(n_17133), .b(FE_OCP_RBN7110_n_44365), .c(delay_xor_ln22_unr12_stage5_stallmux_q_4_), .o(n_17188) );
oa12f08 g763309 ( .a(n_17025), .b(n_17125), .c(n_17226), .o(n_17472) );
in01s03 g763310 ( .a(n_17005), .o(n_17006) );
no02s08 g763311 ( .a(n_16910), .b(n_16868), .o(n_17005) );
no02f08 g763312 ( .a(n_17578), .b(n_17432), .o(n_17736) );
oa22f02 g763313 ( .a(n_16916), .b(FE_OCP_RBN3193_n_15599), .c(n_16872), .d(n_16339), .o(n_17004) );
in01f02 g763314 ( .a(n_46974), .o(n_17003) );
in01s02 g763316 ( .a(n_16917), .o(n_16918) );
in01s02 g763317 ( .a(n_16884), .o(n_16917) );
ao12s06 g763318 ( .a(n_16762), .b(n_16793), .c(n_16706), .o(n_16884) );
in01s01 g763319 ( .a(n_17386), .o(n_17387) );
na02m02 TIMEBOOST_cell_1182 ( .a(n_23500), .b(TIMEBOOST_net_205), .o(n_23516) );
in01s01 g763321 ( .a(n_17384), .o(n_17385) );
no02f08 TIMEBOOST_cell_1190 ( .a(TIMEBOOST_net_209), .b(n_7332), .o(n_47176) );
in01s01 g763323 ( .a(n_17382), .o(n_17383) );
na02s02 g763324 ( .a(n_17178), .b(n_17215), .o(n_17382) );
in01f02 g763325 ( .a(n_46973), .o(n_17187) );
in01m02 g763327 ( .a(n_17001), .o(n_17002) );
no02f08 g763328 ( .a(n_16883), .b(n_16876), .o(n_17001) );
no02m08 g763329 ( .a(n_16882), .b(n_16843), .o(n_16951) );
no02s06 g763333 ( .a(n_17132), .b(n_17033), .o(n_17233) );
oa22f02 g763334 ( .a(n_17128), .b(FE_OCP_RBN3193_n_15599), .c(n_17061), .d(n_16339), .o(n_17224) );
no02s01 TIMEBOOST_cell_3406 ( .a(n_27204), .b(FE_RN_1535_0), .o(TIMEBOOST_net_994) );
in01s02 g763337 ( .a(n_17380), .o(n_17381) );
na02s02 g763338 ( .a(n_17185), .b(n_17223), .o(n_17380) );
in01s01 g763339 ( .a(n_17378), .o(n_17379) );
no02s01 TIMEBOOST_cell_5580 ( .a(n_39590), .b(n_40247), .o(TIMEBOOST_net_1738) );
in01s01 g763341 ( .a(n_17376), .o(n_17377) );
na02s02 g763342 ( .a(n_17180), .b(n_17217), .o(n_17376) );
in01s01 g763344 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_17_), .o(n_16921) );
in01s01 g763348 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_18_), .o(n_17186) );
na02s01 g763350 ( .a(n_17708), .b(n_17665), .o(n_17710) );
in01m03 g763351 ( .a(n_17040), .o(n_17244) );
na02s10 g763353 ( .a(FE_OCP_RBN7111_n_44365), .b(delay_xor_ln21_unr12_stage5_stallmux_q_3_), .o(n_16915) );
no02s20 g763356 ( .a(FE_OCP_RBN7104_n_44365), .b(delay_xor_ln22_unr12_stage5_stallmux_q_4_), .o(n_17133) );
na02f08 g763357 ( .a(n_17632), .b(n_17532), .o(n_17633) );
na02s01 g763358 ( .a(n_17708), .b(n_17467), .o(n_17709) );
no02s01 g763359 ( .a(n_17026), .b(n_17125), .o(n_17227) );
na02f02 g763361 ( .a(n_16938), .b(n_16753), .o(n_16999) );
in01s03 g763363 ( .a(n_17083), .o(n_17123) );
in01s06 g763364 ( .a(n_17039), .o(n_17083) );
na02s06 g763365 ( .a(n_16905), .b(n_16998), .o(n_17039) );
na02f02 g763367 ( .a(n_16811), .b(n_16785), .o(n_16840) );
no02m06 g763368 ( .a(n_16836), .b(FE_OCP_RBN3084_n_15314), .o(n_16952) );
in01m02 g763370 ( .a(n_17331), .o(n_17390) );
no02s01 TIMEBOOST_cell_1175 ( .a(n_37750), .b(n_37749), .o(TIMEBOOST_net_202) );
na02s06 g763372 ( .a(FE_OCP_RBN6175_n_16923), .b(n_15479), .o(n_17331) );
in01s01 g763373 ( .a(n_17081), .o(n_17082) );
na02s02 g763374 ( .a(n_16948), .b(n_16986), .o(n_17081) );
na02s02 g763375 ( .a(FE_OCP_RBN6174_n_16923), .b(FE_OCP_RBN3072_n_15433), .o(n_17332) );
no02s03 g763376 ( .a(FE_OCPN900_n_16923), .b(n_15479), .o(n_17391) );
na02s02 g763377 ( .a(FE_OCP_RBN6175_n_16923), .b(FE_OCP_RBN4370_n_46982), .o(n_17185) );
na02s02 g763378 ( .a(FE_OCP_RBN6174_n_16923), .b(FE_OCP_RBN3134_n_46982), .o(n_17223) );
in01s01 g763379 ( .a(n_17329), .o(n_17326) );
na02s01 g763380 ( .a(FE_OCPN900_n_16923), .b(FE_OCPN1274_n_15708), .o(n_17329) );
no02s01 g763381 ( .a(FE_OCP_RBN6175_n_16923), .b(FE_OCPN1274_n_15708), .o(n_17325) );
na02s01 g763382 ( .a(FE_OCP_RBN6174_n_16923), .b(n_15762), .o(n_17328) );
no02f06 TIMEBOOST_cell_5579 ( .a(TIMEBOOST_net_1737), .b(FE_RN_1180_0), .o(n_46978) );
na02s01 g763384 ( .a(FE_OCP_RBN6174_n_16923), .b(n_15983), .o(n_17221) );
in01s01 g763386 ( .a(n_16957), .o(n_17037) );
no02s02 g763387 ( .a(n_16919), .b(n_15939), .o(n_16957) );
in01s01 g763390 ( .a(n_17036), .o(n_17135) );
no02s02 g763391 ( .a(n_16912), .b(FE_OCP_RBN3204_n_15900), .o(n_17036) );
na02s04 TIMEBOOST_cell_1181 ( .a(FE_RN_1571_0), .b(n_23515), .o(TIMEBOOST_net_205) );
no02s01 g763393 ( .a(n_16923), .b(FE_OCP_RBN3235_n_16041), .o(n_17137) );
in01s01 g763397 ( .a(n_16996), .o(n_17035) );
no02s06 g763398 ( .a(n_16919), .b(FE_OCP_RBN3220_n_15992), .o(n_16996) );
na02s01 g763399 ( .a(FE_OCP_RBN6172_n_16923), .b(FE_OCP_RBN3220_n_15992), .o(n_17323) );
no02m01 g763400 ( .a(FE_OCPN900_n_16923), .b(n_15992), .o(n_17388) );
na02s01 g763401 ( .a(FE_OCP_RBN6175_n_16923), .b(FE_OCP_RBN6078_n_16084), .o(n_17180) );
na02s01 g763402 ( .a(FE_OCP_RBN6172_n_16923), .b(n_16084), .o(n_17217) );
no02s01 g763403 ( .a(FE_OCP_RBN6176_n_16923), .b(n_16146), .o(n_17216) );
na02m06 TIMEBOOST_cell_1187 ( .a(FE_RN_1994_0), .b(FE_RN_650_0), .o(TIMEBOOST_net_208) );
no02s02 TIMEBOOST_cell_1189 ( .a(FE_RN_1840_0), .b(FE_RN_2825_0), .o(TIMEBOOST_net_209) );
na02s01 g763406 ( .a(FE_OCP_RBN6175_n_16923), .b(n_16003), .o(n_17178) );
na02s01 g763407 ( .a(FE_OCP_RBN6172_n_16923), .b(n_16038), .o(n_17215) );
na02s06 g763408 ( .a(n_16941), .b(n_16902), .o(n_17033) );
in01s06 g763409 ( .a(n_17072), .o(n_17073) );
na02s02 g763411 ( .a(n_16838), .b(n_16874), .o(n_16950) );
no02m01 g763412 ( .a(n_16876), .b(n_16837), .o(n_16995) );
in01s02 g763413 ( .a(n_17213), .o(n_17214) );
no02m02 g763414 ( .a(n_17118), .b(n_16839), .o(n_17213) );
in01m02 g763415 ( .a(n_16910), .o(n_16911) );
na02m08 g763416 ( .a(n_16838), .b(n_16758), .o(n_16910) );
in01s01 g763418 ( .a(n_17132), .o(n_17121) );
na02s06 g763419 ( .a(n_17032), .b(n_16976), .o(n_17132) );
na02s01 g763420 ( .a(n_16902), .b(n_16944), .o(n_17031) );
no02s02 g763421 ( .a(n_16942), .b(n_16903), .o(n_17071) );
ao12f08 g763422 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n_17577), .c(n_17496), .o(n_17578) );
no02f04 g763423 ( .a(n_16837), .b(n_16759), .o(n_16883) );
no03s02 TIMEBOOST_cell_7650 ( .a(FE_OCP_RBN4163_n_3390), .b(n_2958), .c(FE_OCP_RBN4164_n_3390), .o(TIMEBOOST_net_2456) );
in01s01 g763425 ( .a(n_17176), .o(n_17177) );
na02s01 g763426 ( .a(n_16986), .b(n_16943), .o(n_17176) );
no02s02 g763428 ( .a(n_16903), .b(n_16867), .o(n_16920) );
no02m06 g763429 ( .a(n_16839), .b(n_15651), .o(n_16882) );
in01s02 g763430 ( .a(n_17268), .o(n_17269) );
no02s02 g763431 ( .a(n_17454), .b(n_17022), .o(n_17268) );
ao12s01 g763433 ( .a(n_17366), .b(n_17576), .c(n_17614), .o(n_17615) );
oa22f02 g763434 ( .a(n_46975), .b(FE_OCP_RBN3193_n_15599), .c(n_16895), .d(n_17753), .o(n_17029) );
no02s06 g763435 ( .a(n_16923), .b(n_15694), .o(n_16993) );
in01s02 g763436 ( .a(n_17069), .o(n_17070) );
in01s01 g763438 ( .a(n_17027), .o(n_17069) );
no02s01 g763439 ( .a(n_16912), .b(n_15995), .o(n_17027) );
in01s01 g763440 ( .a(FE_OCPN919_n_17042), .o(n_16991) );
no02s01 g763441 ( .a(n_16836), .b(n_15949), .o(n_17042) );
in01s01 g763443 ( .a(n_17120), .o(n_17174) );
in01s02 g763446 ( .a(n_17321), .o(n_17322) );
in01s01 TIMEBOOST_cell_5912 ( .a(TIMEBOOST_net_1800), .o(TIMEBOOST_net_1801) );
in01s01 g763448 ( .a(n_17319), .o(n_17320) );
na02s02 g763449 ( .a(n_17170), .b(n_17113), .o(n_17319) );
in01s01 g763450 ( .a(n_17317), .o(n_17318) );
na02s01 g763451 ( .a(n_17119), .b(n_17169), .o(n_17317) );
in01s01 g763452 ( .a(n_17315), .o(n_17316) );
na02s02 g763453 ( .a(n_17115), .b(n_17167), .o(n_17315) );
ao22s01 g763454 ( .a(n_17577), .b(n_17527), .c(n_17503), .d(n_17526), .o(n_18419) );
in01s01 g763455 ( .a(n_17313), .o(n_17314) );
no02s02 TIMEBOOST_cell_3408 ( .a(n_27204), .b(FE_OCP_RBN3078_n_25816), .o(TIMEBOOST_net_995) );
in01s02 g763457 ( .a(n_17311), .o(n_17312) );
na02s06 g763458 ( .a(n_17171), .b(n_17114), .o(n_17311) );
in01s01 g763463 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_17_), .o(n_16990) );
no02s10 g763468 ( .a(n_17129), .b(n_16973), .o(n_17247) );
no02s40 g763469 ( .a(FE_OCP_RBN7110_n_44365), .b(delay_xor_ln22_unr12_stage5_stallmux_q_3_), .o(n_17084) );
no02m08 g763470 ( .a(n_16987), .b(delay_add_ln22_unr11_stage5_stallmux_q_1_), .o(n_17125) );
in01s01 g763471 ( .a(n_17025), .o(n_17026) );
na02f06 g763472 ( .a(n_16987), .b(delay_add_ln22_unr11_stage5_stallmux_q_1_), .o(n_17025) );
na02s01 g763474 ( .a(n_17541), .b(n_17302), .o(n_17543) );
in01s02 g763475 ( .a(n_16908), .o(n_16909) );
na02s04 g763476 ( .a(n_16880), .b(n_16879), .o(n_16908) );
no02m06 g763480 ( .a(n_16814), .b(FE_OCPN1278_n_15656), .o(n_16839) );
na02s01 g763481 ( .a(n_16843), .b(FE_OCP_RBN3179_n_16088), .o(n_16948) );
na02s01 g763482 ( .a(n_17108), .b(FE_OCP_RBN3179_n_16088), .o(n_17119) );
in01s01 g763483 ( .a(n_17734), .o(n_17708) );
na04s02 TIMEBOOST_cell_7168 ( .a(n_2460), .b(n_2858), .c(n_2433), .d(n_2102), .o(n_2607) );
in01s01 g763486 ( .a(n_17118), .o(n_17172) );
no02s08 g763487 ( .a(n_16977), .b(n_15549), .o(n_17118) );
in01s04 g763490 ( .a(n_16838), .o(n_16876) );
na02m08 g763491 ( .a(n_16814), .b(FE_OCP_DRV_N3524_FE_OCP_RBN3021_n_15319), .o(n_16838) );
in01s01 g763495 ( .a(n_16986), .o(n_17023) );
na02s03 g763496 ( .a(n_16843), .b(n_15948), .o(n_16986) );
na02m01 TIMEBOOST_cell_5024 ( .a(n_41324), .b(n_41525), .o(TIMEBOOST_net_1460) );
in01s02 g763499 ( .a(n_16904), .o(n_16905) );
ao12s06 g763500 ( .a(n_16777), .b(n_16784), .c(n_16752), .o(n_16904) );
in01s01 g763502 ( .a(n_16837), .o(n_16874) );
no02m04 g763503 ( .a(n_16814), .b(FE_OCP_DRV_N3524_FE_OCP_RBN3021_n_15319), .o(n_16837) );
na02s02 g763504 ( .a(n_16977), .b(n_15651), .o(n_17171) );
no02s06 g763505 ( .a(n_17108), .b(n_16940), .o(n_17454) );
in01s01 g763507 ( .a(n_16903), .o(n_16944) );
no02s02 g763508 ( .a(n_16814), .b(FE_OCP_RBN2111_n_15911), .o(n_16903) );
na02s01 g763509 ( .a(n_16977), .b(n_16118), .o(n_17170) );
na02s02 g763512 ( .a(n_16796), .b(n_15993), .o(n_16943) );
na02s01 g763513 ( .a(n_16977), .b(n_16088), .o(n_17169) );
no02s01 g763514 ( .a(n_17108), .b(n_16086), .o(n_17117) );
na02s01 g763515 ( .a(n_16977), .b(n_16011), .o(n_17167) );
oa12m06 g763516 ( .a(n_17541), .b(n_17424), .c(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17542) );
no02f08 g763517 ( .a(n_17576), .b(n_17429), .o(n_17632) );
in01s01 g763522 ( .a(n_16902), .o(n_16942) );
na02s06 g763523 ( .a(n_16843), .b(FE_OCP_RBN2111_n_15911), .o(n_16902) );
na02s01 g763524 ( .a(n_17108), .b(FE_OCP_RBN6057_n_16011), .o(n_17115) );
na02s02 g763525 ( .a(n_16814), .b(n_15912), .o(n_17032) );
no02m04 TIMEBOOST_cell_1303 ( .a(n_24175), .b(n_21852), .o(TIMEBOOST_net_266) );
no02s02 TIMEBOOST_cell_3407 ( .a(TIMEBOOST_net_994), .b(n_27390), .o(n_27494) );
no02f04 TIMEBOOST_cell_3409 ( .a(TIMEBOOST_net_995), .b(n_27392), .o(n_27498) );
na02s02 g763529 ( .a(n_17108), .b(FE_OCP_RBN3060_n_15595), .o(n_17114) );
na02s06 g763530 ( .a(n_16843), .b(n_16089), .o(n_16941) );
na02s01 g763531 ( .a(n_16089), .b(n_17108), .o(n_17113) );
in01s01 g763534 ( .a(n_16976), .o(n_17022) );
na02s02 g763535 ( .a(n_16814), .b(n_16940), .o(n_16976) );
ao12f04 g763537 ( .a(n_16751), .b(n_16827), .c(n_16726), .o(n_16938) );
oa22f02 g763538 ( .a(n_16810), .b(FE_OCP_RBN3193_n_15599), .c(n_16781), .d(n_16339), .o(n_16873) );
in01f02 g763539 ( .a(n_16916), .o(n_16872) );
no02s06 TIMEBOOST_cell_4203 ( .a(FE_RN_768_0), .b(n_6641), .o(TIMEBOOST_net_1192) );
in01f01 g763542 ( .a(n_16793), .o(n_16811) );
ao12f08 g763543 ( .a(n_16667), .b(n_16690), .c(n_16708), .o(n_16793) );
in01s01 g763545 ( .a(n_16912), .o(n_16919) );
in01m08 g763546 ( .a(n_16836), .o(n_16912) );
in01m06 g763566 ( .a(n_16836), .o(n_16923) );
no02m10 g763570 ( .a(n_16764), .b(n_16717), .o(n_16836) );
in01f02 g763571 ( .a(n_17128), .o(n_17061) );
no02s01 TIMEBOOST_cell_1510 ( .a(TIMEBOOST_net_369), .b(n_3212), .o(n_3213) );
in01s03 g763573 ( .a(n_16868), .o(n_16869) );
no02m08 g763574 ( .a(n_16796), .b(n_15657), .o(n_16868) );
no02s01 g763575 ( .a(n_16814), .b(n_16866), .o(n_16867) );
no02s02 g763576 ( .a(n_17108), .b(FE_OCPN1644_n_16866), .o(n_17451) );
na02s20 g763579 ( .a(n_16988), .b(n_16900), .o(n_17129) );
na02s02 g763581 ( .a(n_17535), .b(n_17609), .o(n_17613) );
no02s06 g763583 ( .a(n_17575), .b(n_17574), .o(n_17611) );
in01s06 g763585 ( .a(n_16899), .o(n_16973) );
na02s20 g763589 ( .a(n_44365), .b(n_16807), .o(n_16899) );
na02s02 TIMEBOOST_cell_5023 ( .a(TIMEBOOST_net_1459), .b(n_44867), .o(n_38001) );
in01s10 g763591 ( .a(n_17192), .o(n_17020) );
no02m04 TIMEBOOST_cell_5042 ( .a(n_37884), .b(n_44867), .o(TIMEBOOST_net_1469) );
no02s06 g763593 ( .a(n_17539), .b(n_17465), .o(n_17540) );
no02s02 g763594 ( .a(n_17374), .b(n_17496), .o(n_17432) );
in01s01 g763595 ( .a(n_17577), .o(n_17503) );
no02f10 g763596 ( .a(n_17375), .b(n_17156), .o(n_17577) );
na02s01 g763597 ( .a(n_17610), .b(n_17609), .o(n_18326) );
no02s01 g763598 ( .a(n_17607), .b(n_17604), .o(n_17608) );
na02s01 g763599 ( .a(n_17430), .b(n_17421), .o(n_17431) );
no02s08 g763600 ( .a(n_16712), .b(n_16716), .o(n_16717) );
no02m08 g763601 ( .a(n_16713), .b(n_16735), .o(n_16764) );
no02s01 TIMEBOOST_cell_1509 ( .a(n_2706), .b(n_2661), .o(TIMEBOOST_net_369) );
no02m08 TIMEBOOST_cell_8582 ( .a(FE_OCP_RBN5898_n_35005), .b(n_30546), .o(TIMEBOOST_net_2778) );
na02m02 g763604 ( .a(n_16731), .b(n_16736), .o(n_16763) );
no02s06 TIMEBOOST_cell_4202 ( .a(TIMEBOOST_net_1191), .b(FE_RN_690_0), .o(FE_RN_692_0) );
in01s02 g763606 ( .a(n_16833), .o(n_16834) );
na02m04 g763607 ( .a(n_16809), .b(n_16761), .o(n_16833) );
in01s02 g763608 ( .a(n_16808), .o(n_16880) );
no02s04 g763609 ( .a(n_16791), .b(FE_OCP_RBN3048_n_15200), .o(n_16808) );
ao12s01 g763610 ( .a(n_17575), .b(n_17423), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_29_), .o(n_18382) );
na02m04 g763611 ( .a(FE_OCP_RBN3048_n_15200), .b(n_16791), .o(n_16879) );
in01f02 g763615 ( .a(n_16864), .o(n_16865) );
na02m04 g763616 ( .a(n_16758), .b(n_16832), .o(n_16864) );
in01m04 g763617 ( .a(n_17471), .o(n_17541) );
oa12m04 g763618 ( .a(n_17430), .b(n_17208), .c(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17471) );
in01f06 g763619 ( .a(n_17502), .o(n_17576) );
oa12f08 g763620 ( .a(n_17470), .b(n_17469), .c(n_17262), .o(n_17502) );
ao12s01 g763621 ( .a(n_17663), .b(n_17732), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_30_), .o(n_18385) );
oa12s06 g763622 ( .a(n_17498), .b(n_17573), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_29_), .o(n_17665) );
ao12s01 g763623 ( .a(n_17373), .b(n_17372), .c(n_17371), .o(n_18417) );
oa22f02 g763624 ( .a(n_46977), .b(FE_OCP_RBN3193_n_15599), .c(n_16705), .d(n_17753), .o(n_16789) );
oa22f02 g763625 ( .a(n_46976), .b(FE_OCP_RBN3193_n_15599), .c(n_16774), .d(n_16339), .o(n_16863) );
in01s06 g763634 ( .a(n_16977), .o(n_17108) );
in01s10 g763643 ( .a(n_16843), .o(n_16977) );
in01m10 g763646 ( .a(n_16796), .o(n_16843) );
in01m08 g763647 ( .a(n_16814), .o(n_16796) );
na02m10 g763648 ( .a(n_16714), .b(n_16671), .o(n_16814) );
in01f02 g763650 ( .a(n_46975), .o(n_16895) );
in01s01 g763652 ( .a(n_18404), .o(n_16931) );
oa12s01 g763653 ( .a(n_16828), .b(n_16829), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_0_), .o(n_18404) );
in01s01 g763654 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_15_), .o(n_18159) );
in01s20 g763656 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_2_), .o(n_16807) );
in01s01 g763658 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_16_), .o(n_16830) );
in01s10 g763661 ( .a(n_16893), .o(n_16894) );
in01s10 g763662 ( .a(n_16900), .o(n_16893) );
na02s40 g763663 ( .a(n_44365), .b(n_44720), .o(n_16900) );
in01s01 g763665 ( .a(n_16857), .o(n_17437) );
na02s04 TIMEBOOST_cell_5041 ( .a(TIMEBOOST_net_1468), .b(n_24500), .o(TIMEBOOST_net_1059) );
na02s06 g763668 ( .a(n_17212), .b(FE_OFN736_n_17093), .o(n_17609) );
na02s06 g763669 ( .a(n_17614), .b(n_17468), .o(n_17539) );
in01f08 g763670 ( .a(n_17374), .o(n_17375) );
na02f10 g763671 ( .a(n_17372), .b(n_17257), .o(n_17374) );
no02s02 g763672 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_30_), .b(n_17423), .o(n_17663) );
no02s06 g763673 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_29_), .b(n_17423), .o(n_17575) );
no02s01 g763674 ( .a(n_17372), .b(n_17371), .o(n_17373) );
na02s01 g763675 ( .a(n_16829), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_0_), .o(n_16828) );
na02s02 g763676 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_27_), .b(n_17423), .o(n_17610) );
na02m08 g763677 ( .a(n_17365), .b(n_17428), .o(n_17429) );
no02s01 g763678 ( .a(n_17605), .b(n_17604), .o(n_18293) );
na02s01 g763679 ( .a(n_17306), .b(n_17055), .o(n_17370) );
na02s01 g763680 ( .a(n_17367), .b(n_17098), .o(n_17369) );
na02s06 g763681 ( .a(n_16649), .b(n_16397), .o(n_16671) );
na02m08 g763682 ( .a(n_16650), .b(n_16396), .o(n_16714) );
na02f03 g763684 ( .a(n_16755), .b(n_16728), .o(n_16787) );
in01f01 g763686 ( .a(n_16827), .o(n_16855) );
na02f08 g763687 ( .a(n_16750), .b(n_16734), .o(n_16827) );
no02f02 g763689 ( .a(n_16762), .b(n_16707), .o(n_16785) );
na02s06 g763690 ( .a(n_16739), .b(FE_OCP_RBN3037_n_15079), .o(n_16809) );
in01m02 g763691 ( .a(n_16760), .o(n_16761) );
no02m06 g763692 ( .a(n_16739), .b(FE_OCP_RBN3037_n_15079), .o(n_16760) );
na02s04 g763693 ( .a(n_16749), .b(n_16726), .o(n_16784) );
in01f02 g763694 ( .a(n_16759), .o(n_16832) );
no02f02 g763695 ( .a(n_16719), .b(FE_OCP_RBN3007_n_15206), .o(n_16759) );
no02s04 g763696 ( .a(n_17266), .b(n_17210), .o(n_17430) );
na02s06 g763698 ( .a(n_17265), .b(n_17367), .o(n_17368) );
in01s01 g763699 ( .a(n_17706), .o(n_17707) );
ao12s01 g763700 ( .a(n_17533), .b(n_17423), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_25_), .o(n_17706) );
in01s02 g763702 ( .a(n_16758), .o(n_16782) );
na02m04 g763703 ( .a(FE_OCP_RBN3007_n_15206), .b(n_16719), .o(n_16758) );
in01s01 g763704 ( .a(n_17537), .o(n_17607) );
oa12s02 g763705 ( .a(n_17498), .b(n_17497), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_25_), .o(n_17537) );
in01m04 g763706 ( .a(n_16712), .o(n_16713) );
ao12m08 g763707 ( .a(n_46426), .b(n_16643), .c(n_47268), .o(n_16712) );
na02s06 g763708 ( .a(n_16733), .b(n_16778), .o(n_16998) );
oa22f02 g763709 ( .a(n_16757), .b(n_17336), .c(n_16725), .d(n_17753), .o(n_16804) );
in01f02 g763710 ( .a(n_16810), .o(n_16781) );
no02f04 TIMEBOOST_cell_1522 ( .a(TIMEBOOST_net_375), .b(n_8462), .o(n_8540) );
in01f02 g763712 ( .a(n_16736), .o(n_16737) );
in01f01 g763713 ( .a(n_16690), .o(n_16736) );
ao12f08 g763714 ( .a(n_16603), .b(n_16646), .c(n_16641), .o(n_16690) );
ao22s01 g763716 ( .a(n_17259), .b(n_17427), .c(n_17258), .d(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_18418) );
in01s02 g763723 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_27_), .o(n_17212) );
in01s01 g763725 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_15_), .o(n_16779) );
no02s06 g763730 ( .a(n_17309), .b(n_17310), .o(n_17614) );
no02f10 g763731 ( .a(n_17260), .b(n_17211), .o(n_17470) );
in01s01 g763732 ( .a(n_17536), .o(n_17604) );
na02s02 g763733 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_26_), .b(n_17423), .o(n_17536) );
in01s01 g763734 ( .a(n_17605), .o(n_17535) );
no02s06 g763735 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_26_), .b(n_17423), .o(n_17605) );
no02m01 g763737 ( .a(n_17498), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_25_), .o(n_17533) );
na02s01 g763738 ( .a(n_17428), .b(n_17468), .o(n_18234) );
no02s01 g763739 ( .a(n_17574), .b(n_17573), .o(n_18350) );
na02s01 g763740 ( .a(n_17532), .b(n_17466), .o(n_18255) );
no02f04 g763742 ( .a(n_16685), .b(n_16600), .o(n_16755) );
in01f04 g763743 ( .a(n_16733), .o(n_16734) );
no02f08 g763744 ( .a(n_16684), .b(FE_OCP_RBN4459_FE_RN_1190_0), .o(n_16733) );
na02s02 TIMEBOOST_cell_5571 ( .a(TIMEBOOST_net_1733), .b(n_6369), .o(n_6500) );
no02f04 TIMEBOOST_cell_1521 ( .a(FE_OCP_RBN4141_n_7743), .b(n_8455), .o(TIMEBOOST_net_375) );
in01m02 g763747 ( .a(n_16731), .o(n_16732) );
na02m02 g763748 ( .a(n_16708), .b(n_16668), .o(n_16731) );
no02s06 g763749 ( .a(n_46978), .b(FE_OCP_RBN3012_n_14985), .o(n_16762) );
in01f01 g763750 ( .a(n_16706), .o(n_16707) );
na02f06 g763751 ( .a(n_46978), .b(FE_OCP_RBN3012_n_14985), .o(n_16706) );
in01f06 g763752 ( .a(n_16801), .o(n_16802) );
in01s01 g763754 ( .a(n_16825), .o(n_16826) );
na02f04 g763755 ( .a(n_16727), .b(n_16726), .o(n_16825) );
no02f02 g763757 ( .a(n_16777), .b(n_16715), .o(n_16753) );
no02s01 TIMEBOOST_cell_1546 ( .a(TIMEBOOST_net_387), .b(n_42782), .o(n_42821) );
oa12f10 g763759 ( .a(n_17202), .b(n_17096), .c(n_17427), .o(n_17372) );
ao12s06 g763760 ( .a(n_17308), .b(n_17207), .c(n_17152), .o(n_17469) );
in01s01 g763761 ( .a(n_17704), .o(n_17705) );
ao12s01 g763762 ( .a(n_17310), .b(n_17423), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_21_), .o(n_17704) );
in01s01 g763763 ( .a(n_17702), .o(n_17703) );
ao12s01 g763764 ( .a(n_17211), .b(n_17423), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_19_), .o(n_17702) );
no02s06 g763765 ( .a(n_16715), .b(n_16751), .o(n_16752) );
no02s06 g763766 ( .a(n_16748), .b(n_16777), .o(n_16778) );
in01s01 g763768 ( .a(n_17266), .o(n_17306) );
no02s03 g763769 ( .a(n_17107), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17266) );
in01s01 g763771 ( .a(n_17367), .o(n_17305) );
no03m02 TIMEBOOST_cell_2248 ( .a(TIMEBOOST_net_93), .b(n_17971), .c(n_18004), .o(n_18093) );
oa12s06 g763773 ( .a(n_17015), .b(n_17263), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_7_), .o(n_17265) );
in01s01 g763774 ( .a(n_17365), .o(n_17366) );
oa12m08 g763775 ( .a(n_17101), .b(n_17304), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_21_), .o(n_17365) );
ao12f10 g763776 ( .a(FE_OFN736_n_17093), .b(n_17261), .c(n_17057), .o(n_17262) );
in01s04 g763777 ( .a(n_16649), .o(n_16650) );
oa12m08 g763778 ( .a(n_16373), .b(n_16609), .c(n_16232), .o(n_16649) );
oa22f02 g763779 ( .a(n_16686), .b(FE_OCP_RBN3193_n_15599), .c(n_16658), .d(n_16339), .o(n_16730) );
in01m02 g763780 ( .a(n_46977), .o(n_16705) );
na02m06 g763782 ( .a(n_16648), .b(n_16629), .o(n_16739) );
ao22s10 g763783 ( .a(FE_OCP_RBN7107_n_44365), .b(FE_OCP_RBN4590_n_44847), .c(FE_OCP_RBN7109_n_44365), .d(n_44847), .o(n_16829) );
in01m02 g763784 ( .a(n_46976), .o(n_16774) );
in01f04 g763786 ( .a(n_16749), .o(n_16750) );
na02m06 TIMEBOOST_cell_8815 ( .a(TIMEBOOST_net_2894), .b(n_11251), .o(TIMEBOOST_net_2290) );
in01s01 g763789 ( .a(n_18483), .o(n_16968) );
ao12s01 g763790 ( .a(n_16854), .b(n_16853), .c(delay_add_ln22_unr11_stage5_stallmux_q_0_), .o(n_18483) );
no02s06 g763794 ( .a(n_17362), .b(n_17363), .o(n_17364) );
no02s20 g763796 ( .a(FE_OCP_RBN7112_n_44365), .b(n_44847), .o(n_16936) );
na02m20 g763797 ( .a(n_44365), .b(FE_OCP_RBN4590_n_44847), .o(n_16988) );
na02s06 g763798 ( .a(n_16799), .b(delay_add_ln22_unr11_stage5_stallmux_q_0_), .o(n_17226) );
in01s01 g763799 ( .a(n_17467), .o(n_17573) );
na02s02 g763800 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_28_), .b(n_17101), .o(n_17467) );
in01s01 g763801 ( .a(n_17465), .o(n_17466) );
no02s06 g763802 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_23_), .b(n_17423), .o(n_17465) );
in01s06 g763803 ( .a(n_17358), .o(n_17468) );
no02s03 g763804 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_22_), .b(n_17101), .o(n_17358) );
no02s06 g763805 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_21_), .b(n_17101), .o(n_17310) );
no02s20 g763806 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_19_), .b(n_17101), .o(n_17211) );
no02s06 g763807 ( .a(n_17422), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_15_), .o(n_17424) );
no02s06 g763808 ( .a(n_17100), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_13_), .o(n_17208) );
no02s04 g763809 ( .a(n_17106), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_), .o(n_17107) );
na02m06 TIMEBOOST_cell_3997 ( .a(n_14511), .b(FE_OCP_RBN5803_FE_RN_2224_0), .o(TIMEBOOST_net_1089) );
no02s02 TIMEBOOST_cell_5956 ( .a(TIMEBOOST_net_1829), .b(n_32534), .o(n_32604) );
na02s06 g763812 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_23_), .b(n_17423), .o(n_17532) );
na02s02 g763813 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_22_), .b(n_17101), .o(n_17428) );
in01s01 g763814 ( .a(n_17574), .o(n_17531) );
no02m01 g763815 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_28_), .b(n_17498), .o(n_17574) );
no02s01 g763816 ( .a(n_16853), .b(delay_add_ln22_unr11_stage5_stallmux_q_0_), .o(n_16854) );
no02s01 g763817 ( .a(n_17153), .b(n_17308), .o(n_18083) );
no02s01 g763818 ( .a(n_17154), .b(n_17260), .o(n_18141) );
no02s01 g763819 ( .a(n_17572), .b(n_17497), .o(n_18211) );
in01s01 g763820 ( .a(n_17356), .o(n_17357) );
no02s01 g763821 ( .a(n_17309), .b(n_17304), .o(n_17356) );
no02s01 g763822 ( .a(n_17464), .b(n_17463), .o(n_17992) );
no02s01 g763823 ( .a(n_17362), .b(n_17422), .o(n_17958) );
no02s01 g763824 ( .a(n_17355), .b(n_17263), .o(n_17818) );
no02s01 g763825 ( .a(n_17354), .b(n_17104), .o(n_17961) );
no02s01 g763826 ( .a(n_17530), .b(n_17106), .o(n_17902) );
no02s01 g763827 ( .a(n_17462), .b(n_17099), .o(n_17711) );
in01s01 g763828 ( .a(n_17258), .o(n_17259) );
na02s01 g763829 ( .a(n_17097), .b(n_17202), .o(n_17258) );
na02s01 g763830 ( .a(n_17157), .b(n_17257), .o(n_17371) );
na02s01 g763831 ( .a(n_17421), .b(n_17300), .o(n_17980) );
na02s04 g763832 ( .a(n_16612), .b(n_16464), .o(n_16648) );
na02s04 g763833 ( .a(n_16611), .b(n_16465), .o(n_16629) );
in01f02 g763834 ( .a(n_16684), .o(n_16685) );
na02f08 g763835 ( .a(n_16637), .b(n_16640), .o(n_16684) );
na02f01 g763837 ( .a(n_16640), .b(n_16656), .o(n_16703) );
na02f02 g763839 ( .a(n_16607), .b(n_16585), .o(n_16628) );
in01s02 g763840 ( .a(n_16669), .o(n_16670) );
in01s01 g763841 ( .a(n_16646), .o(n_16669) );
na02m06 g763843 ( .a(n_16645), .b(FE_OCP_RBN3006_n_14905), .o(n_16708) );
in01s02 g763844 ( .a(n_16667), .o(n_16668) );
no02f06 g763845 ( .a(n_16645), .b(FE_OCP_RBN3006_n_14905), .o(n_16667) );
no02f02 g763847 ( .a(n_16682), .b(FE_OCP_RBN4459_FE_RN_1190_0), .o(n_16728) );
in01m02 g763848 ( .a(n_16751), .o(n_16727) );
no02f08 g763849 ( .a(n_16702), .b(FE_OCP_RBN2092_n_14991), .o(n_16751) );
in01s02 g763851 ( .a(n_16726), .o(n_16748) );
na02m08 g763852 ( .a(FE_OCP_RBN2092_n_14991), .b(n_16702), .o(n_16726) );
no02s04 g763853 ( .a(n_16638), .b(FE_OCP_RBN2102_n_15083), .o(n_16715) );
no02f04 g763854 ( .a(n_16639), .b(n_15083), .o(n_16777) );
ao12s01 g763855 ( .a(n_17425), .b(n_17256), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_11_), .o(n_17986) );
ao12s01 g763856 ( .a(n_17360), .b(n_17256), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_13_), .o(n_18033) );
ao12s01 g763857 ( .a(n_17363), .b(n_17256), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_15_), .o(n_17989) );
in01s01 g763858 ( .a(n_17602), .o(n_17603) );
ao12s01 g763859 ( .a(n_17297), .b(n_17256), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_7_), .o(n_17602) );
no02f06 TIMEBOOST_cell_3401 ( .a(n_36552), .b(TIMEBOOST_net_991), .o(n_36655) );
oa22m02 g763861 ( .a(n_46979), .b(n_17584), .c(n_16634), .d(FE_OCP_RBN3196_n_15599), .o(n_16700) );
oa22m02 g763862 ( .a(n_16699), .b(n_17336), .c(n_16681), .d(n_16339), .o(n_16747) );
in01s02 g763865 ( .a(n_16643), .o(n_16665) );
na02s06 g763866 ( .a(n_16590), .b(n_16534), .o(n_16643) );
in01m02 g763867 ( .a(n_16757), .o(n_16725) );
no02s01 TIMEBOOST_cell_4095 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(FE_RN_1873_0), .o(TIMEBOOST_net_1138) );
oa22s01 g763869 ( .a(n_16928), .b(n_16310), .c(n_16929), .d(n_16311), .o(n_17058) );
oa22s01 g763870 ( .a(FE_OCP_RBN6212_n_16962), .b(n_16260), .c(n_16962), .d(n_16259), .o(n_17103) );
oa22s01 g763871 ( .a(n_16961), .b(n_16308), .c(n_16960), .d(n_16309), .o(n_17102) );
oa22s01 g763872 ( .a(n_17256), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_), .c(n_16618), .d(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17983) );
oa22s01 g763873 ( .a(n_17158), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .c(n_17256), .d(delay_sub_ln23_0_unr12_stage5_stallmux_q_5_), .o(n_17788) );
in01s01 g763874 ( .a(n_17526), .o(n_17527) );
oa22s01 g763875 ( .a(n_17256), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_3_), .c(n_17496), .d(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17526) );
in01s01 g763876 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_13_), .o(n_18048) );
in01s20 g763889 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_19_), .o(n_17057) );
in01s02 g763891 ( .a(n_17353), .o(n_17497) );
na02s01 g763892 ( .a(n_17101), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_24_), .o(n_17353) );
no02m03 g763893 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_20_), .b(n_17101), .o(n_17309) );
no02s20 g763894 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_18_), .b(n_17101), .o(n_17260) );
no02s06 g763895 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_17_), .b(n_17498), .o(n_17308) );
no02m01 g763896 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_16_), .b(n_17256), .o(n_17464) );
in01s01 g763897 ( .a(n_17302), .o(n_17422) );
na02s06 g763898 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_14_), .b(n_17255), .o(n_17302) );
in01s02 g763899 ( .a(n_17421), .o(n_17100) );
na02s01 g763900 ( .a(n_17054), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_12_), .o(n_17421) );
in01s01 g763901 ( .a(n_17106), .o(n_17056) );
no02s03 g763902 ( .a(n_16591), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17106) );
in01s01 g763903 ( .a(n_17104), .o(n_17055) );
no02s02 g763904 ( .a(n_16617), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17104) );
no02s01 g763905 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_15_), .b(n_17256), .o(n_17363) );
in01s01 g763906 ( .a(n_17362), .o(n_17301) );
no02m01 g763907 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_14_), .b(n_17256), .o(n_17362) );
no02s01 g763908 ( .a(n_17255), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_13_), .o(n_17360) );
in01s01 g763909 ( .a(n_17359), .o(n_17300) );
no02s01 g763910 ( .a(n_17054), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_12_), .o(n_17359) );
no02s02 g763911 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_11_), .b(n_17015), .o(n_17425) );
in01s01 g763912 ( .a(n_17354), .o(n_17299) );
no02s02 g763913 ( .a(n_17255), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_10_), .o(n_17354) );
in01s01 g763914 ( .a(n_17159), .o(n_17099) );
na02s02 g763915 ( .a(n_17054), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_4_), .o(n_17159) );
in01s02 g763916 ( .a(n_17098), .o(n_17263) );
na02s06 g763917 ( .a(n_17054), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_6_), .o(n_17098) );
in01s02 g763918 ( .a(n_17297), .o(n_17298) );
no02s01 g763919 ( .a(n_17255), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_7_), .o(n_17297) );
no02m01 g763920 ( .a(n_17054), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_6_), .o(n_17355) );
na02f20 g763921 ( .a(FE_OCP_RBN3845_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_1_), .o(n_17202) );
in01s01 g763922 ( .a(n_17096), .o(n_17097) );
no02f20 g763923 ( .a(FE_OCP_RBN3844_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_1_), .o(n_17096) );
na02s10 g763924 ( .a(n_17018), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17257) );
in01s01 g763925 ( .a(n_17156), .o(n_17157) );
no02s06 g763926 ( .a(n_17018), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17156) );
in01s10 g763927 ( .a(n_17155), .o(n_17304) );
na02s40 g763928 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_20_), .b(n_17101), .o(n_17155) );
in01s01 g763929 ( .a(n_17261), .o(n_17154) );
na02m40 g763930 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_18_), .b(n_17101), .o(n_17261) );
in01s01 g763931 ( .a(n_17207), .o(n_17463) );
na02s06 g763932 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_16_), .b(n_17015), .o(n_17207) );
in01s01 g763933 ( .a(n_17152), .o(n_17153) );
na02s06 g763934 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_17_), .b(n_17101), .o(n_17152) );
no02s01 g763936 ( .a(n_17423), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_24_), .o(n_17572) );
no02s01 g763937 ( .a(n_17256), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_4_), .o(n_17462) );
no02s01 g763938 ( .a(n_17256), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_8_), .o(n_17530) );
no03f04 TIMEBOOST_cell_8375 ( .a(FE_RN_2472_0), .b(n_45101), .c(n_20615), .o(n_20641) );
no02m10 TIMEBOOST_cell_8489 ( .a(TIMEBOOST_net_2731), .b(n_17972), .o(n_18077) );
in01s01 g763941 ( .a(n_16611), .o(n_16612) );
no02s04 g763942 ( .a(n_16570), .b(n_16533), .o(n_16611) );
na02s06 g763943 ( .a(n_16570), .b(n_16441), .o(n_16590) );
in01m02 g763944 ( .a(n_16661), .o(n_16662) );
na02f02 g763945 ( .a(n_16604), .b(n_16641), .o(n_16661) );
na02s02 TIMEBOOST_cell_4905 ( .a(TIMEBOOST_net_1400), .b(n_23027), .o(n_23088) );
ao12f08 g763951 ( .a(n_16583), .b(n_16560), .c(n_16562), .o(n_16640) );
ao12s02 g763953 ( .a(n_17255), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_8_), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_), .o(n_17426) );
no02s06 TIMEBOOST_cell_1548 ( .a(TIMEBOOST_net_388), .b(n_38650), .o(n_38683) );
in01s01 g763956 ( .a(n_16609), .o(n_16626) );
oa12s06 g763957 ( .a(n_16399), .b(n_16532), .c(n_16431), .o(n_16609) );
in01m02 g763958 ( .a(n_16686), .o(n_16658) );
no02s04 TIMEBOOST_cell_6730 ( .a(TIMEBOOST_net_2122), .b(n_24808), .o(n_24830) );
oa12f01 g763961 ( .a(n_16564), .b(n_16565), .c(n_16535), .o(n_16607) );
na02m06 g763962 ( .a(n_16569), .b(n_16537), .o(n_16645) );
in01s01 g763964 ( .a(n_16799), .o(n_16853) );
oa22s01 g763966 ( .a(n_16851), .b(n_16300), .c(n_16850), .d(n_16301), .o(n_16967) );
oa22s01 g763967 ( .a(n_16889), .b(n_16064), .c(n_16890), .d(n_16063), .o(n_17017) );
in01f02 g763968 ( .a(n_16638), .o(n_16639) );
in01s01 g763976 ( .a(n_17783), .o(n_17815) );
in01s02 g763977 ( .a(FE_OFN739_n_17093), .o(n_17783) );
in01s01 g763978 ( .a(FE_OFN739_n_17093), .o(n_19222) );
in01s02 g764009 ( .a(n_18140), .o(n_18230) );
in01s06 g764012 ( .a(n_18119), .o(n_18140) );
in01s01 g764013 ( .a(n_19418), .o(n_19645) );
in01s06 g764015 ( .a(n_19418), .o(n_18119) );
in01s06 g764016 ( .a(n_18032), .o(n_19418) );
in01s01 g764024 ( .a(n_18099), .o(n_18117) );
in01s02 g764026 ( .a(n_18032), .o(n_18099) );
in01s06 g764033 ( .a(n_18032), .o(n_18010) );
in01s06 g764034 ( .a(n_17900), .o(n_18032) );
in01s01 g764039 ( .a(n_19170), .o(FE_RN_1458_0) );
in01s01 g764040 ( .a(n_17900), .o(n_19170) );
in01s06 g764043 ( .a(n_17881), .o(n_17900) );
in01m06 g764044 ( .a(FE_OFN738_n_17093), .o(n_17881) );
in01s02 g764051 ( .a(FE_OFN736_n_17093), .o(n_17732) );
in01s03 g764055 ( .a(FE_OFN737_n_17093), .o(n_17661) );
in01s02 g764064 ( .a(FE_OFN736_n_17093), .o(n_17498) );
in01s03 g764067 ( .a(FE_OFN736_n_17093), .o(n_17423) );
in01s40 g764075 ( .a(FE_OFN736_n_17093), .o(n_17101) );
in01s02 g764087 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17256) );
in01s02 g764090 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17255) );
in01s02 g764097 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17015) );
in01s06 g764099 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17054) );
na02s02 TIMEBOOST_cell_8823 ( .a(TIMEBOOST_net_2898), .b(n_3685), .o(n_3890) );
na02s04 g764105 ( .a(n_16500), .b(n_16370), .o(n_16537) );
na02s03 g764107 ( .a(n_16518), .b(n_16495), .o(n_16567) );
no02f04 TIMEBOOST_cell_5569 ( .a(n_31060), .b(TIMEBOOST_net_1732), .o(n_31165) );
no02s02 TIMEBOOST_cell_1401 ( .a(n_7864), .b(n_7925), .o(TIMEBOOST_net_315) );
na02f06 g764110 ( .a(n_16565), .b(n_16564), .o(n_16566) );
in01f01 g764111 ( .a(n_16603), .o(n_16604) );
no02f06 g764112 ( .a(n_16588), .b(FE_OCP_RBN2983_n_14814), .o(n_16603) );
na02s06 g764113 ( .a(n_16588), .b(FE_OCP_RBN2983_n_14814), .o(n_16641) );
na02f02 g764115 ( .a(n_16620), .b(n_16637), .o(n_16656) );
in01m02 g764116 ( .a(n_16624), .o(n_16625) );
ao12m04 g764117 ( .a(n_16524), .b(n_16552), .c(n_16580), .o(n_16624) );
oa12s01 g764119 ( .a(n_16017), .b(n_16930), .c(n_16099), .o(n_16962) );
in01s01 g764120 ( .a(n_16960), .o(n_16961) );
ao12s01 g764121 ( .a(n_16134), .b(n_16930), .c(n_16261), .o(n_16960) );
in01s01 g764122 ( .a(n_16928), .o(n_16929) );
oa12s01 g764123 ( .a(n_16065), .b(n_16852), .c(n_16021), .o(n_16928) );
oa22f02 g764124 ( .a(n_16601), .b(n_17584), .c(n_16578), .d(FE_OCP_RBN3196_n_15599), .o(n_16636) );
in01s02 g764125 ( .a(n_46979), .o(n_16634) );
no02s01 g764128 ( .a(n_16563), .b(n_16475), .o(n_16585) );
no02s02 TIMEBOOST_cell_1142 ( .a(TIMEBOOST_net_185), .b(n_37586), .o(n_37611) );
in01m02 g764130 ( .a(n_16699), .o(n_16681) );
oa22m02 g764131 ( .a(n_16576), .b(n_16594), .c(n_16552), .d(n_16595), .o(n_16699) );
oa22s01 g764134 ( .a(n_16821), .b(n_15962), .c(n_16820), .d(n_15963), .o(n_16927) );
oa22s01 g764135 ( .a(n_16886), .b(n_16132), .c(n_16885), .d(n_16131), .o(n_17014) );
oa22m02 g764136 ( .a(n_16602), .b(n_17584), .c(n_16579), .d(FE_OCP_RBN3196_n_15599), .o(n_16633) );
oa22s01 g764137 ( .a(n_16819), .b(n_16250), .c(n_16818), .d(n_16249), .o(n_16926) );
oa22s01 g764138 ( .a(n_16817), .b(n_16304), .c(n_16816), .d(n_16305), .o(n_16925) );
oa22s01 g764139 ( .a(n_16823), .b(n_16257), .c(n_16822), .d(n_16256), .o(n_16924) );
in01s01 g764146 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_13_), .o(n_18152) );
na02s01 TIMEBOOST_cell_7017 ( .a(FE_RN_1275_0), .b(FE_RN_1606_0), .o(TIMEBOOST_net_2267) );
no02s02 g764152 ( .a(n_16499), .b(n_16446), .o(n_16500) );
na02s06 g764153 ( .a(n_16499), .b(n_46421), .o(n_16518) );
no02s06 g764154 ( .a(n_16533), .b(n_16332), .o(n_16534) );
no02f06 g764155 ( .a(n_16561), .b(n_16516), .o(n_16562) );
na02f08 g764156 ( .a(n_16526), .b(n_16515), .o(n_16560) );
in01s01 g764157 ( .a(n_16889), .o(n_16890) );
na02s01 g764158 ( .a(n_16852), .b(n_16102), .o(n_16889) );
na02s02 g764160 ( .a(n_16527), .b(n_16486), .o(n_16559) );
in01s01 g764161 ( .a(n_16557), .o(n_16558) );
in01s01 g764162 ( .a(n_16565), .o(n_16557) );
ao12f06 g764163 ( .a(n_16461), .b(n_16439), .c(n_16437), .o(n_16565) );
in01m01 g764164 ( .a(n_16555), .o(n_16556) );
na02m01 g764165 ( .a(n_16494), .b(n_16564), .o(n_16555) );
no02s01 g764166 ( .a(n_16474), .b(FE_OCP_RBN4319_n_14768), .o(n_16475) );
no02m08 g764167 ( .a(n_16468), .b(FE_OCP_RBN2973_n_14768), .o(n_16563) );
no02s02 TIMEBOOST_cell_7075 ( .a(n_39910), .b(n_39965), .o(TIMEBOOST_net_2296) );
in01f01 g764170 ( .a(n_16600), .o(n_16620) );
no02f06 g764171 ( .a(n_16582), .b(FE_OCPN1642_FE_OCP_RBN1596_n_14823), .o(n_16600) );
in01s01 g764172 ( .a(n_16598), .o(n_16599) );
no02s02 g764173 ( .a(n_16583), .b(n_16561), .o(n_16598) );
na02m06 g764174 ( .a(n_16582), .b(FE_OCPN1642_FE_OCP_RBN1596_n_14823), .o(n_16637) );
in01m02 g764176 ( .a(n_16532), .o(n_16553) );
na02f08 g764177 ( .a(n_16469), .b(n_16445), .o(n_16532) );
na02m08 g764179 ( .a(n_16529), .b(n_16406), .o(n_16596) );
in01s01 g764180 ( .a(n_16850), .o(n_16851) );
ao12s01 g764181 ( .a(n_16173), .b(n_16824), .c(n_16255), .o(n_16850) );
in01m01 g764182 ( .a(n_16887), .o(n_16888) );
oa12m02 g764183 ( .a(n_16313), .b(FE_OCP_RBN6186_n_16824), .c(n_16262), .o(n_16887) );
no02f08 TIMEBOOST_cell_1134 ( .a(TIMEBOOST_net_181), .b(n_37579), .o(n_37755) );
oa22s01 g764185 ( .a(n_16824), .b(n_16306), .c(FE_OCP_RBN6186_n_16824), .d(n_16307), .o(n_16849) );
in01s01 g764187 ( .a(n_16499), .o(n_16472) );
na02m08 TIMEBOOST_cell_7705 ( .a(TIMEBOOST_net_2483), .b(n_24532), .o(n_24648) );
no02f04 g764189 ( .a(n_16443), .b(n_16435), .o(n_16497) );
no02f06 TIMEBOOST_cell_1133 ( .a(n_37602), .b(n_37659), .o(TIMEBOOST_net_181) );
na02s06 g764191 ( .a(n_16495), .b(n_16442), .o(n_16533) );
in01m02 g764192 ( .a(n_16594), .o(n_16595) );
na02s02 g764193 ( .a(n_16580), .b(n_16515), .o(n_16594) );
in01f02 g764194 ( .a(n_16530), .o(n_16531) );
na02f06 g764195 ( .a(n_16401), .b(n_16490), .o(n_16530) );
na02m08 g764196 ( .a(n_16491), .b(n_16368), .o(n_16529) );
na02s01 g764197 ( .a(n_16824), .b(n_15927), .o(n_16852) );
in01m01 g764198 ( .a(n_16535), .o(n_16494) );
no02f06 g764199 ( .a(n_16471), .b(FE_OCP_RBN2927_n_14684), .o(n_16535) );
na02s04 g764200 ( .a(n_16471), .b(FE_OCP_RBN2927_n_14684), .o(n_16564) );
no02f06 g764201 ( .a(n_16484), .b(FE_OCP_RBN1599_n_14763), .o(n_16583) );
no02f04 g764202 ( .a(n_47340), .b(FE_OCP_RBN1600_n_14763), .o(n_16561) );
in01s01 g764204 ( .a(n_16822), .o(n_16823) );
ao12s01 g764205 ( .a(n_16022), .b(n_16798), .c(n_15880), .o(n_16822) );
in01s01 g764206 ( .a(n_16820), .o(n_16821) );
ao12s01 g764207 ( .a(n_16210), .b(n_16798), .c(n_15929), .o(n_16820) );
in01s01 g764208 ( .a(n_16885), .o(n_16886) );
in01s01 g764209 ( .a(n_16930), .o(n_16885) );
na02s01 g764210 ( .a(n_16772), .b(n_16385), .o(n_16930) );
in01s01 g764211 ( .a(n_16818), .o(n_16819) );
ao12s01 g764212 ( .a(n_15834), .b(n_16741), .c(n_15778), .o(n_16818) );
in01s01 g764213 ( .a(n_16816), .o(n_16817) );
ao12s01 g764214 ( .a(n_15928), .b(n_16798), .c(n_15922), .o(n_16816) );
in01s02 g764215 ( .a(n_16602), .o(n_16579) );
no02s01 TIMEBOOST_cell_1396 ( .a(TIMEBOOST_net_312), .b(n_29708), .o(n_29742) );
in01m04 g764217 ( .a(n_16474), .o(n_16468) );
na02s02 g764220 ( .a(n_16462), .b(n_16436), .o(n_16527) );
in01m02 g764221 ( .a(n_16601), .o(n_16578) );
na02f08 TIMEBOOST_cell_1294 ( .a(TIMEBOOST_net_261), .b(FE_OCP_RBN7023_n_18650), .o(n_18829) );
in01s01 g764224 ( .a(n_16552), .o(n_16576) );
in01m02 g764225 ( .a(n_16526), .o(n_16552) );
na02f06 g764227 ( .a(n_16460), .b(n_16485), .o(n_16582) );
oa22s01 g764228 ( .a(n_16742), .b(n_16253), .c(n_16743), .d(n_16254), .o(n_16815) );
oa22s01 g764229 ( .a(n_16741), .b(n_15872), .c(n_16768), .d(n_15871), .o(n_16847) );
oa22s01 g764230 ( .a(n_16798), .b(n_15959), .c(n_16770), .d(n_15960), .o(n_16846) );
oa22s01 g764231 ( .a(n_16575), .b(n_17584), .c(n_16551), .d(FE_OCP_RBN3196_n_15599), .o(n_16619) );
in01s01 g764232 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_11_), .o(n_17995) );
in01m01 g764237 ( .a(n_16516), .o(n_16580) );
no02m04 g764238 ( .a(n_16493), .b(FE_OCPN6285_FE_OCP_RBN1602_n_14638), .o(n_16516) );
in01s01 g764240 ( .a(n_16515), .o(n_16524) );
na02s06 g764241 ( .a(FE_OCPN6285_FE_OCP_RBN1602_n_14638), .b(n_16493), .o(n_16515) );
no02s06 g764242 ( .a(n_16376), .b(n_16405), .o(n_16445) );
in01f02 g764243 ( .a(n_16443), .o(n_16444) );
no02f04 g764244 ( .a(n_16296), .b(n_16336), .o(n_16443) );
na02f04 TIMEBOOST_cell_6312 ( .a(n_36457), .b(TIMEBOOST_net_2007), .o(TIMEBOOST_net_1710) );
in01s02 g764247 ( .a(n_16464), .o(n_16465) );
na02s04 g764248 ( .a(n_16377), .b(n_16441), .o(n_16464) );
na02m06 g764249 ( .a(n_16295), .b(n_47268), .o(n_16735) );
no02m06 g764250 ( .a(n_16293), .b(n_46426), .o(n_16716) );
in01m04 g764251 ( .a(n_16490), .o(n_16491) );
na02f08 g764252 ( .a(FE_OCP_RBN6868_n_16392), .b(FE_OCP_RBN4401_n_16321), .o(n_16490) );
na02s03 g764253 ( .a(n_16402), .b(n_16374), .o(n_16440) );
no02f02 g764254 ( .a(n_16376), .b(n_16375), .o(n_16463) );
na02m02 g764255 ( .a(n_16458), .b(n_16429), .o(n_16489) );
no02m02 g764256 ( .a(n_16431), .b(FE_OCP_RBN4409_n_16429), .o(n_16514) );
na02m04 g764258 ( .a(n_16722), .b(n_16263), .o(n_16824) );
na02s01 g764259 ( .a(n_16723), .b(n_16384), .o(n_16772) );
no02s02 TIMEBOOST_cell_5563 ( .a(TIMEBOOST_net_1729), .b(n_22098), .o(n_22233) );
na02s02 g764261 ( .a(n_16424), .b(n_16364), .o(n_16462) );
no02s01 g764263 ( .a(n_16438), .b(n_16461), .o(n_16486) );
no02f04 g764264 ( .a(n_16438), .b(n_16272), .o(n_16439) );
na02f06 g764265 ( .a(n_16394), .b(n_16436), .o(n_16437) );
na02s03 g764266 ( .a(n_16432), .b(FE_OCP_RBN6867_n_16392), .o(n_16460) );
na02m02 g764267 ( .a(n_16452), .b(n_16455), .o(n_16513) );
na02f08 TIMEBOOST_cell_1293 ( .a(n_18718), .b(n_18554), .o(TIMEBOOST_net_261) );
na02f02 g764269 ( .a(n_16433), .b(n_16392), .o(n_16485) );
no02s01 TIMEBOOST_cell_1395 ( .a(n_44045), .b(n_28922), .o(TIMEBOOST_net_312) );
in01f02 g764271 ( .a(n_16434), .o(n_16435) );
in01f02 g764272 ( .a(n_16407), .o(n_16434) );
no02f06 g764273 ( .a(n_16290), .b(n_16237), .o(n_16407) );
na02s01 TIMEBOOST_cell_1128 ( .a(TIMEBOOST_net_178), .b(n_33275), .o(n_33346) );
in01m02 g764275 ( .a(n_47340), .o(n_16484) );
oa22s01 g764277 ( .a(n_16675), .b(n_16303), .c(n_16676), .d(n_16302), .o(n_16744) );
na02s01 TIMEBOOST_cell_1127 ( .a(n_33276), .b(n_32895), .o(TIMEBOOST_net_178) );
no02f04 g764280 ( .a(n_16234), .b(n_16207), .o(n_16337) );
in01s02 g764281 ( .a(n_16405), .o(n_16406) );
na02s06 g764282 ( .a(n_16286), .b(n_16221), .o(n_16405) );
no02m04 g764283 ( .a(n_16321), .b(n_16273), .o(n_16379) );
in01s01 g764284 ( .a(n_16446), .o(n_16404) );
no02m02 g764285 ( .a(n_16230), .b(n_14588), .o(n_16296) );
no02s03 g764286 ( .a(n_16230), .b(FE_OCPN1733_n_14524), .o(n_16446) );
no02f04 g764287 ( .a(FE_OCP_RBN4391_n_16230), .b(n_14618), .o(n_16336) );
na02s03 TIMEBOOST_cell_4521 ( .a(n_39844), .b(n_39816), .o(TIMEBOOST_net_1351) );
na02s06 g764289 ( .a(n_16333), .b(FE_OCPN1705_n_14730), .o(n_16442) );
na02s02 TIMEBOOST_cell_5401 ( .a(TIMEBOOST_net_1648), .b(n_43128), .o(n_43282) );
no02s06 g764292 ( .a(n_16330), .b(n_14588), .o(n_16332) );
na02s04 g764293 ( .a(n_16278), .b(FE_OCPN1705_n_14730), .o(n_16377) );
na02s06 g764294 ( .a(n_16330), .b(n_14588), .o(n_16441) );
in01m02 g764295 ( .a(n_46426), .o(n_16295) );
in01m02 g764298 ( .a(n_47268), .o(n_16293) );
in01s01 g764302 ( .a(n_16376), .o(n_16402) );
no02s03 g764303 ( .a(n_16328), .b(n_14588), .o(n_16376) );
in01m02 g764304 ( .a(n_16432), .o(n_16433) );
na02f04 g764305 ( .a(n_16401), .b(FE_OCP_RBN4401_n_16321), .o(n_16432) );
in01m01 g764306 ( .a(n_16374), .o(n_16375) );
no02s01 TIMEBOOST_cell_6985 ( .a(n_4528), .b(n_3641), .o(TIMEBOOST_net_2251) );
na02f01 g764308 ( .a(n_16328), .b(n_14805), .o(n_16374) );
in01s01 g764310 ( .a(n_16431), .o(n_16458) );
no02m08 g764311 ( .a(n_16398), .b(n_14588), .o(n_16431) );
na02s06 g764313 ( .a(n_16398), .b(n_14805), .o(n_16399) );
na02s02 g764314 ( .a(n_16398), .b(n_14805), .o(n_16429) );
in01f04 g764317 ( .a(n_16397), .o(n_16396) );
na02f08 g764318 ( .a(n_16283), .b(n_16373), .o(n_16397) );
in01s01 g764320 ( .a(n_16798), .o(n_16770) );
na02s01 g764321 ( .a(n_16678), .b(n_16103), .o(n_16798) );
in01s01 g764322 ( .a(n_16722), .o(n_16723) );
na02m04 g764323 ( .a(n_15973), .b(n_16677), .o(n_16722) );
no02f02 g764324 ( .a(n_16319), .b(FE_OCP_RBN2905_n_14590), .o(n_16438) );
na02f02 g764326 ( .a(n_16322), .b(n_16274), .o(n_16372) );
no02f06 g764327 ( .a(n_16418), .b(n_16422), .o(n_16426) );
oa12m04 g764329 ( .a(n_16206), .b(n_16234), .c(n_16233), .o(n_16291) );
no02m08 TIMEBOOST_cell_1126 ( .a(TIMEBOOST_net_177), .b(n_40942), .o(n_40979) );
na02m04 g764332 ( .a(n_16289), .b(n_16363), .o(n_16493) );
in01s01 g764334 ( .a(n_16742), .o(n_16743) );
oa12s01 g764335 ( .a(n_16018), .b(n_16673), .c(n_15967), .o(n_16742) );
in01s01 g764337 ( .a(n_16741), .o(n_16768) );
oa12s01 g764338 ( .a(n_15930), .b(n_16673), .c(n_16059), .o(n_16741) );
oa12s01 g764339 ( .a(n_16367), .b(n_16366), .c(n_16365), .o(n_16425) );
in01s01 g764341 ( .a(n_16424), .o(n_16456) );
in01s01 g764342 ( .a(n_16394), .o(n_16424) );
oa12f06 g764343 ( .a(n_16181), .b(n_16366), .c(n_16271), .o(n_16394) );
in01s02 g764344 ( .a(n_16575), .o(n_16551) );
no02m02 TIMEBOOST_cell_1288 ( .a(n_18602), .b(TIMEBOOST_net_258), .o(n_18683) );
in01m01 g764346 ( .a(n_16454), .o(n_16455) );
oa22m01 g764347 ( .a(n_16317), .b(n_14598), .c(n_16423), .d(FE_OCPN1324_n_14577), .o(n_16454) );
in01s01 g764348 ( .a(n_16452), .o(n_16453) );
oa12s01 g764349 ( .a(n_16314), .b(n_16361), .c(n_16422), .o(n_16452) );
in01m04 g764353 ( .a(n_16371), .o(n_16392) );
ao12f08 g764354 ( .a(n_16203), .b(n_16288), .c(n_16224), .o(n_16371) );
oa22s01 g764355 ( .a(n_16653), .b(n_16060), .c(n_16673), .d(n_16061), .o(n_16767) );
no02f06 g764356 ( .a(n_16418), .b(n_16318), .o(n_16419) );
in01s01 g764357 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_11_), .o(n_18055) );
no03m08 TIMEBOOST_cell_1125 ( .a(n_40941), .b(n_40963), .c(n_40824), .o(TIMEBOOST_net_177) );
na02s02 g764361 ( .a(n_16288), .b(n_16157), .o(n_16289) );
na02f04 g764362 ( .a(n_16206), .b(n_16205), .o(n_16207) );
no02m04 g764363 ( .a(n_16236), .b(n_16233), .o(n_16204) );
na02s04 g764364 ( .a(n_16200), .b(n_16226), .o(n_16287) );
no02s04 g764365 ( .a(n_16201), .b(n_16168), .o(n_16324) );
in01s02 g764366 ( .a(n_16369), .o(n_16370) );
na02m04 g764367 ( .a(n_16225), .b(n_46421), .o(n_16369) );
no02f02 g764369 ( .a(n_16288), .b(n_16188), .o(n_16322) );
na02s04 g764370 ( .a(n_16285), .b(n_14730), .o(n_16286) );
na02f04 g764371 ( .a(n_16285), .b(FE_OCPN1705_n_14730), .o(n_16401) );
in01m02 g764372 ( .a(n_16390), .o(n_16391) );
na02m04 g764373 ( .a(n_16219), .b(n_16368), .o(n_16390) );
no02m06 g764374 ( .a(n_16231), .b(FE_OCPN1705_n_14730), .o(n_16232) );
na02f06 g764375 ( .a(n_16190), .b(n_14805), .o(n_16283) );
na02m08 g764376 ( .a(n_16231), .b(FE_OCPN1705_n_14730), .o(n_16373) );
no02f08 g764378 ( .a(n_16285), .b(n_14730), .o(n_16321) );
na02s01 g764379 ( .a(n_16366), .b(n_16365), .o(n_16367) );
in01s01 g764380 ( .a(n_16388), .o(n_16389) );
na02s01 g764381 ( .a(n_16364), .b(n_16436), .o(n_16388) );
no02f08 g764382 ( .a(n_16316), .b(n_16266), .o(n_16418) );
na02s01 g764383 ( .a(n_16417), .b(n_16361), .o(n_16482) );
no02s02 TIMEBOOST_cell_1287 ( .a(n_18263), .b(n_18316), .o(TIMEBOOST_net_258) );
in01s01 g764385 ( .a(n_16677), .o(n_16678) );
no02m04 g764386 ( .a(n_16632), .b(n_16062), .o(n_16677) );
in01s01 g764387 ( .a(n_16675), .o(n_16676) );
ao12s02 g764388 ( .a(n_15866), .b(n_16615), .c(n_15925), .o(n_16675) );
no02f02 g764390 ( .a(n_16193), .b(n_16161), .o(n_16319) );
na02s01 TIMEBOOST_cell_4485 ( .a(n_5584), .b(n_5583), .o(TIMEBOOST_net_1333) );
in01f02 g764395 ( .a(n_16333), .o(n_16279) );
in01s02 g764397 ( .a(n_16330), .o(n_16278) );
na02f04 TIMEBOOST_cell_4520 ( .a(TIMEBOOST_net_1350), .b(n_11295), .o(n_11356) );
na02s08 TIMEBOOST_cell_904 ( .a(n_206), .b(TIMEBOOST_net_66), .o(n_207) );
na02m02 g764400 ( .a(n_16277), .b(n_16194), .o(n_16363) );
no02s10 TIMEBOOST_cell_972 ( .a(TIMEBOOST_net_100), .b(n_17698), .o(n_17954) );
na02f06 TIMEBOOST_cell_1060 ( .a(TIMEBOOST_net_144), .b(FE_RN_1018_0), .o(n_23270) );
no02s01 TIMEBOOST_cell_6383 ( .a(n_23339), .b(n_23317), .o(TIMEBOOST_net_2043) );
in01s01 g764406 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_), .o(n_16618) );
in01s01 g764409 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_10_), .o(n_16617) );
in01m02 g764412 ( .a(n_16234), .o(n_16228) );
na02f08 g764413 ( .a(n_16172), .b(n_16171), .o(n_16234) );
na02f08 g764414 ( .a(n_16202), .b(n_16157), .o(n_16203) );
na02f04 g764416 ( .a(n_16095), .b(n_14618), .o(n_16205) );
no02f06 g764417 ( .a(n_16095), .b(n_14420), .o(n_16236) );
in01s02 g764419 ( .a(n_16200), .o(n_16201) );
na02f04 g764420 ( .a(n_16169), .b(n_14420), .o(n_16170) );
na02s04 g764421 ( .a(n_16169), .b(FE_OCP_DRV_N3514_n_14650), .o(n_16200) );
in01s02 g764423 ( .a(n_16168), .o(n_16226) );
no02s04 g764424 ( .a(n_16169), .b(n_14420), .o(n_16168) );
no02f04 g764425 ( .a(n_16169), .b(FE_OCP_DRV_N3514_n_14650), .o(n_16166) );
no02m04 TIMEBOOST_cell_4484 ( .a(TIMEBOOST_net_1332), .b(n_5555), .o(TIMEBOOST_net_1156) );
no02s04 g764427 ( .a(n_16053), .b(n_14419), .o(n_16094) );
na02m04 g764429 ( .a(n_16151), .b(FE_OCPN1705_n_14730), .o(n_16225) );
na02s02 TIMEBOOST_cell_4517 ( .a(n_10892), .b(n_10747), .o(TIMEBOOST_net_1349) );
no02s01 TIMEBOOST_cell_8473 ( .a(TIMEBOOST_net_2723), .b(n_7515), .o(TIMEBOOST_net_255) );
no02m04 TIMEBOOST_cell_6257 ( .a(TIMEBOOST_net_1669), .b(n_5813), .o(TIMEBOOST_net_1980) );
na02s01 TIMEBOOST_cell_903 ( .a(beta_31), .b(beta_11), .o(TIMEBOOST_net_66) );
no02s04 g764438 ( .a(n_16084), .b(n_14524), .o(n_16125) );
na02m02 g764439 ( .a(n_16159), .b(n_16157), .o(n_16277) );
na02f02 g764441 ( .a(n_16224), .b(n_16202), .o(n_16274) );
in01m03 g764442 ( .a(n_16273), .o(n_16368) );
no02m06 g764443 ( .a(n_16220), .b(n_14730), .o(n_16273) );
na02f06 TIMEBOOST_cell_1059 ( .a(FE_RN_1019_0), .b(n_23196), .o(TIMEBOOST_net_144) );
no02f08 g764445 ( .a(n_16158), .b(n_16194), .o(n_16288) );
no02m08 g764446 ( .a(FE_OCP_RBN4394_n_16146), .b(FE_OCPN1705_n_14730), .o(n_16223) );
na02s04 g764447 ( .a(n_16220), .b(n_14730), .o(n_16221) );
na02s02 g764448 ( .a(n_16220), .b(FE_OCPN1705_n_14730), .o(n_16219) );
no02s08 TIMEBOOST_cell_3297 ( .a(TIMEBOOST_net_939), .b(n_10620), .o(n_10711) );
no02s03 TIMEBOOST_cell_971 ( .a(n_17758), .b(n_17825), .o(TIMEBOOST_net_100) );
no02f08 TIMEBOOST_cell_3179 ( .a(n_25734), .b(TIMEBOOST_net_880), .o(n_25816) );
in01s01 g764452 ( .a(n_16272), .o(n_16364) );
na02s06 TIMEBOOST_cell_1118 ( .a(TIMEBOOST_net_173), .b(n_17954), .o(n_18061) );
no02m02 g764455 ( .a(n_16124), .b(n_45331), .o(n_16193) );
in01s01 g764456 ( .a(n_16416), .o(n_16417) );
no02s01 g764457 ( .a(n_16422), .b(n_16266), .o(n_16416) );
no02s01 g764458 ( .a(n_16084), .b(FE_OCP_RBN3220_n_15992), .o(n_16192) );
na02f04 g764459 ( .a(n_16267), .b(FE_OCP_RBN2082_n_14554), .o(n_16318) );
in01s01 g764463 ( .a(n_16653), .o(n_16673) );
in01s01 g764465 ( .a(n_16632), .o(n_16653) );
no02s01 TIMEBOOST_cell_4860 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_36540), .o(TIMEBOOST_net_1378) );
no02f08 g764467 ( .a(n_16155), .b(n_16112), .o(n_16366) );
in01m01 g764468 ( .a(n_16423), .o(n_16317) );
na02f04 g764469 ( .a(n_16160), .b(n_16189), .o(n_16423) );
oa12s01 g764470 ( .a(n_16270), .b(n_16269), .c(n_16268), .o(n_16362) );
in01s01 g764472 ( .a(n_16361), .o(n_16386) );
in01s01 g764473 ( .a(n_16316), .o(n_16361) );
ao12f06 g764474 ( .a(n_16180), .b(n_16179), .c(n_16107), .o(n_16316) );
na02f08 g764475 ( .a(n_16119), .b(n_16090), .o(n_16285) );
in01m02 g764476 ( .a(n_16231), .o(n_16190) );
na04s01 TIMEBOOST_cell_8394 ( .a(n_5174), .b(n_6051), .c(n_5175), .d(n_6052), .o(n_6159) );
oa12s01 g764478 ( .a(n_16574), .b(n_16573), .c(n_16572), .o(n_16616) );
na02s01 TIMEBOOST_cell_5411 ( .a(TIMEBOOST_net_1653), .b(FE_OCP_RBN6191_n_43103), .o(n_43605) );
na02m02 g764481 ( .a(n_16113), .b(n_16037), .o(n_16160) );
na02f02 g764482 ( .a(FE_OCP_RBN3256_n_16113), .b(n_16036), .o(n_16189) );
in01s02 g764483 ( .a(n_16123), .o(n_16124) );
no02f04 g764484 ( .a(n_16010), .b(n_15954), .o(n_16123) );
na02f08 g764485 ( .a(n_45332), .b(n_16008), .o(n_16171) );
in01s01 g764486 ( .a(n_16158), .o(n_16159) );
no02m08 g764487 ( .a(n_16122), .b(FE_OCPN1733_n_14524), .o(n_16158) );
in01s02 g764489 ( .a(n_16157), .o(n_16188) );
na02m08 g764490 ( .a(n_16122), .b(FE_OCPN1733_n_14524), .o(n_16157) );
na02f08 g764491 ( .a(n_16075), .b(n_14618), .o(n_16224) );
na02f04 g764492 ( .a(n_16074), .b(FE_OCPN1733_n_14524), .o(n_16202) );
na02f08 g764493 ( .a(FE_OCP_RBN6070_n_16041), .b(FE_OCP_DRV_N3514_n_14650), .o(n_16119) );
no02s02 TIMEBOOST_cell_7615 ( .a(TIMEBOOST_net_2438), .b(n_19417), .o(n_20265) );
na02s03 g764495 ( .a(n_16003), .b(n_14730), .o(n_16056) );
na02m04 g764496 ( .a(n_16041), .b(n_14524), .o(n_16090) );
na02s01 g764497 ( .a(n_16573), .b(n_16572), .o(n_16574) );
in01s01 g764499 ( .a(n_16615), .o(n_16630) );
no02s01 g764500 ( .a(n_16542), .b(n_15878), .o(n_16615) );
no02s01 g764501 ( .a(n_16182), .b(n_16271), .o(n_16365) );
na02s01 g764502 ( .a(n_16269), .b(n_16268), .o(n_16270) );
in01s04 g764503 ( .a(n_16267), .o(n_16422) );
na02m06 g764504 ( .a(n_16216), .b(FE_OCP_RBN2814_n_14441), .o(n_16267) );
in01s01 g764506 ( .a(n_16266), .o(n_16314) );
no02m06 g764507 ( .a(n_16216), .b(FE_OCP_RBN2814_n_14441), .o(n_16266) );
na02s01 TIMEBOOST_cell_7846 ( .a(TIMEBOOST_net_1311), .b(FE_OCP_RBN3052_n_10100), .o(TIMEBOOST_net_2554) );
ao12f06 g764509 ( .a(n_46980), .b(n_16154), .c(FE_OCPN5126_n_16111), .o(n_16155) );
no02s02 TIMEBOOST_cell_1120 ( .a(TIMEBOOST_net_174), .b(FE_OCP_RBN2505_n_33226), .o(n_33394) );
na02f08 g764513 ( .a(n_15918), .b(n_15860), .o(n_16095) );
no02s06 TIMEBOOST_cell_4513 ( .a(n_39969), .b(FE_OCP_RBN6853_n_39793), .o(TIMEBOOST_net_1347) );
in01s01 g764517 ( .a(n_16089), .o(n_16118) );
in01s01 g764518 ( .a(n_16053), .o(n_16089) );
in01f02 g764519 ( .a(n_16053), .o(n_16052) );
in01s02 g764521 ( .a(n_16197), .o(n_16151) );
no02m08 g764522 ( .a(n_16046), .b(n_16004), .o(n_16197) );
na02f08 g764538 ( .a(n_16049), .b(n_16047), .o(n_16194) );
na02s02 TIMEBOOST_cell_8704 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_11_), .b(FE_OCP_RBN6540_n_44083), .o(TIMEBOOST_net_2839) );
oa12s01 g764551 ( .a(n_16110), .b(n_16154), .c(n_16109), .o(n_16183) );
oa12s01 g764552 ( .a(n_16507), .b(n_16506), .c(n_16505), .o(n_16550) );
oa12s01 g764553 ( .a(n_16548), .b(n_16547), .c(n_16546), .o(n_16593) );
oa12s01 g764554 ( .a(n_16545), .b(n_16544), .c(n_16543), .o(n_16592) );
oa12s01 g764555 ( .a(n_16510), .b(n_16509), .c(n_16508), .o(n_16549) );
in01s01 g764556 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_9_), .o(n_17886) );
in01s02 g764558 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_8_), .o(n_16591) );
na02f08 g764560 ( .a(n_16001), .b(n_16048), .o(n_16049) );
no02m10 TIMEBOOST_cell_1144 ( .a(n_37412), .b(TIMEBOOST_net_186), .o(n_37515) );
na03s08 TIMEBOOST_cell_1117 ( .a(n_17930), .b(n_17893), .c(n_18002), .o(TIMEBOOST_net_173) );
no02f04 g764564 ( .a(n_16007), .b(n_14524), .o(n_16010) );
na02s04 TIMEBOOST_cell_6886 ( .a(TIMEBOOST_net_2201), .b(n_18113), .o(TIMEBOOST_net_1426) );
no02f02 g764566 ( .a(n_15915), .b(n_14419), .o(n_15954) );
na02s06 g764567 ( .a(n_16007), .b(n_14452), .o(n_16008) );
na02f06 g764568 ( .a(FE_OCP_RBN3109_n_15817), .b(n_14650), .o(n_15918) );
na02s04 g764569 ( .a(n_15817), .b(n_14588), .o(n_15860) );
na02m04 g764570 ( .a(n_15911), .b(n_14419), .o(n_15953) );
no02f06 TIMEBOOST_cell_4512 ( .a(TIMEBOOST_net_1346), .b(n_39719), .o(n_39733) );
no02s06 g764572 ( .a(n_15948), .b(FE_OCPN1733_n_14524), .o(n_16004) );
no02m08 g764573 ( .a(n_15993), .b(FE_OCP_DRV_N3514_n_14650), .o(n_16046) );
na02m02 TIMEBOOST_cell_4556 ( .a(TIMEBOOST_net_1368), .b(n_17350), .o(FE_RN_341_0) );
na02s03 g764577 ( .a(n_15992), .b(FE_OCP_DRV_N3514_n_14650), .o(n_16044) );
na02s01 g764578 ( .a(n_16509), .b(n_16508), .o(n_16510) );
na02s01 g764579 ( .a(n_16547), .b(n_16546), .o(n_16548) );
na02s01 g764580 ( .a(n_16506), .b(n_16505), .o(n_16507) );
na02s01 g764581 ( .a(n_16544), .b(n_16543), .o(n_16545) );
no02s06 g764582 ( .a(n_16154), .b(FE_OCPN5126_n_16111), .o(n_16112) );
in01s01 g764583 ( .a(n_16181), .o(n_16182) );
na02s06 g764584 ( .a(n_16144), .b(FE_OCPN4929_n_16143), .o(n_16181) );
no02s06 g764585 ( .a(n_16144), .b(FE_OCPN4929_n_16143), .o(n_16271) );
no02f04 g764586 ( .a(n_15998), .b(n_15985), .o(n_16077) );
no02s01 TIMEBOOST_cell_1119 ( .a(n_33317), .b(n_33316), .o(TIMEBOOST_net_174) );
na02s01 g764588 ( .a(n_16109), .b(n_16154), .o(n_16110) );
no02s01 g764589 ( .a(n_16180), .b(n_16108), .o(n_16268) );
no02s01 g764590 ( .a(FE_OCP_RBN3111_n_15817), .b(FE_OCP_RBN3075_n_15706), .o(n_16866) );
in01s01 g764591 ( .a(n_16541), .o(n_16542) );
na02m04 g764592 ( .a(n_16504), .b(n_15877), .o(n_16541) );
ao12s01 g764593 ( .a(n_16025), .b(n_16448), .c(n_15821), .o(n_16573) );
in01m02 g764594 ( .a(n_16074), .o(n_16075) );
in01s01 g764596 ( .a(FE_OCP_RBN3234_n_16041), .o(n_17139) );
in01m02 g764601 ( .a(n_16003), .o(n_16038) );
oa22f02 g764603 ( .a(n_15802), .b(n_15567), .c(n_15803), .d(n_15568), .o(n_16003) );
oa12s01 g764604 ( .a(n_16141), .b(n_16142), .c(n_16140), .o(n_16212) );
in01s01 g764605 ( .a(n_16179), .o(n_16269) );
oa12f06 g764606 ( .a(n_15980), .b(n_16142), .c(n_16067), .o(n_16179) );
no02s01 TIMEBOOST_cell_1152 ( .a(TIMEBOOST_net_190), .b(n_41171), .o(n_41231) );
na02m08 TIMEBOOST_cell_3220 ( .a(n_20767), .b(n_20464), .o(TIMEBOOST_net_901) );
in01s01 g764609 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_9_), .o(n_17931) );
in01s01 g764611 ( .a(n_16036), .o(n_16037) );
no02m01 g764612 ( .a(n_16001), .b(n_15946), .o(n_16036) );
no02s01 TIMEBOOST_cell_1151 ( .a(n_40908), .b(n_40944), .o(TIMEBOOST_net_190) );
no02m04 g764614 ( .a(n_15988), .b(n_15893), .o(n_16072) );
na02m02 g764615 ( .a(FE_OCP_RBN3125_n_15856), .b(n_15999), .o(n_16000) );
no02m02 g764616 ( .a(n_16080), .b(n_15856), .o(n_15998) );
no02s10 TIMEBOOST_cell_1143 ( .a(FE_RN_185_0), .b(n_36998), .o(TIMEBOOST_net_186) );
no02m08 TIMEBOOST_cell_4551 ( .a(n_16953), .b(n_17045), .o(TIMEBOOST_net_1366) );
na02f08 g764621 ( .a(n_15951), .b(n_14588), .o(n_16048) );
na02f06 TIMEBOOST_cell_3219 ( .a(n_1238), .b(TIMEBOOST_net_900), .o(n_1248) );
no02s04 g764623 ( .a(n_15861), .b(n_14588), .o(n_15917) );
in01s01 g764624 ( .a(n_16504), .o(n_16544) );
na02m04 g764625 ( .a(n_16447), .b(n_16024), .o(n_16504) );
in01s04 g764626 ( .a(n_15818), .o(n_15819) );
oa12s06 g764627 ( .a(n_15639), .b(n_15810), .c(n_15661), .o(n_15818) );
no02s01 g764628 ( .a(n_15983), .b(n_15762), .o(n_15995) );
no02s01 g764629 ( .a(n_15901), .b(n_15708), .o(n_15949) );
na02s01 g764630 ( .a(n_16142), .b(n_16140), .o(n_16141) );
no02m04 g764631 ( .a(n_16071), .b(n_16070), .o(n_16180) );
in01s01 g764632 ( .a(n_16107), .o(n_16108) );
na02f04 g764633 ( .a(n_16071), .b(n_16070), .o(n_16107) );
ao12s01 g764634 ( .a(n_15787), .b(n_16450), .c(n_15783), .o(n_16509) );
no02s01 g764635 ( .a(n_16449), .b(n_15883), .o(n_16547) );
ao12s01 g764636 ( .a(n_15932), .b(n_16450), .c(n_15881), .o(n_16506) );
no02f08 g764637 ( .a(n_15945), .b(n_15937), .o(n_16154) );
ao12s01 g764638 ( .a(n_15944), .b(n_46980), .c(FE_OCPN5126_n_16111), .o(n_16109) );
in01m06 g764640 ( .a(n_15915), .o(n_16007) );
na02f06 TIMEBOOST_cell_5372 ( .a(n_26010), .b(n_23353), .o(TIMEBOOST_net_1634) );
in01s01 g764644 ( .a(FE_OCP_RBN3111_n_15817), .o(n_15912) );
na02s01 TIMEBOOST_cell_3897 ( .a(n_18852), .b(n_18481), .o(TIMEBOOST_net_1039) );
oa12f04 g764651 ( .a(FE_OCP_RBN3016_n_15300), .b(FE_OCP_RBN6006_n_15704), .c(n_15771), .o(n_15815) );
no02s01 TIMEBOOST_cell_894 ( .a(TIMEBOOST_net_61), .b(n_17736), .o(n_17819) );
in01m04 g764654 ( .a(n_15948), .o(n_15993) );
no02s06 TIMEBOOST_cell_896 ( .a(TIMEBOOST_net_62), .b(n_32643), .o(FE_RN_2002_0) );
in01s04 g764657 ( .a(n_15908), .o(n_15909) );
oa12s02 g764659 ( .a(n_15578), .b(FE_OCP_RBN3102_n_15768), .c(n_15810), .o(n_15857) );
na02m04 TIMEBOOST_cell_7567 ( .a(TIMEBOOST_net_2414), .b(FE_RN_860_0), .o(TIMEBOOST_net_1471) );
na02m04 TIMEBOOST_cell_6002 ( .a(TIMEBOOST_net_1852), .b(n_18089), .o(n_18163) );
oa12m04 g764666 ( .a(n_15373), .b(n_15808), .c(n_15806), .o(n_15820) );
na02f08 TIMEBOOST_cell_8569 ( .a(TIMEBOOST_net_2771), .b(n_14943), .o(n_15047) );
in01s04 g764668 ( .a(n_15989), .o(n_15990) );
no02s06 g764669 ( .a(n_15854), .b(n_15455), .o(n_15989) );
oa12s01 g764670 ( .a(n_16032), .b(n_16031), .c(n_16030), .o(n_16106) );
oa12s01 g764671 ( .a(n_16481), .b(n_16480), .c(n_16479), .o(n_16523) );
no02f06 g764674 ( .a(n_15845), .b(n_15905), .o(n_16001) );
no02f08 g764677 ( .a(n_15765), .b(n_14650), .o(n_15856) );
na02s04 TIMEBOOST_cell_5371 ( .a(TIMEBOOST_net_1633), .b(n_46957), .o(TIMEBOOST_net_1312) );
na02m04 g764679 ( .a(n_15706), .b(n_14524), .o(n_15743) );
in01m02 g764680 ( .a(n_15987), .o(n_15988) );
no02m02 g764681 ( .a(n_15946), .b(n_15905), .o(n_15987) );
no02m08 g764682 ( .a(n_15797), .b(n_14452), .o(n_16080) );
na02m02 g764683 ( .a(n_15765), .b(n_14419), .o(n_15999) );
na02s01 g764684 ( .a(n_16480), .b(n_16479), .o(n_16481) );
no02f06 g764685 ( .a(n_16030), .b(n_15938), .o(n_15945) );
no02s01 g764686 ( .a(n_46980), .b(FE_OCPN5126_n_16111), .o(n_15944) );
na02m04 g764687 ( .a(n_15895), .b(n_15736), .o(n_15943) );
na02s02 TIMEBOOST_cell_6968 ( .a(TIMEBOOST_net_2242), .b(n_8404), .o(n_10214) );
in01s01 TIMEBOOST_cell_7379 ( .a(TIMEBOOST_net_2315), .o(TIMEBOOST_net_2314) );
no02s02 TIMEBOOST_cell_3896 ( .a(TIMEBOOST_net_1038), .b(TIMEBOOST_net_242), .o(n_38698) );
no02s01 TIMEBOOST_cell_893 ( .a(n_17713), .b(n_17305), .o(TIMEBOOST_net_61) );
no03s08 TIMEBOOST_cell_895 ( .a(FE_OCP_RBN6520_n_32706), .b(n_32704), .c(FE_OCP_RBN5518_n_32436), .o(TIMEBOOST_net_62) );
no02s04 g764693 ( .a(n_15768), .b(n_15523), .o(n_15770) );
no02f04 TIMEBOOST_cell_6180 ( .a(TIMEBOOST_net_1941), .b(n_10480), .o(TIMEBOOST_net_1610) );
no02s01 g764695 ( .a(n_15981), .b(n_16067), .o(n_16140) );
na02s02 g764696 ( .a(n_15808), .b(n_15375), .o(n_15809) );
na03s04 TIMEBOOST_cell_5713 ( .a(n_12445), .b(n_12364), .c(n_12363), .o(TIMEBOOST_net_1198) );
no02s02 TIMEBOOST_cell_7068 ( .a(TIMEBOOST_net_2292), .b(n_11589), .o(n_11741) );
no02s06 g764699 ( .a(n_15853), .b(n_15404), .o(n_15854) );
na02s01 g764700 ( .a(n_16031), .b(n_16030), .o(n_16032) );
no02s01 g764701 ( .a(n_16415), .b(n_15882), .o(n_16449) );
in01s01 g764702 ( .a(n_16447), .o(n_16448) );
na02m04 g764703 ( .a(n_15838), .b(n_16450), .o(n_16447) );
in01s02 g764704 ( .a(n_15984), .o(n_15985) );
in01s02 g764705 ( .a(n_15942), .o(n_15984) );
no02f08 g764706 ( .a(n_15801), .b(n_15799), .o(n_15942) );
in01s01 g764708 ( .a(n_15901), .o(n_15983) );
in01s01 g764711 ( .a(n_15861), .o(n_15901) );
in01f02 g764712 ( .a(n_15861), .o(n_15862) );
in01s01 g764715 ( .a(FE_OCP_RBN3204_n_15900), .o(n_15939) );
oa12s02 g764718 ( .a(n_15258), .b(n_15804), .c(n_15180), .o(n_15805) );
ao12s06 g764719 ( .a(n_15178), .b(FE_OCP_RBN3154_n_15804), .c(n_15218), .o(n_15852) );
in01m01 g764720 ( .a(n_15802), .o(n_15803) );
oa12f01 g764721 ( .a(n_15604), .b(n_15739), .c(n_15487), .o(n_15802) );
ao12f06 g764722 ( .a(n_15843), .b(n_16029), .c(n_15934), .o(n_16142) );
no02s02 TIMEBOOST_cell_7034 ( .a(TIMEBOOST_net_2275), .b(n_4459), .o(TIMEBOOST_net_1307) );
oa12s01 g764724 ( .a(n_16028), .b(n_16029), .c(n_16027), .o(n_16105) );
in01m01 g764725 ( .a(n_15951), .o(n_15898) );
no02f08 g764726 ( .a(n_15741), .b(n_15767), .o(n_15951) );
no02s01 TIMEBOOST_cell_5130 ( .a(FE_OCP_RBN6671_n_34297), .b(FE_OCP_RBN4920_n_33691), .o(TIMEBOOST_net_1513) );
na02f04 g764730 ( .a(n_15795), .b(FE_OCP_RBN3217_n_15758), .o(n_15850) );
na02f04 TIMEBOOST_cell_4538 ( .a(TIMEBOOST_net_1359), .b(n_11291), .o(n_11369) );
na02f06 g764732 ( .a(n_15701), .b(n_15800), .o(n_15801) );
in01s02 g764733 ( .a(n_15895), .o(n_15896) );
no02f02 TIMEBOOST_cell_3196 ( .a(n_9807), .b(n_9750), .o(TIMEBOOST_net_889) );
na02s01 TIMEBOOST_cell_1016 ( .a(TIMEBOOST_net_122), .b(n_37291), .o(n_37289) );
no02f06 g764736 ( .a(FE_OCP_RBN4377_n_15700), .b(n_14419), .o(n_15767) );
no02f04 g764737 ( .a(n_15847), .b(n_14524), .o(n_15849) );
no02m02 g764738 ( .a(n_15847), .b(n_14588), .o(n_15946) );
no02s04 g764739 ( .a(n_15761), .b(n_14618), .o(n_15905) );
no02s04 g764740 ( .a(n_15700), .b(n_14524), .o(n_15741) );
in01s01 g764741 ( .a(n_16415), .o(n_16480) );
in01s01 g764742 ( .a(n_16450), .o(n_16415) );
na02m04 g764743 ( .a(n_16265), .b(n_16211), .o(n_16450) );
ao12s06 g764744 ( .a(n_15495), .b(n_45135), .c(n_15493), .o(n_15661) );
in01m04 g764745 ( .a(n_15808), .o(n_15853) );
na02s06 g764746 ( .a(n_15739), .b(n_44052), .o(n_15808) );
no02s01 g764747 ( .a(n_15938), .b(n_15937), .o(n_16031) );
in01s01 g764748 ( .a(n_15980), .o(n_15981) );
na02s04 g764749 ( .a(n_46981), .b(n_15935), .o(n_15980) );
na02s01 g764750 ( .a(n_16029), .b(n_16027), .o(n_16028) );
no02f04 g764751 ( .a(n_46981), .b(n_15935), .o(n_16067) );
in01s01 g764753 ( .a(n_15845), .o(n_15893) );
no02f06 g764754 ( .a(n_15732), .b(n_15731), .o(n_15845) );
ao12f06 g764755 ( .a(n_15725), .b(n_15889), .c(n_15793), .o(n_16030) );
in01s01 g764757 ( .a(FE_OCP_RBN3075_n_15706), .o(n_16940) );
na03f06 TIMEBOOST_cell_8324 ( .a(n_9635), .b(FE_RN_319_0), .c(n_9761), .o(FE_RN_320_0) );
oa12m02 g764761 ( .a(n_15273), .b(n_45139), .c(n_15269), .o(n_15629) );
ao12f04 g764762 ( .a(n_15270), .b(FE_OCP_RBN3040_n_45139), .c(n_15272), .o(n_15660) );
ao12f08 g764765 ( .a(n_15461), .b(FE_OCP_RBN3040_n_45139), .c(n_15410), .o(n_15704) );
oa12m10 g764767 ( .a(n_15494), .b(FE_OCP_RBN3041_n_45139), .c(n_15492), .o(n_15768) );
oa12s01 g764768 ( .a(n_15891), .b(n_15890), .c(n_15889), .o(n_15979) );
oa12s01 g764769 ( .a(n_16360), .b(n_16359), .c(n_16358), .o(n_16414) );
in01m04 g764771 ( .a(n_15765), .o(n_15797) );
na02s03 TIMEBOOST_cell_2998 ( .a(n_33816), .b(n_33813), .o(TIMEBOOST_net_790) );
in01s01 g764773 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_7_), .o(n_15892) );
in01s01 g764775 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_5_), .o(n_17158) );
no02m04 g764777 ( .a(n_15649), .b(n_15696), .o(n_15738) );
in01s02 g764779 ( .a(n_15736), .o(n_15737) );
na02s04 g764780 ( .a(n_15702), .b(n_15701), .o(n_15736) );
na02f06 g764781 ( .a(n_15734), .b(FE_RN_1486_0), .o(n_15800) );
na02s04 g764782 ( .a(n_15595), .b(FE_RN_1486_0), .o(n_15628) );
no02f08 TIMEBOOST_cell_2997 ( .a(TIMEBOOST_net_789), .b(n_19172), .o(n_19565) );
na02s04 TIMEBOOST_cell_4255 ( .a(n_29036), .b(n_28704), .o(TIMEBOOST_net_1218) );
na02s01 TIMEBOOST_cell_1015 ( .a(n_37288), .b(n_36970), .o(TIMEBOOST_net_122) );
na03s02 TIMEBOOST_cell_7316 ( .a(n_36750), .b(n_36588), .c(n_36657), .o(n_36658) );
na02s01 g764788 ( .a(n_16359), .b(n_16358), .o(n_16360) );
no02f04 g764789 ( .a(n_15755), .b(n_13879), .o(n_15938) );
no02s10 TIMEBOOST_cell_6861 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_), .o(TIMEBOOST_net_2189) );
no02f02 g764791 ( .a(n_15510), .b(n_15274), .o(n_15559) );
na02s01 g764794 ( .a(n_15844), .b(n_15934), .o(n_16027) );
na02s01 g764795 ( .a(n_15890), .b(n_15889), .o(n_15891) );
no02m06 g764796 ( .a(n_15756), .b(n_13880), .o(n_15937) );
no02s01 g764797 ( .a(FE_OCP_RBN3060_n_15595), .b(n_15656), .o(n_15657) );
no02s06 TIMEBOOST_cell_932 ( .a(TIMEBOOST_net_80), .b(n_23138), .o(n_23237) );
na02f04 g764799 ( .a(n_15730), .b(n_15621), .o(n_15731) );
oa12s04 g764800 ( .a(FE_OCP_RBN6053_n_15514), .b(n_16177), .c(n_16244), .o(n_16265) );
in01s01 g764803 ( .a(n_15708), .o(n_15762) );
in01s01 g764804 ( .a(n_15700), .o(n_15708) );
oa12s04 g764807 ( .a(n_15219), .b(FE_OCP_RBN3099_n_15561), .c(n_15144), .o(n_15698) );
ao12s02 g764808 ( .a(n_46419), .b(FE_OCP_RBN3098_n_15561), .c(n_15182), .o(n_15655) );
oa12f06 g764811 ( .a(n_15723), .b(n_15888), .c(n_15790), .o(n_16029) );
oa12s01 g764812 ( .a(n_15887), .b(n_15888), .c(n_15886), .o(n_15978) );
oa12s01 g764813 ( .a(n_16357), .b(n_16356), .c(n_16355), .o(n_16413) );
in01f02 g764814 ( .a(n_15761), .o(n_15847) );
in01s01 g764816 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_7_), .o(n_17800) );
no02f06 g764818 ( .a(n_15627), .b(n_15622), .o(n_15701) );
no02f04 g764820 ( .a(n_15688), .b(n_15727), .o(n_15728) );
no02m04 g764822 ( .a(n_15627), .b(n_15592), .o(n_15696) );
na02f06 g764823 ( .a(n_15623), .b(n_15591), .o(n_15702) );
na02f04 g764824 ( .a(n_15652), .b(n_14618), .o(n_15730) );
no02s06 TIMEBOOST_cell_931 ( .a(n_23308), .b(FE_RN_248_0), .o(TIMEBOOST_net_80) );
no02f08 TIMEBOOST_cell_3145 ( .a(n_42736), .b(TIMEBOOST_net_863), .o(n_42811) );
na02s01 g764827 ( .a(n_16178), .b(n_16136), .o(n_16359) );
na02s01 g764828 ( .a(n_16356), .b(n_16355), .o(n_16357) );
no02s01 g764829 ( .a(FE_OCP_RBN3134_n_46982), .b(FE_OCP_RBN3072_n_15433), .o(n_15694) );
no02m08 g764831 ( .a(n_15561), .b(FE_OCP_DRV_N4508_n_15099), .o(n_15625) );
na02f04 g764832 ( .a(n_15792), .b(n_15791), .o(n_15934) );
na02s01 g764833 ( .a(n_15726), .b(n_15793), .o(n_15890) );
in01s01 g764834 ( .a(n_15843), .o(n_15844) );
no02m04 g764835 ( .a(n_15792), .b(n_15791), .o(n_15843) );
na02s01 g764836 ( .a(n_15888), .b(n_15886), .o(n_15887) );
ao12f04 g764838 ( .a(n_15553), .b(n_15727), .c(n_15648), .o(n_15758) );
no02s02 g764839 ( .a(n_16139), .b(n_15744), .o(n_16211) );
in01s02 g764841 ( .a(n_15734), .o(n_15692) );
no03f06 TIMEBOOST_cell_8446 ( .a(n_26748), .b(n_26783), .c(n_26827), .o(n_26967) );
in01s01 g764845 ( .a(FE_OCP_RBN3060_n_15595), .o(n_15651) );
no03s06 TIMEBOOST_cell_6623 ( .a(n_32976), .b(n_32961), .c(n_32962), .o(TIMEBOOST_net_2069) );
oa12s01 g764855 ( .a(n_15685), .b(n_15684), .c(n_15683), .o(n_15757) );
in01m02 g764856 ( .a(n_15755), .o(n_15756) );
na02f06 g764857 ( .a(n_15619), .b(n_47333), .o(n_15755) );
oa12s01 g764858 ( .a(n_16354), .b(n_16353), .c(n_16352), .o(n_16412) );
in01s01 g764861 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_4_), .o(n_16503) );
no02s04 g764864 ( .a(n_15623), .b(n_15622), .o(n_15649) );
na02m04 TIMEBOOST_cell_3889 ( .a(n_40890), .b(n_41049), .o(TIMEBOOST_net_1035) );
no02f04 g764866 ( .a(n_15557), .b(n_14452), .o(n_15627) );
in01s02 g764867 ( .a(n_15591), .o(n_15592) );
na02m04 g764868 ( .a(n_15557), .b(FE_OCP_RBN6693_n_13796), .o(n_15591) );
na02f02 g764873 ( .a(n_15551), .b(n_15545), .o(n_15620) );
no02s02 g764874 ( .a(n_16137), .b(n_16138), .o(n_16139) );
na02s01 g764875 ( .a(n_16353), .b(n_16352), .o(n_16354) );
na02f04 g764877 ( .a(n_15687), .b(n_15686), .o(n_15793) );
in01s01 g764878 ( .a(n_15725), .o(n_15726) );
no02f04 g764879 ( .a(n_15687), .b(n_15686), .o(n_15725) );
no02s03 TIMEBOOST_cell_6863 ( .a(n_6708), .b(n_6600), .o(TIMEBOOST_net_2190) );
no02s01 TIMEBOOST_cell_6049 ( .a(FE_OFN738_n_17093), .b(n_18032), .o(TIMEBOOST_net_1876) );
na02s01 g764882 ( .a(n_15684), .b(n_15683), .o(n_15685) );
na02m04 g764883 ( .a(n_15543), .b(n_15586), .o(n_15619) );
no02s01 g764884 ( .a(n_15790), .b(n_15724), .o(n_15886) );
in01s01 g764885 ( .a(n_16177), .o(n_16178) );
na02m04 g764886 ( .a(n_16137), .b(n_15632), .o(n_16177) );
oa12s01 g764887 ( .a(n_16136), .b(n_16026), .c(n_16135), .o(n_16356) );
na02f08 g764896 ( .a(n_15438), .b(n_15390), .o(n_15561) );
no02f06 g764898 ( .a(n_15677), .b(n_15680), .o(n_15888) );
in01s01 g764899 ( .a(n_15652), .o(n_15598) );
no03s04 TIMEBOOST_cell_7542 ( .a(FE_OCP_RBN6600_n_7708), .b(n_9304), .c(FE_OCP_RBN2612_FE_OCPN857_n_7802), .o(TIMEBOOST_net_2402) );
oa12s01 g764901 ( .a(n_15754), .b(n_15753), .c(n_15752), .o(n_15842) );
na02m06 g764903 ( .a(n_15473), .b(n_15502), .o(n_15622) );
na02f08 g764905 ( .a(n_15546), .b(n_15548), .o(n_15727) );
na02f06 TIMEBOOST_cell_2994 ( .a(n_13353), .b(n_13380), .o(TIMEBOOST_net_788) );
no02f04 TIMEBOOST_cell_7541 ( .a(TIMEBOOST_net_2401), .b(n_13559), .o(TIMEBOOST_net_2080) );
no02f08 TIMEBOOST_cell_2124 ( .a(n_43788), .b(TIMEBOOST_net_676), .o(n_43885) );
no02m04 g764911 ( .a(n_15552), .b(n_14588), .o(n_15553) );
na02f02 g764912 ( .a(n_15552), .b(n_14452), .o(n_15551) );
na02s04 g764913 ( .a(n_15552), .b(n_14524), .o(n_15648) );
na02f06 g764915 ( .a(n_15440), .b(n_15437), .o(n_15586) );
na02m02 g764916 ( .a(n_15433), .b(n_14420), .o(n_15476) );
na02m04 g764917 ( .a(n_16066), .b(n_15633), .o(n_16137) );
no02f06 g764918 ( .a(n_15612), .b(n_15611), .o(n_15615) );
no02f04 g764919 ( .a(n_15679), .b(n_15678), .o(n_15790) );
no02m04 TIMEBOOST_cell_6098 ( .a(TIMEBOOST_net_1900), .b(n_14281), .o(n_14441) );
na02m02 g764922 ( .a(n_15434), .b(n_15187), .o(n_15475) );
ao12f06 g764923 ( .a(FE_OCP_DRV_N6895_n_15391), .b(n_15320), .c(FE_OCP_RBN5948_n_14982), .o(n_15438) );
na02f02 g764925 ( .a(n_15584), .b(n_15537), .o(n_15614) );
na02f06 TIMEBOOST_cell_7557 ( .a(TIMEBOOST_net_2409), .b(TIMEBOOST_net_1481), .o(n_13883) );
in01s01 g764927 ( .a(n_15723), .o(n_15724) );
na02m04 g764928 ( .a(n_15679), .b(n_15678), .o(n_15723) );
na02s01 g764929 ( .a(n_15753), .b(n_15752), .o(n_15754) );
in01s02 g764930 ( .a(n_15394), .o(n_15395) );
na02m02 g764931 ( .a(n_15357), .b(n_15113), .o(n_15394) );
ao12s01 g764932 ( .a(n_16066), .b(FE_OCP_RBN3195_n_15599), .c(n_16246), .o(n_16353) );
ao12s01 g764933 ( .a(n_16312), .b(n_16264), .c(n_16384), .o(n_16385) );
no02s02 TIMEBOOST_cell_3274 ( .a(n_15974), .b(n_16019), .o(TIMEBOOST_net_928) );
no02f06 g764935 ( .a(n_15612), .b(n_15536), .o(n_15613) );
in01s01 g764937 ( .a(FE_OCPN1278_n_15656), .o(n_15549) );
in01s01 g764938 ( .a(n_45502), .o(n_15656) );
ao12f06 g764941 ( .a(n_15194), .b(n_15286), .c(FE_OCPN1077_n_13831), .o(n_15356) );
oa12s01 g764942 ( .a(n_15675), .b(n_15674), .c(n_15673), .o(n_15751) );
oa12s01 g764943 ( .a(n_15608), .b(n_15674), .c(n_15611), .o(n_15684) );
ao12s01 g764944 ( .a(n_15541), .b(n_15610), .c(n_15609), .o(n_15683) );
ao12f04 g764945 ( .a(n_15643), .b(n_15676), .c(n_15606), .o(n_15677) );
oa12s01 g764946 ( .a(n_16351), .b(n_16350), .c(n_16349), .o(n_16411) );
in01m04 g764948 ( .a(n_15547), .o(n_15548) );
na02s04 g764950 ( .a(n_15387), .b(FE_OCP_RBN6693_n_13796), .o(n_15437) );
no02m08 TIMEBOOST_cell_2993 ( .a(FE_RN_152_0), .b(TIMEBOOST_net_787), .o(n_45521) );
no02s04 TIMEBOOST_cell_4335 ( .a(n_14613), .b(n_14396), .o(TIMEBOOST_net_1258) );
in01m04 g764956 ( .a(n_15545), .o(n_15546) );
no03s08 TIMEBOOST_cell_2272 ( .a(FE_OCP_RBN4007_n_32860), .b(n_32963), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_23_), .o(FE_RN_656_0) );
na02f04 g764958 ( .a(FE_OCP_RBN5994_n_15387), .b(FE_OCPN1703_n_14210), .o(n_15440) );
na02m04 g764959 ( .a(FE_OCP_RBN5993_n_15387), .b(n_14215), .o(n_15473) );
na02f06 g764961 ( .a(n_15503), .b(n_15502), .o(n_15543) );
na02s01 g764962 ( .a(n_16350), .b(n_16349), .o(n_16351) );
no02s03 g764963 ( .a(n_15385), .b(n_15468), .o(n_15501) );
no02f06 TIMEBOOST_cell_3273 ( .a(TIMEBOOST_net_927), .b(n_5732), .o(n_5893) );
no02f08 g764965 ( .a(n_15498), .b(n_15496), .o(n_15612) );
na02f04 g764967 ( .a(FE_OCP_RBN2103_n_15286), .b(FE_RN_1141_0), .o(n_15353) );
na02m06 g764968 ( .a(n_15242), .b(n_15157), .o(n_15357) );
no02m02 g764970 ( .a(n_15389), .b(n_15391), .o(n_15434) );
na02s06 g764971 ( .a(n_15389), .b(n_13950), .o(n_15390) );
na02s01 g764972 ( .a(n_15674), .b(n_15673), .o(n_15675) );
no02s01 g764973 ( .a(n_15610), .b(n_15609), .o(n_15541) );
ao12s01 g764974 ( .a(n_16312), .b(n_16176), .c(FE_OCP_RBN3193_n_15599), .o(n_16313) );
in01s01 g764975 ( .a(n_16066), .o(n_16026) );
no02m04 g764976 ( .a(n_15933), .b(n_15563), .o(n_16066) );
in01s01 g764981 ( .a(FE_OCP_RBN3072_n_15433), .o(n_15479) );
oa22f02 g764984 ( .a(n_15321), .b(n_15154), .c(n_15284), .d(n_15153), .o(n_15433) );
no03f04 TIMEBOOST_cell_5346 ( .a(n_20977), .b(n_21012), .c(n_20976), .o(TIMEBOOST_net_1621) );
no02m40 TIMEBOOST_cell_8135 ( .a(TIMEBOOST_net_2698), .b(TIMEBOOST_net_1379), .o(n_16972) );
oa12s01 g764987 ( .a(n_15642), .b(n_15641), .c(n_15640), .o(n_15722) );
na02s01 g764988 ( .a(n_15607), .b(n_15580), .o(n_15753) );
ao12s01 g764989 ( .a(n_15581), .b(n_15644), .c(n_15643), .o(n_15752) );
in01s01 g764990 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_5_), .o(n_17589) );
in01m01 g764992 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_3_), .o(n_17496) );
in01f02 g764994 ( .a(n_15468), .o(n_15469) );
na02f06 g764995 ( .a(n_15427), .b(n_15323), .o(n_15468) );
na02f04 g764996 ( .a(n_15429), .b(n_14419), .o(n_15504) );
in01s01 g764997 ( .a(n_15537), .o(n_15538) );
na02m02 g764998 ( .a(n_15500), .b(n_15426), .o(n_15537) );
no02m02 g764999 ( .a(n_15314), .b(n_14420), .o(n_15352) );
no02m06 TIMEBOOST_cell_7620 ( .a(n_44139), .b(n_29160), .o(TIMEBOOST_net_2441) );
na02f04 TIMEBOOST_cell_5635 ( .a(TIMEBOOST_net_1765), .b(n_40557), .o(n_40577) );
na02s02 TIMEBOOST_cell_6945 ( .a(n_2419), .b(n_2394), .o(TIMEBOOST_net_2231) );
na02f08 g765003 ( .a(n_15385), .b(n_15427), .o(n_15503) );
na02f04 g765004 ( .a(n_15497), .b(n_15609), .o(n_15536) );
no02s01 g765005 ( .a(n_15644), .b(n_15643), .o(n_15581) );
no02m06 g765006 ( .a(n_15321), .b(n_15112), .o(n_15389) );
na02f06 g765007 ( .a(FE_OCP_RBN1821_n_13858), .b(n_15321), .o(n_15320) );
na02s01 g765008 ( .a(n_15497), .b(n_15608), .o(n_15673) );
no02f02 TIMEBOOST_cell_4450 ( .a(TIMEBOOST_net_1315), .b(n_5284), .o(TIMEBOOST_net_1120) );
no02f04 g765010 ( .a(n_15465), .b(n_15420), .o(n_15535) );
na02f06 g765011 ( .a(n_15529), .b(n_15580), .o(n_15676) );
na02s01 g765012 ( .a(n_15641), .b(n_15640), .o(n_15642) );
na02s01 g765013 ( .a(n_15641), .b(n_15606), .o(n_15607) );
in01s01 g765014 ( .a(n_16263), .o(n_16264) );
no02s01 TIMEBOOST_cell_8574 ( .a(FE_OCP_RBN5852_n_3625), .b(FE_OCP_RBN5851_n_3625), .o(TIMEBOOST_net_2774) );
in01s01 g765016 ( .a(n_15933), .o(n_16350) );
no02s04 g765017 ( .a(n_15789), .b(n_15721), .o(n_15933) );
na02s06 TIMEBOOST_cell_8715 ( .a(TIMEBOOST_net_2844), .b(n_17828), .o(n_17932) );
in01s01 g765019 ( .a(n_15498), .o(n_15674) );
ao12f06 g765020 ( .a(n_15380), .b(n_15532), .c(n_15460), .o(n_15498) );
in01f04 g765027 ( .a(n_15242), .o(n_15286) );
ao12f08 g765028 ( .a(n_14987), .b(n_15084), .c(n_14986), .o(n_15242) );
oa12s01 g765029 ( .a(n_15534), .b(n_15533), .c(n_15532), .o(n_15605) );
no02s04 TIMEBOOST_cell_5280 ( .a(n_4405), .b(n_4543), .o(TIMEBOOST_net_1588) );
in01m01 g765033 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_4_), .o(n_17478) );
no02m04 g765036 ( .a(n_15206), .b(FE_OCP_RBN5800_n_13962), .o(n_15241) );
in01f02 g765037 ( .a(n_15464), .o(n_15465) );
na02f04 g765038 ( .a(n_15426), .b(n_15425), .o(n_15464) );
na02m04 g765039 ( .a(n_15382), .b(n_15425), .o(n_15500) );
na02f06 g765040 ( .a(n_15282), .b(n_14215), .o(n_15323) );
na02s06 g765041 ( .a(n_15282), .b(FE_OCP_RBN5801_n_13962), .o(n_15502) );
na02s06 g765042 ( .a(n_15281), .b(FE_OCP_RBN6693_n_13796), .o(n_15427) );
na02s06 TIMEBOOST_cell_6940 ( .a(TIMEBOOST_net_2228), .b(FE_OCP_RBN4191_n_34285), .o(FE_RN_2266_0) );
no02s02 g765044 ( .a(n_16103), .b(n_15972), .o(n_16104) );
oa12s01 g765045 ( .a(n_16102), .b(n_15975), .c(FE_OCP_RBN3190_n_15599), .o(n_16312) );
in01s02 g765047 ( .a(n_15497), .o(n_15611) );
in01s01 g765049 ( .a(n_15496), .o(n_15608) );
na02s01 TIMEBOOST_cell_7876 ( .a(n_4213), .b(n_4087), .o(TIMEBOOST_net_2569) );
na02s01 g765052 ( .a(n_15533), .b(n_15532), .o(n_15534) );
no02f02 g765053 ( .a(n_15530), .b(FE_OFN806_n_13742), .o(n_15531) );
no02s01 g765054 ( .a(n_15490), .b(n_15530), .o(n_15640) );
na02s01 g765055 ( .a(n_16133), .b(n_16175), .o(n_16176) );
in01m02 g765057 ( .a(n_15385), .o(n_15423) );
ao12f08 g765058 ( .a(n_15239), .b(n_15276), .c(n_15205), .o(n_15385) );
no02s01 g765059 ( .a(n_15977), .b(n_15926), .o(n_16384) );
ao12m02 g765060 ( .a(n_15514), .b(n_16347), .c(n_15788), .o(n_15789) );
in01s01 g765065 ( .a(n_15321), .o(n_15284) );
in01f01 g765067 ( .a(n_15429), .o(n_15384) );
no02s01 TIMEBOOST_cell_8537 ( .a(TIMEBOOST_net_2755), .b(n_14081), .o(TIMEBOOST_net_1295) );
na02f04 g765069 ( .a(n_15383), .b(n_15422), .o(n_15644) );
in01s01 g765070 ( .a(n_15529), .o(n_15641) );
oa12f06 g765071 ( .a(n_15378), .b(n_15526), .c(n_15457), .o(n_15529) );
oa12s01 g765072 ( .a(n_15528), .b(n_15527), .c(n_15526), .o(n_15603) );
oa12s01 g765073 ( .a(n_16348), .b(n_16347), .c(n_16346), .o(n_16410) );
in01s40 g765075 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_2_), .o(n_17018) );
na02f02 g765077 ( .a(n_15344), .b(n_15305), .o(n_15383) );
na02f04 g765078 ( .a(n_15345), .b(n_15306), .o(n_15422) );
na02f02 g765079 ( .a(n_15237), .b(n_15278), .o(n_15313) );
no02m02 g765080 ( .a(n_15239), .b(n_15238), .o(n_15349) );
na02m02 g765081 ( .a(n_15200), .b(n_14215), .o(n_15240) );
no02m04 TIMEBOOST_cell_5335 ( .a(TIMEBOOST_net_1615), .b(n_20736), .o(n_20889) );
na02s04 g765083 ( .a(FE_OCP_RBN2833_n_13962), .b(n_15275), .o(n_15425) );
na02f04 g765085 ( .a(FE_OCP_RBN3070_n_15275), .b(n_14419), .o(n_15426) );
na02s01 g765086 ( .a(n_15976), .b(n_15923), .o(n_15977) );
na02s01 g765087 ( .a(n_16024), .b(n_15837), .o(n_16025) );
no02s01 g765088 ( .a(n_16101), .b(n_16098), .o(n_16261) );
in01s01 g765089 ( .a(n_15494), .o(n_15495) );
ao12m06 g765090 ( .a(n_15461), .b(FE_OCP_RBN6798_n_15156), .c(n_15341), .o(n_15494) );
no02s02 g765091 ( .a(n_15492), .b(n_15491), .o(n_15493) );
in01s01 g765092 ( .a(n_15580), .o(n_15490) );
na02m04 g765093 ( .a(n_15459), .b(n_15458), .o(n_15580) );
na02s01 g765095 ( .a(n_15381), .b(n_15460), .o(n_15533) );
in01s02 g765096 ( .a(n_15530), .o(n_15606) );
no02f04 g765097 ( .a(n_15459), .b(n_15458), .o(n_15530) );
na02s01 g765098 ( .a(n_15527), .b(n_15526), .o(n_15528) );
na02s01 g765099 ( .a(n_16347), .b(n_16346), .o(n_16348) );
in01s02 g765100 ( .a(n_15420), .o(n_15421) );
in01s02 g765101 ( .a(n_15382), .o(n_15420) );
ao12f04 g765102 ( .a(n_15233), .b(n_15243), .c(n_15311), .o(n_15382) );
na02s01 g765103 ( .a(n_15931), .b(n_16023), .o(n_16103) );
in01s01 g765104 ( .a(n_16310), .o(n_16311) );
oa12s01 g765105 ( .a(n_15976), .b(n_15884), .c(FE_OCP_RBN3190_n_15599), .o(n_16310) );
in01s01 g765106 ( .a(n_16259), .o(n_16260) );
ao12s01 g765107 ( .a(n_16101), .b(n_16100), .c(n_16245), .o(n_16259) );
in01s01 g765108 ( .a(n_16308), .o(n_16309) );
oa12s01 g765109 ( .a(n_16258), .b(n_16175), .c(FE_OCP_RBN3190_n_15599), .o(n_16308) );
in01s01 g765110 ( .a(n_16133), .o(n_16134) );
oa12s01 g765111 ( .a(FE_OCP_RBN3193_n_15599), .b(n_16100), .c(n_16099), .o(n_16133) );
na02f06 g765112 ( .a(n_15277), .b(n_15310), .o(n_15463) );
in01m02 g765113 ( .a(n_15163), .o(n_15164) );
in01m01 g765114 ( .a(n_15084), .o(n_15163) );
oa12f08 g765115 ( .a(n_14908), .b(n_15026), .c(n_14909), .o(n_15084) );
oa12f06 g765116 ( .a(n_15264), .b(n_15415), .c(n_15339), .o(n_15532) );
no02s02 TIMEBOOST_cell_8697 ( .a(TIMEBOOST_net_2835), .b(n_37514), .o(TIMEBOOST_net_1432) );
oa12s01 g765118 ( .a(n_15417), .b(n_15416), .c(n_15415), .o(n_15489) );
oa12s01 g765119 ( .a(n_15414), .b(n_15413), .c(n_15412), .o(n_15488) );
in01f04 g765120 ( .a(n_15281), .o(n_15282) );
na02m06 TIMEBOOST_cell_2988 ( .a(n_13201), .b(n_13209), .o(TIMEBOOST_net_785) );
in01s06 g765127 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_3_), .o(n_17347) );
in01f01 g765130 ( .a(n_15239), .o(n_15278) );
no02f06 g765131 ( .a(n_15204), .b(n_14215), .o(n_15239) );
no02f06 TIMEBOOST_cell_5142 ( .a(FE_OCP_RBN4177_n_38586), .b(FE_OFN5092_delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(TIMEBOOST_net_1519) );
in01m02 g765133 ( .a(n_15237), .o(n_15238) );
na02m06 g765134 ( .a(n_15204), .b(FE_OCP_RBN5790_n_13962), .o(n_15205) );
na02m02 g765135 ( .a(n_15204), .b(n_14215), .o(n_15237) );
in01f02 g765136 ( .a(n_15344), .o(n_15345) );
na02f02 g765137 ( .a(n_15311), .b(n_15234), .o(n_15344) );
no02s02 TIMEBOOST_cell_7461 ( .a(TIMEBOOST_net_2361), .b(n_33146), .o(TIMEBOOST_net_1419) );
na02s01 g765139 ( .a(FE_OCP_RBN3190_n_15599), .b(n_15884), .o(n_15976) );
na02s01 g765140 ( .a(n_15836), .b(n_15830), .o(n_15883) );
no02s01 g765141 ( .a(n_16020), .b(n_15634), .o(n_15975) );
na02s01 g765142 ( .a(n_15971), .b(n_15969), .o(n_16022) );
no02s02 g765143 ( .a(n_15638), .b(n_15788), .o(n_15721) );
no02s01 g765144 ( .a(n_16100), .b(FE_OCP_RBN3194_n_15599), .o(n_16101) );
na02s01 g765145 ( .a(n_16175), .b(FE_OCP_RBN3190_n_15599), .o(n_16258) );
na02s04 g765146 ( .a(n_15151), .b(n_15235), .o(n_15277) );
na02f04 g765147 ( .a(n_15189), .b(FE_OCP_RBN5970_n_15235), .o(n_15310) );
na02s06 g765148 ( .a(n_15343), .b(n_15342), .o(n_15460) );
in01s01 g765149 ( .a(n_15380), .o(n_15381) );
no02f04 g765150 ( .a(n_15343), .b(n_15342), .o(n_15380) );
no02s01 g765151 ( .a(n_15457), .b(n_15379), .o(n_15527) );
no02s01 TIMEBOOST_cell_6227 ( .a(n_3706), .b(FE_OCP_RBN4274_n_3700), .o(TIMEBOOST_net_1965) );
na02s01 g765155 ( .a(n_15416), .b(n_15415), .o(n_15417) );
na02s01 g765156 ( .a(n_15413), .b(n_15412), .o(n_15414) );
oa12s02 g765157 ( .a(n_15879), .b(n_15827), .c(FE_OCP_RBN6845_n_15599), .o(n_15974) );
no02s01 g765158 ( .a(n_15832), .b(n_15932), .o(n_16024) );
na02s01 g765159 ( .a(n_15930), .b(n_15835), .o(n_15931) );
in01s02 g765160 ( .a(n_15308), .o(n_15309) );
in01s02 g765161 ( .a(n_15276), .o(n_15308) );
in01s01 g765163 ( .a(n_15972), .o(n_15973) );
na02s02 g765164 ( .a(n_15841), .b(n_15929), .o(n_15972) );
no02m04 g765165 ( .a(n_15637), .b(n_15515), .o(n_16347) );
no02f04 g765167 ( .a(n_15123), .b(n_15159), .o(n_15275) );
no02s01 TIMEBOOST_cell_2926 ( .a(n_28672), .b(n_28673), .o(TIMEBOOST_net_754) );
in01s01 g765174 ( .a(n_15124), .o(n_15160) );
oa12f08 g765175 ( .a(n_14927), .b(n_15023), .c(n_14877), .o(n_15124) );
ao12f06 g765177 ( .a(n_15340), .b(n_15296), .c(n_15256), .o(n_15526) );
oa12s01 g765178 ( .a(n_16345), .b(n_16344), .c(FE_OCP_RBN5394_cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n_16409) );
oa12s01 g765179 ( .a(n_16343), .b(n_16342), .c(n_16341), .o(n_16408) );
in01s06 g765180 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_2_), .o(n_17229) );
na02s01 g765182 ( .a(n_16344), .b(FE_OCP_RBN5394_cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n_16345) );
na02f04 g765184 ( .a(n_15082), .b(n_15118), .o(n_15235) );
no02f04 g765185 ( .a(FE_OCP_RBN5984_n_15079), .b(FE_OCP_RBN5800_n_13962), .o(n_15159) );
no02m02 g765186 ( .a(n_15079), .b(FE_OCP_RBN2837_n_13962), .o(n_15123) );
in01f01 g765187 ( .a(n_15233), .o(n_15234) );
no02f04 g765188 ( .a(n_15198), .b(FE_OCPN1703_n_14210), .o(n_15233) );
na02m04 g765189 ( .a(n_15198), .b(FE_OCPN1703_n_14210), .o(n_15311) );
no02s01 g765190 ( .a(n_15840), .b(n_15839), .o(n_15841) );
no02s01 g765191 ( .a(n_16020), .b(n_16016), .o(n_16065) );
na02s01 g765192 ( .a(n_15881), .b(n_15749), .o(n_15882) );
no02s01 g765193 ( .a(n_15828), .b(n_15839), .o(n_15880) );
in01s01 g765194 ( .a(n_16063), .o(n_16064) );
no02s01 g765195 ( .a(n_16021), .b(n_16020), .o(n_16063) );
in01s01 g765196 ( .a(n_16131), .o(n_16132) );
no02s01 g765197 ( .a(n_16099), .b(n_16098), .o(n_16131) );
na02f02 g765199 ( .a(n_15081), .b(n_15157), .o(n_15196) );
na02s02 g765200 ( .a(n_15272), .b(n_15273), .o(n_15274) );
no02f02 g765201 ( .a(n_15269), .b(n_15270), .o(n_15271) );
in01s02 g765202 ( .a(n_15408), .o(n_15409) );
no02s06 g765203 ( .a(n_15771), .b(n_15300), .o(n_15408) );
na02m02 g765204 ( .a(n_15302), .b(n_15299), .o(n_15341) );
no02s04 TIMEBOOST_cell_2925 ( .a(TIMEBOOST_net_753), .b(n_19184), .o(n_19280) );
no02s01 g765206 ( .a(n_15257), .b(n_15340), .o(n_15413) );
in01s01 g765207 ( .a(n_15378), .o(n_15379) );
na02m04 g765208 ( .a(n_15338), .b(n_15337), .o(n_15378) );
na02s01 g765209 ( .a(n_15405), .b(n_15403), .o(n_15487) );
no02s01 g765210 ( .a(n_15265), .b(n_15339), .o(n_15416) );
no02f04 g765213 ( .a(n_15338), .b(n_15337), .o(n_15457) );
na02s01 g765214 ( .a(n_16342), .b(n_16341), .o(n_16343) );
in01m02 g765215 ( .a(n_15305), .o(n_15306) );
in01m01 g765216 ( .a(n_15243), .o(n_15305) );
ao12f04 g765217 ( .a(n_15110), .b(n_15136), .c(n_15195), .o(n_15243) );
na02s01 g765218 ( .a(n_15968), .b(n_16023), .o(n_16062) );
in01s01 g765219 ( .a(n_16256), .o(n_16257) );
ao12s01 g765220 ( .a(n_15840), .b(n_16245), .c(n_15748), .o(n_16256) );
no02s01 g765221 ( .a(n_15785), .b(n_15750), .o(n_15838) );
in01s01 g765222 ( .a(n_15878), .o(n_15879) );
ao12s01 g765223 ( .a(FE_OCP_RBN6845_n_15599), .b(n_15837), .c(n_14779), .o(n_15878) );
na02f06 TIMEBOOST_cell_6270 ( .a(TIMEBOOST_net_1986), .b(n_10591), .o(n_10709) );
in01s01 g765225 ( .a(n_15836), .o(n_15932) );
oa12s01 g765226 ( .a(n_15719), .b(n_15787), .c(n_15786), .o(n_15836) );
in01s01 g765227 ( .a(n_15637), .o(n_15638) );
na02s02 TIMEBOOST_cell_6894 ( .a(TIMEBOOST_net_2205), .b(FE_OCP_RBN2507_n_37720), .o(n_37769) );
in01s01 g765229 ( .a(n_15971), .o(n_16210) );
oa12s01 g765230 ( .a(n_15664), .b(n_15928), .c(n_15360), .o(n_15971) );
ao12s01 g765231 ( .a(FE_OCP_RBN3190_n_15599), .b(n_15969), .c(n_15512), .o(n_15970) );
oa12s01 g765232 ( .a(n_15664), .b(n_15834), .c(n_15833), .o(n_15835) );
ao12s01 g765233 ( .a(n_15664), .b(n_15830), .c(n_15666), .o(n_15832) );
in01m02 g765238 ( .a(n_15059), .o(n_15060) );
in01s02 g765239 ( .a(n_15026), .o(n_15059) );
ao12f08 g765240 ( .a(n_14854), .b(n_14944), .c(n_14906), .o(n_15026) );
no02s02 TIMEBOOST_cell_4469 ( .a(n_39479), .b(n_39250), .o(TIMEBOOST_net_1325) );
in01s01 g765242 ( .a(n_15453), .o(n_15454) );
na02s02 g765243 ( .a(n_15407), .b(n_15335), .o(n_15453) );
in01s01 g765244 ( .a(n_15635), .o(n_15636) );
no02s01 TIMEBOOST_cell_2924 ( .a(n_18425), .b(n_18426), .o(TIMEBOOST_net_753) );
no02s01 g765247 ( .a(n_15142), .b(n_15297), .o(n_15455) );
oa12s01 g765248 ( .a(n_15227), .b(n_15226), .c(n_15225), .o(n_15303) );
oa12s01 g765250 ( .a(n_15333), .b(n_15332), .c(n_15331), .o(n_15406) );
na02f06 g765251 ( .a(n_15025), .b(n_15058), .o(n_15204) );
in01s01 g765252 ( .a(n_15884), .o(n_15634) );
ao12s01 g765253 ( .a(n_15522), .b(n_15521), .c(n_15520), .o(n_15884) );
ao12s01 g765254 ( .a(n_15577), .b(n_15576), .c(n_15575), .o(n_16175) );
oa12s01 g765255 ( .a(n_15574), .b(n_15573), .c(n_15572), .o(n_16100) );
in01s02 g765256 ( .a(n_15601), .o(n_15602) );
na02s02 g765257 ( .a(n_15486), .b(n_15452), .o(n_15601) );
in01s01 g765258 ( .a(n_15266), .o(n_15267) );
in01s02 g765260 ( .a(n_15376), .o(n_15377) );
na02s04 g765261 ( .a(n_15230), .b(n_15263), .o(n_15376) );
in01s01 g765262 ( .a(n_15671), .o(n_15672) );
na02s02 g765263 ( .a(n_15517), .b(n_15571), .o(n_15671) );
in01s01 g765264 ( .a(n_15523), .o(n_15524) );
no02s01 g765266 ( .a(n_15521), .b(n_15520), .o(n_15522) );
no02s01 g765267 ( .a(n_15576), .b(n_15575), .o(n_15577) );
na02s01 g765268 ( .a(n_15573), .b(n_15572), .o(n_15574) );
na02m02 g765269 ( .a(n_15047), .b(FE_OCP_RBN5790_n_13962), .o(n_15082) );
na02f02 g765271 ( .a(n_14991), .b(FE_OCP_RBN5800_n_13962), .o(n_15025) );
na02f04 g765272 ( .a(FE_OCP_RBN2093_n_14991), .b(FE_OCP_RBN2834_n_13962), .o(n_15058) );
na02f04 g765273 ( .a(FE_OCP_RBN5328_n_15047), .b(FE_OCP_RBN2834_n_13962), .o(n_15118) );
na02f04 g765276 ( .a(n_15195), .b(FE_OCP_RBN6807_n_15110), .o(n_15231) );
in01s01 g765277 ( .a(n_15785), .o(n_15881) );
na02s01 g765278 ( .a(n_15668), .b(n_15783), .o(n_15785) );
na02s01 g765279 ( .a(n_15714), .b(n_15749), .o(n_15750) );
no02s01 g765280 ( .a(n_15826), .b(n_15829), .o(n_16023) );
no02s01 g765281 ( .a(n_15876), .b(n_15873), .o(n_15877) );
na02s01 g765282 ( .a(n_15921), .b(n_15924), .o(n_16019) );
in01s01 g765283 ( .a(n_15828), .o(n_15929) );
na02s01 g765284 ( .a(n_15922), .b(n_15784), .o(n_15828) );
in01s01 g765285 ( .a(n_15926), .o(n_15927) );
na02s01 g765286 ( .a(n_15875), .b(n_16255), .o(n_15926) );
no02s01 g765287 ( .a(n_15967), .b(n_15868), .o(n_15968) );
in01s01 g765288 ( .a(n_16306), .o(n_16307) );
na02s01 g765289 ( .a(n_16255), .b(n_16174), .o(n_16306) );
na02f04 TIMEBOOST_cell_6269 ( .a(FE_OCP_RBN6049_n_10570), .b(FE_OCPN1067_n_44461), .o(TIMEBOOST_net_1986) );
in01s01 g765291 ( .a(n_16060), .o(n_16061) );
na02s01 g765292 ( .a(n_15919), .b(n_16018), .o(n_16060) );
no02s01 g765293 ( .a(n_15961), .b(FE_OCP_RBN3190_n_15599), .o(n_16099) );
no02s01 g765294 ( .a(n_15781), .b(n_15869), .o(n_15827) );
in01s01 g765295 ( .a(n_15964), .o(n_15965) );
na02s01 g765296 ( .a(n_15925), .b(n_15924), .o(n_15964) );
in01s01 g765297 ( .a(n_15923), .o(n_16021) );
na02s01 g765298 ( .a(FE_OCP_RBN3190_n_15599), .b(n_15870), .o(n_15923) );
na02s01 g765299 ( .a(n_15716), .b(n_15783), .o(n_16479) );
no02s01 g765300 ( .a(n_15709), .b(n_15717), .o(n_16505) );
no02s01 g765301 ( .a(n_15745), .b(n_15873), .o(n_16543) );
in01s01 g765302 ( .a(n_15871), .o(n_15872) );
no02s01 g765303 ( .a(n_15826), .b(n_15834), .o(n_15871) );
in01s01 g765304 ( .a(n_15962), .o(n_15963) );
na02s01 g765305 ( .a(n_15710), .b(n_15969), .o(n_15962) );
no02s01 g765306 ( .a(FE_OCP_RBN6846_n_15599), .b(n_15748), .o(n_15840) );
no02s01 g765307 ( .a(n_15719), .b(n_15870), .o(n_16020) );
in01s01 g765308 ( .a(n_16017), .o(n_16098) );
na02s01 g765309 ( .a(FE_OCP_RBN3190_n_15599), .b(n_15961), .o(n_16017) );
in01s01 g765310 ( .a(n_15959), .o(n_15960) );
na02s01 g765311 ( .a(n_15922), .b(n_15822), .o(n_15959) );
no02f04 g765312 ( .a(n_15208), .b(n_15207), .o(n_15339) );
in01s01 g765313 ( .a(n_15264), .o(n_15265) );
na02f04 g765314 ( .a(n_15208), .b(n_15207), .o(n_15264) );
na02s02 g765315 ( .a(n_15021), .b(FE_OCP_DRV_N4499_n_13785), .o(n_15157) );
na02s02 g765316 ( .a(n_15194), .b(FE_OCPN1250_n_13882), .o(n_15273) );
no02f01 g765317 ( .a(n_15156), .b(n_13912), .o(n_15270) );
na02s02 g765318 ( .a(n_15156), .b(n_13912), .o(n_15272) );
no02s02 g765319 ( .a(n_15194), .b(FE_OCPN1250_n_13882), .o(n_15269) );
na02s02 g765320 ( .a(FE_OCP_RBN5711_n_13984), .b(FE_OCP_RBN4324_n_15156), .o(n_15230) );
na02s02 g765321 ( .a(FE_OCP_RBN4322_n_15156), .b(FE_OCP_RBN5710_n_13984), .o(n_15263) );
in01m01 g765322 ( .a(n_15302), .o(n_15771) );
na02s06 g765324 ( .a(FE_OCP_RBN4322_n_15156), .b(FE_OCP_RBN2727_n_14018), .o(n_15302) );
in01s01 g765325 ( .a(FE_OCP_RBN3015_n_15300), .o(n_15336) );
no02s04 g765327 ( .a(FE_OCP_RBN4322_n_15156), .b(FE_OCP_RBN2727_n_14018), .o(n_15300) );
in01s04 g765328 ( .a(n_15113), .o(n_15114) );
na02m01 g765329 ( .a(n_15048), .b(FE_OCP_DRV_N4500_n_13785), .o(n_15081) );
na02s06 g765330 ( .a(n_15048), .b(FE_OCP_DRV_N4500_n_13785), .o(n_15113) );
na02s02 g765331 ( .a(FE_OCP_RBN6799_n_15156), .b(FE_OCP_RBN2731_n_14072), .o(n_15335) );
na02s04 g765332 ( .a(FE_OCP_RBN4323_n_15156), .b(n_15299), .o(n_15407) );
na02s01 g765333 ( .a(FE_OCP_RBN6801_n_15156), .b(n_14157), .o(n_15486) );
na02s02 g765334 ( .a(FE_OCP_RBN6802_n_15156), .b(FE_OCP_RBN2750_n_14157), .o(n_15452) );
na02f08 TIMEBOOST_cell_2923 ( .a(TIMEBOOST_net_752), .b(n_13513), .o(n_13633) );
no02s01 g765338 ( .a(FE_OCP_RBN6798_n_15156), .b(n_14397), .o(n_15491) );
na02s01 g765339 ( .a(FE_OCP_RBN5987_n_15135), .b(n_14225), .o(n_15517) );
na02s01 g765340 ( .a(FE_OCP_RBN6798_n_15156), .b(n_14265), .o(n_15571) );
in01m02 g765341 ( .a(n_15153), .o(n_15154) );
no02f02 g765342 ( .a(n_15112), .b(n_15049), .o(n_15153) );
no02s02 g765345 ( .a(n_15127), .b(n_15180), .o(n_15298) );
na02s03 g765346 ( .a(n_15258), .b(n_15218), .o(n_15259) );
no02s03 g765347 ( .a(n_15180), .b(FE_OCP_RBN2079_n_14149), .o(n_15228) );
in01s01 g765349 ( .a(n_15374), .o(n_15375) );
no02s02 g765350 ( .a(n_15806), .b(n_15293), .o(n_15374) );
no02f04 g765351 ( .a(n_15224), .b(n_15223), .o(n_15340) );
in01s01 TIMEBOOST_cell_5914 ( .a(TIMEBOOST_net_1802), .o(TIMEBOOST_net_1803) );
in01s01 g765353 ( .a(n_15404), .o(n_15405) );
na02s02 g765354 ( .a(n_15373), .b(n_15330), .o(n_15404) );
na02s01 g765355 ( .a(n_15226), .b(n_15225), .o(n_15227) );
no02m04 TIMEBOOST_cell_5423 ( .a(TIMEBOOST_net_1659), .b(FE_OCP_RBN3237_n_5130), .o(n_5308) );
in01s01 g765357 ( .a(n_15256), .o(n_15257) );
na02f04 g765358 ( .a(n_15224), .b(n_15223), .o(n_15256) );
na02s01 g765359 ( .a(n_15332), .b(n_15331), .o(n_15333) );
no02m04 TIMEBOOST_cell_4468 ( .a(TIMEBOOST_net_1324), .b(FE_OCP_RBN6092_n_5531), .o(n_5700) );
in01s01 g765362 ( .a(n_15569), .o(n_16341) );
na02m06 TIMEBOOST_cell_6809 ( .a(FE_OCP_RBN3287_n_5656), .b(n_4759), .o(TIMEBOOST_net_2162) );
in01s01 g765364 ( .a(n_16253), .o(n_16254) );
oa12s01 g765365 ( .a(n_15867), .b(n_16245), .c(n_15823), .o(n_16253) );
in01s01 g765366 ( .a(n_16304), .o(n_16305) );
oa12s01 g765367 ( .a(n_15784), .b(FE_OCP_RBN6847_n_15599), .c(n_15711), .o(n_16304) );
ao12s01 g765368 ( .a(n_15715), .b(FE_OCP_RBN6847_n_15599), .c(n_14652), .o(n_16546) );
in01s01 g765369 ( .a(n_16249), .o(n_16250) );
ao12s01 g765370 ( .a(n_15829), .b(n_16245), .c(n_15833), .o(n_16249) );
ao12s01 g765371 ( .a(n_15667), .b(FE_OCP_RBN6847_n_15599), .c(n_15786), .o(n_16508) );
ao12s01 g765372 ( .a(n_16135), .b(FE_OCP_RBN3195_n_15599), .c(n_15564), .o(n_16352) );
ao12s01 g765373 ( .a(n_15876), .b(FE_OCP_RBN6847_n_15599), .c(n_15779), .o(n_16572) );
in01s01 g765374 ( .a(n_16302), .o(n_16303) );
ao12s01 g765375 ( .a(n_15920), .b(FE_OCP_RBN6847_n_15599), .c(n_15869), .o(n_16302) );
in01s01 g765376 ( .a(n_16300), .o(n_16301) );
oa12s01 g765377 ( .a(n_15875), .b(FE_OCP_RBN3190_n_15599), .c(n_15958), .o(n_16300) );
no02s01 g765378 ( .a(n_16135), .b(n_15566), .o(n_15633) );
in01s01 g765379 ( .a(n_16016), .o(n_16102) );
ao12s01 g765380 ( .a(FE_OCP_RBN3190_n_15599), .b(n_15958), .c(n_15957), .o(n_16016) );
na02s08 g765381 ( .a(FE_OCP_RBN4324_n_15156), .b(n_14056), .o(n_15410) );
in01s01 g765383 ( .a(n_15578), .o(n_15516) );
na02m01 g765384 ( .a(FE_OCP_RBN6801_n_15156), .b(n_14277), .o(n_15578) );
no02s06 g765385 ( .a(FE_OCP_RBN6801_n_15156), .b(n_14276), .o(n_15810) );
in01s01 g765390 ( .a(n_15023), .o(n_15055) );
ao12f08 g765391 ( .a(n_14789), .b(n_14942), .c(n_14845), .o(n_15023) );
in01s01 g765392 ( .a(n_15371), .o(n_15372) );
no02s02 TIMEBOOST_cell_5070 ( .a(n_13781), .b(n_13690), .o(TIMEBOOST_net_1483) );
in01s02 g765394 ( .a(n_15369), .o(n_15370) );
na02s02 g765395 ( .a(n_15330), .b(n_15252), .o(n_15369) );
oa12s01 g765396 ( .a(n_15141), .b(n_15140), .c(n_15139), .o(n_15221) );
in01s01 g765397 ( .a(n_15449), .o(n_15450) );
no02s01 TIMEBOOST_cell_3062 ( .a(n_7577), .b(n_8742), .o(TIMEBOOST_net_822) );
no02s02 TIMEBOOST_cell_8557 ( .a(TIMEBOOST_net_2765), .b(n_38131), .o(n_38153) );
no02s02 TIMEBOOST_cell_4383 ( .a(n_20062), .b(n_19583), .o(TIMEBOOST_net_1282) );
in01s01 g765401 ( .a(n_15296), .o(n_15412) );
na02f08 g765402 ( .a(n_15177), .b(n_15170), .o(n_15296) );
oa22s01 g765403 ( .a(FE_OCP_RBN3195_n_15599), .b(n_15482), .c(n_16245), .d(n_15513), .o(n_16342) );
in01f02 g765405 ( .a(n_15151), .o(n_15189) );
na02f08 g765406 ( .a(n_15054), .b(n_15050), .o(n_15151) );
oa22s01 g765407 ( .a(FE_OCP_RBN3195_n_15599), .b(n_16246), .c(n_16245), .d(n_14433), .o(n_16349) );
ao22s01 g765408 ( .a(n_16245), .b(n_15788), .c(FE_OCP_RBN3195_n_15599), .d(n_14112), .o(n_16346) );
ao22s01 g765409 ( .a(n_16245), .b(n_14081), .c(FE_OCP_RBN3195_n_15599), .d(n_14044), .o(n_16344) );
oa22s01 g765410 ( .a(FE_OCP_RBN3195_n_15599), .b(n_15631), .c(n_16245), .d(n_14391), .o(n_16355) );
oa22s01 g765411 ( .a(FE_OCP_RBN3195_n_15599), .b(n_16244), .c(n_16245), .d(n_16138), .o(n_16358) );
oa22s02 g765413 ( .a(FE_OCP_RBN5946_n_14982), .b(FE_OCP_RBN1821_n_13858), .c(FE_OCP_RBN5948_n_14982), .d(n_13950), .o(n_15187) );
in01s02 g765414 ( .a(n_15294), .o(n_15295) );
na02m04 g765415 ( .a(n_15181), .b(n_15143), .o(n_15294) );
in01s01 g765416 ( .a(n_15567), .o(n_15568) );
na02s01 g765417 ( .a(n_15402), .b(n_15448), .o(n_15567) );
no02m04 TIMEBOOST_cell_4382 ( .a(TIMEBOOST_net_1281), .b(n_26233), .o(n_26313) );
no02m04 g765477 ( .a(n_15042), .b(n_15097), .o(n_15149) );
no02s06 g765478 ( .a(n_15053), .b(n_15017), .o(n_15054) );
na02m04 g765480 ( .a(n_15077), .b(FE_OCP_RBN2834_n_13962), .o(n_15195) );
no02f04 g765482 ( .a(n_15077), .b(FE_OCP_RBN2834_n_13962), .o(n_15110) );
in01f02 g765483 ( .a(n_15108), .o(n_15109) );
no02s02 TIMEBOOST_cell_4271 ( .a(n_44866), .b(n_37901), .o(TIMEBOOST_net_1226) );
na02f06 g765485 ( .a(n_15018), .b(n_14989), .o(n_15050) );
na02f02 g765486 ( .a(n_14985), .b(FE_OCPN1703_n_14210), .o(n_15022) );
in01s01 g765487 ( .a(n_16173), .o(n_16174) );
no02s01 g765488 ( .a(FE_OCP_RBN3190_n_15599), .b(n_15957), .o(n_16173) );
in01s01 g765489 ( .a(n_15920), .o(n_15921) );
no02s01 g765490 ( .a(FE_OCP_RBN6828_n_15514), .b(n_15869), .o(n_15920) );
no02s02 g765491 ( .a(n_15514), .b(n_15513), .o(n_15515) );
na02s01 g765492 ( .a(FE_OCP_RBN6846_n_15599), .b(n_15665), .o(n_15969) );
na02s01 g765493 ( .a(n_15719), .b(n_15957), .o(n_16255) );
no02s01 g765494 ( .a(FE_OCP_RBN6846_n_15599), .b(n_15833), .o(n_15829) );
in01s01 g765495 ( .a(n_15781), .o(n_15925) );
no02s01 g765496 ( .a(n_15664), .b(n_15747), .o(n_15781) );
in01s01 g765497 ( .a(n_15867), .o(n_15868) );
na02s01 g765498 ( .a(n_15664), .b(n_15823), .o(n_15867) );
na02s01 g765499 ( .a(n_15719), .b(n_15958), .o(n_15875) );
in01s01 g765500 ( .a(n_15928), .o(n_15822) );
no02s01 g765501 ( .a(FE_OCP_RBN6829_n_15514), .b(n_15712), .o(n_15928) );
na02s01 g765502 ( .a(FE_OCP_RBN3185_n_15599), .b(n_15669), .o(n_15783) );
no02s01 g765503 ( .a(n_15565), .b(n_15631), .o(n_15566) );
no02s01 g765504 ( .a(n_15719), .b(n_15779), .o(n_15876) );
in01s01 g765505 ( .a(n_15826), .o(n_15778) );
no02s01 g765506 ( .a(FE_OCP_RBN6846_n_15599), .b(n_15087), .o(n_15826) );
in01s01 g765507 ( .a(n_15837), .o(n_15745) );
na02s01 g765508 ( .a(n_15719), .b(n_15718), .o(n_15837) );
na02s01 g765509 ( .a(FE_OCP_RBN6053_n_15514), .b(n_15631), .o(n_15632) );
na02s02 TIMEBOOST_cell_6893 ( .a(n_37671), .b(n_37692), .o(TIMEBOOST_net_2205) );
in01s01 g765511 ( .a(n_15749), .o(n_15717) );
na02s01 g765512 ( .a(FE_OCP_RBN3185_n_15599), .b(n_15663), .o(n_15749) );
in01s01 g765513 ( .a(n_15787), .o(n_15716) );
no02s01 g765514 ( .a(n_15514), .b(n_15669), .o(n_15787) );
no02s01 g765515 ( .a(n_15565), .b(n_15564), .o(n_16135) );
no02s01 g765516 ( .a(n_15565), .b(n_16246), .o(n_15563) );
in01s01 g765517 ( .a(n_15667), .o(n_15668) );
no02s01 g765518 ( .a(n_15565), .b(n_15786), .o(n_15667) );
in01s01 g765519 ( .a(n_15714), .o(n_15715) );
na02s01 g765520 ( .a(FE_OCP_RBN3185_n_15599), .b(n_15666), .o(n_15714) );
in01s01 g765521 ( .a(n_15924), .o(n_15866) );
na02s01 g765522 ( .a(n_15664), .b(n_15747), .o(n_15924) );
na02s01 g765523 ( .a(n_15565), .b(n_15865), .o(n_16018) );
in01s01 g765524 ( .a(n_15967), .o(n_15919) );
no02s01 g765525 ( .a(FE_OCP_RBN6847_n_15599), .b(n_15865), .o(n_15967) );
no02s01 g765526 ( .a(FE_OCP_RBN6829_n_15514), .b(n_15086), .o(n_15834) );
na02s01 g765527 ( .a(FE_OCP_RBN6829_n_15514), .b(n_15712), .o(n_15922) );
na02s01 g765528 ( .a(n_15719), .b(n_15711), .o(n_15784) );
in01s01 g765529 ( .a(n_15873), .o(n_15821) );
no02s01 g765530 ( .a(FE_OCP_RBN6053_n_15514), .b(n_15718), .o(n_15873) );
in01s01 g765531 ( .a(n_15839), .o(n_15710) );
no02s01 g765532 ( .a(n_15664), .b(n_15665), .o(n_15839) );
in01s01 g765533 ( .a(n_15709), .o(n_15830) );
no02s01 g765534 ( .a(n_15664), .b(n_15663), .o(n_15709) );
na02m02 g765535 ( .a(n_15014), .b(n_14986), .o(n_15076) );
no02m02 g765536 ( .a(n_15012), .b(n_14987), .o(n_15075) );
no02f02 g765537 ( .a(FE_OCP_RBN2056_n_13784), .b(n_14982), .o(n_15112) );
no02m02 g765538 ( .a(n_14983), .b(FE_OCP_RBN2057_n_13784), .o(n_15049) );
no02m06 g765539 ( .a(FE_OCP_RBN5946_n_14982), .b(FE_OCP_RBN2058_n_13784), .o(n_15391) );
in01s02 g765542 ( .a(n_46419), .o(n_15219) );
in01s01 g765547 ( .a(n_15144), .o(n_15182) );
no02s06 g765549 ( .a(FE_OCP_RBN3032_n_15150), .b(FE_OCPN1244_n_13992), .o(n_15144) );
na02s01 g765550 ( .a(n_15103), .b(FE_OCP_RBN5728_n_14120), .o(n_15181) );
na02s02 g765551 ( .a(n_15142), .b(FE_OCP_RBN2073_n_14120), .o(n_15143) );
in01s01 g765555 ( .a(n_15180), .o(n_15218) );
no02m03 g765556 ( .a(FE_OCP_RBN5947_n_14982), .b(FE_OCP_RBN2068_n_14069), .o(n_15180) );
in01s01 g765558 ( .a(n_15258), .o(n_15178) );
in01s02 g765559 ( .a(n_15127), .o(n_15258) );
no02s02 g765560 ( .a(FE_OCP_RBN2069_n_14069), .b(FE_OCP_RBN3032_n_15150), .o(n_15127) );
no02s02 TIMEBOOST_cell_3063 ( .a(TIMEBOOST_net_822), .b(n_8747), .o(n_8788) );
no02s06 g765564 ( .a(n_15142), .b(FE_OCPN4857_n_14317), .o(n_15806) );
na02s06 TIMEBOOST_cell_4387 ( .a(n_20311), .b(FE_RN_109_0), .o(TIMEBOOST_net_1284) );
in01s01 g765567 ( .a(n_15293), .o(n_15373) );
no02m01 g765568 ( .a(n_15103), .b(n_14396), .o(n_15293) );
na02s01 g765569 ( .a(n_15103), .b(n_15250), .o(n_15252) );
na02s01 g765570 ( .a(n_15142), .b(n_14364), .o(n_15330) );
na02s01 g765571 ( .a(n_15140), .b(n_15139), .o(n_15141) );
no02s01 TIMEBOOST_cell_4029 ( .a(n_30790), .b(FE_OCPN5130_FE_OFN1198_n_27014), .o(TIMEBOOST_net_1105) );
na02s01 g765573 ( .a(n_15142), .b(n_14821), .o(n_15403) );
na02s01 g765574 ( .a(n_15103), .b(FE_OCP_RBN5759_n_14444), .o(n_15402) );
na02s01 g765575 ( .a(n_15142), .b(FE_OCP_RBN5758_n_14444), .o(n_15448) );
no02s01 g765576 ( .a(n_45523), .b(n_15137), .o(n_15226) );
no02s01 g765577 ( .a(n_15171), .b(n_15133), .o(n_15332) );
na02f06 g765578 ( .a(n_15132), .b(n_15091), .o(n_15177) );
no02s20 TIMEBOOST_cell_6881 ( .a(n_32818), .b(n_32820), .o(TIMEBOOST_net_2199) );
oa12s01 g765580 ( .a(n_14488), .b(n_15446), .c(n_14456), .o(n_15521) );
oa12s01 g765581 ( .a(n_14526), .b(n_15481), .c(n_14528), .o(n_15576) );
ao12s01 g765582 ( .a(n_14426), .b(n_15481), .c(n_14388), .o(n_15573) );
in01f02 g765584 ( .a(n_15136), .o(n_15175) );
na02f04 g765585 ( .a(n_15044), .b(n_15045), .o(n_15136) );
in01s01 g765586 ( .a(n_16136), .o(n_15744) );
na02s01 g765587 ( .a(FE_OCP_RBN6053_n_15514), .b(n_14434), .o(n_16136) );
ao12s01 g765588 ( .a(FE_OCP_RBN6847_n_15599), .b(n_15085), .c(n_15865), .o(n_16059) );
in01s01 g765589 ( .a(n_15748), .o(n_15512) );
na02s01 g765590 ( .a(n_15366), .b(n_15397), .o(n_15748) );
no02s06 TIMEBOOST_cell_6954 ( .a(TIMEBOOST_net_2235), .b(n_8315), .o(n_8445) );
in01f02 g765610 ( .a(n_15021), .o(n_15156) );
in01s04 g765611 ( .a(n_15048), .o(n_15194) );
in01m06 g765616 ( .a(n_15021), .o(n_15048) );
no02s06 g765619 ( .a(FE_OCP_RBN3032_n_15150), .b(n_14192), .o(n_15099) );
ao12s01 g765626 ( .a(n_15443), .b(n_15481), .c(n_15442), .o(n_15961) );
in01m02 g765628 ( .a(n_14944), .o(n_14964) );
oa12f08 g765629 ( .a(n_14851), .b(n_14830), .c(n_14794), .o(n_14944) );
na02m06 TIMEBOOST_cell_5141 ( .a(TIMEBOOST_net_1518), .b(n_9254), .o(n_9450) );
ao12f04 g765633 ( .a(n_15070), .b(n_15003), .c(n_14916), .o(n_15225) );
ao12s01 g765634 ( .a(n_15399), .b(n_15446), .c(n_15398), .o(n_15870) );
no02s01 g765636 ( .a(n_15446), .b(n_15398), .o(n_15399) );
no02s01 g765637 ( .a(n_15481), .b(n_15442), .o(n_15443) );
na02f08 TIMEBOOST_cell_7555 ( .a(TIMEBOOST_net_2408), .b(n_13859), .o(n_14059) );
na02s01 g765639 ( .a(n_15324), .b(n_14424), .o(n_15366) );
na02f02 g765641 ( .a(n_15019), .b(n_15043), .o(n_15044) );
in01s02 g765642 ( .a(n_15041), .o(n_15042) );
no02m02 g765643 ( .a(n_15019), .b(n_47262), .o(n_15041) );
na02f02 g765644 ( .a(n_15005), .b(n_14920), .o(n_15040) );
na02s01 g765645 ( .a(n_15325), .b(n_14423), .o(n_15397) );
in01s02 g765646 ( .a(n_15038), .o(n_15039) );
no02f06 g765647 ( .a(n_15018), .b(n_15017), .o(n_15038) );
no02s08 g765648 ( .a(n_14988), .b(FE_OCP_RBN4234_n_13962), .o(n_15053) );
na02s04 g765650 ( .a(n_14911), .b(FE_OCP_RBN5790_n_13962), .o(n_14943) );
no02s06 TIMEBOOST_cell_4270 ( .a(TIMEBOOST_net_1225), .b(n_33804), .o(n_33937) );
na02s02 g765652 ( .a(n_14988), .b(FE_OCP_RBN4234_n_13962), .o(n_14989) );
in01m02 g765653 ( .a(n_15097), .o(n_15098) );
na02f04 g765654 ( .a(n_15008), .b(n_15043), .o(n_15097) );
no02s06 TIMEBOOST_cell_6953 ( .a(FE_OCP_RBN6645_n_8342), .b(FE_OCP_RBN2739_n_8300), .o(TIMEBOOST_net_2235) );
na02f04 g765657 ( .a(n_15009), .b(n_14923), .o(n_15037) );
in01s01 g765659 ( .a(n_14987), .o(n_15014) );
no02f04 g765660 ( .a(n_14962), .b(FE_OCP_RBN2644_n_13667), .o(n_14987) );
in01s01 g765662 ( .a(n_14986), .o(n_15012) );
na02f04 g765663 ( .a(n_14962), .b(FE_OCP_RBN2644_n_13667), .o(n_14986) );
na02f02 g765666 ( .a(n_15036), .b(n_15035), .o(n_15071) );
in01s01 g765667 ( .a(n_15170), .o(n_15171) );
na02m06 g765668 ( .a(n_15067), .b(n_13479), .o(n_15170) );
no02s01 g765669 ( .a(n_15004), .b(n_15070), .o(n_15140) );
in01s01 g765670 ( .a(n_15132), .o(n_15133) );
na02f04 g765671 ( .a(n_15066), .b(n_13478), .o(n_15132) );
in01s02 g765676 ( .a(n_15664), .o(n_15719) );
in01s02 g765677 ( .a(n_15565), .o(n_15664) );
in01s01 g765685 ( .a(FE_OCP_RBN6847_n_15599), .o(n_16245) );
in01s03 g765690 ( .a(FE_OCP_RBN3196_n_15599), .o(n_17336) );
in01s02 g765697 ( .a(FE_OCP_RBN3196_n_15599), .o(n_17584) );
in01s03 g765706 ( .a(FE_OCP_RBN3193_n_15599), .o(n_16339) );
in01s03 g765711 ( .a(FE_OCP_RBN3193_n_15599), .o(n_17753) );
in01s02 g765737 ( .a(n_15514), .o(n_15565) );
in01s06 g765738 ( .a(n_15441), .o(n_15514) );
in01m04 g765739 ( .a(n_15396), .o(n_15441) );
oa12m04 g765740 ( .a(n_14619), .b(n_15287), .c(n_14563), .o(n_15396) );
in01s02 g765744 ( .a(n_14959), .o(n_14960) );
in01s01 g765745 ( .a(n_14942), .o(n_14959) );
oa12f08 g765746 ( .a(n_14718), .b(n_14862), .c(n_14717), .o(n_14942) );
in01s01 g765747 ( .a(n_14982), .o(n_14983) );
in01s08 g765762 ( .a(n_15103), .o(n_15142) );
in01m06 g765763 ( .a(FE_OCP_RBN5947_n_14982), .o(n_15103) );
no03s04 TIMEBOOST_cell_8272 ( .a(n_8069), .b(n_8002), .c(n_8022), .o(n_8175) );
oa12s01 g765774 ( .a(n_15094), .b(n_15093), .c(n_15092), .o(n_15168) );
ao12s01 g765775 ( .a(n_15363), .b(n_15362), .c(n_15361), .o(n_15958) );
in01s06 g765776 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_1_), .o(n_17193) );
no02s01 g765778 ( .a(n_15362), .b(n_15361), .o(n_15363) );
no02s01 g765779 ( .a(n_15288), .b(n_14490), .o(n_15481) );
no02f02 g765780 ( .a(n_14958), .b(n_14903), .o(n_15019) );
in01m02 g765781 ( .a(n_15009), .o(n_15010) );
na02s06 TIMEBOOST_cell_6870 ( .a(TIMEBOOST_net_581), .b(TIMEBOOST_net_2193), .o(n_32583) );
na02s02 TIMEBOOST_cell_5646 ( .a(n_6238), .b(n_6170), .o(TIMEBOOST_net_1771) );
na02f02 g765785 ( .a(n_14950), .b(FE_OCPN1703_n_14210), .o(n_15008) );
in01s02 g765786 ( .a(n_15005), .o(n_15006) );
no02f02 g765787 ( .a(n_47262), .b(n_14958), .o(n_15005) );
na02f04 g765788 ( .a(n_14979), .b(FE_OCP_RBN5796_n_13962), .o(n_15043) );
no02f08 g765790 ( .a(n_14923), .b(n_14956), .o(n_15018) );
in01s01 g765791 ( .a(n_15003), .o(n_15004) );
na02f04 g765792 ( .a(n_14978), .b(FE_OCPN5264_n_14977), .o(n_15003) );
na02m06 g765794 ( .a(n_14921), .b(FE_OCP_RBN5021_n_13726), .o(n_15035) );
no02f04 g765795 ( .a(n_14978), .b(FE_OCPN5264_n_14977), .o(n_15070) );
na02s01 g765796 ( .a(n_15093), .b(n_15092), .o(n_15094) );
na02f02 g765797 ( .a(FE_OCP_RBN2091_n_14909), .b(n_14908), .o(n_14976) );
no02f02 g765798 ( .a(FE_OCP_RBN2090_n_14908), .b(n_14909), .o(n_14975) );
oa12s01 g765799 ( .a(n_14353), .b(n_15289), .c(n_14491), .o(n_15446) );
in01m04 g765800 ( .a(n_14912), .o(n_14913) );
oa12f08 g765801 ( .a(n_14646), .b(n_14891), .c(n_14647), .o(n_14912) );
in01s01 g765802 ( .a(n_15324), .o(n_15325) );
oa12s01 g765803 ( .a(n_14390), .b(n_15290), .c(n_14345), .o(n_15324) );
in01m02 g765806 ( .a(n_14889), .o(n_14890) );
in01m01 g765807 ( .a(n_14830), .o(n_14889) );
ao12s06 g765808 ( .a(n_14697), .b(n_14775), .c(n_14754), .o(n_14830) );
oa12s01 g765810 ( .a(n_14973), .b(n_14972), .c(n_14971), .o(n_15033) );
in01m02 g765811 ( .a(n_15066), .o(n_15067) );
no02s01 TIMEBOOST_cell_5352 ( .a(n_3786), .b(n_3727), .o(TIMEBOOST_net_1624) );
in01s01 g765813 ( .a(n_15091), .o(n_15331) );
oa12f04 g765814 ( .a(n_14970), .b(n_14969), .c(n_15032), .o(n_15091) );
in01f02 g765819 ( .a(n_14988), .o(n_14955) );
no02s01 TIMEBOOST_cell_7430 ( .a(n_6752), .b(n_6609), .o(TIMEBOOST_net_2346) );
oa12s01 g765821 ( .a(n_15248), .b(n_15290), .c(n_15247), .o(n_15665) );
na02s01 g765822 ( .a(n_15289), .b(n_14561), .o(n_15362) );
na02f02 g765823 ( .a(n_14917), .b(n_14808), .o(n_14954) );
no02s01 TIMEBOOST_cell_8556 ( .a(FE_OCP_RBN4060_n_44875), .b(n_37653), .o(TIMEBOOST_net_2765) );
no02f02 g765827 ( .a(FE_OCP_RBN5791_n_13962), .b(n_14873), .o(n_14958) );
no02s06 g765828 ( .a(n_14872), .b(FE_OCP_RBN4210_n_13796), .o(n_14956) );
no02s06 g765830 ( .a(n_14932), .b(FE_OCP_RBN4229_n_13962), .o(n_15017) );
no02s04 g765831 ( .a(n_14823), .b(FE_OCP_RBN4209_n_13796), .o(n_14864) );
na02s02 TIMEBOOST_cell_5261 ( .a(TIMEBOOST_net_1578), .b(FE_OCP_RBN5958_n_4165), .o(n_4391) );
na02s01 g765833 ( .a(n_15290), .b(n_15247), .o(n_15248) );
no02f06 g765836 ( .a(n_14865), .b(FE_OCP_RBN4152_n_13616), .o(n_14909) );
na02s01 g765837 ( .a(n_14972), .b(n_14971), .o(n_14973) );
na02f01 g765838 ( .a(n_14927), .b(n_14899), .o(n_14928) );
no02f01 g765839 ( .a(n_14878), .b(n_14877), .o(n_14953) );
na02f06 g765842 ( .a(n_14865), .b(FE_OCP_RBN4152_n_13616), .o(n_14908) );
na02f02 g765843 ( .a(n_14906), .b(n_14875), .o(n_14907) );
no02f02 g765844 ( .a(n_14853), .b(n_14854), .o(n_14924) );
in01s01 g765845 ( .a(n_15287), .o(n_15288) );
na02m04 g765846 ( .a(n_15212), .b(n_14492), .o(n_15287) );
in01m04 g765847 ( .a(n_14886), .o(n_14887) );
no02s04 TIMEBOOST_cell_6653 ( .a(TIMEBOOST_net_1877), .b(n_14144), .o(TIMEBOOST_net_2084) );
no02f08 g765851 ( .a(n_14857), .b(n_14860), .o(n_14923) );
no02s02 TIMEBOOST_cell_3164 ( .a(n_30246), .b(n_30296), .o(TIMEBOOST_net_873) );
in01s02 g765856 ( .a(n_14884), .o(n_14885) );
in01s01 g765857 ( .a(n_14862), .o(n_14884) );
ao12f08 g765858 ( .a(n_14662), .b(n_14771), .c(n_14719), .o(n_14862) );
no02f06 g765860 ( .a(n_14827), .b(n_14861), .o(n_14921) );
in01m02 g765861 ( .a(n_14979), .o(n_14950) );
na02s01 TIMEBOOST_cell_5316 ( .a(n_43106), .b(FE_OCP_RBN3306_n_43022), .o(TIMEBOOST_net_1606) );
oa12s01 g765863 ( .a(n_14967), .b(n_15032), .c(n_14966), .o(n_15093) );
in01s01 g765864 ( .a(n_15711), .o(n_15360) );
ao12s01 g765865 ( .a(n_15246), .b(n_15245), .c(n_15244), .o(n_15711) );
ao12s01 g765866 ( .a(n_15211), .b(n_15210), .c(n_15209), .o(n_15957) );
oa12s01 g765867 ( .a(n_15000), .b(n_14999), .c(n_14998), .o(n_15065) );
no02s04 g765868 ( .a(n_14792), .b(n_14225), .o(n_14827) );
no02f04 g765869 ( .a(n_14793), .b(n_14265), .o(n_14861) );
in01s01 g765870 ( .a(n_15212), .o(n_15289) );
no02m04 g765871 ( .a(n_15128), .b(n_14486), .o(n_15212) );
no02s01 g765872 ( .a(n_15210), .b(n_15209), .o(n_15211) );
na02s04 g765873 ( .a(n_14796), .b(n_14859), .o(n_14860) );
no03s02 TIMEBOOST_cell_8528 ( .a(n_2449), .b(n_2448), .c(n_2390), .o(TIMEBOOST_net_2751) );
na02m04 g765876 ( .a(n_14856), .b(n_14859), .o(n_14881) );
in01f02 g765877 ( .a(n_14919), .o(n_14920) );
in01f02 g765878 ( .a(n_14903), .o(n_14919) );
na02m04 g765879 ( .a(n_14880), .b(n_14808), .o(n_14903) );
no02f02 g765880 ( .a(n_14818), .b(n_14801), .o(n_14858) );
in01f02 g765882 ( .a(n_14901), .o(n_14902) );
in01s01 TIMEBOOST_cell_8909 ( .a(TIMEBOOST_net_2952), .o(TIMEBOOST_net_2953) );
in01s01 TIMEBOOST_cell_8906 ( .a(n_1334), .o(TIMEBOOST_net_2950) );
no02f02 g765885 ( .a(n_14814), .b(n_14215), .o(n_14855) );
no02s01 g765886 ( .a(n_15245), .b(n_15244), .o(n_15246) );
in01f01 g765887 ( .a(n_14927), .o(n_14878) );
na02f04 g765888 ( .a(n_14829), .b(n_13659), .o(n_14927) );
in01m01 g765890 ( .a(n_14877), .o(n_14899) );
no02m04 g765891 ( .a(n_14829), .b(n_13659), .o(n_14877) );
na02s04 g765892 ( .a(n_15092), .b(n_14968), .o(n_14970) );
no02f02 g765893 ( .a(n_15092), .b(n_14968), .o(n_14969) );
na02s01 g765894 ( .a(n_14999), .b(n_14998), .o(n_15000) );
na02s01 g765895 ( .a(n_15032), .b(n_14966), .o(n_14967) );
in01m01 g765897 ( .a(n_14854), .o(n_14875) );
no02f06 g765898 ( .a(n_14826), .b(FE_OCPN4937_n_13570), .o(n_14854) );
in01m01 g765899 ( .a(n_14906), .o(n_14853) );
na02f06 g765900 ( .a(n_14826), .b(FE_OCPN4937_n_13570), .o(n_14906) );
na02s02 g765901 ( .a(n_14815), .b(n_14851), .o(n_14852) );
no02f02 g765902 ( .a(n_14795), .b(n_14816), .o(n_14874) );
no02s04 TIMEBOOST_cell_2097 ( .a(n_20616), .b(n_20338), .o(TIMEBOOST_net_663) );
in01m01 g765904 ( .a(n_14891), .o(n_14824) );
no02s06 TIMEBOOST_cell_2093 ( .a(n_26318), .b(n_23564), .o(TIMEBOOST_net_661) );
in01s02 g765906 ( .a(n_14917), .o(n_14918) );
no02s02 TIMEBOOST_cell_3058 ( .a(n_38182), .b(n_38218), .o(TIMEBOOST_net_820) );
oa12s01 g765908 ( .a(n_14348), .b(n_15088), .c(n_14389), .o(n_15290) );
in01s01 g765912 ( .a(n_14916), .o(n_15139) );
oa12f04 g765913 ( .a(n_14744), .b(n_14898), .c(n_14743), .o(n_14916) );
oa12s01 g765914 ( .a(n_14870), .b(n_14898), .c(n_14869), .o(n_14972) );
in01f02 g765915 ( .a(n_14873), .o(n_14935) );
in01f02 g765917 ( .a(n_14872), .o(n_14932) );
in01m02 g765920 ( .a(n_14802), .o(n_14803) );
in01m02 g765921 ( .a(n_14775), .o(n_14802) );
oa12m06 g765922 ( .a(n_14664), .b(n_14696), .c(n_14611), .o(n_14775) );
no02s01 g765924 ( .a(n_15089), .b(n_14347), .o(n_15245) );
no02m08 TIMEBOOST_cell_3057 ( .a(n_24802), .b(TIMEBOOST_net_819), .o(n_24823) );
na02s06 g765926 ( .a(n_14785), .b(FE_OCP_RBN5795_n_13962), .o(n_14880) );
in01s02 g765927 ( .a(n_14818), .o(n_14819) );
no02s01 TIMEBOOST_cell_4303 ( .a(n_24620), .b(FE_OCPN1920_n_22393), .o(TIMEBOOST_net_1242) );
no02f08 TIMEBOOST_cell_7585 ( .a(TIMEBOOST_net_2423), .b(n_24464), .o(n_24614) );
na03s03 TIMEBOOST_cell_8179 ( .a(n_1393), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_1_), .c(n_1452), .o(TIMEBOOST_net_2336) );
na02m02 g765931 ( .a(n_14798), .b(FE_OCP_RBN4198_n_13796), .o(n_14799) );
na02s04 g765932 ( .a(n_14798), .b(FE_OCP_RBN4206_n_13796), .o(n_14796) );
na02s02 g765933 ( .a(n_14811), .b(n_14845), .o(n_14846) );
no02f02 g765934 ( .a(n_14812), .b(n_14788), .o(n_14871) );
na02s01 g765935 ( .a(n_14898), .b(n_14869), .o(n_14870) );
in01m01 g765936 ( .a(n_14851), .o(n_14795) );
na02f08 g765937 ( .a(n_14774), .b(FE_OCP_RBN4120_n_13483), .o(n_14851) );
in01f02 g765938 ( .a(n_14815), .o(n_14816) );
in01m02 g765939 ( .a(n_14794), .o(n_14815) );
no02f08 g765940 ( .a(n_14774), .b(FE_OCP_RBN2602_n_13483), .o(n_14794) );
na02f02 g765941 ( .a(n_14754), .b(FE_OCP_RBN4249_n_14697), .o(n_14755) );
no02f02 g765942 ( .a(n_14697), .b(n_14698), .o(n_14773) );
in01m02 g765943 ( .a(n_14792), .o(n_14793) );
in01m04 g765944 ( .a(n_14772), .o(n_14792) );
oa12m08 g765945 ( .a(n_14656), .b(n_14750), .c(n_14626), .o(n_14772) );
no03s10 TIMEBOOST_cell_2221 ( .a(n_40749), .b(n_40750), .c(n_40738), .o(n_40751) );
in01s01 g765947 ( .a(n_15128), .o(n_15210) );
ao12m04 g765948 ( .a(n_14431), .b(n_15090), .c(n_14430), .o(n_15128) );
in01m02 g765952 ( .a(n_14790), .o(n_14791) );
in01m01 g765953 ( .a(n_14771), .o(n_14790) );
oa12f08 g765954 ( .a(n_14573), .b(n_14673), .c(n_14572), .o(n_14771) );
na02s01 TIMEBOOST_cell_6190 ( .a(TIMEBOOST_net_1946), .b(n_16018), .o(n_15930) );
oa12f04 g765956 ( .a(n_14734), .b(n_14915), .c(n_14735), .o(n_15092) );
oa22f02 g765957 ( .a(n_14842), .b(n_14738), .c(n_14841), .d(n_14706), .o(n_15032) );
ao12s01 g765958 ( .a(n_15064), .b(n_15090), .c(n_15063), .o(n_15712) );
oa12s01 g765959 ( .a(n_14897), .b(n_14915), .c(n_14896), .o(n_14999) );
na02f06 g765960 ( .a(n_14699), .b(n_14727), .o(n_14826) );
na02f04 g765962 ( .a(n_14670), .b(n_14633), .o(n_14727) );
na02s03 g765963 ( .a(n_14669), .b(n_14632), .o(n_14699) );
na02s01 TIMEBOOST_cell_6189 ( .a(n_15823), .b(n_15719), .o(TIMEBOOST_net_1946) );
na02m04 g765965 ( .a(n_14750), .b(n_14679), .o(n_14751) );
no02s01 TIMEBOOST_cell_6823 ( .a(n_43351), .b(FE_RN_1620_0), .o(TIMEBOOST_net_2169) );
na02s02 g765967 ( .a(n_45520), .b(FE_OCP_RBN4198_n_13796), .o(n_14859) );
in01s01 g765968 ( .a(n_15088), .o(n_15089) );
na02s01 g765969 ( .a(n_15090), .b(n_14385), .o(n_15088) );
no02s01 g765972 ( .a(n_15090), .b(n_15063), .o(n_15064) );
in01m01 g765973 ( .a(n_14811), .o(n_14812) );
in01f01 g765974 ( .a(n_14789), .o(n_14811) );
no02m06 g765975 ( .a(n_14770), .b(FE_OCPN6279_FE_OCP_RBN1594_n_13557), .o(n_14789) );
in01s01 g765976 ( .a(n_14845), .o(n_14788) );
na02s06 g765977 ( .a(n_14770), .b(FE_OCPN6279_FE_OCP_RBN1594_n_13557), .o(n_14845) );
in01f01 g765978 ( .a(n_14754), .o(n_14698) );
na02s01 g765980 ( .a(n_14915), .b(n_14896), .o(n_14897) );
in01f02 g765985 ( .a(n_14696), .o(n_14722) );
oa12f06 g765986 ( .a(n_14636), .b(n_14451), .c(n_14584), .o(n_14696) );
in01f04 g765987 ( .a(n_14746), .o(n_14747) );
in01m04 g765988 ( .a(n_14721), .o(n_14746) );
na02s01 TIMEBOOST_cell_4243 ( .a(n_18915), .b(n_18914), .o(TIMEBOOST_net_1212) );
no02f04 g765990 ( .a(n_14761), .b(n_14745), .o(n_14898) );
na02f04 g765994 ( .a(n_14666), .b(n_14694), .o(n_14768) );
in01f01 g765995 ( .a(n_14809), .o(n_14810) );
oa22f01 g765996 ( .a(n_14716), .b(n_13563), .c(n_14707), .d(n_13562), .o(n_14809) );
in01s01 g765997 ( .a(n_15086), .o(n_15087) );
ao12s01 g765998 ( .a(n_14997), .b(n_14996), .c(n_14995), .o(n_15086) );
in01f02 g765999 ( .a(n_14785), .o(n_14786) );
in01f02 g766001 ( .a(n_14798), .o(n_14764) );
na02s01 TIMEBOOST_cell_5260 ( .a(n_4134), .b(n_4133), .o(TIMEBOOST_net_1578) );
oa12s01 g766007 ( .a(n_15031), .b(n_15030), .c(n_15029), .o(n_15833) );
no02m02 TIMEBOOST_cell_2906 ( .a(n_18377), .b(n_18200), .o(TIMEBOOST_net_744) );
na03f04 TIMEBOOST_cell_8417 ( .a(n_10795), .b(n_10773), .c(n_10847), .o(n_10950) );
in01s02 g766010 ( .a(n_14669), .o(n_14670) );
na02f04 g766011 ( .a(n_14616), .b(n_14634), .o(n_14669) );
na02s02 TIMEBOOST_cell_2905 ( .a(TIMEBOOST_net_743), .b(n_29018), .o(n_29064) );
na02m02 TIMEBOOST_cell_8496 ( .a(FE_RN_1584_0), .b(n_12542), .o(TIMEBOOST_net_2735) );
no02m02 g766014 ( .a(n_14709), .b(n_47256), .o(n_14745) );
no02f04 g766015 ( .a(n_14575), .b(n_14710), .o(n_14761) );
na02s01 g766016 ( .a(n_15030), .b(n_15029), .o(n_15031) );
in01s01 g766018 ( .a(n_14808), .o(n_14843) );
no02m06 g766019 ( .a(n_14782), .b(n_14706), .o(n_14808) );
na02s04 g766020 ( .a(n_14638), .b(FE_OCP_RBN4206_n_13796), .o(n_14667) );
no02f08 TIMEBOOST_cell_5259 ( .a(TIMEBOOST_net_1577), .b(n_39063), .o(n_39109) );
no02s01 g766022 ( .a(n_14996), .b(n_14995), .o(n_14997) );
na02f04 g766023 ( .a(n_14971), .b(FE_OCPN1398_n_14742), .o(n_14744) );
no02f04 g766024 ( .a(n_14971), .b(n_14742), .o(n_14743) );
na02f04 g766025 ( .a(n_14642), .b(n_14601), .o(n_14666) );
na02f02 g766026 ( .a(n_14600), .b(n_14643), .o(n_14694) );
na02f01 g766027 ( .a(n_14687), .b(n_14719), .o(n_14720) );
no02m01 g766028 ( .a(n_14662), .b(n_14661), .o(n_14741) );
na02s06 g766029 ( .a(n_14716), .b(n_13563), .o(n_14718) );
no02s06 g766030 ( .a(n_14716), .b(n_13563), .o(n_14717) );
na02f02 g766031 ( .a(FE_OCP_RBN2083_n_14611), .b(n_14664), .o(n_14665) );
no02f02 g766032 ( .a(FE_OCP_RBN1834_n_14664), .b(n_14611), .o(n_14693) );
na02m08 g766034 ( .a(n_14615), .b(n_14472), .o(n_14750) );
in01f02 g766035 ( .a(n_14841), .o(n_14842) );
no02f02 g766036 ( .a(n_14782), .b(n_14759), .o(n_14841) );
na02f04 g766037 ( .a(n_14760), .b(n_14781), .o(n_14915) );
in01s02 g766038 ( .a(n_14714), .o(n_14715) );
in01f01 g766039 ( .a(n_14673), .o(n_14714) );
oa12s01 g766041 ( .a(n_14686), .b(n_14689), .c(n_14685), .o(n_14740) );
no02s03 TIMEBOOST_cell_3026 ( .a(n_8173), .b(n_8200), .o(TIMEBOOST_net_804) );
in01s01 g766043 ( .a(n_15823), .o(n_15085) );
ao12s01 g766044 ( .a(n_14994), .b(n_14993), .c(n_14992), .o(n_15823) );
no02s06 TIMEBOOST_cell_8784 ( .a(n_3106), .b(FE_OCP_RBN5940_n_4238), .o(TIMEBOOST_net_2879) );
no02f06 TIMEBOOST_cell_4306 ( .a(TIMEBOOST_net_1243), .b(n_20065), .o(n_20164) );
na02m04 TIMEBOOST_cell_4153 ( .a(n_17005), .b(n_16904), .o(TIMEBOOST_net_1167) );
na02m06 g766053 ( .a(n_14582), .b(n_14473), .o(n_14615) );
in01f02 g766054 ( .a(n_14613), .o(n_14614) );
na02f04 g766055 ( .a(n_14516), .b(n_14503), .o(n_14613) );
no02f06 g766056 ( .a(n_14645), .b(n_14376), .o(n_14647) );
na02m06 g766057 ( .a(n_14645), .b(n_14376), .o(n_14646) );
na02f02 g766058 ( .a(n_14736), .b(n_14681), .o(n_14760) );
na02f04 g766059 ( .a(n_14737), .b(n_14569), .o(n_14781) );
na02s01 TIMEBOOST_cell_4985 ( .a(TIMEBOOST_net_1440), .b(n_37855), .o(TIMEBOOST_net_1030) );
in01s02 g766061 ( .a(n_14801), .o(n_14711) );
in01s01 TIMEBOOST_cell_8889 ( .a(TIMEBOOST_net_2932), .o(TIMEBOOST_net_2933) );
no02f02 g766064 ( .a(FE_OCP_RBN6785_n_14704), .b(FE_OCP_RBN6696_n_13796), .o(n_14759) );
no02m06 g766065 ( .a(n_14704), .b(FE_OCP_RBN2830_n_13962), .o(n_14782) );
na02s04 g766066 ( .a(n_14554), .b(FE_OCP_RBN2762_n_13796), .o(n_14586) );
no02s01 g766067 ( .a(n_14993), .b(n_14992), .o(n_14994) );
no02f06 g766068 ( .a(n_14689), .b(FE_OCPN5136_n_12795), .o(n_14971) );
in01f01 g766069 ( .a(n_14642), .o(n_14643) );
na02f01 g766070 ( .a(FE_OCP_RBN5803_FE_RN_2224_0), .b(n_14587), .o(n_14642) );
in01f01 g766072 ( .a(n_14662), .o(n_14687) );
no02f06 g766073 ( .a(n_14641), .b(n_13487), .o(n_14662) );
in01m01 g766074 ( .a(n_14719), .o(n_14661) );
na02m06 g766075 ( .a(n_13487), .b(n_14641), .o(n_14719) );
na02s01 g766076 ( .a(n_14685), .b(n_14689), .o(n_14686) );
na02f06 g766081 ( .a(n_14585), .b(FE_OCP_DRV_N3508_n_13329), .o(n_14664) );
na02m08 g766082 ( .a(n_14515), .b(n_14471), .o(n_14616) );
no02s04 TIMEBOOST_cell_1925 ( .a(n_11578), .b(FE_OCP_RBN3289_n_10915), .o(TIMEBOOST_net_577) );
in01m02 g766084 ( .a(n_14709), .o(n_14710) );
na02m04 TIMEBOOST_cell_5614 ( .a(n_16625), .b(n_16598), .o(TIMEBOOST_net_1755) );
ao12s01 g766086 ( .a(n_14947), .b(n_14894), .c(n_14386), .o(n_14996) );
na02f04 g766089 ( .a(n_14580), .b(n_14602), .o(n_14684) );
in01f01 g766091 ( .a(n_14716), .o(n_14707) );
no02m08 TIMEBOOST_cell_8725 ( .a(TIMEBOOST_net_2849), .b(n_28331), .o(n_28422) );
na02f06 TIMEBOOST_cell_2105 ( .a(n_35214), .b(n_30633), .o(TIMEBOOST_net_667) );
oa12f02 g766096 ( .a(n_14379), .b(FE_OCP_RBN5045_n_14450), .c(n_14479), .o(n_14485) );
in01s01 TIMEBOOST_cell_5907 ( .a(FE_OFN1_n_43918), .o(TIMEBOOST_net_1796) );
oa12f04 g766098 ( .a(n_14415), .b(n_14556), .c(n_14555), .o(n_14584) );
in01f02 g766099 ( .a(n_14659), .o(n_14660) );
na02f04 g766100 ( .a(n_14636), .b(n_14579), .o(n_14659) );
na03f06 TIMEBOOST_cell_8398 ( .a(n_39598), .b(FE_RN_1873_0), .c(n_39637), .o(n_39648) );
na02m04 g766104 ( .a(n_14552), .b(FE_OCP_RBN2743_n_14114), .o(n_14583) );
in01s02 g766105 ( .a(n_14607), .o(n_14608) );
in01s02 g766106 ( .a(n_14582), .o(n_14607) );
ao12m06 g766107 ( .a(n_14407), .b(n_14483), .c(n_14368), .o(n_14582) );
na02f06 g766110 ( .a(n_14605), .b(n_14634), .o(n_14635) );
na02s04 TIMEBOOST_cell_8783 ( .a(TIMEBOOST_net_2878), .b(n_3263), .o(n_3362) );
no02s02 TIMEBOOST_cell_5219 ( .a(TIMEBOOST_net_1557), .b(n_47261), .o(n_15371) );
in01m02 g766113 ( .a(n_14632), .o(n_14633) );
na02f02 g766114 ( .a(n_14605), .b(n_14550), .o(n_14632) );
in01s01 g766116 ( .a(n_14706), .o(n_14738) );
na02s04 g766117 ( .a(n_14682), .b(n_14681), .o(n_14706) );
na02m02 TIMEBOOST_cell_2931 ( .a(TIMEBOOST_net_756), .b(n_19365), .o(n_19476) );
na02s01 g766119 ( .a(n_14895), .b(n_14296), .o(n_14993) );
no02s04 TIMEBOOST_cell_5978 ( .a(TIMEBOOST_net_1840), .b(n_23312), .o(n_23377) );
no02s06 TIMEBOOST_cell_5979 ( .a(n_18040), .b(n_17951), .o(TIMEBOOST_net_1841) );
na02s02 g766122 ( .a(n_14545), .b(n_44850), .o(n_14580) );
na02f02 g766123 ( .a(n_14546), .b(n_44849), .o(n_14602) );
na02f02 g766126 ( .a(n_14519), .b(n_13272), .o(n_14587) );
na02f01 g766127 ( .a(n_14573), .b(n_14593), .o(n_14658) );
no02f01 g766128 ( .a(FE_OCP_RBN4248_n_14573), .b(n_14572), .o(n_14657) );
no02f06 g766129 ( .a(n_14450), .b(n_14416), .o(n_14451) );
na02f02 g766130 ( .a(n_14476), .b(n_14450), .o(n_14557) );
no02f06 TIMEBOOST_cell_4973 ( .a(TIMEBOOST_net_1434), .b(n_1958), .o(FE_RN_2082_0) );
na02f02 g766132 ( .a(n_14507), .b(n_13293), .o(n_14579) );
na02s06 g766133 ( .a(n_14556), .b(FE_OCPN1685_n_14555), .o(n_14636) );
na02f08 TIMEBOOST_cell_2106 ( .a(n_35365), .b(TIMEBOOST_net_667), .o(n_35405) );
in01m02 g766135 ( .a(n_14515), .o(n_14516) );
na02s06 TIMEBOOST_cell_8714 ( .a(FE_OCPN1358_n_17778), .b(n_17721), .o(TIMEBOOST_net_2844) );
in01f02 g766137 ( .a(n_14736), .o(n_14737) );
no02s01 TIMEBOOST_cell_4343 ( .a(FE_OFN4763_n_3029), .b(n_2913), .o(TIMEBOOST_net_1262) );
no02m04 g766139 ( .a(n_14868), .b(n_14387), .o(n_14948) );
in01f02 g766140 ( .a(n_14600), .o(n_14601) );
oa12f04 g766141 ( .a(n_14510), .b(n_14467), .c(n_44850), .o(n_14600) );
na02f04 g766144 ( .a(n_14576), .b(n_14549), .o(n_14689) );
oa22f04 g766146 ( .a(n_14590), .b(FE_OCP_RBN4209_n_13796), .c(FE_OCP_RBN2904_n_14590), .d(FE_OCP_RBN4229_n_13962), .o(n_14704) );
oa12s01 g766147 ( .a(n_14840), .b(n_14839), .c(n_14838), .o(n_15869) );
in01s01 g766150 ( .a(FE_OCPN1324_n_14577), .o(n_14598) );
oa12s01 g766155 ( .a(n_14837), .b(n_14836), .c(n_14835), .o(n_15865) );
in01s02 g766159 ( .a(n_14550), .o(n_14551) );
na02s04 g766160 ( .a(n_14462), .b(n_13469), .o(n_14550) );
na02s03 g766161 ( .a(n_14444), .b(n_13514), .o(n_14477) );
no02s01 TIMEBOOST_cell_1992 ( .a(TIMEBOOST_net_610), .b(FE_OCP_RBN5032_n_18951), .o(n_19059) );
in01m01 g766163 ( .a(n_14678), .o(n_14679) );
na02m08 g766164 ( .a(n_14656), .b(n_14625), .o(n_14678) );
na02s01 g766166 ( .a(n_14839), .b(n_14838), .o(n_14840) );
no02s01 TIMEBOOST_cell_5250 ( .a(n_25693), .b(n_25749), .o(TIMEBOOST_net_1573) );
na02m02 g766168 ( .a(n_14498), .b(FE_OCP_RBN4200_n_13796), .o(n_14576) );
na02s02 g766169 ( .a(n_14547), .b(FE_OCP_RBN2759_n_13796), .o(n_14549) );
na02f04 g766170 ( .a(n_14591), .b(FE_OCP_RBN4228_n_13962), .o(n_14682) );
na02s01 g766171 ( .a(n_14836), .b(n_14835), .o(n_14837) );
in01s01 g766172 ( .a(n_14894), .o(n_14895) );
in01s01 g766173 ( .a(n_14868), .o(n_14894) );
na02m04 g766174 ( .a(n_14836), .b(n_14295), .o(n_14868) );
in01s01 g766175 ( .a(n_47256), .o(n_14575) );
in01m01 g766178 ( .a(n_14545), .o(n_14546) );
na02f01 g766179 ( .a(n_14511), .b(n_14510), .o(n_14545) );
in01m01 g766185 ( .a(n_14572), .o(n_14593) );
no02f06 g766186 ( .a(n_14543), .b(n_14544), .o(n_14572) );
no02f04 g766187 ( .a(n_14998), .b(n_14733), .o(n_14735) );
na02f02 g766188 ( .a(n_14998), .b(n_14733), .o(n_14734) );
in01f02 g766189 ( .a(n_14475), .o(n_14476) );
in01s01 TIMEBOOST_cell_7382 ( .a(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_2318) );
na02m08 g766192 ( .a(n_14250), .b(n_14380), .o(n_14478) );
no02f08 g766193 ( .a(n_14504), .b(n_14469), .o(n_14634) );
in01s04 g766194 ( .a(n_14571), .o(n_14628) );
oa12s01 g766197 ( .a(n_14998), .b(n_14677), .c(n_14676), .o(n_14732) );
in01f01 g766200 ( .a(n_14556), .o(n_14507) );
na02f06 g766201 ( .a(n_14414), .b(n_14377), .o(n_14556) );
in01s03 g766202 ( .a(n_14539), .o(n_14540) );
na02s04 g766204 ( .a(n_14447), .b(n_14315), .o(n_14448) );
no02f06 g766205 ( .a(n_14408), .b(n_14270), .o(n_14474) );
no02m08 g766206 ( .a(n_14447), .b(n_14369), .o(n_14483) );
in01m04 g766207 ( .a(n_14505), .o(n_14506) );
na02m08 g766208 ( .a(n_14473), .b(n_14472), .o(n_14505) );
na02s08 g766209 ( .a(n_14535), .b(n_14376), .o(n_14656) );
in01s02 g766210 ( .a(n_14625), .o(n_14626) );
na02m08 g766211 ( .a(n_14536), .b(n_13515), .o(n_14625) );
na02f08 g766214 ( .a(n_14204), .b(n_14251), .o(n_14380) );
na02m04 g766215 ( .a(n_14468), .b(n_13469), .o(n_14471) );
no02f04 g766216 ( .a(n_14468), .b(FE_OCP_RBN4108_n_12880), .o(n_14469) );
no02m04 g766217 ( .a(n_14731), .b(n_14205), .o(n_14836) );
in01s03 g766220 ( .a(n_14379), .o(n_14416) );
na02m04 g766221 ( .a(n_14283), .b(n_13141), .o(n_14379) );
in01s01 g766222 ( .a(n_14511), .o(n_14467) );
na02m04 g766224 ( .a(n_14372), .b(n_13098), .o(n_14510) );
na02f06 g766225 ( .a(n_14677), .b(n_14676), .o(n_14998) );
in01m01 g766226 ( .a(n_14415), .o(n_14479) );
in01s01 TIMEBOOST_cell_7381 ( .a(TIMEBOOST_net_2316), .o(TIMEBOOST_net_2317) );
na02m04 g766228 ( .a(n_14254), .b(FE_OCP_RBN2557_n_13141), .o(n_14415) );
na02f04 g766229 ( .a(n_14335), .b(FE_OCP_RBN5725_n_14120), .o(n_14414) );
na02f02 g766230 ( .a(n_14334), .b(FE_OCP_RBN2071_n_14120), .o(n_14377) );
in01m04 g766231 ( .a(n_14503), .o(n_14504) );
ao12s01 g766233 ( .a(n_14171), .b(n_14780), .c(n_14213), .o(n_14839) );
oa12f06 g766244 ( .a(n_14400), .b(n_14365), .c(n_14318), .o(n_14508) );
in01m01 g766246 ( .a(n_14547), .o(n_14498) );
no02m06 TIMEBOOST_cell_8127 ( .a(TIMEBOOST_net_2694), .b(TIMEBOOST_net_1322), .o(n_21897) );
in01f02 g766248 ( .a(n_14591), .o(n_14592) );
no03f04 TIMEBOOST_cell_8328 ( .a(n_30511), .b(n_30510), .c(TIMEBOOST_net_1105), .o(n_30622) );
in01m02 g766256 ( .a(n_14412), .o(n_14413) );
na02f06 TIMEBOOST_cell_5188 ( .a(FE_OCP_RBN3058_n_15595), .b(n_14524), .o(TIMEBOOST_net_1542) );
ao12s01 g766258 ( .a(n_14757), .b(n_14780), .c(n_14756), .o(n_15747) );
na02s06 g766259 ( .a(n_14323), .b(n_14376), .o(n_14473) );
na02s08 g766260 ( .a(n_14324), .b(n_13515), .o(n_14472) );
na02s02 TIMEBOOST_cell_5191 ( .a(TIMEBOOST_net_1543), .b(n_2646), .o(n_2795) );
no03s01 TIMEBOOST_cell_8438 ( .a(n_36063), .b(n_36062), .c(FE_OCPN950_n_44180), .o(TIMEBOOST_net_2670) );
no02s04 g766264 ( .a(n_14249), .b(n_13418), .o(n_14466) );
na02m04 g766266 ( .a(n_14249), .b(n_13437), .o(n_14250) );
in01s01 TIMEBOOST_cell_8898 ( .a(n_1009), .o(TIMEBOOST_net_2942) );
no02s01 g766268 ( .a(n_14780), .b(n_14756), .o(n_14757) );
no02s04 TIMEBOOST_cell_7734 ( .a(n_4221), .b(FE_OCP_RBN5959_n_4165), .o(TIMEBOOST_net_2498) );
no02s01 TIMEBOOST_cell_6853 ( .a(FE_OCP_DRV_N1434_n_21283), .b(n_22292), .o(TIMEBOOST_net_2184) );
na02f06 g766271 ( .a(n_14245), .b(FE_OCP_RBN6375_n_14154), .o(n_14248) );
na03s02 TIMEBOOST_cell_8327 ( .a(n_4399), .b(n_4495), .c(n_4565), .o(n_4792) );
no02f04 TIMEBOOST_cell_5187 ( .a(TIMEBOOST_net_1541), .b(FE_OCP_RBN3022_n_15319), .o(n_15557) );
na02f02 g766274 ( .a(n_14197), .b(n_13048), .o(n_14247) );
na02m02 g766275 ( .a(n_14436), .b(n_14398), .o(n_14461) );
in01m02 g766276 ( .a(n_14447), .o(n_14408) );
na02f06 g766277 ( .a(n_14329), .b(n_14235), .o(n_14447) );
na02m04 g766278 ( .a(n_14370), .b(n_14332), .o(n_14407) );
na02f06 g766279 ( .a(n_14165), .b(n_14203), .o(n_14204) );
ao12m02 g766280 ( .a(n_14121), .b(n_14240), .c(n_14286), .o(n_14287) );
na02f02 g766281 ( .a(n_14241), .b(n_14091), .o(n_14336) );
in01f02 g766282 ( .a(n_14334), .o(n_14335) );
no03m04 TIMEBOOST_cell_7156 ( .a(n_41367), .b(n_41366), .c(n_41361), .o(n_41390) );
na02f06 g766284 ( .a(n_14245), .b(n_14155), .o(n_14246) );
ao12s02 g766285 ( .a(n_14181), .b(n_14199), .c(FE_OCP_RBN6376_n_14154), .o(n_14244) );
na02m02 g766286 ( .a(n_14200), .b(n_14117), .o(n_14285) );
in01s04 g766289 ( .a(n_14535), .o(n_14536) );
na02s02 TIMEBOOST_cell_4105 ( .a(n_39640), .b(n_39743), .o(TIMEBOOST_net_1143) );
no02f04 g766291 ( .a(n_14534), .b(n_14568), .o(n_14677) );
in01s01 TIMEBOOST_cell_5922 ( .a(TIMEBOOST_net_1810), .o(TIMEBOOST_net_1811) );
in01s01 g766295 ( .a(n_14779), .o(n_15779) );
ao12s01 g766296 ( .a(n_14702), .b(n_14701), .c(n_14700), .o(n_14779) );
in01f02 g766297 ( .a(n_14283), .o(n_14254) );
in01s02 g766301 ( .a(n_14439), .o(n_14821) );
in01s01 g766302 ( .a(n_45521), .o(n_14439) );
ao12m02 g766305 ( .a(n_14214), .b(n_14703), .c(n_14136), .o(n_14731) );
no02s01 TIMEBOOST_cell_1960 ( .a(TIMEBOOST_net_594), .b(n_12662), .o(n_12741) );
no02m04 g766310 ( .a(n_14333), .b(n_14270), .o(n_14370) );
no02m06 g766311 ( .a(n_14201), .b(n_14120), .o(n_14165) );
na02s01 TIMEBOOST_cell_6860 ( .a(TIMEBOOST_net_2188), .b(TIMEBOOST_net_1377), .o(n_1478) );
na02f02 g766313 ( .a(n_14286), .b(n_14240), .o(n_14241) );
in01f04 g766314 ( .a(n_14403), .o(n_14404) );
no02f04 g766315 ( .a(n_14333), .b(n_14369), .o(n_14403) );
na02m02 g766316 ( .a(n_14271), .b(FE_OFN1181_n_13195), .o(n_14332) );
na02s06 g766317 ( .a(n_14272), .b(n_13515), .o(n_14368) );
na02s04 TIMEBOOST_cell_5432 ( .a(n_26118), .b(FE_OCPN3578_n_23354), .o(TIMEBOOST_net_1664) );
na02s06 g766319 ( .a(n_14359), .b(n_13515), .o(n_14402) );
no02s01 g766320 ( .a(n_14703), .b(n_14076), .o(n_14780) );
in01f01 g766321 ( .a(n_14681), .o(n_14569) );
na02m02 g766322 ( .a(n_14533), .b(FE_OCP_RBN4228_n_13962), .o(n_14681) );
no02m02 g766323 ( .a(n_14533), .b(FE_OCP_RBN6695_n_13796), .o(n_14534) );
no02f02 g766324 ( .a(n_14496), .b(FE_OCP_RBN4228_n_13962), .o(n_14568) );
no02m02 g766325 ( .a(n_14182), .b(n_14199), .o(n_14281) );
na02f08 g766326 ( .a(n_14117), .b(n_14133), .o(n_14245) );
in01s01 TIMEBOOST_cell_5923 ( .a(FE_OFN1_n_43918), .o(TIMEBOOST_net_1812) );
no02s01 g766328 ( .a(n_14701), .b(n_14700), .o(n_14702) );
in01s02 g766329 ( .a(n_14436), .o(n_14437) );
na02m02 g766330 ( .a(n_14400), .b(n_14319), .o(n_14436) );
na02m02 g766331 ( .a(n_14199), .b(FE_OCP_RBN6376_n_14154), .o(n_14200) );
no02m08 TIMEBOOST_cell_3936 ( .a(TIMEBOOST_net_1058), .b(n_29339), .o(n_29401) );
in01f02 g766334 ( .a(n_14366), .o(n_14367) );
in01f02 g766335 ( .a(n_14329), .o(n_14366) );
na02f04 g766336 ( .a(n_14185), .b(n_14184), .o(n_14329) );
no02s04 g766337 ( .a(n_14161), .b(n_14135), .o(n_14251) );
in01s01 g766338 ( .a(n_14398), .o(n_14399) );
in01s01 g766339 ( .a(n_14365), .o(n_14398) );
ao12f06 g766340 ( .a(n_14146), .b(n_14228), .c(n_14230), .o(n_14365) );
in01s01 g766341 ( .a(n_15250), .o(n_14364) );
in01s01 g766342 ( .a(n_14328), .o(n_15250) );
in01f02 g766343 ( .a(n_14328), .o(n_14327) );
no02f06 g766344 ( .a(n_14162), .b(n_14193), .o(n_14328) );
no02f06 TIMEBOOST_cell_7763 ( .a(TIMEBOOST_net_2512), .b(n_19597), .o(n_19802) );
in01s04 g766351 ( .a(n_14326), .o(n_16070) );
na02s01 TIMEBOOST_cell_7806 ( .a(n_16261), .b(n_16258), .o(TIMEBOOST_net_2534) );
in01s04 g766355 ( .a(n_14323), .o(n_14324) );
in01s01 g766359 ( .a(n_14362), .o(n_14363) );
ao22m02 g766360 ( .a(n_14176), .b(n_13514), .c(n_14225), .d(n_13515), .o(n_14362) );
no03m03 TIMEBOOST_cell_8389 ( .a(n_34954), .b(FE_OCP_RBN6074_n_44256), .c(n_35984), .o(n_36032) );
na02s06 g766363 ( .a(n_14163), .b(n_13322), .o(n_14194) );
no02s04 g766364 ( .a(n_14123), .b(n_13131), .o(n_14162) );
no02f04 g766365 ( .a(n_14124), .b(n_13130), .o(n_14193) );
no02s04 g766366 ( .a(n_14177), .b(n_13469), .o(n_14333) );
no02f06 g766367 ( .a(n_14178), .b(n_13514), .o(n_14369) );
no02s02 g766368 ( .a(n_14099), .b(FE_OCP_RBN4102_n_12880), .o(n_14135) );
in01s02 g766369 ( .a(n_14160), .o(n_14161) );
na02s02 g766370 ( .a(n_14096), .b(n_13916), .o(n_14160) );
na02s01 g766372 ( .a(n_14653), .b(n_14040), .o(n_14701) );
no02m04 g766373 ( .a(n_14137), .b(n_14653), .o(n_14703) );
na02f04 g766374 ( .a(n_14278), .b(FE_OCP_DRV_N4502_FE_OCP_RBN1807_n_13010), .o(n_14400) );
na02m08 TIMEBOOST_cell_8548 ( .a(TIMEBOOST_net_1233), .b(n_19264), .o(TIMEBOOST_net_2761) );
in01m01 g766376 ( .a(n_14318), .o(n_14319) );
no02m04 g766377 ( .a(FE_OCP_DRV_N3504_FE_OCP_RBN1807_n_13010), .b(n_14278), .o(n_14318) );
na02s01 g766378 ( .a(n_14274), .b(FE_OCP_RBN2750_n_14157), .o(n_14277) );
no02s01 g766379 ( .a(FE_RN_1606_0), .b(FE_OCP_RBN2750_n_14157), .o(n_14276) );
no02s01 g766380 ( .a(FE_OCP_RBN2073_n_14120), .b(n_14190), .o(n_14192) );
in01s01 g766381 ( .a(n_14238), .o(n_14239) );
na02s01 g766382 ( .a(FE_OCP_RBN2073_n_14120), .b(n_14190), .o(n_14238) );
na02f06 TIMEBOOST_cell_7483 ( .a(TIMEBOOST_net_2372), .b(n_37312), .o(n_37461) );
na02m04 g766384 ( .a(n_14268), .b(n_14267), .o(n_14360) );
no02s02 TIMEBOOST_cell_2911 ( .a(TIMEBOOST_net_746), .b(n_12983), .o(n_13062) );
na02s02 TIMEBOOST_cell_8751 ( .a(TIMEBOOST_net_2862), .b(n_2539), .o(n_47026) );
in01m01 g766389 ( .a(n_14199), .o(n_14187) );
in01s02 g766390 ( .a(n_14133), .o(n_14199) );
ao12f06 g766391 ( .a(n_14028), .b(n_14026), .c(n_14101), .o(n_14133) );
in01m02 g766392 ( .a(n_14286), .o(n_14186) );
no02f08 g766393 ( .a(n_14103), .b(n_14105), .o(n_14286) );
na03f04 TIMEBOOST_cell_8186 ( .a(TIMEBOOST_net_1826), .b(n_37366), .c(n_37353), .o(TIMEBOOST_net_2372) );
na02f02 g766395 ( .a(n_14122), .b(n_14128), .o(n_14184) );
in01s01 g766396 ( .a(n_14397), .o(n_15518) );
in01s01 g766397 ( .a(n_14359), .o(n_14397) );
in01s04 g766398 ( .a(n_14359), .o(n_14358) );
no02s06 TIMEBOOST_cell_5479 ( .a(TIMEBOOST_net_1687), .b(n_11001), .o(n_11118) );
in01f01 g766400 ( .a(n_14533), .o(n_14496) );
ao22f02 g766401 ( .a(n_14355), .b(FE_OCP_RBN4229_n_13962), .c(n_16143), .d(FE_OCP_RBN4209_n_13796), .o(n_14533) );
in01s01 g766402 ( .a(n_15666), .o(n_14652) );
ao12s01 g766403 ( .a(n_14567), .b(n_14566), .c(n_14565), .o(n_15666) );
oa12s01 g766404 ( .a(n_14622), .b(n_14621), .c(n_14620), .o(n_15718) );
in01s01 g766405 ( .a(n_14317), .o(n_14396) );
in01s02 g766408 ( .a(n_14273), .o(n_14317) );
in01m02 g766409 ( .a(n_14273), .o(n_14252) );
na02f08 g766410 ( .a(n_14156), .b(n_14132), .o(n_14273) );
in01s02 g766411 ( .a(n_14271), .o(n_14272) );
na02m04 g766413 ( .a(FE_OCP_RBN2075_n_14093), .b(n_13132), .o(n_14156) );
na02s04 g766414 ( .a(n_14093), .b(n_13133), .o(n_14132) );
na02m02 g766415 ( .a(n_14032), .b(n_14000), .o(n_14034) );
no02f04 g766416 ( .a(n_14002), .b(n_13958), .o(n_14071) );
na02s01 TIMEBOOST_cell_6184 ( .a(TIMEBOOST_net_1943), .b(n_43248), .o(n_43405) );
na02s02 TIMEBOOST_cell_8883 ( .a(TIMEBOOST_net_2928), .b(n_22266), .o(n_22379) );
na02s02 g766419 ( .a(n_14102), .b(n_14240), .o(n_14129) );
na02f02 g766420 ( .a(n_14127), .b(n_13437), .o(n_14128) );
na02m06 g766421 ( .a(n_14233), .b(n_13469), .o(n_14235) );
in01s02 g766423 ( .a(n_14270), .o(n_14315) );
no02m06 g766424 ( .a(FE_OCP_RBN4109_n_12880), .b(n_14233), .o(n_14270) );
na02m04 g766425 ( .a(n_14564), .b(n_14108), .o(n_14653) );
no02m08 TIMEBOOST_cell_5173 ( .a(TIMEBOOST_net_1534), .b(n_34287), .o(n_34342) );
na02s01 TIMEBOOST_cell_6355 ( .a(n_16086), .b(n_16977), .o(TIMEBOOST_net_2029) );
no02f06 g766428 ( .a(n_14104), .b(n_13887), .o(n_14105) );
na02f06 g766429 ( .a(n_14102), .b(n_13886), .o(n_14103) );
in01f02 g766430 ( .a(n_14268), .o(n_14269) );
na02f02 g766431 ( .a(n_14147), .b(n_14230), .o(n_14268) );
no02s01 g766432 ( .a(n_14566), .b(n_14565), .o(n_14567) );
in01s01 g766433 ( .a(n_14125), .o(n_14126) );
na02m02 g766434 ( .a(n_14029), .b(n_14101), .o(n_14125) );
na02s04 g766435 ( .a(n_14100), .b(n_13122), .o(n_14163) );
na02s01 g766436 ( .a(n_14621), .b(n_14620), .o(n_14622) );
in01m02 g766437 ( .a(n_14123), .o(n_14124) );
no02f04 g766439 ( .a(n_14154), .b(n_14153), .o(n_14155) );
na02s02 g766440 ( .a(FE_OCP_RBN6376_n_14154), .b(n_14117), .o(n_14229) );
no02m02 g766441 ( .a(n_14181), .b(n_14154), .o(n_14182) );
in01s02 g766447 ( .a(n_14099), .o(n_14120) );
in01f02 g766450 ( .a(n_14177), .o(n_14178) );
in01m02 g766452 ( .a(n_14266), .o(n_14267) );
in01s01 g766453 ( .a(n_14228), .o(n_14266) );
no02f06 g766454 ( .a(n_14089), .b(n_14116), .o(n_14228) );
in01s01 g766464 ( .a(n_14225), .o(n_14265) );
in01s03 g766465 ( .a(n_14176), .o(n_14225) );
no02s01 TIMEBOOST_cell_3822 ( .a(TIMEBOOST_net_1001), .b(n_46200), .o(TIMEBOOST_net_185) );
oa12s01 g766468 ( .a(n_14066), .b(n_14065), .c(n_14064), .o(n_15935) );
oa12s01 g766469 ( .a(n_14495), .b(n_14494), .c(n_14493), .o(n_15786) );
no02m06 g766476 ( .a(n_14030), .b(n_14067), .o(n_14149) );
ao12s01 g766482 ( .a(n_14532), .b(n_14531), .c(n_14530), .o(n_15663) );
na02f04 g766484 ( .a(n_13959), .b(n_14005), .o(n_14096) );
na02s02 g766485 ( .a(n_14023), .b(n_13441), .o(n_14068) );
na02s02 TIMEBOOST_cell_6611 ( .a(n_12233), .b(n_11900), .o(TIMEBOOST_net_2063) );
no02s04 g766489 ( .a(n_13995), .b(n_13029), .o(n_14030) );
no02f04 g766490 ( .a(n_13997), .b(n_12968), .o(n_14100) );
no02m04 g766491 ( .a(n_13996), .b(n_13028), .o(n_14067) );
na02m02 g766492 ( .a(n_13927), .b(n_13195), .o(n_13959) );
na02f04 g766493 ( .a(FE_OCP_RBN5038_n_13927), .b(FE_OCP_RBN4102_n_12880), .o(n_14005) );
no02s01 g766494 ( .a(n_14531), .b(n_14530), .o(n_14532) );
na02s01 g766495 ( .a(n_14494), .b(n_14493), .o(n_14495) );
na02m04 g766496 ( .a(n_14118), .b(FE_OCP_RBN2045_n_12907), .o(n_14230) );
in01f01 g766497 ( .a(n_14146), .o(n_14147) );
no02f04 g766498 ( .a(FE_OCP_RBN2045_n_12907), .b(n_14118), .o(n_14146) );
in01s02 g766499 ( .a(n_14144), .o(n_14145) );
no02s06 TIMEBOOST_cell_6624 ( .a(TIMEBOOST_net_2069), .b(n_33023), .o(FE_RN_428_0) );
na02s01 g766501 ( .a(n_14065), .b(n_14064), .o(n_14066) );
na02f04 g766502 ( .a(n_14004), .b(FE_OCP_RBN2512_n_12800), .o(n_14101) );
in01m01 g766503 ( .a(n_14028), .o(n_14029) );
no02f04 g766504 ( .a(n_14004), .b(FE_OCP_RBN2512_n_12800), .o(n_14028) );
no02f06 g766506 ( .a(n_14092), .b(n_12877), .o(n_14154) );
in01m01 g766509 ( .a(n_14117), .o(n_14181) );
na02m08 g766510 ( .a(n_14092), .b(n_12877), .o(n_14117) );
in01m01 g766511 ( .a(n_14032), .o(n_14002) );
oa12f06 g766512 ( .a(n_13883), .b(n_13930), .c(FE_OFN4792_n_13195), .o(n_14032) );
oa12f04 g766513 ( .a(n_13948), .b(n_14027), .c(FE_OFN4793_n_13195), .o(n_14104) );
ao12f04 g766514 ( .a(n_13947), .b(n_14027), .c(FE_OFN4793_n_13195), .o(n_14102) );
na02f06 g766515 ( .a(n_14000), .b(n_13891), .o(n_14001) );
ao12s01 g766516 ( .a(n_14080), .b(n_14457), .c(n_14078), .o(n_14566) );
in01s02 g766517 ( .a(n_16143), .o(n_14355) );
na02f04 g766518 ( .a(n_14172), .b(n_14222), .o(n_16143) );
ao12f04 g766519 ( .a(n_46984), .b(n_14115), .c(n_12868), .o(n_14116) );
in01s01 g766526 ( .a(FE_OCP_RBN2744_n_14114), .o(n_14274) );
na02m06 TIMEBOOST_cell_5671 ( .a(TIMEBOOST_net_1783), .b(n_11511), .o(n_11731) );
in01s01 g766530 ( .a(n_14062), .o(n_14063) );
in01s01 g766531 ( .a(n_14026), .o(n_14062) );
ao12f06 g766532 ( .a(n_13922), .b(n_13994), .c(n_14064), .o(n_14026) );
in01s01 g766533 ( .a(n_14564), .o(n_14621) );
oa12m04 g766534 ( .a(n_14111), .b(n_14432), .c(n_14079), .o(n_14564) );
no02m08 g766535 ( .a(n_14057), .b(n_14090), .o(n_14233) );
no02s01 TIMEBOOST_cell_6801 ( .a(n_6250), .b(n_5341), .o(TIMEBOOST_net_2158) );
na02m04 g766538 ( .a(FE_OCP_RBN5701_n_13954), .b(n_13376), .o(n_14025) );
na03m06 TIMEBOOST_cell_6457 ( .a(n_2627), .b(n_2626), .c(n_2688), .o(n_2778) );
na02m08 g766541 ( .a(n_13014), .b(n_13957), .o(n_13997) );
in01s01 g766542 ( .a(n_14121), .o(n_14091) );
no02f06 g766543 ( .a(n_14059), .b(FE_OFN4793_n_13195), .o(n_14121) );
na02s06 g766544 ( .a(n_14059), .b(FE_OFN4793_n_13195), .o(n_14240) );
no02s03 g766545 ( .a(n_14018), .b(n_13437), .o(n_14057) );
no02s06 g766546 ( .a(FE_OCP_RBN2724_n_14018), .b(FE_OFN4796_n_13195), .o(n_14090) );
na02f04 g766547 ( .a(n_13858), .b(FE_OCP_RBN4096_n_12880), .o(n_13891) );
in01s01 g766548 ( .a(n_14000), .o(n_13958) );
na02f06 g766549 ( .a(n_13930), .b(FE_OFN4792_n_13195), .o(n_14000) );
no02s01 g766550 ( .a(n_14457), .b(n_14110), .o(n_14531) );
in01m02 g766551 ( .a(n_13995), .o(n_13996) );
na02f01 g766553 ( .a(n_14115), .b(n_14140), .o(n_14172) );
na02m02 g766554 ( .a(n_14049), .b(n_14141), .o(n_14222) );
no02s04 g766555 ( .a(n_14115), .b(n_12868), .o(n_14089) );
na02s01 g766556 ( .a(FE_OCP_RBN5710_n_13984), .b(FE_OCPN1250_n_13882), .o(n_14056) );
no02s01 g766557 ( .a(FE_OCP_RBN5710_n_13984), .b(FE_OCPN1250_n_13882), .o(n_14055) );
in01s01 g766558 ( .a(n_14023), .o(n_14024) );
na02f08 TIMEBOOST_cell_2032 ( .a(TIMEBOOST_net_630), .b(n_33835), .o(n_33946) );
in01s02 g766560 ( .a(n_13928), .o(n_13929) );
oa12m04 g766561 ( .a(n_46415), .b(n_13866), .c(n_13138), .o(n_13928) );
in01m04 g766562 ( .a(n_13955), .o(n_13956) );
na02s01 g766564 ( .a(n_13923), .b(n_13994), .o(n_14065) );
oa12f02 g766565 ( .a(n_13981), .b(n_14019), .c(n_14051), .o(n_14052) );
no02f02 g766566 ( .a(n_14020), .b(n_13982), .o(n_14088) );
oa12s01 g766567 ( .a(n_13967), .b(n_14435), .c(n_14039), .o(n_14494) );
in01s04 g766568 ( .a(n_14021), .o(n_14022) );
na02m04 TIMEBOOST_cell_5445 ( .a(TIMEBOOST_net_1670), .b(n_5717), .o(TIMEBOOST_net_1342) );
ao12s01 g766570 ( .a(n_14393), .b(n_14435), .c(n_14392), .o(n_15669) );
in01s02 g766576 ( .a(FE_OCP_RBN5039_n_13927), .o(n_14190) );
no02f04 g766580 ( .a(n_13989), .b(n_13952), .o(n_14118) );
no02m06 TIMEBOOST_cell_8517 ( .a(TIMEBOOST_net_2745), .b(n_38121), .o(n_38141) );
in01s01 g766583 ( .a(FE_OCP_RBN2730_n_14072), .o(n_15299) );
no02f06 g766585 ( .a(n_13953), .b(n_13926), .o(n_14072) );
no02m08 g766588 ( .a(n_13924), .b(n_13470), .o(n_13954) );
no02m04 g766589 ( .a(FE_OCP_RBN6660_n_13884), .b(n_13363), .o(n_13953) );
no02s03 g766590 ( .a(n_13884), .b(n_13364), .o(n_13926) );
no02f02 TIMEBOOST_cell_4086 ( .a(TIMEBOOST_net_1133), .b(n_30963), .o(n_30987) );
no02f02 g766593 ( .a(n_13988), .b(n_14019), .o(n_14020) );
no02s02 g766594 ( .a(n_13931), .b(FE_OCP_DRV_N4499_n_13785), .o(n_13952) );
no02m04 g766595 ( .a(n_13988), .b(FE_OCP_DRV_N4500_n_13785), .o(n_13989) );
na02s01 TIMEBOOST_cell_8719 ( .a(TIMEBOOST_net_2846), .b(n_7359), .o(n_7425) );
in01s01 g766597 ( .a(n_13922), .o(n_13923) );
no02m04 g766598 ( .a(n_13890), .b(FE_OCPN5222_FE_OFN753_n_13889), .o(n_13922) );
no02s01 g766599 ( .a(n_14435), .b(n_14392), .o(n_14393) );
na02s01 g766600 ( .a(n_14354), .b(n_14433), .o(n_14434) );
na02f04 g766602 ( .a(n_13890), .b(FE_OCPN5222_FE_OFN753_n_13889), .o(n_13994) );
no02s01 g766603 ( .a(n_14015), .b(n_13944), .o(n_14050) );
no02s04 TIMEBOOST_cell_8090 ( .a(FE_OCPN5226_n_25509), .b(FE_OCP_RBN6815_n_25753), .o(TIMEBOOST_net_2676) );
in01m02 g766605 ( .a(n_14457), .o(n_14432) );
no02m04 g766606 ( .a(n_14435), .b(n_14007), .o(n_14457) );
in01s01 g766607 ( .a(n_14115), .o(n_14049) );
na02f08 g766608 ( .a(n_13946), .b(n_13980), .o(n_14115) );
in01m01 g766609 ( .a(n_14140), .o(n_14141) );
oa22f01 g766610 ( .a(n_46984), .b(n_12868), .c(n_14013), .d(n_12846), .o(n_14140) );
na02f04 TIMEBOOST_cell_1981 ( .a(n_41348), .b(FE_OCP_RBN4045_n_41298), .o(TIMEBOOST_net_605) );
in01s01 g766616 ( .a(n_16138), .o(n_16244) );
ao12s01 g766617 ( .a(n_14309), .b(n_14308), .c(n_14307), .o(n_16138) );
in01s01 g766618 ( .a(n_15631), .o(n_14391) );
oa12s01 g766619 ( .a(n_14262), .b(n_14261), .c(n_14260), .o(n_15631) );
in01s01 g766626 ( .a(FE_OCP_RBN1821_n_13858), .o(n_13950) );
na02f06 g766630 ( .a(n_13817), .b(n_13783), .o(n_13930) );
na02f06 g766631 ( .a(n_13862), .b(n_13842), .o(n_14027) );
no02f02 TIMEBOOST_cell_6124 ( .a(TIMEBOOST_net_1913), .b(n_14905), .o(TIMEBOOST_net_1555) );
in01s01 g766637 ( .a(n_13960), .o(n_13984) );
in01f02 g766638 ( .a(n_13960), .o(n_13949) );
no02m08 g766640 ( .a(n_13857), .b(n_13319), .o(n_13924) );
na02s01 g766641 ( .a(n_14261), .b(n_14260), .o(n_14262) );
no02s01 g766642 ( .a(n_14308), .b(n_14307), .o(n_14309) );
in01s01 g766643 ( .a(n_13948), .o(n_14019) );
na02m06 g766644 ( .a(n_13918), .b(FE_OCP_RBN4104_n_12880), .o(n_13948) );
in01s01 g766645 ( .a(n_13981), .o(n_13982) );
in01s01 g766646 ( .a(n_13947), .o(n_13981) );
no02f06 g766647 ( .a(n_13918), .b(FE_OCP_RBN4104_n_12880), .o(n_13947) );
na02f04 g766648 ( .a(FE_OCP_RBN2683_n_13818), .b(FE_OFN4793_n_13195), .o(n_13862) );
na02s04 g766649 ( .a(n_13818), .b(FE_OCP_RBN4102_n_12880), .o(n_13842) );
no02s01 TIMEBOOST_cell_6123 ( .a(n_14215), .b(FE_OCP_RBN2834_n_13962), .o(TIMEBOOST_net_1913) );
no02m06 TIMEBOOST_cell_8843 ( .a(TIMEBOOST_net_2908), .b(n_10435), .o(n_10559) );
na02m02 g766652 ( .a(n_13756), .b(FE_OCPN929_n_12880), .o(n_13783) );
na02f04 g766653 ( .a(n_13784), .b(FE_OCP_RBN4099_n_12880), .o(n_13817) );
na02f06 g766654 ( .a(n_13945), .b(n_13944), .o(n_13946) );
in01s01 g766655 ( .a(n_14015), .o(n_14016) );
na02s01 g766656 ( .a(n_13980), .b(n_13945), .o(n_14015) );
in01s02 g766657 ( .a(n_13931), .o(n_14051) );
in01f02 g766658 ( .a(n_13931), .o(n_13988) );
na02f06 g766659 ( .a(n_13887), .b(n_13886), .o(n_13931) );
na02f04 TIMEBOOST_cell_2031 ( .a(FE_OCP_RBN4914_n_33833), .b(n_33697), .o(TIMEBOOST_net_630) );
no02s01 TIMEBOOST_cell_8770 ( .a(n_14016), .b(n_13909), .o(TIMEBOOST_net_2872) );
na02s04 g766663 ( .a(n_13857), .b(n_13282), .o(n_13884) );
in01s06 g766665 ( .a(n_13815), .o(n_13866) );
in01m02 g766666 ( .a(n_13815), .o(n_13816) );
no03f02 TIMEBOOST_cell_8270 ( .a(n_3673), .b(n_3155), .c(FE_OCP_RBN2804_n_3261), .o(TIMEBOOST_net_2110) );
oa12m02 g766668 ( .a(n_13707), .b(n_13813), .c(n_13781), .o(n_13814) );
no02s02 TIMEBOOST_cell_6680 ( .a(TIMEBOOST_net_2097), .b(n_3982), .o(n_4252) );
in01f02 g766671 ( .a(n_13883), .o(n_13913) );
ao12s01 g766674 ( .a(n_13855), .b(n_13854), .c(n_13853), .o(n_15791) );
in01s01 g766675 ( .a(n_15564), .o(n_14354) );
oa12s01 g766676 ( .a(n_14221), .b(n_14220), .c(n_14219), .o(n_15564) );
no02m04 g766677 ( .a(n_14009), .b(n_14218), .o(n_14435) );
na02f08 TIMEBOOST_cell_1958 ( .a(n_37353), .b(TIMEBOOST_net_593), .o(n_37399) );
na02s02 g766679 ( .a(n_13806), .b(n_13381), .o(n_13839) );
na02m06 TIMEBOOST_cell_4957 ( .a(TIMEBOOST_net_1426), .b(FE_RN_349_0), .o(n_46972) );
na02m08 g766681 ( .a(n_13774), .b(n_13279), .o(n_13857) );
no02m04 g766683 ( .a(n_13729), .b(n_12869), .o(n_13757) );
na02s01 g766684 ( .a(n_14220), .b(n_14219), .o(n_14221) );
no02m04 g766685 ( .a(n_14217), .b(n_13899), .o(n_14218) );
na02m06 TIMEBOOST_cell_5960 ( .a(TIMEBOOST_net_1831), .b(FE_RN_1400_0), .o(FE_RN_1399_0) );
oa12s01 g766687 ( .a(n_14562), .b(n_14529), .c(n_14527), .o(n_14619) );
ao12m04 g766688 ( .a(n_13124), .b(n_13778), .c(n_13777), .o(n_13812) );
na02m04 g766689 ( .a(n_13779), .b(n_13238), .o(n_13838) );
na02f04 g766690 ( .a(n_13849), .b(n_12798), .o(n_13945) );
na02m06 g766691 ( .a(n_13850), .b(FE_OCPN847_n_12799), .o(n_13980) );
no02s01 g766692 ( .a(n_13853), .b(n_13854), .o(n_13855) );
ao12s01 g766693 ( .a(n_13976), .b(n_14139), .c(n_13876), .o(n_14261) );
na02s01 g766694 ( .a(n_14217), .b(n_13977), .o(n_14308) );
no02f04 TIMEBOOST_cell_4108 ( .a(TIMEBOOST_net_1144), .b(n_15620), .o(n_15732) );
in01f01 g766699 ( .a(n_46984), .o(n_14013) );
in01s01 g766704 ( .a(n_13882), .o(n_13912) );
in01s01 g766705 ( .a(n_13860), .o(n_13882) );
in01s04 g766706 ( .a(n_13860), .o(n_13859) );
na03s04 TIMEBOOST_cell_6538 ( .a(n_31029), .b(n_27536), .c(n_31007), .o(n_31103) );
oa12f08 g766708 ( .a(n_13753), .b(n_13853), .c(n_13805), .o(n_14064) );
in01f02 g766714 ( .a(n_13756), .o(n_13784) );
no02f02 TIMEBOOST_cell_4085 ( .a(n_30910), .b(FE_OCPN1404_n_30823), .o(TIMEBOOST_net_1133) );
na02s04 g766724 ( .a(n_13778), .b(n_13777), .o(n_13779) );
no02s04 g766725 ( .a(n_13732), .b(n_13261), .o(n_13759) );
na02m04 TIMEBOOST_cell_8745 ( .a(TIMEBOOST_net_2859), .b(n_33960), .o(n_34059) );
no02f08 g766727 ( .a(n_13694), .b(n_12870), .o(n_13729) );
no02s01 g766728 ( .a(n_14139), .b(n_13903), .o(n_14220) );
na02f02 g766730 ( .a(n_13829), .b(FE_OCP_RBN2640_n_13667), .o(n_13851) );
na02s06 TIMEBOOST_cell_6790 ( .a(TIMEBOOST_net_2152), .b(n_43282), .o(n_43332) );
no02f04 TIMEBOOST_cell_4084 ( .a(TIMEBOOST_net_1132), .b(FE_RN_2439_0), .o(n_15700) );
no02f02 g766733 ( .a(n_13725), .b(n_13690), .o(n_13731) );
no02s02 TIMEBOOST_cell_1901 ( .a(n_11439), .b(n_45300), .o(TIMEBOOST_net_565) );
in01s02 g766736 ( .a(n_13806), .o(n_13807) );
in01s02 g766737 ( .a(n_13774), .o(n_13806) );
no02s01 g766739 ( .a(n_13805), .b(n_13754), .o(n_13854) );
no02f06 g766741 ( .a(n_13724), .b(n_13725), .o(n_13813) );
na02m04 g766742 ( .a(n_14139), .b(n_13905), .o(n_14217) );
in01s01 g766743 ( .a(n_13944), .o(n_13909) );
na02f04 g766744 ( .a(n_13828), .b(n_13801), .o(n_13944) );
in01m02 g766745 ( .a(n_13849), .o(n_13850) );
in01s01 g766747 ( .a(n_13879), .o(n_13880) );
oa12s01 g766748 ( .a(n_13804), .b(n_13803), .c(n_13827), .o(n_13879) );
in01s01 g766749 ( .a(n_15788), .o(n_14112) );
ao12s01 g766750 ( .a(n_14012), .b(n_14011), .c(n_14010), .o(n_15788) );
in01s01 g766751 ( .a(n_16246), .o(n_14433) );
oa12s01 g766752 ( .a(n_14084), .b(n_14085), .c(n_14083), .o(n_16246) );
no02s01 g766753 ( .a(n_14011), .b(n_14010), .o(n_14012) );
no02m04 g766754 ( .a(n_14085), .b(n_13902), .o(n_14139) );
na02s01 g766755 ( .a(n_14085), .b(n_14083), .o(n_14084) );
no02f02 g766757 ( .a(n_13789), .b(n_13788), .o(n_13829) );
no02s01 g766758 ( .a(n_14489), .b(n_14528), .o(n_14529) );
in01s06 g766759 ( .a(n_13732), .o(n_13778) );
no02m06 g766762 ( .a(n_13722), .b(FE_OCPN1306_n_13721), .o(n_13805) );
in01s01 g766763 ( .a(n_13753), .o(n_13754) );
na02s01 g766765 ( .a(n_13803), .b(n_13827), .o(n_13804) );
ao12m02 g766766 ( .a(n_13173), .b(n_13645), .c(n_13213), .o(n_13695) );
oa12f04 g766767 ( .a(n_13099), .b(n_13664), .c(n_13083), .o(n_13709) );
oa12f08 g766769 ( .a(FE_OCPN1695_n_12836), .b(n_13601), .c(n_12766), .o(n_13694) );
oa12f04 g766770 ( .a(n_13573), .b(FE_OCP_RBN4092_n_12880), .c(n_13693), .o(n_13725) );
oa12s01 g766777 ( .a(n_13749), .b(n_13748), .c(n_13747), .o(n_15678) );
oa12f02 g766778 ( .a(n_13743), .b(n_13827), .c(n_13800), .o(n_13828) );
in01s01 g766782 ( .a(n_13751), .o(n_13785) );
in01s03 g766783 ( .a(n_13751), .o(n_13750) );
no02s06 TIMEBOOST_cell_6044 ( .a(TIMEBOOST_net_1873), .b(n_24163), .o(n_24288) );
na02s01 TIMEBOOST_cell_5225 ( .a(TIMEBOOST_net_1560), .b(n_34927), .o(n_34990) );
no02s40 TIMEBOOST_cell_8134 ( .a(FE_OCP_RBN7101_n_44365), .b(delay_xor_ln22_unr12_stage5_stallmux_q_0_), .o(TIMEBOOST_net_2698) );
no02f04 TIMEBOOST_cell_4080 ( .a(TIMEBOOST_net_1130), .b(n_5693), .o(TIMEBOOST_net_927) );
in01s01 g766790 ( .a(n_13690), .o(n_13707) );
no02m02 g766791 ( .a(n_13661), .b(FE_OCP_RBN4092_n_12880), .o(n_13690) );
no02m04 TIMEBOOST_cell_8597 ( .a(TIMEBOOST_net_2785), .b(n_30858), .o(n_30875) );
na02s06 TIMEBOOST_cell_8754 ( .a(n_14358), .b(n_14376), .o(TIMEBOOST_net_2864) );
no02s02 g766794 ( .a(n_13661), .b(FE_OCPN929_n_12880), .o(n_13781) );
na02s01 g766795 ( .a(n_14526), .b(n_14525), .o(n_14527) );
na02s01 g766796 ( .a(n_14429), .b(n_14562), .o(n_14563) );
na02s01 g766797 ( .a(n_14525), .b(n_14562), .o(n_15575) );
na02s01 g766798 ( .a(n_13747), .b(n_13748), .o(n_13749) );
na02s02 g766799 ( .a(n_13827), .b(n_13800), .o(n_13801) );
na02f04 g766800 ( .a(FE_OCP_RBN6661_n_13702), .b(FE_OCP_RBN2697_n_13703), .o(n_13746) );
no02s03 g766801 ( .a(n_13703), .b(n_13702), .o(n_13713) );
oa12s01 g766802 ( .a(n_13864), .b(n_13943), .c(n_13939), .o(n_14011) );
no02m04 g766803 ( .a(n_13940), .b(n_13865), .o(n_14085) );
no02f06 g766804 ( .a(FE_OCP_RBN2696_n_13703), .b(n_13644), .o(n_13789) );
na02f08 g766805 ( .a(FE_OCP_RBN6662_n_13702), .b(n_13635), .o(n_13788) );
no02s01 TIMEBOOST_cell_7099 ( .a(n_27308), .b(n_27309), .o(TIMEBOOST_net_2308) );
in01s01 g766807 ( .a(n_14489), .o(n_14490) );
no03s10 TIMEBOOST_cell_5721 ( .a(TIMEBOOST_net_1438), .b(n_28030), .c(n_28251), .o(n_28347) );
ao12f08 g766810 ( .a(n_13657), .b(n_13747), .c(n_13705), .o(n_13853) );
oa12s01 g766811 ( .a(n_13704), .b(n_13743), .c(n_13800), .o(n_13803) );
in01s01 g766812 ( .a(n_15482), .o(n_15513) );
oa12s01 g766813 ( .a(n_13942), .b(n_13943), .c(n_13941), .o(n_15482) );
na02s01 g766814 ( .a(n_14346), .b(n_14351), .o(n_14431) );
no02s01 g766815 ( .a(n_14349), .b(n_14382), .o(n_14430) );
na02s01 g766816 ( .a(n_13943), .b(n_13941), .o(n_13942) );
no02s01 g766817 ( .a(n_14342), .b(n_14425), .o(n_14526) );
in01s01 g766818 ( .a(n_14352), .o(n_14353) );
na02s01 g766819 ( .a(n_14306), .b(n_14561), .o(n_14352) );
no02s01 g766820 ( .a(n_14350), .b(n_14300), .o(n_14351) );
in01s01 g766821 ( .a(n_14429), .o(n_14528) );
no02s01 g766822 ( .a(n_14426), .b(n_14343), .o(n_14429) );
na02s01 g766823 ( .a(n_14381), .b(n_14297), .o(n_14382) );
na02s01 g766824 ( .a(n_14488), .b(n_14339), .o(n_15398) );
no02s01 g766825 ( .a(n_14455), .b(n_14454), .o(n_15520) );
na02s01 g766826 ( .a(n_14341), .b(n_14344), .o(n_15572) );
na02s01 g766827 ( .a(n_14422), .b(n_14306), .o(n_15361) );
na02s01 g766828 ( .a(n_13908), .b(n_14452), .o(n_14562) );
oa12s01 g766829 ( .a(n_14427), .b(n_14947), .c(n_14299), .o(n_14428) );
no02s01 g766830 ( .a(n_14426), .b(n_14425), .o(n_15442) );
in01s01 g766831 ( .a(n_14423), .o(n_14424) );
na02s01 g766832 ( .a(n_14381), .b(n_14301), .o(n_14423) );
na02s01 g766833 ( .a(n_13907), .b(n_14215), .o(n_14525) );
na02s01 g766834 ( .a(n_13658), .b(n_13705), .o(n_13748) );
na02s01 g766835 ( .a(n_13743), .b(n_13800), .o(n_13704) );
in01m06 g766836 ( .a(n_13645), .o(n_13711) );
in01m04 g766837 ( .a(n_13664), .o(n_13665) );
in01m04 g766838 ( .a(n_13645), .o(n_13664) );
ao12f08 g766839 ( .a(n_13043), .b(n_13633), .c(FE_OCPN4522_n_13015), .o(n_13645) );
ao12f08 g766842 ( .a(n_12722), .b(n_13560), .c(n_12773), .o(n_13601) );
no03s10 TIMEBOOST_cell_6410 ( .a(n_17192), .b(n_17084), .c(n_17188), .o(TIMEBOOST_net_1828) );
ao12s01 g766848 ( .a(n_13741), .b(n_13740), .c(n_13739), .o(n_15686) );
na02f06 g766854 ( .a(n_13712), .b(n_13669), .o(n_13827) );
in01s01 g766855 ( .a(FE_OFN806_n_13742), .o(n_15643) );
oa12s01 g766856 ( .a(n_13686), .b(n_13685), .c(n_13684), .o(n_13742) );
in01s01 g766857 ( .a(n_14044), .o(n_14081) );
oa22s01 g766858 ( .a(n_13869), .b(FE_OCP_RBN5395_cordic_combinational_sub_ln23_0_unr12_z_0_), .c(n_13870), .d(FE_OCP_RBN5392_cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n_14044) );
in01s02 g766860 ( .a(n_13659), .o(n_13673) );
in01s02 g766861 ( .a(n_13661), .o(n_13659) );
no02f04 g766863 ( .a(n_13595), .b(n_13574), .o(n_13693) );
in01m02 g766864 ( .a(n_13629), .o(n_13630) );
na02m04 g766865 ( .a(n_13599), .b(n_13567), .o(n_13629) );
no02f04 g766866 ( .a(FE_OCP_RBN4151_n_13616), .b(FE_OCP_RBN4100_n_12880), .o(n_13644) );
na02m04 g766867 ( .a(n_13616), .b(FE_OCP_RBN4088_n_12880), .o(n_13635) );
no02f04 g766868 ( .a(FE_OCP_RBN1591_n_13557), .b(FE_OCP_RBN4087_n_12880), .o(n_13595) );
no02m02 g766869 ( .a(n_13557), .b(FE_OCP_RBN2540_n_12880), .o(n_13574) );
no02s01 g766870 ( .a(n_13976), .b(n_13937), .o(n_13977) );
na02s01 g766871 ( .a(n_14390), .b(n_14385), .o(n_14349) );
no02s01 g766872 ( .a(n_14347), .b(n_14350), .o(n_14348) );
no02s01 g766873 ( .a(n_14345), .b(n_14347), .o(n_14346) );
na02s01 g766874 ( .a(n_14008), .b(n_14042), .o(n_14080) );
in01s01 g766875 ( .a(n_14343), .o(n_14344) );
no02s01 g766876 ( .a(FE_OCP_RBN5802_n_13962), .b(n_14304), .o(n_14343) );
na02s01 g766877 ( .a(n_14390), .b(n_14298), .o(n_15247) );
in01s01 g766878 ( .a(n_14491), .o(n_14422) );
no02s01 g766879 ( .a(n_14216), .b(FE_OCP_RBN6699_n_13796), .o(n_14491) );
in01s01 g766880 ( .a(n_14421), .o(n_14488) );
no02s01 g766881 ( .a(n_14303), .b(FE_OCP_RBN6699_n_13796), .o(n_14421) );
no02s01 g766882 ( .a(n_14389), .b(n_14350), .o(n_15244) );
in01s01 g766883 ( .a(n_14341), .o(n_14342) );
na02s01 g766884 ( .a(n_14304), .b(FE_OCP_RBN5802_n_13962), .o(n_14341) );
no02s01 g766885 ( .a(n_13846), .b(n_14340), .o(n_14454) );
in01s01 g766886 ( .a(n_14339), .o(n_14456) );
na02s01 g766887 ( .a(n_14303), .b(n_14215), .o(n_14339) );
na02s01 g766888 ( .a(n_14216), .b(n_14215), .o(n_14306) );
in01s01 g766889 ( .a(n_14300), .o(n_14301) );
no02s01 g766890 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14259), .o(n_14300) );
na02s01 g766891 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14259), .o(n_14381) );
no02s01 g766892 ( .a(FE_OCP_RBN5802_n_13962), .b(n_13847), .o(n_14455) );
in01s01 g766893 ( .a(n_14425), .o(n_14388) );
no02s01 g766894 ( .a(n_13877), .b(FE_OCP_RBN4205_n_13796), .o(n_14425) );
no02s01 g766895 ( .a(n_13878), .b(FE_OCP_RBN5802_n_13962), .o(n_14426) );
no02s01 g766896 ( .a(n_13740), .b(n_13739), .o(n_13741) );
na02f04 g766897 ( .a(n_13642), .b(n_13683), .o(n_13712) );
na02f04 g766898 ( .a(n_13647), .b(FE_OFN5070_n_13646), .o(n_13705) );
na02s01 g766899 ( .a(n_13684), .b(n_13685), .o(n_13686) );
in01s01 g766900 ( .a(n_13657), .o(n_13658) );
no02m04 g766901 ( .a(n_13647), .b(FE_OFN5070_n_13646), .o(n_13657) );
ao12m02 g766902 ( .a(n_13793), .b(n_13848), .c(FE_OCP_RBN5394_cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n_13943) );
no02m03 TIMEBOOST_cell_8728 ( .a(n_45180), .b(n_40679), .o(TIMEBOOST_net_2851) );
no02s01 g766904 ( .a(n_14110), .b(n_14043), .o(n_14111) );
na02s02 g766905 ( .a(n_13906), .b(n_13938), .o(n_14009) );
na02f04 g766906 ( .a(n_13628), .b(n_13615), .o(n_13743) );
oa12f08 g766907 ( .a(n_13618), .b(n_13684), .c(n_13637), .o(n_13747) );
in01s01 g766908 ( .a(n_13907), .o(n_13908) );
oa12s01 g766909 ( .a(n_13826), .b(n_13825), .c(n_13824), .o(n_13907) );
in01m02 g766910 ( .a(n_13575), .o(n_13576) );
in01s02 g766911 ( .a(n_13560), .o(n_13575) );
oa12f08 g766912 ( .a(n_12683), .b(n_13459), .c(n_12658), .o(n_13560) );
na02f04 g766913 ( .a(n_13570), .b(n_13583), .o(n_13628) );
na02s02 g766914 ( .a(n_13582), .b(n_13589), .o(n_13615) );
na02s01 g766915 ( .a(n_14258), .b(n_14296), .o(n_14947) );
in01s01 g766916 ( .a(n_14110), .o(n_14008) );
na02s01 g766917 ( .a(n_13967), .b(n_13966), .o(n_14110) );
na02s01 g766918 ( .a(n_13971), .b(n_14042), .o(n_14043) );
in01s01 g766919 ( .a(n_13906), .o(n_13976) );
no02s01 g766920 ( .a(n_13892), .b(n_13903), .o(n_13906) );
no02s01 g766921 ( .a(n_13937), .b(n_13900), .o(n_13938) );
na02s01 g766922 ( .a(n_13864), .b(n_13863), .o(n_13865) );
no02s01 g766923 ( .a(n_13904), .b(n_13895), .o(n_13905) );
na02s01 g766924 ( .a(n_13973), .b(n_14006), .o(n_14007) );
na02s01 g766925 ( .a(n_14035), .b(n_14078), .o(n_14079) );
na02s01 g766926 ( .a(n_14292), .b(n_14386), .o(n_14387) );
in01s01 g766927 ( .a(n_14076), .o(n_14077) );
na02s01 g766928 ( .a(n_14041), .b(n_14040), .o(n_14076) );
no02s01 g766929 ( .a(n_13892), .b(n_13895), .o(n_14219) );
no02s01 g766930 ( .a(n_13970), .b(n_14036), .o(n_14565) );
na02s01 g766931 ( .a(n_13901), .b(n_13898), .o(n_14307) );
na02s01 g766932 ( .a(n_14041), .b(n_14138), .o(n_14700) );
na02s01 g766933 ( .a(n_13863), .b(n_13822), .o(n_14010) );
no02s01 g766934 ( .a(n_13972), .b(n_14109), .o(n_14620) );
na02s01 g766935 ( .a(n_14385), .b(n_14294), .o(n_15063) );
na02s01 g766936 ( .a(n_14258), .b(n_14386), .o(n_14992) );
na02s01 g766937 ( .a(n_13966), .b(n_14006), .o(n_14493) );
no02s01 g766938 ( .a(n_14293), .b(n_14208), .o(n_15029) );
na02s01 g766939 ( .a(n_14487), .b(n_14561), .o(n_15209) );
na02s01 g766940 ( .a(n_14212), .b(n_14206), .o(n_14838) );
no02s01 g766941 ( .a(n_13823), .b(n_13939), .o(n_13941) );
no02s01 g766942 ( .a(n_13974), .b(n_14037), .o(n_14530) );
no02s01 g766943 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14257), .o(n_14350) );
na02s01 g766944 ( .a(n_14209), .b(n_14211), .o(n_14299) );
in01s01 g766945 ( .a(n_13869), .o(n_13870) );
na02s01 g766946 ( .a(n_13794), .b(n_13848), .o(n_13869) );
no02s01 g766947 ( .a(n_13937), .b(n_13904), .o(n_14260) );
in01s01 g766948 ( .a(n_14345), .o(n_14298) );
no02s01 g766949 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14253), .o(n_14345) );
in01s01 g766950 ( .a(n_14297), .o(n_14389) );
na02s01 g766951 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14257), .o(n_14297) );
na02s01 g766952 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14253), .o(n_14390) );
no02s01 g766953 ( .a(n_14338), .b(n_14291), .o(n_14995) );
no02s01 g766954 ( .a(n_13903), .b(n_13902), .o(n_14083) );
no02s01 g766955 ( .a(n_13897), .b(n_14039), .o(n_14392) );
no02s01 g766956 ( .a(n_14075), .b(n_14171), .o(n_14756) );
na02s01 g766957 ( .a(n_14296), .b(n_14295), .o(n_14835) );
no02s01 g766958 ( .a(n_13670), .b(n_13643), .o(n_13740) );
no02s01 g766959 ( .a(n_13637), .b(n_13619), .o(n_13685) );
na02s01 g766960 ( .a(n_13825), .b(n_13824), .o(n_13826) );
in01s02 g766961 ( .a(n_13633), .o(n_13594) );
in01s01 g766971 ( .a(n_13683), .o(n_13739) );
no02s02 g766973 ( .a(n_13668), .b(n_13682), .o(n_15609) );
ao12s01 g766974 ( .a(n_13614), .b(n_13613), .c(n_13612), .o(n_15458) );
in01s01 g766975 ( .a(n_13846), .o(n_13847) );
ao12s01 g766976 ( .a(n_13768), .b(n_13767), .c(n_13766), .o(n_13846) );
oa12s01 g766983 ( .a(n_13799), .b(n_13798), .c(n_13797), .o(n_14304) );
in01s01 g766984 ( .a(n_13877), .o(n_13878) );
ao12s01 g766985 ( .a(n_13792), .b(n_13791), .c(n_13790), .o(n_13877) );
oa12s01 g766986 ( .a(n_13763), .b(n_13762), .c(n_13761), .o(n_14303) );
oa12s01 g766987 ( .a(n_13738), .b(n_13737), .c(n_13736), .o(n_14216) );
ao12s01 g766988 ( .a(n_13771), .b(n_13770), .c(n_13769), .o(n_14259) );
na02s06 TIMEBOOST_cell_4916 ( .a(n_1744), .b(n_1745), .o(TIMEBOOST_net_1406) );
no02s01 g766991 ( .a(n_13770), .b(n_13769), .o(n_13771) );
no02s01 g766992 ( .a(n_13767), .b(n_13766), .o(n_13768) );
in01f02 g766993 ( .a(n_13582), .o(n_13583) );
no02s01 TIMEBOOST_cell_2980 ( .a(n_28735), .b(n_28736), .o(TIMEBOOST_net_781) );
na02s01 g766995 ( .a(n_13737), .b(n_13736), .o(n_13738) );
na02s01 g766996 ( .a(n_13798), .b(n_13797), .o(n_13799) );
no02s02 TIMEBOOST_cell_4052 ( .a(TIMEBOOST_net_1116), .b(n_25418), .o(n_25454) );
na02s02 g766998 ( .a(n_13497), .b(FE_OCP_RBN2540_n_12880), .o(n_13573) );
na02s02 g766999 ( .a(n_13497), .b(FE_OCP_RBN2540_n_12880), .o(n_13567) );
no02s04 TIMEBOOST_cell_1918 ( .a(TIMEBOOST_net_573), .b(n_17452), .o(n_17513) );
in01s01 g767002 ( .a(n_14211), .o(n_14338) );
na02s01 g767003 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14170), .o(n_14211) );
na02m01 g767004 ( .a(n_13765), .b(n_13764), .o(n_13848) );
in01s01 g767005 ( .a(n_14213), .o(n_14075) );
na02s01 g767006 ( .a(FE_OCPN924_n_13962), .b(n_14038), .o(n_14213) );
in01s01 g767007 ( .a(n_14486), .o(n_14487) );
no02s01 g767008 ( .a(FE_RN_1486_0), .b(n_14207), .o(n_14486) );
na02s01 g767009 ( .a(FE_OCP_RBN5802_n_13962), .b(n_13715), .o(n_14386) );
in01s01 g767010 ( .a(n_14137), .o(n_14138) );
no02s01 g767011 ( .a(FE_OCPN924_n_13962), .b(n_13975), .o(n_14137) );
in01s01 g767012 ( .a(n_14078), .o(n_14037) );
na02s01 g767013 ( .a(FE_OCP_RBN4200_n_13796), .b(n_13936), .o(n_14078) );
no02s01 g767014 ( .a(FE_OCP_RBN4188_n_13765), .b(n_13325), .o(n_13904) );
in01s01 g767015 ( .a(n_14171), .o(n_14136) );
no02s01 g767016 ( .a(FE_OCPN924_n_13962), .b(n_14038), .o(n_14171) );
na02s01 g767017 ( .a(FE_OCP_RBN5802_n_13962), .b(n_13650), .o(n_14295) );
in01s01 g767018 ( .a(n_13864), .o(n_13823) );
na02s02 g767019 ( .a(n_13760), .b(n_13795), .o(n_13864) );
na02s02 g767020 ( .a(FE_OCP_RBN4188_n_13765), .b(n_13787), .o(n_13863) );
no02s01 g767021 ( .a(FE_OCP_RBN4188_n_13765), .b(n_13135), .o(n_13902) );
in01s01 g767022 ( .a(n_14108), .o(n_14109) );
na02s01 g767023 ( .a(FE_OCP_RBN6694_n_13796), .b(n_13961), .o(n_14108) );
in01s01 g767024 ( .a(n_14347), .o(n_14294) );
no02s01 g767025 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14256), .o(n_14347) );
in01s01 g767026 ( .a(n_14427), .o(n_14293) );
na02s01 g767027 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14168), .o(n_14427) );
in01s01 g767028 ( .a(n_14208), .o(n_14209) );
no02s01 g767029 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14168), .o(n_14208) );
na02s01 g767030 ( .a(FE_OCP_RBN2835_n_13962), .b(n_13714), .o(n_14258) );
na02s01 g767031 ( .a(FE_OCP_RBN2835_n_13962), .b(n_13649), .o(n_14296) );
na02s01 g767032 ( .a(FE_OCP_RBN2759_n_13796), .b(n_13975), .o(n_14041) );
na02s01 g767033 ( .a(FE_OCP_RBN2759_n_13796), .b(n_13501), .o(n_13966) );
in01s01 g767034 ( .a(n_13974), .o(n_14042) );
no02s01 g767035 ( .a(FE_OCP_RBN4189_n_13765), .b(n_13936), .o(n_13974) );
no02s01 g767036 ( .a(FE_OCP_RBN2756_n_13796), .b(n_13134), .o(n_13903) );
in01s01 g767037 ( .a(n_13900), .o(n_13901) );
no02s01 g767038 ( .a(FE_OCP_RBN2756_n_13796), .b(n_13875), .o(n_13900) );
no02m01 g767039 ( .a(FE_OCP_RBN4188_n_13765), .b(n_13795), .o(n_13939) );
in01s01 g767040 ( .a(n_13821), .o(n_13822) );
no02s01 g767041 ( .a(FE_OCP_RBN4188_n_13765), .b(n_13787), .o(n_13821) );
in01s01 g767042 ( .a(n_13973), .o(n_14039) );
na02s01 g767043 ( .a(FE_OCP_RBN4200_n_13796), .b(n_13893), .o(n_13973) );
in01s01 g767044 ( .a(n_14035), .o(n_14036) );
na02s01 g767045 ( .a(FE_OCP_RBN4200_n_13796), .b(n_13934), .o(n_14035) );
in01s01 g767046 ( .a(n_14291), .o(n_14292) );
no02s01 g767047 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14170), .o(n_14291) );
in01s01 g767048 ( .a(n_13895), .o(n_13876) );
no02s01 g767049 ( .a(FE_OCP_RBN4188_n_13765), .b(n_13289), .o(n_13895) );
na02s01 g767050 ( .a(FE_OCP_RBN4200_n_13796), .b(n_13502), .o(n_14006) );
in01s01 g767051 ( .a(n_13898), .o(n_13899) );
na02s01 g767052 ( .a(FE_OCP_RBN2756_n_13796), .b(n_13875), .o(n_13898) );
na02s01 g767053 ( .a(n_14215), .b(n_14207), .o(n_14561) );
in01s01 g767054 ( .a(n_13972), .o(n_14040) );
no02s01 g767055 ( .a(FE_OCP_RBN4200_n_13796), .b(n_13961), .o(n_13972) );
na02s01 g767056 ( .a(FE_OCPN924_n_13962), .b(n_14107), .o(n_14212) );
in01s01 g767057 ( .a(n_13970), .o(n_13971) );
no02s01 g767058 ( .a(FE_OCP_RBN4189_n_13765), .b(n_13934), .o(n_13970) );
no02s01 g767059 ( .a(FE_OCP_RBN2756_n_13796), .b(n_13324), .o(n_13937) );
na02s01 g767060 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14256), .o(n_14385) );
no02s01 g767061 ( .a(FE_OCP_RBN2756_n_13796), .b(n_13288), .o(n_13892) );
in01s01 g767062 ( .a(n_14205), .o(n_14206) );
no02s01 g767063 ( .a(FE_OCP_RBN2835_n_13962), .b(n_14107), .o(n_14205) );
in01s01 g767064 ( .a(n_13897), .o(n_13967) );
no02s01 g767065 ( .a(FE_OCP_RBN4189_n_13765), .b(n_13893), .o(n_13897) );
in01s01 g767066 ( .a(n_13793), .o(n_13794) );
no02m01 g767067 ( .a(n_13765), .b(n_13764), .o(n_13793) );
no02s01 g767068 ( .a(n_13624), .b(n_13639), .o(n_13668) );
no02s01 g767069 ( .a(n_13623), .b(n_13640), .o(n_13682) );
no02s01 g767070 ( .a(n_13612), .b(n_13613), .o(n_13614) );
in01s01 g767071 ( .a(n_13618), .o(n_13619) );
na02m04 g767072 ( .a(n_13591), .b(FE_OCPN5258_n_13590), .o(n_13618) );
in01s01 g767073 ( .a(n_13669), .o(n_13670) );
na02m06 g767074 ( .a(n_13598), .b(n_12586), .o(n_13669) );
no02m06 g767075 ( .a(n_13591), .b(FE_OCPN5258_n_13590), .o(n_13637) );
na02s01 g767076 ( .a(n_13762), .b(n_13761), .o(n_13763) );
in01s01 g767077 ( .a(n_13642), .o(n_13643) );
na02f04 g767078 ( .a(n_13597), .b(FE_OCP_DRV_N1452_n_12585), .o(n_13642) );
no02s01 g767079 ( .a(n_13791), .b(n_13790), .o(n_13792) );
oa12s01 g767080 ( .a(n_13611), .b(n_13610), .c(n_13609), .o(n_15462) );
oa12f08 g767081 ( .a(n_13578), .b(n_13612), .c(n_13517), .o(n_13684) );
oa12s01 g767082 ( .a(n_13287), .b(n_13699), .c(n_13378), .o(n_13825) );
ao12s01 g767083 ( .a(n_13719), .b(n_13718), .c(n_13717), .o(n_14257) );
ao12s01 g767084 ( .a(n_13735), .b(n_13734), .c(n_13733), .o(n_14253) );
no02s01 g767085 ( .a(n_13718), .b(n_13717), .o(n_13719) );
na02s01 g767086 ( .a(n_13610), .b(n_13609), .o(n_13611) );
na02s01 g767087 ( .a(n_13578), .b(n_13518), .o(n_13613) );
no02s01 g767089 ( .a(n_13734), .b(n_13733), .o(n_13735) );
in01m02 g767090 ( .a(n_13532), .o(n_13533) );
in01m01 g767091 ( .a(n_13513), .o(n_13532) );
no03m04 TIMEBOOST_cell_2646 ( .a(FE_OCP_RBN4338_n_9521), .b(n_9399), .c(n_9562), .o(n_9785) );
ao12f04 g767094 ( .a(FE_OCPN1240_n_13412), .b(n_13413), .c(FE_OCPN1242_n_12633), .o(n_13460) );
no02s02 TIMEBOOST_cell_1885 ( .a(n_39803), .b(n_39878), .o(TIMEBOOST_net_557) );
in01s06 g767145 ( .a(n_14524), .o(n_14618) );
in01f03 g767148 ( .a(n_14420), .o(n_14524) );
in01s40 g767153 ( .a(FE_OCP_RBN2837_n_13962), .o(n_14420) );
in01f01 g767161 ( .a(n_14452), .o(n_14650) );
in01s06 g767192 ( .a(n_14730), .o(n_14805) );
in01s06 g767195 ( .a(n_14588), .o(n_14730) );
in01s10 g767200 ( .a(FE_RN_1486_0), .o(n_14588) );
in01s06 g767204 ( .a(FE_RN_1486_0), .o(n_14452) );
in01s06 g767205 ( .a(FE_OCP_RBN2832_n_13962), .o(FE_RN_1486_0) );
in01s03 g767213 ( .a(n_14215), .o(n_14340) );
in01s06 g767214 ( .a(FE_OCP_RBN2833_n_13962), .o(n_14215) );
in01s01 g767231 ( .a(n_13765), .o(n_13760) );
na03m08 TIMEBOOST_cell_7365 ( .a(FE_RN_1554_0), .b(FE_RN_1555_0), .c(n_18178), .o(n_18224) );
oa12s01 g767233 ( .a(n_13252), .b(n_13696), .c(n_13249), .o(n_13770) );
ao12s01 g767234 ( .a(n_13157), .b(n_13716), .c(n_13284), .o(n_13767) );
no02s02 TIMEBOOST_cell_1867 ( .a(n_40009), .b(FE_OCP_RBN6154_n_39816), .o(TIMEBOOST_net_548) );
no02s01 g767236 ( .a(n_13701), .b(n_13285), .o(n_13791) );
ao12s01 g767237 ( .a(n_13210), .b(n_13697), .c(n_13248), .o(n_13737) );
no02m06 TIMEBOOST_cell_4089 ( .a(n_39193), .b(n_39104), .o(TIMEBOOST_net_1135) );
na02m02 g767239 ( .a(n_13535), .b(n_13530), .o(n_13536) );
no02s04 TIMEBOOST_cell_8126 ( .a(n_21538), .b(n_21731), .o(TIMEBOOST_net_2694) );
in01m02 g767243 ( .a(n_13597), .o(n_13598) );
no03m06 TIMEBOOST_cell_6542 ( .a(n_35274), .b(FE_OCP_RBN5973_n_35231), .c(n_35352), .o(TIMEBOOST_net_1998) );
in01s01 g767245 ( .a(n_13639), .o(n_13640) );
oa12s01 g767246 ( .a(n_13588), .b(n_13626), .c(FE_RN_1759_0), .o(n_13639) );
in01s01 g767247 ( .a(n_13623), .o(n_13624) );
oa12s01 g767248 ( .a(n_13525), .b(n_13568), .c(n_13608), .o(n_13623) );
oa22s01 g767249 ( .a(n_13697), .b(n_13274), .c(n_13716), .d(n_13275), .o(n_14207) );
ao12s01 g767250 ( .a(n_13681), .b(n_13680), .c(n_13679), .o(n_14168) );
oa12s01 g767251 ( .a(n_13542), .b(n_13541), .c(n_13540), .o(n_15337) );
in01s01 g767254 ( .a(n_13562), .o(n_13563) );
in01m01 g767258 ( .a(n_13497), .o(n_13562) );
no02m04 g767263 ( .a(n_13512), .b(n_13488), .o(n_13591) );
oa12s01 g767264 ( .a(n_13202), .b(n_13716), .c(n_13088), .o(n_13762) );
in01s01 g767266 ( .a(n_13570), .o(n_13589) );
in01s01 g767267 ( .a(n_13559), .o(n_13570) );
in01s02 g767268 ( .a(n_13559), .o(n_13558) );
na02f06 g767269 ( .a(n_13490), .b(n_13458), .o(n_13559) );
na02f04 g767270 ( .a(n_13430), .b(n_12891), .o(n_13458) );
na03m40 TIMEBOOST_cell_8195 ( .a(FE_RN_1566_0), .b(delay_xor_ln22_unr15_stage6_stallmux_q_13_), .c(FE_OCP_RBN6540_n_44083), .o(FE_RN_1567_0) );
no02s06 TIMEBOOST_cell_1886 ( .a(TIMEBOOST_net_557), .b(n_39937), .o(n_39938) );
na02f04 g767273 ( .a(n_13431), .b(n_12890), .o(n_13490) );
no02s01 g767274 ( .a(n_13716), .b(n_13700), .o(n_13701) );
na02f02 g767275 ( .a(n_13489), .b(FE_OCP_RBN4112_n_12880), .o(n_13530) );
in01s01 g767278 ( .a(n_13698), .o(n_13699) );
no02s01 g767279 ( .a(n_13697), .b(n_13379), .o(n_13698) );
no02m02 g767281 ( .a(n_13436), .b(n_13429), .o(n_13512) );
no02m02 g767282 ( .a(n_13456), .b(n_13388), .o(n_13488) );
na02s01 g767283 ( .a(n_13541), .b(n_13540), .o(n_13542) );
no02s01 g767284 ( .a(n_13608), .b(n_13569), .o(n_13610) );
na02s01 g767285 ( .a(n_13626), .b(FE_RN_1759_0), .o(n_13588) );
na02s01 TIMEBOOST_cell_2974 ( .a(n_13422), .b(n_13391), .o(TIMEBOOST_net_778) );
na02m06 g767287 ( .a(n_13511), .b(FE_OCPN1372_n_13510), .o(n_13578) );
no02f06 g767288 ( .a(n_13569), .b(n_13547), .o(n_13606) );
in01s01 g767289 ( .a(n_13517), .o(n_13518) );
no02m06 g767290 ( .a(n_13511), .b(FE_OCPN1372_n_13510), .o(n_13517) );
no02s01 g767291 ( .a(n_13680), .b(n_13679), .o(n_13681) );
no02m06 TIMEBOOST_cell_4943 ( .a(TIMEBOOST_net_1419), .b(n_33072), .o(n_33191) );
ao12s01 g767294 ( .a(n_13080), .b(n_13678), .c(n_13115), .o(n_13718) );
na02f08 TIMEBOOST_cell_4997 ( .a(TIMEBOOST_net_1446), .b(n_41353), .o(n_41355) );
na02s01 g767296 ( .a(n_13696), .b(n_13036), .o(n_13734) );
ao12f01 g767297 ( .a(n_13550), .b(n_13549), .c(n_13548), .o(n_15342) );
oa12f06 g767298 ( .a(n_13500), .b(n_13468), .c(n_13451), .o(n_13612) );
oa12s01 g767299 ( .a(n_13676), .b(n_13675), .c(n_13674), .o(n_14170) );
in01s01 g767300 ( .a(n_13714), .o(n_13715) );
oa12s01 g767301 ( .a(n_13653), .b(n_13652), .c(n_13651), .o(n_13714) );
ao12s01 g767302 ( .a(n_13672), .b(n_13678), .c(n_13671), .o(n_14256) );
na02s01 g767303 ( .a(n_13675), .b(n_13674), .o(n_13676) );
no02s01 g767304 ( .a(n_13678), .b(n_13671), .o(n_13672) );
na02s01 g767305 ( .a(n_13652), .b(n_13651), .o(n_13653) );
na02s01 g767306 ( .a(n_13452), .b(n_13500), .o(n_13541) );
no02s01 g767307 ( .a(n_13549), .b(n_13548), .o(n_13550) );
in01m02 g767308 ( .a(n_13538), .o(n_13608) );
na02f04 g767309 ( .a(n_13496), .b(FE_OCP_DRV_N5360_n_13495), .o(n_13538) );
in01s01 g767310 ( .a(n_13569), .o(n_13525) );
no02f06 g767311 ( .a(n_13496), .b(FE_OCP_DRV_N5360_n_13495), .o(n_13569) );
in01m02 g767312 ( .a(n_13410), .o(n_13411) );
in01m02 g767313 ( .a(n_13413), .o(n_13410) );
in01f02 g767315 ( .a(n_13430), .o(n_13431) );
in01m02 g767316 ( .a(n_13409), .o(n_13430) );
oa12f06 g767317 ( .a(n_12809), .b(n_13336), .c(n_12731), .o(n_13409) );
in01s01 g767318 ( .a(n_13697), .o(n_13716) );
oa12f08 g767319 ( .a(n_13347), .b(n_13636), .c(n_13316), .o(n_13697) );
no02s04 TIMEBOOST_cell_2006 ( .a(TIMEBOOST_net_617), .b(n_7990), .o(n_9304) );
oa12s01 g767321 ( .a(n_13039), .b(n_13638), .c(n_13312), .o(n_13680) );
in01m02 g767323 ( .a(n_13436), .o(n_13456) );
oa12m04 g767325 ( .a(FE_OCP_RBN4112_n_12880), .b(n_13407), .c(n_13453), .o(n_13535) );
na02f02 TIMEBOOST_cell_8761 ( .a(TIMEBOOST_net_2867), .b(n_8270), .o(n_8390) );
no02f04 g767327 ( .a(n_13508), .b(n_13482), .o(n_13626) );
ao12s01 g767328 ( .a(n_13493), .b(n_13492), .c(n_13491), .o(n_15223) );
in01s01 g767329 ( .a(n_13429), .o(n_13487) );
in01m01 g767333 ( .a(n_13388), .o(n_13429) );
in01s01 g767335 ( .a(n_13568), .o(n_13609) );
in01s01 g767336 ( .a(n_13547), .o(n_13568) );
no02s01 TIMEBOOST_cell_1985 ( .a(n_6704), .b(n_6765), .o(TIMEBOOST_net_607) );
no02s02 TIMEBOOST_cell_6756 ( .a(TIMEBOOST_net_2135), .b(n_39097), .o(n_39209) );
in01m02 g767345 ( .a(n_13489), .o(n_13483) );
na02s01 g767348 ( .a(n_13636), .b(n_13256), .o(n_13678) );
no02s06 TIMEBOOST_cell_2007 ( .a(n_33827), .b(n_33855), .o(TIMEBOOST_net_618) );
no02m02 g767350 ( .a(n_13446), .b(n_13453), .o(n_13482) );
na02m03 TIMEBOOST_cell_1947 ( .a(FE_OCP_RBN3980_n_32436), .b(n_32439), .o(TIMEBOOST_net_588) );
no02m04 g767353 ( .a(n_13447), .b(FE_OCP_RBN4083_n_13453), .o(n_13508) );
no02s01 g767354 ( .a(n_13507), .b(n_13480), .o(n_13549) );
no02s01 g767355 ( .a(n_13492), .b(n_13491), .o(n_13493) );
na02m04 g767356 ( .a(n_13435), .b(n_13434), .o(n_13500) );
na02m04 g767357 ( .a(n_13390), .b(n_13385), .o(n_13408) );
no02s01 TIMEBOOST_cell_1986 ( .a(n_7527), .b(TIMEBOOST_net_607), .o(n_7603) );
no02s02 TIMEBOOST_cell_6755 ( .a(n_38608), .b(FE_OCP_RBN4328_n_38878), .o(TIMEBOOST_net_2135) );
in01s01 g767360 ( .a(n_13451), .o(n_13452) );
no02f04 g767361 ( .a(n_13435), .b(n_13434), .o(n_13451) );
no02s02 TIMEBOOST_cell_1861 ( .a(n_40011), .b(FE_OCP_RBN6154_n_39816), .o(TIMEBOOST_net_545) );
oa12s01 g767363 ( .a(n_13621), .b(n_13620), .c(n_13150), .o(n_13652) );
in01s01 g767364 ( .a(n_13649), .o(n_13650) );
oa12s01 g767365 ( .a(n_13603), .b(n_13620), .c(n_13602), .o(n_13649) );
oa12s01 g767366 ( .a(n_13450), .b(n_13449), .c(n_13448), .o(n_15207) );
in01s01 g767367 ( .a(n_13468), .o(n_13540) );
ao12f06 g767368 ( .a(n_13417), .b(n_13397), .c(n_13383), .o(n_13468) );
no02m04 TIMEBOOST_cell_7488 ( .a(n_12499), .b(n_12238), .o(TIMEBOOST_net_2375) );
oa12s01 g767370 ( .a(n_13586), .b(n_13585), .c(n_13584), .o(n_14107) );
na02s01 g767371 ( .a(n_13587), .b(n_13164), .o(n_13638) );
na02s01 g767372 ( .a(n_13620), .b(n_13602), .o(n_13603) );
no02f06 g767373 ( .a(n_13399), .b(n_12437), .o(n_13507) );
na03f06 TIMEBOOST_cell_8317 ( .a(n_14918), .b(n_14843), .c(n_14954), .o(n_15066) );
na02s01 g767375 ( .a(n_13449), .b(n_13448), .o(n_13450) );
no02s01 g767376 ( .a(n_13417), .b(n_13384), .o(n_13492) );
no02m04 g767377 ( .a(n_13398), .b(FE_OCP_DRV_N5358_n_12436), .o(n_13480) );
na02f04 g767378 ( .a(n_13361), .b(n_13301), .o(n_13386) );
na02s01 g767379 ( .a(n_13585), .b(n_13584), .o(n_13586) );
in01s02 g767380 ( .a(n_13298), .o(n_13299) );
in01m01 g767381 ( .a(n_13270), .o(n_13298) );
ao12f06 g767382 ( .a(n_12558), .b(n_13139), .c(n_12576), .o(n_13270) );
in01s02 g767383 ( .a(n_13343), .o(n_13344) );
in01s02 g767384 ( .a(n_13336), .o(n_13343) );
ao12f08 g767385 ( .a(n_12695), .b(n_13235), .c(n_12733), .o(n_13336) );
in01m02 g767386 ( .a(n_13446), .o(n_13447) );
in01m02 g767387 ( .a(n_13433), .o(n_13446) );
na02m04 g767388 ( .a(n_13406), .b(n_13405), .o(n_13407) );
na02m04 g767389 ( .a(n_13406), .b(n_13405), .o(n_13433) );
in01s02 g767390 ( .a(n_13390), .o(n_13362) );
na02m08 g767391 ( .a(n_13310), .b(n_13244), .o(n_13390) );
na02f08 g767392 ( .a(n_13587), .b(n_13313), .o(n_13636) );
in01s01 g767397 ( .a(n_13478), .o(n_13479) );
ao12s01 g767398 ( .a(n_13402), .b(n_13401), .c(n_13400), .o(n_13478) );
oa12s01 g767399 ( .a(n_13522), .b(n_13521), .c(n_13520), .o(n_13975) );
in01s01 g767400 ( .a(n_13385), .o(n_14543) );
in01s02 g767401 ( .a(n_13365), .o(n_13385) );
in01s02 g767402 ( .a(n_13335), .o(n_13365) );
no02s06 TIMEBOOST_cell_6301 ( .a(n_35591), .b(n_36075), .o(TIMEBOOST_net_2002) );
ao12f06 g767405 ( .a(n_13358), .b(n_13448), .c(n_13403), .o(n_13548) );
oa12s01 g767406 ( .a(n_13546), .b(n_13545), .c(n_13544), .o(n_14038) );
na02s01 g767407 ( .a(n_13545), .b(n_13544), .o(n_13546) );
na02s04 g767408 ( .a(n_13334), .b(FE_OCP_RBN4110_n_12880), .o(n_13405) );
no02s02 TIMEBOOST_cell_5127 ( .a(TIMEBOOST_net_1511), .b(FE_RN_893_0), .o(FE_RN_894_0) );
na03m06 TIMEBOOST_cell_4747 ( .a(n_20795), .b(n_20761), .c(n_20793), .o(n_20878) );
na02s04 g767411 ( .a(n_13232), .b(FE_OCP_RBN2519_n_12721), .o(n_13244) );
na02s01 g767412 ( .a(n_13359), .b(n_13403), .o(n_13449) );
no02s04 g767413 ( .a(n_13367), .b(n_13366), .o(n_13417) );
no02s01 g767414 ( .a(n_13401), .b(n_13400), .o(n_13402) );
in01s01 g767415 ( .a(n_13383), .o(n_13384) );
na02m04 g767416 ( .a(n_13367), .b(n_13366), .o(n_13383) );
na02s01 g767417 ( .a(n_13521), .b(n_13520), .o(n_13522) );
in01s06 g767418 ( .a(n_13361), .o(n_13406) );
na02f08 g767420 ( .a(n_13268), .b(n_13332), .o(n_13361) );
oa12s01 g767421 ( .a(n_13171), .b(n_13472), .c(n_13200), .o(n_13585) );
oa12s01 g767423 ( .a(n_13396), .b(n_13395), .c(n_13394), .o(n_13476) );
ao12s01 g767424 ( .a(n_13475), .b(n_13474), .c(n_13473), .o(n_13934) );
in01s01 g767425 ( .a(n_13587), .o(n_13620) );
no02s02 TIMEBOOST_cell_1998 ( .a(n_44869), .b(TIMEBOOST_net_613), .o(n_37911) );
in01f02 g767427 ( .a(n_13398), .o(n_13399) );
ao12s01 g767429 ( .a(n_13506), .b(n_13505), .c(n_13504), .o(n_13961) );
in01s01 g767430 ( .a(n_13397), .o(n_13491) );
no02s01 g767432 ( .a(n_13494), .b(n_13208), .o(n_13545) );
na02m04 g767433 ( .a(n_13228), .b(n_12910), .o(n_13268) );
na02s01 g767434 ( .a(n_13360), .b(n_13338), .o(n_13401) );
na02s01 g767436 ( .a(n_13395), .b(n_13394), .o(n_13396) );
no02s01 g767437 ( .a(n_13505), .b(n_13504), .o(n_13506) );
na02m04 g767438 ( .a(n_13331), .b(FE_OCP_DRV_N6273_n_13330), .o(n_13403) );
in01s01 g767439 ( .a(n_13358), .o(n_13359) );
no02s04 g767440 ( .a(n_13331), .b(FE_OCP_DRV_N6273_n_13330), .o(n_13358) );
no02s01 g767441 ( .a(n_13474), .b(n_13473), .o(n_13475) );
in01m02 g767442 ( .a(n_13175), .o(n_13176) );
in01s01 g767443 ( .a(n_13139), .o(n_13175) );
oa12m08 g767444 ( .a(n_12563), .b(n_13009), .c(n_12549), .o(n_13139) );
in01m02 g767445 ( .a(n_13266), .o(n_13267) );
in01s01 g767446 ( .a(n_13235), .o(n_13266) );
oa12m08 g767447 ( .a(n_12697), .b(n_13097), .c(n_12656), .o(n_13235) );
no02s01 TIMEBOOST_cell_1995 ( .a(n_37871), .b(n_37882), .o(TIMEBOOST_net_612) );
in01s02 g767449 ( .a(n_13310), .o(n_13269) );
no02m08 g767450 ( .a(n_13229), .b(n_13153), .o(n_13310) );
oa12s01 g767451 ( .a(n_12951), .b(n_13462), .c(n_13033), .o(n_13521) );
in01m02 g767452 ( .a(n_13334), .o(n_13301) );
in01s01 g767453 ( .a(n_13301), .o(n_13329) );
no02s01 TIMEBOOST_cell_5120 ( .a(n_14421), .b(n_14491), .o(TIMEBOOST_net_1508) );
in01s01 g767458 ( .a(n_14968), .o(n_14966) );
oa12s01 g767459 ( .a(n_13297), .b(n_13296), .c(n_13295), .o(n_14968) );
in01m02 g767461 ( .a(n_13272), .o(n_13273) );
in01m02 g767462 ( .a(n_13232), .o(n_13272) );
oa12f06 g767464 ( .a(n_13302), .b(n_13394), .c(n_13357), .o(n_13448) );
ao12s01 g767465 ( .a(n_13445), .b(n_13444), .c(n_13443), .o(n_13936) );
in01s01 g767466 ( .a(n_13501), .o(n_13502) );
oa12s01 g767467 ( .a(n_13427), .b(n_13426), .c(n_13425), .o(n_13501) );
no02s01 g767468 ( .a(n_13444), .b(n_13443), .o(n_13445) );
na02s01 g767469 ( .a(n_13426), .b(n_13425), .o(n_13427) );
no02s06 g767470 ( .a(n_13098), .b(n_12790), .o(n_13153) );
na02s01 g767471 ( .a(n_13296), .b(n_13295), .o(n_13297) );
no02s01 g767472 ( .a(n_13303), .b(n_13357), .o(n_13395) );
na02s06 g767473 ( .a(n_13226), .b(n_12322), .o(n_13360) );
na02s01 g767474 ( .a(n_13462), .b(n_12999), .o(n_13505) );
no02s20 TIMEBOOST_cell_6862 ( .a(FE_OCP_RBN3963_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(TIMEBOOST_net_2189), .o(FE_RN_158_0) );
na02m02 g767476 ( .a(n_13229), .b(n_13098), .o(n_13230) );
na02m02 g767477 ( .a(n_13225), .b(n_12321), .o(n_13338) );
in01s01 g767478 ( .a(n_13494), .o(n_13472) );
no02f08 g767479 ( .a(n_13462), .b(n_13166), .o(n_13494) );
ao12f08 g767480 ( .a(FE_OCP_RBN2580_n_13154), .b(FE_OCP_RBN2555_n_13141), .c(n_12881), .o(n_13332) );
na02f04 g767481 ( .a(n_13234), .b(n_13154), .o(n_13294) );
ao12s01 g767482 ( .a(n_12844), .b(n_13393), .c(n_12963), .o(n_13474) );
in01s01 g767484 ( .a(n_13293), .o(n_14555) );
in01m04 g767485 ( .a(n_13245), .o(n_13293) );
in01m04 g767486 ( .a(n_13228), .o(n_13245) );
ao12s01 g767489 ( .a(n_13292), .b(n_13291), .c(n_13290), .o(n_14977) );
oa12m04 g767490 ( .a(n_13142), .b(n_13227), .c(n_13295), .o(n_13400) );
in01m02 g767492 ( .a(n_13097), .o(n_13151) );
oa12m08 g767493 ( .a(n_12640), .b(n_12948), .c(n_12622), .o(n_13097) );
no02s01 g767494 ( .a(n_13393), .b(n_12788), .o(n_13444) );
na02f04 g767495 ( .a(FE_OCP_RBN2556_n_13141), .b(n_12910), .o(n_13234) );
no02s01 g767496 ( .a(n_13291), .b(n_13290), .o(n_13292) );
in01s01 g767497 ( .a(n_13302), .o(n_13303) );
na02s04 g767498 ( .a(n_13265), .b(FE_OCP_DRV_N6271_n_13264), .o(n_13302) );
no02s01 g767499 ( .a(n_13143), .b(n_13227), .o(n_13296) );
no02m04 g767500 ( .a(n_13265), .b(FE_OCP_DRV_N6271_n_13264), .o(n_13357) );
in01m02 g767501 ( .a(n_13059), .o(n_13060) );
in01m01 g767502 ( .a(n_13009), .o(n_13059) );
ao12m08 g767503 ( .a(n_12502), .b(n_12904), .c(n_12522), .o(n_13009) );
na02f08 g767504 ( .a(n_13393), .b(n_13037), .o(n_13462) );
oa12s01 g767505 ( .a(n_12774), .b(n_13382), .c(n_12982), .o(n_13426) );
na02m06 g767506 ( .a(n_13146), .b(n_13057), .o(n_13229) );
no02m02 g767507 ( .a(n_13144), .b(n_13058), .o(n_13145) );
ao12s01 g767508 ( .a(n_13355), .b(n_13382), .c(n_13354), .o(n_13893) );
in01s01 g767509 ( .a(n_14733), .o(n_14896) );
oa12s01 g767510 ( .a(n_13223), .b(n_13222), .c(n_13221), .o(n_14733) );
in01s02 g767514 ( .a(n_13098), .o(n_13148) );
in01s02 g767517 ( .a(n_13225), .o(n_13226) );
in01s01 g767519 ( .a(n_13057), .o(n_13058) );
na02m04 g767520 ( .a(n_12981), .b(FE_OCP_RBN2519_n_12721), .o(n_13057) );
in01s01 g767521 ( .a(n_13142), .o(n_13143) );
na02s02 g767522 ( .a(n_13096), .b(n_13095), .o(n_13142) );
no02s01 g767523 ( .a(n_13224), .b(n_13183), .o(n_13291) );
na02s01 g767524 ( .a(n_13222), .b(n_13221), .o(n_13223) );
no02s01 g767526 ( .a(n_13382), .b(n_13354), .o(n_13355) );
no02m02 g767527 ( .a(n_13096), .b(n_13095), .o(n_13227) );
oa12m02 g767528 ( .a(n_12617), .b(n_12983), .c(n_12975), .o(n_13008) );
no03s40 TIMEBOOST_cell_2177 ( .a(n_32635), .b(n_32731), .c(n_32754), .o(n_32772) );
no02f08 g767530 ( .a(n_13382), .b(n_12995), .o(n_13393) );
no02f08 g767534 ( .a(n_13006), .b(FE_OCP_RBN6577_n_13011), .o(n_13154) );
ao12s01 g767535 ( .a(n_13307), .b(n_13306), .c(n_13305), .o(n_13875) );
na02m04 g767536 ( .a(n_13094), .b(n_13063), .o(n_13265) );
in01s01 g767537 ( .a(FE_OCPN1398_n_14742), .o(n_14869) );
na02s01 g767538 ( .a(n_13140), .b(n_13093), .o(n_14742) );
in01s01 g767545 ( .a(n_13324), .o(n_13325) );
ao12s01 g767546 ( .a(n_13217), .b(n_13216), .c(n_13215), .o(n_13324) );
na02s01 g767547 ( .a(n_13322), .b(n_13193), .o(n_13323) );
no02s08 g767550 ( .a(n_12875), .b(n_12947), .o(n_12948) );
no02s02 TIMEBOOST_cell_1902 ( .a(TIMEBOOST_net_565), .b(n_11478), .o(n_11498) );
no02s01 g767552 ( .a(n_13306), .b(n_13305), .o(n_13307) );
no02s01 g767553 ( .a(n_13216), .b(n_13215), .o(n_13217) );
na02m02 g767554 ( .a(n_13011), .b(n_12987), .o(n_13063) );
na02m02 g767555 ( .a(FE_OCP_RBN6576_n_13011), .b(n_13005), .o(n_13094) );
no02f06 g767556 ( .a(n_13005), .b(n_13004), .o(n_13006) );
na02s01 g767557 ( .a(n_13053), .b(n_12796), .o(n_13140) );
na02s01 g767558 ( .a(n_13052), .b(n_12768), .o(n_13093) );
no02f02 g767559 ( .a(n_13050), .b(n_12283), .o(n_13183) );
no02s06 g767560 ( .a(n_13051), .b(n_12284), .o(n_13224) );
oa12m08 g767563 ( .a(n_12512), .b(n_12805), .c(n_12483), .o(n_12904) );
oa12s02 g767564 ( .a(n_12940), .b(FE_OCP_RBN2046_n_12907), .c(n_13004), .o(n_13144) );
no02m06 g767565 ( .a(n_12978), .b(n_12941), .o(n_13146) );
no02f08 g767566 ( .a(n_13239), .b(n_12924), .o(n_13382) );
in01m02 g767571 ( .a(n_12981), .o(n_13010) );
oa22m02 g767572 ( .a(n_12830), .b(n_12533), .c(n_12831), .d(n_12534), .o(n_12981) );
oa12s01 g767573 ( .a(n_13056), .b(n_13055), .c(n_13054), .o(n_13222) );
no02m04 g767574 ( .a(n_13002), .b(n_12826), .o(n_13295) );
in01s01 g767576 ( .a(n_13288), .o(n_13289) );
ao12s01 g767577 ( .a(n_13179), .b(n_13178), .c(n_13177), .o(n_13288) );
no02s01 g767578 ( .a(n_13470), .b(n_13377), .o(n_13424) );
no02f08 g767580 ( .a(n_13137), .b(n_12958), .o(n_13239) );
no02s01 g767581 ( .a(n_13178), .b(n_13177), .o(n_13179) );
no02m06 g767582 ( .a(FE_OCP_RBN2046_n_12907), .b(FE_OCP_RBN2522_n_12721), .o(n_12978) );
no02s02 g767583 ( .a(n_13087), .b(n_13262), .o(n_13322) );
no02s01 g767584 ( .a(n_13423), .b(n_13470), .o(n_13471) );
na02s01 g767585 ( .a(n_13055), .b(n_13054), .o(n_13056) );
in01m03 g767587 ( .a(n_12875), .o(n_12983) );
ao12f08 g767588 ( .a(n_12555), .b(n_12802), .c(n_12583), .o(n_12875) );
no02f08 TIMEBOOST_cell_8484 ( .a(FE_RN_2466_0), .b(FE_RN_2463_0), .o(TIMEBOOST_net_2729) );
oa12s01 g767590 ( .a(n_12923), .b(n_13100), .c(n_12776), .o(n_13216) );
no03m03 TIMEBOOST_cell_4587 ( .a(n_17339), .b(FE_OCP_RBN5511_n_44365), .c(delay_xor_ln22_unr12_stage5_stallmux_q_6_), .o(TIMEBOOST_net_68) );
no02s01 TIMEBOOST_cell_5937 ( .a(n_24105), .b(n_22788), .o(TIMEBOOST_net_1820) );
in01s01 g767595 ( .a(n_13052), .o(n_13053) );
oa12s01 g767596 ( .a(n_12943), .b(n_12949), .c(n_12942), .o(n_13052) );
in01s02 g767597 ( .a(n_13050), .o(n_13051) );
oa22f02 g767598 ( .a(n_12977), .b(n_12902), .c(n_12845), .d(n_12879), .o(n_13050) );
no02m02 g767599 ( .a(n_12784), .b(n_12980), .o(n_13002) );
in01s01 g767601 ( .a(n_14153), .o(n_13048) );
in01m01 g767602 ( .a(n_13005), .o(n_14153) );
in01m01 g767603 ( .a(n_13005), .o(n_12987) );
na02s01 g767605 ( .a(n_13422), .b(n_13421), .o(n_13423) );
no03m10 TIMEBOOST_cell_8212 ( .a(n_18075), .b(n_18226), .c(n_18204), .o(n_18302) );
in01s01 g767607 ( .a(n_13190), .o(n_13262) );
no02s01 g767608 ( .a(n_13047), .b(n_13138), .o(n_13190) );
na02s01 g767609 ( .a(n_13100), .b(n_12832), .o(n_13178) );
no02s01 g767610 ( .a(n_13700), .b(n_13286), .o(n_13287) );
no02m01 TIMEBOOST_cell_1895 ( .a(FE_OCP_RBN3226_n_39575), .b(FE_OCP_RBN3342_n_39942), .o(TIMEBOOST_net_562) );
na02s01 g767612 ( .a(n_12949), .b(n_12942), .o(n_12943) );
in01s02 g767613 ( .a(n_12830), .o(n_12831) );
in01s01 g767614 ( .a(n_12805), .o(n_12830) );
ao12m08 g767615 ( .a(n_12479), .b(n_12713), .c(n_12506), .o(n_12805) );
in01f06 g767616 ( .a(n_13136), .o(n_13137) );
na02s06 TIMEBOOST_cell_8035 ( .a(TIMEBOOST_net_2648), .b(n_20482), .o(n_20713) );
na02m02 TIMEBOOST_cell_5658 ( .a(n_11294), .b(n_11260), .o(TIMEBOOST_net_1777) );
in01m02 g767620 ( .a(n_12940), .o(n_12941) );
in01m02 g767621 ( .a(n_12888), .o(n_12940) );
in01m01 g767622 ( .a(n_12888), .o(n_12889) );
na02m04 g767623 ( .a(n_12803), .b(n_12849), .o(n_12888) );
ao12m06 g767624 ( .a(n_13253), .b(n_13346), .c(n_13315), .o(n_13347) );
in01s01 g767625 ( .a(n_12980), .o(n_13055) );
na02m02 g767626 ( .a(n_12866), .b(n_12829), .o(n_12980) );
na02s02 TIMEBOOST_cell_6337 ( .a(FE_OCP_RBN6880_n_31819), .b(FE_OCP_RBN6008_n_30608), .o(TIMEBOOST_net_2020) );
in01s01 g767628 ( .a(n_13134), .o(n_13135) );
ao12s01 g767629 ( .a(n_13020), .b(n_13019), .c(n_13018), .o(n_13134) );
oa12s01 g767630 ( .a(n_12939), .b(n_12938), .c(n_12937), .o(n_13787) );
na02m06 g767637 ( .a(n_12804), .b(n_12772), .o(n_12907) );
no02s01 g767638 ( .a(n_13369), .b(n_13392), .o(n_13442) );
na02m02 g767639 ( .a(n_12745), .b(n_12521), .o(n_12772) );
na02m04 g767640 ( .a(n_12746), .b(n_12520), .o(n_12804) );
na02f08 g767641 ( .a(n_13019), .b(n_12815), .o(n_13100) );
no02s01 g767642 ( .a(n_13019), .b(n_13018), .o(n_13020) );
na02s01 g767643 ( .a(n_12938), .b(n_12937), .o(n_12939) );
na02s01 g767644 ( .a(n_13284), .b(n_13243), .o(n_13285) );
na02s04 g767645 ( .a(n_13156), .b(n_13192), .o(n_13700) );
na02m02 g767646 ( .a(n_12771), .b(n_12753), .o(n_12803) );
na02s02 g767647 ( .a(n_12825), .b(n_12849), .o(n_12866) );
na02s02 g767648 ( .a(n_12770), .b(n_12808), .o(n_12829) );
oa12f08 g767651 ( .a(n_12564), .b(n_12727), .c(n_12539), .o(n_12802) );
na02m04 g767652 ( .a(n_13284), .b(n_13242), .o(n_13379) );
in01f04 g767653 ( .a(n_12879), .o(n_12977) );
na02f10 TIMEBOOST_cell_8631 ( .a(TIMEBOOST_net_2802), .b(n_39165), .o(n_39290) );
no03f10 TIMEBOOST_cell_7111 ( .a(TIMEBOOST_net_1830), .b(FE_RN_946_0), .c(FE_RN_945_0), .o(n_46964) );
oa12s01 g767657 ( .a(FE_OCP_RBN2561_n_13084), .b(n_13377), .c(delay_sub_ln21_0_unr8_stage4_stallmux_q_29_), .o(n_13422) );
ao12s01 g767658 ( .a(n_12823), .b(n_13000), .c(n_13013), .o(n_13047) );
in01s01 g767661 ( .a(n_12845), .o(n_12877) );
in01m01 g767663 ( .a(n_12902), .o(n_12845) );
no02s01 g767667 ( .a(n_13281), .b(n_13280), .o(n_13282) );
in01s01 g767668 ( .a(n_13391), .o(n_13392) );
no02s01 g767669 ( .a(n_13356), .b(n_13371), .o(n_13391) );
in01s01 g767672 ( .a(n_13260), .o(n_13261) );
na02m01 g767673 ( .a(n_13238), .b(n_13777), .o(n_13260) );
in01s01 g767674 ( .a(n_13351), .o(n_13352) );
no02s01 g767675 ( .a(n_13281), .b(n_13278), .o(n_13351) );
in01s01 g767676 ( .a(n_13375), .o(n_13376) );
no02s01 g767677 ( .a(n_13377), .b(n_13356), .o(n_13375) );
na02s01 g767678 ( .a(n_13203), .b(n_12271), .o(n_13259) );
in01s01 g767679 ( .a(n_13463), .o(n_13464) );
na02s01 g767680 ( .a(n_13421), .b(n_13370), .o(n_13463) );
no02s02 g767681 ( .a(n_13083), .b(n_13173), .o(n_13180) );
na02s03 g767682 ( .a(n_13213), .b(n_13099), .o(n_13172) );
in01s01 g767683 ( .a(n_13022), .o(n_13023) );
na02s01 g767684 ( .a(n_12956), .b(n_13000), .o(n_13022) );
na02s01 g767686 ( .a(n_13193), .b(n_13121), .o(n_13257) );
in01s01 g767687 ( .a(n_13132), .o(n_13133) );
na02s01 g767688 ( .a(n_12969), .b(n_13101), .o(n_13132) );
in01s01 g767689 ( .a(n_12961), .o(n_12962) );
na02s02 g767690 ( .a(n_12867), .b(n_47250), .o(n_12961) );
na02s01 g767692 ( .a(n_12824), .b(n_12900), .o(n_12935) );
no02s02 g767693 ( .a(n_12807), .b(n_12869), .o(n_12864) );
no02s06 g767694 ( .a(n_13256), .b(n_13255), .o(n_13346) );
na02s02 g767695 ( .a(n_13168), .b(n_13236), .o(n_13286) );
no02s02 g767696 ( .a(n_13160), .b(n_13241), .o(n_13242) );
in01s01 g767697 ( .a(n_13156), .o(n_13157) );
no02s03 g767698 ( .a(n_13088), .b(n_13040), .o(n_13156) );
no02s01 g767699 ( .a(n_13208), .b(n_13197), .o(n_13171) );
no02s01 TIMEBOOST_cell_5513 ( .a(TIMEBOOST_net_1704), .b(n_43470), .o(n_43609) );
na02s01 g767701 ( .a(n_13243), .b(n_13192), .o(n_13766) );
na02s01 g767702 ( .a(n_13314), .b(n_13236), .o(n_13797) );
no02s01 g767703 ( .a(n_13350), .b(n_13349), .o(n_13824) );
in01s01 g767704 ( .a(n_12898), .o(n_12899) );
no02s02 g767705 ( .a(n_12870), .b(n_12869), .o(n_12898) );
in01s01 g767706 ( .a(n_13028), .o(n_13029) );
oa12s01 g767707 ( .a(n_13014), .b(n_12823), .c(n_13013), .o(n_13028) );
na02s01 g767708 ( .a(n_13129), .b(n_13126), .o(n_13212) );
no02s01 g767709 ( .a(n_46414), .b(n_13127), .o(n_13211) );
in01s01 g767710 ( .a(n_13320), .o(n_13321) );
ao12s01 g767711 ( .a(n_13204), .b(n_13084), .c(delay_sub_ln21_0_unr8_stage4_stallmux_q_25_), .o(n_13320) );
in01s01 g767712 ( .a(n_13363), .o(n_13364) );
ao12s01 g767713 ( .a(n_13319), .b(FE_OCP_RBN2562_n_13084), .c(delay_sub_ln21_0_unr8_stage4_stallmux_q_27_), .o(n_13363) );
in01s01 g767714 ( .a(n_13419), .o(n_13420) );
ao12m01 g767715 ( .a(n_13371), .b(FE_OCP_RBN2561_n_13084), .c(delay_sub_ln21_0_unr8_stage4_stallmux_q_29_), .o(n_13419) );
no02s01 g767716 ( .a(n_13221), .b(n_13054), .o(n_12784) );
no02s01 g767717 ( .a(n_12767), .b(n_12245), .o(n_12826) );
in01s02 g767718 ( .a(n_12745), .o(n_12746) );
in01s01 g767719 ( .a(n_12713), .o(n_12745) );
oa12m08 g767720 ( .a(n_12491), .b(n_12655), .c(n_12438), .o(n_12713) );
oa12s01 g767721 ( .a(n_13101), .b(n_12823), .c(n_13086), .o(n_13087) );
na02f08 g767722 ( .a(n_12861), .b(n_12750), .o(n_13019) );
ao12s01 g767723 ( .a(n_12748), .b(n_12863), .c(n_12860), .o(n_12938) );
no02s04 g767724 ( .a(n_13066), .b(n_13210), .o(n_13284) );
no02f02 TIMEBOOST_cell_8741 ( .a(TIMEBOOST_net_2857), .b(n_24896), .o(n_24966) );
in01s01 g767726 ( .a(n_13206), .o(n_13207) );
ao12s01 g767727 ( .a(n_13082), .b(FE_RN_1447_0), .c(delay_add_ln22_unr8_stage4_stallmux_q_31_), .o(n_13206) );
in01s01 g767728 ( .a(n_13440), .o(n_13441) );
ao22s01 g767729 ( .a(FE_OCP_RBN2563_n_13084), .b(n_12229), .c(FE_OCP_RBN2561_n_13084), .d(delay_sub_ln21_0_unr8_stage4_stallmux_q_31_), .o(n_13440) );
oa22s01 g767730 ( .a(FE_OCPN847_n_12799), .b(n_11943), .c(n_12798), .d(n_12747), .o(n_14676) );
oa12s01 g767731 ( .a(n_12822), .b(n_12863), .c(n_12821), .o(n_13795) );
in01s01 g767732 ( .a(n_12846), .o(n_12868) );
in01s01 g767736 ( .a(n_12825), .o(n_12846) );
in01s02 g767737 ( .a(n_12808), .o(n_12825) );
in01s01 g767738 ( .a(n_12771), .o(n_12808) );
in01s01 g767740 ( .a(n_13130), .o(n_13131) );
oa22s01 g767741 ( .a(FE_RN_1447_0), .b(delay_add_ln22_unr8_stage4_stallmux_q_29_), .c(n_12823), .d(n_13086), .o(n_13130) );
in01s01 g767742 ( .a(n_13045), .o(n_13046) );
ao12s01 g767743 ( .a(n_12932), .b(n_12929), .c(delay_add_ln22_unr8_stage4_stallmux_q_25_), .o(n_13045) );
in01s01 g767744 ( .a(n_46414), .o(n_13129) );
in01s01 g767747 ( .a(n_13126), .o(n_13127) );
na02s01 g767748 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_23_), .o(n_13126) );
na02s03 g767749 ( .a(FE_OCP_RBN2559_n_13084), .b(n_12254), .o(n_13777) );
in01s01 g767750 ( .a(n_13238), .o(n_13124) );
na02s06 g767751 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_24_), .o(n_13238) );
no02s01 g767753 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_25_), .o(n_13204) );
in01s02 g767754 ( .a(n_13203), .o(n_13281) );
na02s06 g767755 ( .a(FE_OCP_RBN2562_n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_26_), .o(n_13203) );
in01s01 g767756 ( .a(n_13278), .o(n_13279) );
no02s01 g767757 ( .a(FE_OCP_RBN2562_n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_26_), .o(n_13278) );
in01s02 g767760 ( .a(n_13099), .o(n_13173) );
na02s03 g767761 ( .a(n_13025), .b(n_13024), .o(n_13099) );
no02m01 g767762 ( .a(FE_OCP_RBN2562_n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_27_), .o(n_13319) );
in01s01 g767763 ( .a(n_13356), .o(n_13277) );
no02s01 g767764 ( .a(FE_OCP_RBN2562_n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_28_), .o(n_13356) );
no02s01 g767765 ( .a(FE_OCP_RBN2563_n_13084), .b(n_12188), .o(n_13377) );
no02s01 g767766 ( .a(FE_OCP_RBN2562_n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_29_), .o(n_13371) );
in01s01 g767767 ( .a(n_13369), .o(n_13370) );
no02s01 g767768 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_30_), .b(FE_OCP_RBN2561_n_13084), .o(n_13369) );
na02s01 g767769 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_30_), .b(FE_OCP_RBN2561_n_13084), .o(n_13421) );
in01s03 g767772 ( .a(n_13083), .o(n_13213) );
no02s02 g767773 ( .a(n_13025), .b(n_13024), .o(n_13083) );
no02s01 g767774 ( .a(FE_RN_1447_0), .b(delay_add_ln22_unr8_stage4_stallmux_q_31_), .o(n_13082) );
na02s01 g767775 ( .a(n_13015), .b(n_12986), .o(n_13016) );
no02s02 g767776 ( .a(n_13043), .b(FE_OCPN4521_n_13015), .o(n_13044) );
na02s01 g767779 ( .a(n_46933), .b(delay_add_ln22_unr8_stage4_stallmux_q_26_), .o(n_13000) );
no02s01 g767780 ( .a(n_46933), .b(delay_add_ln22_unr8_stage4_stallmux_q_23_), .o(n_12807) );
na02s01 g767781 ( .a(n_12823), .b(n_11886), .o(n_12824) );
na02s01 g767782 ( .a(n_12823), .b(n_13086), .o(n_13122) );
na02s01 g767783 ( .a(FE_RN_1447_0), .b(delay_add_ln22_unr8_stage4_stallmux_q_28_), .o(n_13101) );
no02s01 g767786 ( .a(n_46933), .b(delay_add_ln22_unr8_stage4_stallmux_q_25_), .o(n_12932) );
na02s01 g767787 ( .a(n_46933), .b(delay_add_ln22_unr8_stage4_stallmux_q_23_), .o(n_12900) );
na02s01 g767788 ( .a(n_46933), .b(delay_add_ln22_unr8_stage4_stallmux_q_24_), .o(n_12867) );
in01s01 g767790 ( .a(n_13120), .o(n_13121) );
no02s01 g767791 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_30_), .b(FE_RN_1447_0), .o(n_13120) );
no02s02 g767792 ( .a(n_12743), .b(delay_add_ln22_unr8_stage4_stallmux_q_22_), .o(n_12869) );
no02s03 g767793 ( .a(n_12744), .b(n_11868), .o(n_12870) );
na02s02 g767794 ( .a(n_12823), .b(n_13013), .o(n_13014) );
in01s01 g767795 ( .a(n_12968), .o(n_12969) );
no02s01 g767796 ( .a(FE_RN_1447_0), .b(delay_add_ln22_unr8_stage4_stallmux_q_28_), .o(n_12968) );
na02s01 g767797 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_30_), .b(FE_RN_1447_0), .o(n_13193) );
na02s01 g767798 ( .a(n_12823), .b(n_12215), .o(n_12956) );
na02s01 g767799 ( .a(n_12863), .b(n_12821), .o(n_12822) );
na02s06 g767800 ( .a(n_13167), .b(n_13315), .o(n_13316) );
na02s04 g767801 ( .a(n_13252), .b(n_13251), .o(n_13253) );
no02s04 g767802 ( .a(n_13038), .b(n_13113), .o(n_13256) );
na02s02 g767803 ( .a(n_12925), .b(n_13248), .o(n_13088) );
no02s01 g767804 ( .a(n_13064), .b(n_13210), .o(n_13202) );
na02s04 g767805 ( .a(n_13065), .b(n_12996), .o(n_13066) );
na02s01 g767806 ( .a(FE_OCP_RBN4095_n_12880), .b(n_13119), .o(n_13236) );
no02s04 g767807 ( .a(n_12764), .b(FE_OCP_RBN4094_n_12880), .o(n_13350) );
na02s02 g767808 ( .a(FE_OCP_RBN4093_n_12880), .b(n_13118), .o(n_13192) );
no02s01 g767809 ( .a(n_12873), .b(n_12918), .o(n_12951) );
no02s02 g767810 ( .a(FE_OCP_RBN4088_n_12880), .b(n_12763), .o(n_13349) );
in01s01 g767811 ( .a(n_13378), .o(n_13314) );
no02s02 g767812 ( .a(n_13119), .b(FE_OCP_RBN4095_n_12880), .o(n_13378) );
in01s01 g767813 ( .a(n_13160), .o(n_13243) );
no02s01 g767814 ( .a(n_13118), .b(FE_OCPN926_n_12914), .o(n_13160) );
no02s01 g767815 ( .a(n_13241), .b(n_13271), .o(n_13790) );
in01s01 g767816 ( .a(n_12849), .o(n_12770) );
na02m02 g767817 ( .a(n_12799), .b(n_12753), .o(n_12849) );
na02s01 g767818 ( .a(n_13065), .b(n_13041), .o(n_13761) );
no02s01 g767819 ( .a(n_13064), .b(n_12926), .o(n_13736) );
na02s02 TIMEBOOST_cell_8852 ( .a(n_5727), .b(n_5728), .o(TIMEBOOST_net_2913) );
in01s01 g767821 ( .a(n_13381), .o(n_13280) );
na02s02 g767822 ( .a(n_13084), .b(n_12255), .o(n_13381) );
in01s01 g767825 ( .a(n_13221), .o(n_12767) );
na02s02 g767826 ( .a(n_12799), .b(n_12747), .o(n_13221) );
in01s01 g767827 ( .a(n_12967), .o(n_13138) );
oa12s01 g767828 ( .a(n_46933), .b(delay_add_ln22_unr8_stage4_stallmux_q_24_), .c(delay_add_ln22_unr8_stage4_stallmux_q_25_), .o(n_12967) );
no02s06 TIMEBOOST_cell_6880 ( .a(TIMEBOOST_net_2198), .b(n_40828), .o(n_40910) );
ao12f08 g767832 ( .a(n_12475), .b(n_12668), .c(n_12507), .o(n_12727) );
no02s01 TIMEBOOST_cell_1775 ( .a(n_42980), .b(FE_OCP_RBN3307_n_43022), .o(TIMEBOOST_net_502) );
na02m08 g767834 ( .a(n_12999), .b(n_12919), .o(n_13208) );
ao22s01 g767835 ( .a(n_12787), .b(FE_OCP_RBN5395_cordic_combinational_sub_ln23_0_unr12_z_0_), .c(n_12786), .d(FE_OCP_RBN5392_cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n_13764) );
in01s01 g767836 ( .a(FE_OCPN5136_n_12795), .o(n_14685) );
ao12s01 g767837 ( .a(n_12725), .b(FE_OFN754_n_13889), .c(n_12724), .o(n_12795) );
in01s01 g767840 ( .a(n_12997), .o(n_12998) );
na02s01 g767841 ( .a(n_12955), .b(n_12954), .o(n_12997) );
na02s02 g767843 ( .a(n_12852), .b(n_11663), .o(n_13015) );
in01s04 g767844 ( .a(n_12986), .o(n_13043) );
na02s04 g767845 ( .a(n_12853), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_21_), .o(n_12986) );
no02m10 g767861 ( .a(FE_OCP_RBN2542_n_12921), .b(n_12435), .o(n_13084) );
in01s02 g767862 ( .a(n_12793), .o(n_12794) );
na02s02 g767863 ( .a(n_12773), .b(n_12723), .o(n_12793) );
na02s02 g767865 ( .a(n_12728), .b(delay_add_ln22_unr8_stage4_stallmux_q_21_), .o(n_12836) );
in01s01 g767874 ( .a(n_12823), .o(n_12929) );
in01s02 g767880 ( .a(n_46933), .o(n_12823) );
no02s06 g767885 ( .a(n_12728), .b(delay_add_ln22_unr8_stage4_stallmux_q_21_), .o(n_12766) );
no02s06 g767886 ( .a(n_13249), .b(n_13198), .o(n_13315) );
na02s01 g767887 ( .a(n_12843), .b(n_12759), .o(n_12844) );
no02f08 g767889 ( .a(FE_OCP_RBN6563_n_12753), .b(FE_OFN754_n_13889), .o(n_12865) );
no02s02 g767890 ( .a(n_13116), .b(FE_OCP_RBN4093_n_12880), .o(n_13241) );
in01s01 g767891 ( .a(n_12925), .o(n_12926) );
na02s02 g767892 ( .a(n_12905), .b(n_12910), .o(n_12925) );
in01s01 g767893 ( .a(n_13064), .o(n_12996) );
no02s02 g767894 ( .a(n_12905), .b(FE_OCPN926_n_12914), .o(n_13064) );
in01s01 g767895 ( .a(n_13040), .o(n_13041) );
no02s02 g767896 ( .a(n_12990), .b(FE_OCP_RBN2539_n_12880), .o(n_13040) );
in01s01 g767897 ( .a(n_13168), .o(n_13271) );
na02s02 g767898 ( .a(FE_OCP_RBN4093_n_12880), .b(n_13116), .o(n_13168) );
na02s01 g767899 ( .a(n_12990), .b(FE_OCP_RBN2539_n_12880), .o(n_13065) );
na02s01 g767900 ( .a(n_13199), .b(n_13251), .o(n_13769) );
in01s01 g767901 ( .a(n_12768), .o(n_12796) );
no02s02 g767902 ( .a(FE_OFN754_n_13889), .b(n_11944), .o(n_12768) );
na02m01 g767903 ( .a(n_12921), .b(n_46985), .o(n_13025) );
no02s01 g767904 ( .a(FE_OFN754_n_13889), .b(n_12724), .o(n_12725) );
in01s02 g767905 ( .a(n_12743), .o(n_12744) );
na03f04 TIMEBOOST_cell_7372 ( .a(FE_OCP_RBN3356_FE_RN_1058_0), .b(n_26498), .c(n_26878), .o(n_27019) );
in01s02 g767907 ( .a(n_12690), .o(n_12691) );
in01s01 g767908 ( .a(n_12655), .o(n_12690) );
ao12m08 g767909 ( .a(n_12392), .b(n_12615), .c(n_12420), .o(n_12655) );
oa12f06 g767910 ( .a(n_12765), .b(n_12700), .c(FE_OCP_RBN5395_cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n_12863) );
no03s04 g767911 ( .a(n_12992), .b(n_13080), .c(n_13079), .o(n_13252) );
in01s01 g767912 ( .a(n_13038), .o(n_13039) );
na02s04 g767913 ( .a(n_12920), .b(n_13621), .o(n_13038) );
in01m04 g767914 ( .a(n_12873), .o(n_12999) );
na02s06 g767915 ( .a(n_12843), .b(n_12783), .o(n_12873) );
na02s06 g767916 ( .a(n_12923), .b(n_12856), .o(n_12924) );
na02f04 TIMEBOOST_cell_8658 ( .a(n_16732), .b(n_16737), .o(TIMEBOOST_net_2816) );
ao12s01 g767918 ( .a(n_12742), .b(n_12741), .c(n_12740), .o(n_13118) );
in01s02 g767919 ( .a(n_12763), .o(n_12764) );
oa12s01 g767920 ( .a(n_12708), .b(n_12707), .c(n_12706), .o(n_12763) );
in01s01 g767921 ( .a(FE_OCPN847_n_12799), .o(n_12798) );
no02m08 TIMEBOOST_cell_4514 ( .a(TIMEBOOST_net_1347), .b(n_39934), .o(n_40107) );
ao12s01 g767923 ( .a(n_12712), .b(n_12711), .c(n_12710), .o(n_13119) );
no02s02 TIMEBOOST_cell_1838 ( .a(TIMEBOOST_net_533), .b(FE_OCPN6901_FE_OCP_RBN4472_n_31819), .o(FE_RN_2882_0) );
na02s04 g767928 ( .a(n_12651), .b(n_12455), .o(n_12686) );
no03f06 TIMEBOOST_cell_7371 ( .a(n_20920), .b(n_20855), .c(n_20942), .o(n_21094) );
na02m06 g767930 ( .a(n_12817), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_20_), .o(n_12954) );
na02s02 g767931 ( .a(n_12816), .b(n_11524), .o(n_12955) );
na02s01 g767932 ( .a(n_12707), .b(n_12706), .o(n_12708) );
na02s02 g767933 ( .a(n_12664), .b(n_12683), .o(n_12684) );
no02s02 g767934 ( .a(n_12635), .b(n_12658), .o(n_12705) );
no02s01 g767935 ( .a(n_12741), .b(n_12740), .o(n_12742) );
in01s01 g767936 ( .a(n_12722), .o(n_12723) );
no02s06 g767937 ( .a(n_12694), .b(n_12693), .o(n_12722) );
na02m02 g767938 ( .a(n_12627), .b(n_12448), .o(n_12654) );
in01m02 g767939 ( .a(n_12890), .o(n_12891) );
na02m02 g767940 ( .a(n_12848), .b(n_12847), .o(n_12890) );
no02s01 g767941 ( .a(n_12711), .b(n_12710), .o(n_12712) );
na02s06 g767942 ( .a(n_12694), .b(n_12693), .o(n_12773) );
na02s04 TIMEBOOST_cell_7032 ( .a(TIMEBOOST_net_2274), .b(n_3950), .o(n_4168) );
no02s02 g767944 ( .a(n_12885), .b(n_12911), .o(n_12920) );
in01s01 g767945 ( .a(n_13255), .o(n_13167) );
na02s02 g767946 ( .a(n_13115), .b(n_13075), .o(n_13255) );
no02s03 g767947 ( .a(n_12782), .b(n_12781), .o(n_12783) );
in01s02 g767948 ( .a(n_12788), .o(n_12843) );
na02s01 g767949 ( .a(n_12775), .b(n_12774), .o(n_12788) );
no02s03 g767950 ( .a(n_12918), .b(n_12882), .o(n_12919) );
na02s02 g767951 ( .a(n_13078), .b(n_13159), .o(n_13166) );
no02s06 g767952 ( .a(n_13034), .b(n_13035), .o(n_13037) );
no02s06 g767954 ( .a(n_12749), .b(n_12748), .o(n_12750) );
in01s02 g767955 ( .a(n_12857), .o(n_12923) );
na02s02 g767956 ( .a(n_12811), .b(n_12832), .o(n_12857) );
no02s02 g767957 ( .a(n_12855), .b(n_12854), .o(n_12856) );
na02s06 g767958 ( .a(n_12994), .b(n_12916), .o(n_12995) );
no02m01 g767959 ( .a(n_13104), .b(n_13200), .o(n_13201) );
in01s01 g767960 ( .a(n_13164), .o(n_13165) );
no02s01 g767961 ( .a(n_13032), .b(n_13150), .o(n_13164) );
no02s01 g767962 ( .a(n_13079), .b(n_13080), .o(n_13036) );
no02s01 g767963 ( .a(n_13150), .b(n_12917), .o(n_13602) );
no02s01 g767964 ( .a(n_12737), .b(n_12982), .o(n_13354) );
na02s01 g767965 ( .a(n_12832), .b(n_12815), .o(n_13018) );
na02s01 g767966 ( .a(FE_OCP_RBN2539_n_12880), .b(n_13163), .o(n_13251) );
in01s01 g767967 ( .a(n_13274), .o(n_13275) );
na02s01 g767968 ( .a(n_13248), .b(n_13161), .o(n_13274) );
no02s01 g767969 ( .a(n_13079), .b(n_13076), .o(n_13717) );
in01s01 g767970 ( .a(n_13198), .o(n_13199) );
no02s02 g767971 ( .a(FE_OCP_RBN2539_n_12880), .b(n_13163), .o(n_13198) );
na02s01 g767972 ( .a(n_12886), .b(n_13196), .o(n_13674) );
na02s01 g767973 ( .a(n_12883), .b(n_13159), .o(n_13520) );
na02s01 g767974 ( .a(n_12775), .b(n_12994), .o(n_13425) );
na02s01 g767975 ( .a(n_12811), .b(n_12810), .o(n_13177) );
no02s01 g767976 ( .a(n_13035), .b(n_12781), .o(n_13473) );
no02s01 g767977 ( .a(n_13034), .b(n_12782), .o(n_13443) );
na02s01 g767978 ( .a(n_12717), .b(n_12860), .o(n_12821) );
na02s01 g767979 ( .a(n_13162), .b(n_12993), .o(n_13733) );
in01s01 g767980 ( .a(n_12786), .o(n_12787) );
na02s01 g767981 ( .a(n_12765), .b(n_12701), .o(n_12786) );
no02s01 g767982 ( .a(n_12749), .b(n_12719), .o(n_12937) );
na02s01 g767983 ( .a(n_13115), .b(n_12988), .o(n_13671) );
na02s01 g767984 ( .a(n_13114), .b(n_13109), .o(n_13679) );
no02s01 g767985 ( .a(n_12958), .b(n_12855), .o(n_13305) );
na02s01 g767986 ( .a(n_12884), .b(n_13078), .o(n_13504) );
na02s01 g767987 ( .a(n_13077), .b(n_13031), .o(n_13651) );
no02s01 g767988 ( .a(n_13200), .b(n_13197), .o(n_13544) );
na02s01 g767989 ( .a(n_13112), .b(n_13103), .o(n_13584) );
na02s01 g767990 ( .a(n_12813), .b(n_12841), .o(n_13215) );
in01m02 g767991 ( .a(n_12688), .o(n_12689) );
in01m01 g767992 ( .a(n_12668), .o(n_12688) );
oa12m08 g767993 ( .a(n_12474), .b(n_12629), .c(n_12432), .o(n_12668) );
in01m01 g767994 ( .a(n_12852), .o(n_12853) );
oa12m01 g767995 ( .a(n_12762), .b(n_12761), .c(n_12760), .o(n_12852) );
no02s01 TIMEBOOST_cell_4407 ( .a(n_843), .b(n_885), .o(TIMEBOOST_net_1294) );
ao12s01 g767997 ( .a(n_12680), .b(n_12679), .c(n_12678), .o(n_13116) );
oa12s02 g767998 ( .a(n_12704), .b(n_12703), .c(n_12702), .o(n_12990) );
ao22s02 g768000 ( .a(n_12646), .b(n_12429), .c(n_12645), .d(n_12430), .o(n_12905) );
na02m01 g768001 ( .a(n_12761), .b(n_12760), .o(n_12762) );
na02s02 g768002 ( .a(n_12616), .b(n_12666), .o(n_12667) );
in01m02 g768003 ( .a(n_12819), .o(n_12820) );
na02m02 g768004 ( .a(n_12809), .b(FE_OCP_RBN2529_n_12731), .o(n_12819) );
in01s04 g768005 ( .a(n_12664), .o(n_12658) );
na02s04 g768007 ( .a(n_12613), .b(n_11492), .o(n_12664) );
in01s01 g768008 ( .a(n_12683), .o(n_12635) );
na02m03 g768009 ( .a(n_12612), .b(delay_add_ln22_unr8_stage4_stallmux_q_19_), .o(n_12683) );
no02s02 g768010 ( .a(n_12634), .b(FE_OCPN1240_n_13412), .o(n_12682) );
na02s02 g768011 ( .a(FE_OCPN1242_n_12633), .b(FE_OCPN1239_n_13412), .o(n_12681) );
no02s02 g768012 ( .a(n_12629), .b(n_12498), .o(n_12630) );
no03s02 TIMEBOOST_cell_2164 ( .a(n_32499), .b(n_32391), .c(n_32498), .o(n_32500) );
na02m02 g768015 ( .a(n_12729), .b(n_11528), .o(n_12847) );
no03f04 TIMEBOOST_cell_3720 ( .a(n_26299), .b(n_26306), .c(n_26252), .o(n_26469) );
na02m04 g768017 ( .a(n_12730), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_19_), .o(n_12848) );
in01s01 g768018 ( .a(n_12651), .o(n_12652) );
na02s04 g768019 ( .a(n_12616), .b(n_12431), .o(n_12651) );
na02s01 g768020 ( .a(n_12703), .b(n_12702), .o(n_12704) );
no02s01 g768021 ( .a(n_12679), .b(n_12678), .o(n_12680) );
na02s01 g768022 ( .a(n_12910), .b(n_12887), .o(n_13248) );
in01s01 g768023 ( .a(n_13080), .o(n_12988) );
no02s02 g768024 ( .a(FE_OCPN926_n_12914), .b(n_12965), .o(n_13080) );
in01s01 g768025 ( .a(n_12992), .o(n_12993) );
no02s01 g768026 ( .a(FE_OCPN926_n_12914), .b(n_12964), .o(n_12992) );
no02s01 g768027 ( .a(FE_OCPN926_n_12914), .b(n_12985), .o(n_13079) );
in01s01 g768028 ( .a(n_13621), .o(n_12917) );
na02s02 g768029 ( .a(n_12910), .b(n_12909), .o(n_13621) );
in01s01 g768030 ( .a(n_12885), .o(n_12886) );
no02s01 g768031 ( .a(n_12790), .b(n_12840), .o(n_12885) );
in01s01 g768032 ( .a(n_12911), .o(n_13077) );
no02s01 g768033 ( .a(n_12790), .b(n_12838), .o(n_12911) );
in01s01 g768034 ( .a(n_13113), .o(n_13114) );
no02s01 g768035 ( .a(FE_OCP_RBN2539_n_12880), .b(n_13073), .o(n_13113) );
in01s01 g768036 ( .a(n_13075), .o(n_13076) );
na02s02 g768037 ( .a(FE_OCPN926_n_12914), .b(n_12985), .o(n_13075) );
na02s02 g768038 ( .a(FE_OCPN926_n_12914), .b(n_12965), .o(n_13115) );
in01s01 g768039 ( .a(n_13162), .o(n_13249) );
na02s02 g768040 ( .a(FE_OCPN926_n_12914), .b(n_12964), .o(n_13162) );
in01s01 g768041 ( .a(n_12782), .o(n_12759) );
no02m01 g768042 ( .a(FE_OCP_RBN4047_n_12721), .b(n_12738), .o(n_12782) );
no02s04 g768043 ( .a(FE_OCP_RBN2522_n_12721), .b(n_12256), .o(n_12781) );
na02s01 g768044 ( .a(FE_OCP_RBN5578_n_12753), .b(n_12289), .o(n_12775) );
in01s01 g768045 ( .a(n_12774), .o(n_12737) );
na02s02 g768046 ( .a(FE_OCP_RBN5578_n_12753), .b(n_12720), .o(n_12774) );
in01s01 g768047 ( .a(n_12918), .o(n_12884) );
no02s02 g768048 ( .a(n_12790), .b(n_12871), .o(n_12918) );
in01s01 g768049 ( .a(n_12882), .o(n_12883) );
no02s01 g768050 ( .a(n_12790), .b(n_12850), .o(n_12882) );
in01s01 g768051 ( .a(n_13111), .o(n_13112) );
no02s01 g768052 ( .a(FE_OCP_RBN2539_n_12880), .b(n_13074), .o(n_13111) );
no02m01 g768053 ( .a(FE_OCP_RBN2539_n_12880), .b(n_12325), .o(n_13197) );
in01s01 g768054 ( .a(n_13078), .o(n_13033) );
na02s02 g768055 ( .a(FE_OCP_RBN2539_n_12880), .b(n_12871), .o(n_13078) );
na02s01 g768056 ( .a(FE_OCP_RBN2539_n_12880), .b(n_12850), .o(n_13159) );
in01s01 g768057 ( .a(n_12963), .o(n_13034) );
na02s06 g768058 ( .a(FE_OCP_RBN2539_n_12880), .b(n_12738), .o(n_12963) );
no02s01 g768059 ( .a(FE_OCP_RBN2538_n_12880), .b(n_12257), .o(n_13035) );
no02s06 g768060 ( .a(n_12881), .b(n_12135), .o(n_12958) );
na02s06 g768061 ( .a(n_12790), .b(n_12789), .o(n_12841) );
in01s01 g768062 ( .a(n_12810), .o(n_12776) );
na02s04 g768063 ( .a(n_13004), .b(n_12223), .o(n_12810) );
na02s06 g768064 ( .a(FE_OCP_RBN5581_n_12753), .b(n_12692), .o(n_12860) );
in01s01 g768065 ( .a(n_12718), .o(n_12719) );
na02s06 g768066 ( .a(FE_OCP_RBN5581_n_12753), .b(n_12699), .o(n_12718) );
na02m06 g768067 ( .a(FE_OCP_RBN5578_n_12753), .b(FE_OCPN3554_n_12671), .o(n_12765) );
in01s01 g768068 ( .a(n_12700), .o(n_12701) );
no02f06 g768069 ( .a(FE_OCP_RBN6565_n_12753), .b(FE_OCPN3554_n_12671), .o(n_12700) );
in01s01 g768070 ( .a(n_12748), .o(n_12717) );
no02s04 g768071 ( .a(FE_OCP_RBN5581_n_12753), .b(n_12692), .o(n_12748) );
no02s04 g768072 ( .a(FE_OCP_RBN5581_n_12753), .b(n_12699), .o(n_12749) );
na02s06 g768073 ( .a(n_13004), .b(n_12222), .o(n_12815) );
na02s02 g768074 ( .a(FE_OCP_RBN4048_n_12721), .b(n_12224), .o(n_12811) );
na02s02 g768075 ( .a(FE_OCP_RBN4048_n_12721), .b(n_12221), .o(n_12832) );
no02s02 g768076 ( .a(n_12790), .b(n_12134), .o(n_12855) );
in01s01 g768077 ( .a(n_12854), .o(n_12813) );
no02s02 g768078 ( .a(n_12790), .b(n_12789), .o(n_12854) );
na02s06 g768079 ( .a(FE_OCP_RBN2539_n_12880), .b(n_12290), .o(n_12994) );
in01s01 g768080 ( .a(n_12982), .o(n_12916) );
no02s01 g768081 ( .a(FE_OCP_RBN4048_n_12721), .b(n_12720), .o(n_12982) );
in01s01 g768082 ( .a(n_13103), .o(n_13104) );
na02s02 g768083 ( .a(FE_OCP_RBN2539_n_12880), .b(n_13074), .o(n_13103) );
no02s06 g768084 ( .a(FE_OCPN926_n_12914), .b(n_12326), .o(n_13200) );
in01s01 g768085 ( .a(n_13196), .o(n_13312) );
na02s01 g768086 ( .a(FE_OCP_RBN2539_n_12880), .b(n_12840), .o(n_13196) );
in01s01 g768087 ( .a(n_13109), .o(n_13110) );
na02s01 g768088 ( .a(FE_OCP_RBN2539_n_12880), .b(n_13073), .o(n_13109) );
in01s01 g768089 ( .a(n_13031), .o(n_13032) );
na02s02 g768090 ( .a(FE_OCP_RBN2539_n_12880), .b(n_12838), .o(n_13031) );
no02s02 g768091 ( .a(FE_OCPN926_n_12914), .b(n_12909), .o(n_13150) );
in01s01 g768092 ( .a(n_13210), .o(n_13161) );
no02s01 g768093 ( .a(FE_OCPN926_n_12914), .b(n_12887), .o(n_13210) );
in01s01 g768094 ( .a(n_12627), .o(n_12628) );
in01s01 g768095 ( .a(n_12615), .o(n_12627) );
oa12m08 g768096 ( .a(n_12398), .b(n_12569), .c(n_12353), .o(n_12615) );
no02s06 TIMEBOOST_cell_1891 ( .a(n_39989), .b(FE_OCP_RBN3333_n_39942), .o(TIMEBOOST_net_560) );
ao12s02 g768098 ( .a(n_12220), .b(n_12663), .c(n_12046), .o(n_12711) );
ao12s01 g768099 ( .a(n_12214), .b(n_12663), .c(n_12119), .o(n_12707) );
oa12s01 g768100 ( .a(n_12598), .b(n_12597), .c(n_12596), .o(n_13800) );
in01s02 g768101 ( .a(n_12816), .o(n_12817) );
oa12m04 g768102 ( .a(n_12736), .b(n_12735), .c(n_12734), .o(n_12816) );
oa22s02 g768103 ( .a(n_12602), .b(n_12494), .c(n_12603), .d(n_12493), .o(n_13163) );
ao12s03 g768104 ( .a(n_12632), .b(n_12589), .c(n_12631), .o(n_12694) );
no02m04 TIMEBOOST_cell_1809 ( .a(n_15734), .b(FE_RN_1486_0), .o(TIMEBOOST_net_519) );
na02m04 g768106 ( .a(n_12735), .b(n_12734), .o(n_12736) );
no02m08 g768109 ( .a(n_12698), .b(n_12415), .o(n_12761) );
no02s02 g768110 ( .a(n_12589), .b(n_12631), .o(n_12632) );
in01m02 g768111 ( .a(n_12755), .o(n_12756) );
na02m02 g768112 ( .a(n_12733), .b(n_12696), .o(n_12755) );
in01s02 g768115 ( .a(n_12633), .o(n_12634) );
na02s06 g768116 ( .a(n_12605), .b(delay_add_ln22_unr8_stage4_stallmux_q_18_), .o(n_12633) );
no02s08 g768120 ( .a(n_12589), .b(n_12400), .o(n_12616) );
no02s04 g768123 ( .a(n_12605), .b(delay_add_ln22_unr8_stage4_stallmux_q_18_), .o(n_13412) );
no02m02 g768125 ( .a(n_12716), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_18_), .o(n_12731) );
in01s01 g768126 ( .a(n_12647), .o(n_12648) );
no02s02 g768127 ( .a(n_12620), .b(n_12619), .o(n_12647) );
na02s02 g768128 ( .a(n_12716), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_18_), .o(n_12809) );
na02s01 g768129 ( .a(n_12597), .b(n_12596), .o(n_12598) );
na02s02 g768130 ( .a(n_12662), .b(n_12085), .o(n_12703) );
no02s01 g768131 ( .a(n_12663), .b(n_12281), .o(n_12679) );
in01s01 g768132 ( .a(n_12645), .o(n_12646) );
oa12s01 g768133 ( .a(n_11892), .b(n_12623), .c(n_12083), .o(n_12645) );
in01m01 g768134 ( .a(n_12629), .o(n_12614) );
ao12m08 g768135 ( .a(n_12386), .b(n_12591), .c(n_12424), .o(n_12629) );
in01s02 g768136 ( .a(FE_OCP_RBN5578_n_12753), .o(n_13004) );
in01s02 g768137 ( .a(n_12790), .o(n_12881) );
in01m02 g768139 ( .a(n_12790), .o(n_12910) );
in01m01 g768148 ( .a(FE_OCP_RBN4102_n_12880), .o(n_13916) );
in01m01 g768164 ( .a(n_13195), .o(n_13437) );
in01s02 g768170 ( .a(n_13515), .o(n_14376) );
in01s06 g768177 ( .a(n_13514), .o(n_13515) );
in01s06 g768180 ( .a(n_13418), .o(n_13514) );
in01s02 g768189 ( .a(FE_OFN1181_n_13195), .o(n_13469) );
in01s06 g768191 ( .a(FE_OFN4795_n_13195), .o(n_13418) );
in01m20 g768227 ( .a(FE_OCP_RBN4048_n_12721), .o(n_12880) );
in01m08 g768229 ( .a(FE_OCP_RBN4048_n_12721), .o(n_12790) );
oa12s01 g768239 ( .a(n_12588), .b(n_12591), .c(n_12587), .o(n_13721) );
in01m02 g768240 ( .a(n_12729), .o(n_12730) );
oa12m02 g768241 ( .a(n_12676), .b(n_12675), .c(n_12674), .o(n_12729) );
ao12s01 g768242 ( .a(n_12611), .b(n_12623), .c(n_12610), .o(n_12887) );
in01s02 g768243 ( .a(n_12612), .o(n_12613) );
oa12s04 g768244 ( .a(n_12572), .b(n_12571), .c(FE_OCP_DRV_N1412_n_12570), .o(n_12612) );
na02m02 g768245 ( .a(n_12675), .b(n_12674), .o(n_12676) );
na02s03 g768246 ( .a(n_12571), .b(FE_OCP_DRV_N1412_n_12570), .o(n_12572) );
in01s04 g768247 ( .a(n_12698), .o(n_12735) );
na02m08 g768248 ( .a(n_12675), .b(n_12384), .o(n_12698) );
no02s02 g768249 ( .a(n_12565), .b(delay_add_ln22_unr8_stage4_stallmux_q_17_), .o(n_12619) );
na02s10 g768253 ( .a(n_12571), .b(FE_OCPN1616_n_12371), .o(n_12589) );
na02s02 g768254 ( .a(n_12604), .b(n_12157), .o(n_12662) );
na02m04 g768256 ( .a(n_12697), .b(n_12657), .o(n_12714) );
in01s02 g768258 ( .a(n_12599), .o(n_12600) );
na02s02 g768259 ( .a(n_12576), .b(n_12559), .o(n_12599) );
na02s01 g768260 ( .a(n_12591), .b(n_12587), .o(n_12588) );
na02m04 g768261 ( .a(n_12673), .b(n_12672), .o(n_12733) );
in01m01 g768262 ( .a(n_12695), .o(n_12696) );
no02f04 g768263 ( .a(n_12673), .b(n_12672), .o(n_12695) );
no02m01 g768264 ( .a(n_12623), .b(n_12279), .o(n_12663) );
no02s01 g768265 ( .a(n_12623), .b(n_12610), .o(n_12611) );
in01s02 g768266 ( .a(n_12602), .o(n_12603) );
ao12s01 g768267 ( .a(n_11974), .b(n_12573), .c(n_11894), .o(n_12602) );
in01s01 g768268 ( .a(n_12569), .o(n_12597) );
ao12m08 g768269 ( .a(n_12300), .b(n_12553), .c(n_12335), .o(n_12569) );
in01s01 g768271 ( .a(FE_OCP_DRV_N1452_n_12585), .o(n_12586) );
ao12s01 g768272 ( .a(n_12552), .b(n_12553), .c(n_12551), .o(n_12585) );
ao12s01 g768273 ( .a(n_12568), .b(n_12573), .c(n_12567), .o(n_12964) );
ao12m01 g768274 ( .a(n_12643), .b(n_12644), .c(n_12642), .o(n_12716) );
oa12s06 g768275 ( .a(n_12562), .b(n_12561), .c(n_12560), .o(n_12605) );
na02s06 g768276 ( .a(n_12621), .b(n_12618), .o(n_12622) );
in01s01 g768277 ( .a(n_12574), .o(n_12575) );
na02s02 g768278 ( .a(n_12550), .b(n_12563), .o(n_12574) );
no02s01 g768279 ( .a(n_12573), .b(n_12567), .o(n_12568) );
na02s06 g768280 ( .a(n_12561), .b(n_12560), .o(n_12562) );
no02s01 g768281 ( .a(n_12553), .b(n_12551), .o(n_12552) );
na02m04 g768282 ( .a(n_12641), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_16_), .o(n_12697) );
in01s01 g768283 ( .a(n_12558), .o(n_12559) );
no02s04 g768284 ( .a(n_12538), .b(n_12537), .o(n_12558) );
no02m08 g768285 ( .a(n_12644), .b(n_12372), .o(n_12675) );
no02m01 g768286 ( .a(n_12644), .b(n_12642), .o(n_12643) );
in01s02 g768287 ( .a(n_12656), .o(n_12657) );
no02m06 g768288 ( .a(n_12641), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_16_), .o(n_12656) );
na02s02 g768290 ( .a(n_12538), .b(n_12537), .o(n_12576) );
in01m02 g768291 ( .a(n_12659), .o(n_12660) );
na02m02 g768292 ( .a(n_12640), .b(n_12621), .o(n_12659) );
in01s01 g768293 ( .a(n_12623), .o(n_12604) );
oa12m08 g768295 ( .a(n_12389), .b(n_44426), .c(n_12346), .o(n_12591) );
oa12m02 g768296 ( .a(n_12608), .b(n_12607), .c(n_12606), .o(n_12673) );
ao12s01 g768297 ( .a(n_12546), .b(n_12545), .c(n_12544), .o(n_12985) );
no03m08 TIMEBOOST_cell_3703 ( .a(n_38885), .b(n_38930), .c(FE_OCP_RBN4327_n_38878), .o(TIMEBOOST_net_887) );
ao22s01 g768300 ( .a(n_44425), .b(n_12408), .c(n_44426), .d(n_12409), .o(n_13646) );
no02s01 g768302 ( .a(n_12535), .b(n_12051), .o(n_12573) );
na02s04 TIMEBOOST_cell_7988 ( .a(n_26014), .b(n_26059), .o(TIMEBOOST_net_2625) );
na02s01 g768304 ( .a(n_12516), .b(n_12388), .o(n_12517) );
na02m02 g768305 ( .a(n_12607), .b(n_12606), .o(n_12608) );
na02m08 g768306 ( .a(n_12607), .b(n_12411), .o(n_12644) );
na02s04 g768307 ( .a(n_12579), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_15_), .o(n_12621) );
no02s10 g768308 ( .a(n_12531), .b(FE_OCPN1657_n_12368), .o(n_12561) );
in01s01 g768310 ( .a(n_12549), .o(n_12550) );
no02s06 g768311 ( .a(n_12530), .b(delay_add_ln22_unr8_stage4_stallmux_q_15_), .o(n_12549) );
na02s06 g768312 ( .a(n_12530), .b(delay_add_ln22_unr8_stage4_stallmux_q_15_), .o(n_12563) );
na02m02 g768314 ( .a(n_12618), .b(n_12617), .o(n_12638) );
na02m06 g768315 ( .a(n_12580), .b(n_11298), .o(n_12640) );
na02m02 g768317 ( .a(n_12522), .b(n_12503), .o(n_12547) );
no02s01 g768318 ( .a(n_12545), .b(n_12544), .o(n_12546) );
oa12m08 g768319 ( .a(FE_OCPN1344_n_12313), .b(n_12519), .c(n_12262), .o(n_12553) );
ao12s01 g768320 ( .a(n_12515), .b(n_12514), .c(n_12513), .o(n_12965) );
ao12s01 g768321 ( .a(n_12487), .b(n_12486), .c(n_12485), .o(n_13073) );
ao22s01 g768322 ( .a(n_12519), .b(n_12329), .c(n_12482), .d(n_12328), .o(n_13625) );
oa12s01 g768323 ( .a(n_12510), .b(n_12509), .c(n_12508), .o(n_13590) );
ao12s04 g768324 ( .a(n_12489), .b(n_12490), .c(FE_OCPN1655_n_12488), .o(n_12538) );
no02s06 g768326 ( .a(n_12490), .b(FE_OCPN1659_n_12488), .o(n_12489) );
in01s01 g768327 ( .a(n_12502), .o(n_12503) );
no02m06 g768328 ( .a(n_12469), .b(n_12468), .o(n_12502) );
no02s01 g768329 ( .a(n_12514), .b(n_12513), .o(n_12515) );
no02s01 g768330 ( .a(n_12486), .b(n_12485), .o(n_12487) );
na02s10 g768331 ( .a(n_12349), .b(n_12465), .o(n_12531) );
no02s06 g768332 ( .a(FE_OCPN1360_n_12370), .b(n_12490), .o(n_12516) );
in01s01 g768333 ( .a(n_12618), .o(n_12975) );
na02s06 g768334 ( .a(n_12584), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_14_), .o(n_12618) );
in01s01 g768335 ( .a(n_12533), .o(n_12534) );
na02s02 g768336 ( .a(n_12484), .b(n_12512), .o(n_12533) );
no02m08 g768339 ( .a(n_12590), .b(n_12355), .o(n_12607) );
na02s01 g768340 ( .a(n_12509), .b(n_12508), .o(n_12510) );
in01m02 g768341 ( .a(n_12592), .o(n_12593) );
na02m02 g768342 ( .a(n_12583), .b(n_12554), .o(n_12592) );
na02s06 g768343 ( .a(n_12469), .b(n_12468), .o(n_12522) );
no02s06 TIMEBOOST_cell_6654 ( .a(TIMEBOOST_net_2084), .b(n_14145), .o(n_14359) );
in01m02 g768345 ( .a(n_12947), .o(n_12617) );
no02m06 g768346 ( .a(n_12584), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_14_), .o(n_12947) );
oa12s01 g768349 ( .a(n_12054), .b(n_12460), .c(n_11896), .o(n_12545) );
ao12s01 g768350 ( .a(n_12472), .b(n_12471), .c(n_12470), .o(n_12840) );
ao12s01 g768351 ( .a(n_12444), .b(n_12443), .c(n_12442), .o(n_12838) );
in01m02 g768352 ( .a(n_12579), .o(n_12580) );
no02s06 TIMEBOOST_cell_7758 ( .a(n_19463), .b(FE_OCP_RBN1829_n_19528), .o(TIMEBOOST_net_2510) );
no02f08 g768355 ( .a(n_12459), .b(n_12053), .o(n_12514) );
na02s01 TIMEBOOST_cell_6053 ( .a(n_7), .b(n_745), .o(TIMEBOOST_net_1878) );
no02m02 g768357 ( .a(n_12542), .b(n_12541), .o(n_12543) );
no02s01 TIMEBOOST_cell_4223 ( .a(FE_OCP_RBN4007_n_32860), .b(n_32991), .o(TIMEBOOST_net_1202) );
in01s02 g768359 ( .a(n_12554), .o(n_12555) );
na02s02 g768360 ( .a(n_12523), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_13_), .o(n_12554) );
in01s03 g768361 ( .a(n_12490), .o(n_12465) );
na02s20 g768362 ( .a(n_12320), .b(n_12445), .o(n_12490) );
in01s01 g768363 ( .a(n_12483), .o(n_12484) );
no02s08 g768364 ( .a(n_12464), .b(delay_add_ln22_unr8_stage4_stallmux_q_13_), .o(n_12483) );
na02s06 g768365 ( .a(n_12464), .b(delay_add_ln22_unr8_stage4_stallmux_q_13_), .o(n_12512) );
na02m08 g768366 ( .a(n_12529), .b(n_12324), .o(n_12590) );
na02m06 g768367 ( .a(n_12524), .b(n_11101), .o(n_12583) );
in01m02 g768368 ( .a(n_12577), .o(n_12578) );
na02m04 g768369 ( .a(n_12540), .b(n_12564), .o(n_12577) );
in01s02 g768370 ( .a(n_12520), .o(n_12521) );
na02m02 g768371 ( .a(n_12506), .b(n_12480), .o(n_12520) );
no02s01 g768372 ( .a(n_12471), .b(n_12470), .o(n_12472) );
no02s01 g768373 ( .a(n_12443), .b(n_12442), .o(n_12444) );
in01s01 g768374 ( .a(n_12519), .o(n_12482) );
ao12m08 g768375 ( .a(n_12192), .b(n_12467), .c(n_12270), .o(n_12519) );
ao12s01 g768376 ( .a(n_12228), .b(n_12481), .c(n_12294), .o(n_12509) );
ao12s01 g768377 ( .a(n_11898), .b(n_12413), .c(n_11960), .o(n_12486) );
ao22s01 g768378 ( .a(n_12481), .b(n_12315), .c(n_12450), .d(n_12314), .o(n_13510) );
oa12s01 g768379 ( .a(n_12441), .b(n_12467), .c(n_12440), .o(n_13495) );
na03f02 TIMEBOOST_cell_5766 ( .a(n_8619), .b(FE_OCPN935_n_7802), .c(n_8595), .o(TIMEBOOST_net_1551) );
no02m02 g768382 ( .a(n_12504), .b(n_12239), .o(n_12505) );
in01m04 g768383 ( .a(n_12542), .o(n_12529) );
na02m08 g768384 ( .a(n_12504), .b(n_12149), .o(n_12542) );
na02s01 g768385 ( .a(n_12467), .b(n_12440), .o(n_12441) );
na02s06 g768387 ( .a(n_12463), .b(n_12462), .o(n_12506) );
in01s01 g768388 ( .a(n_12479), .o(n_12480) );
no02s06 g768389 ( .a(n_12463), .b(n_12462), .o(n_12479) );
in01s01 g768390 ( .a(n_12445), .o(n_12427) );
na02s06 g768392 ( .a(n_12528), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_12_), .o(n_12564) );
in01s02 g768393 ( .a(n_12526), .o(n_12527) );
na02m02 g768394 ( .a(n_12476), .b(n_12507), .o(n_12526) );
na02f04 TIMEBOOST_cell_8813 ( .a(TIMEBOOST_net_2893), .b(n_14799), .o(n_14901) );
in01s02 g768397 ( .a(n_12539), .o(n_12540) );
no02m06 g768398 ( .a(n_12528), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_12_), .o(n_12539) );
in01s02 g768399 ( .a(n_12500), .o(n_12501) );
na02s01 g768401 ( .a(n_12449), .b(n_11976), .o(n_12471) );
oa12s02 g768402 ( .a(n_12414), .b(n_12381), .c(FE_OCP_RBN2402_n_45697), .o(n_12734) );
oa12s01 g768403 ( .a(n_12461), .b(n_12404), .c(FE_OCP_RBN2406_n_45697), .o(n_12760) );
in01s01 g768404 ( .a(n_12459), .o(n_12460) );
oa12s01 g768406 ( .a(n_12115), .b(n_12418), .c(n_12007), .o(n_12443) );
oa22s01 g768407 ( .a(n_12373), .b(n_12165), .c(n_12418), .d(n_12166), .o(n_12909) );
in01m02 g768409 ( .a(n_12523), .o(n_12524) );
no02s02 g768411 ( .a(n_12492), .b(n_12477), .o(n_12478) );
no02m02 TIMEBOOST_cell_3988 ( .a(n_24473), .b(TIMEBOOST_net_1084), .o(n_24581) );
na02s04 g768413 ( .a(n_12361), .b(n_12208), .o(n_12376) );
in01m01 g768414 ( .a(n_12504), .o(n_12499) );
no02m08 g768415 ( .a(n_12492), .b(n_12147), .o(n_12504) );
in01s01 g768416 ( .a(n_12414), .o(n_12415) );
na02s04 g768417 ( .a(n_12381), .b(FE_OCP_RBN2402_n_45697), .o(n_12414) );
na02s01 g768419 ( .a(FE_OCP_RBN2406_n_45697), .b(n_12404), .o(n_12461) );
na02s02 g768420 ( .a(n_12361), .b(n_12059), .o(n_12362) );
no02s06 g768422 ( .a(n_12428), .b(delay_add_ln22_unr8_stage4_stallmux_q_11_), .o(n_12438) );
na02s06 g768423 ( .a(n_12453), .b(n_12452), .o(n_12507) );
in01s02 g768424 ( .a(n_12447), .o(n_12448) );
na02m01 g768425 ( .a(n_12391), .b(n_12420), .o(n_12447) );
in01s01 g768426 ( .a(n_12475), .o(n_12476) );
no02m04 g768427 ( .a(n_12453), .b(n_12452), .o(n_12475) );
in01s01 g768428 ( .a(n_12497), .o(n_12498) );
na02s03 g768429 ( .a(n_12474), .b(n_12433), .o(n_12497) );
na02s06 g768430 ( .a(n_12428), .b(delay_add_ln22_unr8_stage4_stallmux_q_11_), .o(n_12491) );
in01f06 g768431 ( .a(n_12413), .o(n_12449) );
in01s01 g768433 ( .a(n_12495), .o(n_12496) );
oa12s02 g768434 ( .a(n_12434), .b(FE_OCP_RBN2404_n_45697), .c(delay_xor_ln21_unr9_stage4_stallmux_q_22_), .o(n_12495) );
na02s06 g768436 ( .a(n_12374), .b(FE_RN_1387_0), .o(n_12560) );
ao12s02 g768437 ( .a(n_12400), .b(FE_OCP_RBN2404_n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_20_), .o(n_12631) );
in01s01 g768438 ( .a(n_12450), .o(n_12481) );
oa12m08 g768440 ( .a(n_12251), .b(n_12412), .c(n_12186), .o(n_12467) );
in01s01 g768441 ( .a(FE_OCP_DRV_N5358_n_12436), .o(n_12437) );
oa22s01 g768442 ( .a(n_12366), .b(n_12287), .c(n_12412), .d(n_12288), .o(n_12436) );
oa12s01 g768443 ( .a(n_12379), .b(n_12378), .c(n_12377), .o(n_13434) );
ao12m04 g768445 ( .a(n_12458), .b(n_12457), .c(n_12456), .o(n_12528) );
in01s03 g768446 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_20_), .o(n_12381) );
in01s01 g768448 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_21_), .o(n_12404) );
na02s01 g768451 ( .a(n_12398), .b(n_12354), .o(n_12596) );
no02s06 g768453 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_18_), .b(FE_OCP_RBN2399_n_45697), .o(n_12396) );
na02s01 g768455 ( .a(n_12378), .b(n_12377), .o(n_12379) );
in01s02 g768456 ( .a(n_12391), .o(n_12392) );
na02s02 g768457 ( .a(n_12350), .b(delay_add_ln22_unr8_stage4_stallmux_q_10_), .o(n_12391) );
in01m10 g768458 ( .a(n_12361), .o(n_12401) );
no02s02 TIMEBOOST_cell_1659 ( .a(n_44594), .b(n_8781), .o(TIMEBOOST_net_444) );
no02s02 TIMEBOOST_cell_5667 ( .a(TIMEBOOST_net_1781), .b(n_17216), .o(n_17384) );
no02m04 g768461 ( .a(n_12457), .b(n_12456), .o(n_12458) );
in01s01 g768463 ( .a(n_12434), .o(n_12435) );
na02s06 g768464 ( .a(FE_OCP_RBN2404_n_45697), .b(delay_xor_ln21_unr9_stage4_stallmux_q_22_), .o(n_12434) );
na02s06 g768465 ( .a(n_12419), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_10_), .o(n_12474) );
in01s02 g768466 ( .a(n_12432), .o(n_12433) );
no02s06 g768467 ( .a(n_12419), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_10_), .o(n_12432) );
na02s01 g768468 ( .a(n_12424), .b(n_12385), .o(n_12587) );
na02s01 g768469 ( .a(FE_OCP_RBN2406_n_45697), .b(n_12318), .o(n_12431) );
no02s02 g768470 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_20_), .b(FE_OCP_RBN2404_n_45697), .o(n_12400) );
na02s01 g768471 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_18_), .b(FE_OCP_RBN2399_n_45697), .o(n_12374) );
in01s01 g768473 ( .a(n_12418), .o(n_12373) );
ao12f08 g768474 ( .a(n_12298), .b(n_12302), .c(n_11707), .o(n_12418) );
ao12s06 g768475 ( .a(n_12355), .b(FE_OCP_RBN2399_n_45697), .c(delay_xor_ln21_unr9_stage4_stallmux_q_16_), .o(n_12581) );
oa12s01 g768476 ( .a(n_12384), .b(n_12338), .c(FE_OCP_RBN2402_n_45697), .o(n_12674) );
in01s01 g768477 ( .a(n_12454), .o(n_12455) );
oa12s01 g768478 ( .a(n_12406), .b(FE_OCP_RBN2404_n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_22_), .o(n_12454) );
ao12s02 g768479 ( .a(n_12372), .b(FE_OCP_RBN2399_n_45697), .c(delay_xor_ln21_unr9_stage4_stallmux_q_18_), .o(n_12642) );
oa12s02 g768480 ( .a(n_12411), .b(n_12360), .c(FE_OCP_RBN2402_n_45697), .o(n_12606) );
ao12s01 g768482 ( .a(n_12358), .b(n_12357), .c(n_12356), .o(n_13074) );
in01s01 g768486 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_21_), .o(n_12318) );
in01s02 g768489 ( .a(n_12423), .o(n_12457) );
no02s06 g768490 ( .a(FE_OCP_RBN2461_n_12365), .b(n_12043), .o(n_12423) );
na02s06 g768491 ( .a(n_12336), .b(delay_add_ln22_unr8_stage4_stallmux_q_9_), .o(n_12398) );
in01s01 g768492 ( .a(n_12353), .o(n_12354) );
no02s06 g768493 ( .a(n_12336), .b(delay_add_ln22_unr8_stage4_stallmux_q_9_), .o(n_12353) );
na02s10 g768494 ( .a(n_12352), .b(n_11899), .o(n_12394) );
no02s01 g768495 ( .a(n_12357), .b(n_12356), .o(n_12358) );
in01s01 g768496 ( .a(n_12408), .o(n_12409) );
na02s01 g768497 ( .a(n_12347), .b(n_12389), .o(n_12408) );
na02s03 g768498 ( .a(n_12338), .b(FE_OCP_RBN2402_n_45697), .o(n_12384) );
no02s06 g768499 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_18_), .b(FE_OCP_RBN2399_n_45697), .o(n_12372) );
na02s01 g768500 ( .a(n_12299), .b(n_12335), .o(n_12551) );
in01s02 g768501 ( .a(n_12385), .o(n_12386) );
na02s02 g768502 ( .a(n_12342), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_9_), .o(n_12385) );
no02m06 g768503 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_16_), .b(FE_OCP_RBN2399_n_45697), .o(n_12355) );
na02s06 g768504 ( .a(n_12360), .b(FE_OCP_RBN2397_n_45697), .o(n_12411) );
na02s01 g768507 ( .a(FE_OCP_RBN2404_n_45697), .b(delay_xor_ln22_unr9_stage4_stallmux_q_22_), .o(n_12406) );
oa12s01 g768508 ( .a(n_12371), .b(n_12327), .c(FE_OCP_RBN2402_n_45697), .o(n_12570) );
ao12s06 g768509 ( .a(n_12370), .b(FE_OCP_RBN2394_n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_16_), .o(n_12488) );
in01s01 g768510 ( .a(n_12387), .o(n_12388) );
ao12s01 g768511 ( .a(n_12368), .b(FE_OCP_RBN2399_n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_17_), .o(n_12387) );
in01s01 g768512 ( .a(n_12412), .o(n_12366) );
ao12m08 g768513 ( .a(n_12180), .b(n_12341), .c(n_12273), .o(n_12412) );
oa12m06 g768514 ( .a(n_12248), .b(n_12334), .c(n_12182), .o(n_12378) );
ao22s01 g768517 ( .a(n_12286), .b(n_12334), .c(n_12285), .d(n_12291), .o(n_13366) );
ao12s01 g768518 ( .a(n_12332), .b(n_12331), .c(n_12341), .o(n_13330) );
oa22s06 g768520 ( .a(n_12267), .b(n_11939), .c(n_12333), .d(n_11938), .o(n_12350) );
no02s06 g768521 ( .a(n_12345), .b(n_12339), .o(n_12419) );
in01m03 g768522 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_17_), .o(n_12360) );
in01s01 g768525 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_29_), .o(n_13086) );
in01s03 g768527 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_19_), .o(n_12338) );
na02f08 g768532 ( .a(n_12268), .b(n_12164), .o(n_12302) );
no02s01 g768533 ( .a(n_12269), .b(n_12193), .o(n_12357) );
no02s01 g768535 ( .a(n_12331), .b(n_12341), .o(n_12332) );
in01s03 g768536 ( .a(FE_OCPN1360_n_12370), .o(n_12349) );
no02s20 g768537 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_16_), .b(FE_OCP_RBN2394_n_45697), .o(n_12370) );
no02s06 g768539 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_17_), .b(FE_OCP_RBN2399_n_45697), .o(n_12368) );
no02s20 g768541 ( .a(FE_OCPN1717_n_12311), .b(n_12333), .o(n_12352) );
in01s02 g768542 ( .a(n_12299), .o(n_12300) );
na02s02 g768543 ( .a(n_12230), .b(delay_add_ln22_unr8_stage4_stallmux_q_8_), .o(n_12299) );
in01s01 g768544 ( .a(n_12346), .o(n_12347) );
no02s06 g768545 ( .a(n_12316), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_8_), .o(n_12346) );
na02s03 g768546 ( .a(n_12316), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_8_), .o(n_12389) );
no02s06 g768547 ( .a(FE_OCP_RBN2447_n_12312), .b(n_11945), .o(n_12345) );
no02s06 g768548 ( .a(n_12312), .b(n_11946), .o(n_12339) );
no02s10 g768550 ( .a(n_11888), .b(FE_OCP_RBN2447_n_12312), .o(n_12365) );
na02s01 g768551 ( .a(FE_RN_400_0), .b(n_12309), .o(n_12508) );
in01s01 g768552 ( .a(n_12328), .o(n_12329) );
na02s01 g768553 ( .a(n_12313), .b(n_12263), .o(n_12328) );
na02s02 g768554 ( .a(n_12327), .b(FE_OCP_RBN2402_n_45697), .o(n_12371) );
na02s06 g768555 ( .a(n_12231), .b(n_10611), .o(n_12335) );
no02s20 TIMEBOOST_cell_6882 ( .a(FE_OCP_RBN3990_n_32772), .b(TIMEBOOST_net_2199), .o(n_32851) );
ao12m08 g768557 ( .a(n_12323), .b(FE_OCP_RBN2394_n_45697), .c(delay_xor_ln21_unr9_stage4_stallmux_q_15_), .o(n_12541) );
ao12s01 g768562 ( .a(n_12243), .b(n_12242), .c(n_12241), .o(n_12850) );
in01s01 g768563 ( .a(n_12325), .o(n_12326) );
ao12s01 g768564 ( .a(n_12266), .b(n_12265), .c(n_12264), .o(n_12325) );
ao12s02 g768566 ( .a(n_12297), .b(n_12296), .c(n_12295), .o(n_12342) );
no02f06 TIMEBOOST_cell_6744 ( .a(TIMEBOOST_net_2129), .b(TIMEBOOST_net_1098), .o(n_9086) );
in01s01 g768570 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_27_), .o(n_12271) );
in01s02 g768575 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_19_), .o(n_12327) );
na02s02 g768577 ( .a(n_12146), .b(n_11901), .o(n_12161) );
no02m04 TIMEBOOST_cell_6743 ( .a(FE_OCP_RBN2865_n_8850), .b(FE_OCP_RBN5748_n_8637), .o(TIMEBOOST_net_2129) );
na02s01 g768579 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_24_), .b(delay_add_ln22_unr8_stage4_stallmux_q_25_), .o(n_12892) );
no02s01 g768580 ( .a(n_12296), .b(n_12295), .o(n_12297) );
na02s01 g768581 ( .a(n_12191), .b(n_12270), .o(n_12440) );
in01s01 g768582 ( .a(n_12268), .o(n_12269) );
no02f08 g768583 ( .a(n_12234), .b(n_11795), .o(n_12268) );
no02s06 TIMEBOOST_cell_6130 ( .a(TIMEBOOST_net_1916), .b(n_24372), .o(TIMEBOOST_net_1567) );
in01s10 g768585 ( .a(n_12267), .o(n_12333) );
no02s10 g768586 ( .a(n_12233), .b(n_11860), .o(n_12267) );
no02s01 g768587 ( .a(n_12242), .b(n_12241), .o(n_12243) );
no02s01 g768588 ( .a(n_12265), .b(n_12264), .o(n_12266) );
in01s01 g768589 ( .a(n_12262), .o(n_12263) );
no02s06 g768590 ( .a(n_12232), .b(delay_add_ln22_unr8_stage4_stallmux_q_7_), .o(n_12262) );
in01s01 g768591 ( .a(n_12314), .o(n_12315) );
na02s01 g768592 ( .a(n_12294), .b(n_12293), .o(n_12314) );
in01s02 g768593 ( .a(n_12323), .o(n_12324) );
no02s20 g768594 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_15_), .b(FE_OCP_RBN2394_n_45697), .o(n_12323) );
no02s02 g768596 ( .a(n_12261), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_7_), .o(n_12275) );
na02m08 g768598 ( .a(n_12261), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_7_), .o(n_12309) );
no02s10 g768600 ( .a(n_11885), .b(n_12296), .o(n_12312) );
na02s06 g768601 ( .a(n_12232), .b(delay_add_ln22_unr8_stage4_stallmux_q_7_), .o(n_12313) );
in01s02 g768602 ( .a(n_12363), .o(n_12364) );
ao12s06 g768603 ( .a(n_12319), .b(FE_OCP_RBN2394_n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_15_), .o(n_12363) );
oa12m08 g768604 ( .a(n_12130), .b(n_12292), .c(n_12041), .o(n_12341) );
in01s01 g768605 ( .a(n_12334), .o(n_12291) );
oa12m06 g768606 ( .a(n_12179), .b(n_12092), .c(n_12260), .o(n_12334) );
ao12s01 g768612 ( .a(n_12200), .b(n_12199), .c(n_12198), .o(n_12738) );
in01s01 g768613 ( .a(n_12256), .o(n_12257) );
ao12s01 g768614 ( .a(n_12141), .b(n_12140), .c(n_12139), .o(n_12256) );
in01s01 g768615 ( .a(n_12289), .o(n_12290) );
oa12s01 g768616 ( .a(n_12203), .b(n_12202), .c(n_12201), .o(n_12289) );
ao12s01 g768617 ( .a(n_12155), .b(n_12154), .c(n_12153), .o(n_12871) );
in01m02 g768620 ( .a(n_12211), .o(n_12151) );
oa22s01 g768622 ( .a(n_12204), .b(n_12225), .c(n_12205), .d(n_12292), .o(n_13264) );
in01s01 g768623 ( .a(n_12321), .o(n_12322) );
ao12s01 g768624 ( .a(n_12250), .b(n_12249), .c(n_12260), .o(n_12321) );
in01s02 g768626 ( .a(n_12230), .o(n_12231) );
in01s01 g768629 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_31_), .o(n_12229) );
in01s01 g768631 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_27_), .o(n_13013) );
in01s01 g768633 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_26_), .o(n_12215) );
na02s01 g768637 ( .a(n_12254), .b(n_12209), .o(n_12255) );
no02s01 g768638 ( .a(n_12199), .b(n_12198), .o(n_12200) );
no02s01 g768639 ( .a(n_12072), .b(n_12193), .o(n_12265) );
no02s01 g768642 ( .a(n_12140), .b(n_12139), .o(n_12141) );
na02s01 g768643 ( .a(n_12202), .b(n_12201), .o(n_12203) );
in01s06 g768644 ( .a(n_12191), .o(n_12192) );
na02s06 g768645 ( .a(n_12100), .b(delay_add_ln22_unr8_stage4_stallmux_q_6_), .o(n_12191) );
in01s06 g768646 ( .a(n_12319), .o(n_12320) );
no02s20 g768647 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_15_), .b(FE_OCPN1606_n_45697), .o(n_12319) );
in01s06 g768648 ( .a(n_12146), .o(n_12233) );
no02s10 g768649 ( .a(n_12106), .b(n_11840), .o(n_12146) );
na02s01 g768651 ( .a(n_12253), .b(n_12252), .o(n_12377) );
in01s01 g768652 ( .a(n_12287), .o(n_12288) );
na02s01 g768653 ( .a(n_12187), .b(n_12251), .o(n_12287) );
na02s10 g768654 ( .a(n_47211), .b(n_11757), .o(n_12296) );
in01s02 g768655 ( .a(n_12228), .o(n_12293) );
no02s06 g768656 ( .a(n_12195), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_6_), .o(n_12228) );
na02m06 g768658 ( .a(n_12195), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_6_), .o(n_12294) );
no02s01 g768659 ( .a(n_12249), .b(n_12260), .o(n_12250) );
no02s01 g768660 ( .a(n_12154), .b(n_12153), .o(n_12155) );
no02s01 g768661 ( .a(n_12104), .b(n_11825), .o(n_12242) );
in01s02 g768665 ( .a(n_12197), .o(n_12116) );
in01s02 g768668 ( .a(n_12217), .o(n_12190) );
in01m02 g768673 ( .a(n_12240), .o(n_12189) );
in01s01 g768675 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_25_), .o(n_12209) );
in01s01 g768678 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_28_), .o(n_12188) );
no02s01 g768683 ( .a(n_12108), .b(n_11711), .o(n_12104) );
na02s02 g768684 ( .a(n_12098), .b(n_10371), .o(n_12253) );
in01s01 g768685 ( .a(n_12186), .o(n_12187) );
no02s08 g768686 ( .a(n_12137), .b(delay_add_ln22_unr8_stage4_stallmux_q_5_), .o(n_12186) );
na02m06 g768687 ( .a(n_12137), .b(delay_add_ln22_unr8_stage4_stallmux_q_5_), .o(n_12251) );
in01s01 g768688 ( .a(n_47211), .o(n_12185) );
na02s06 g768690 ( .a(n_12099), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_5_), .o(n_12252) );
in01s01 g768691 ( .a(n_12285), .o(n_12286) );
na02s01 g768692 ( .a(n_12183), .b(n_12248), .o(n_12285) );
na02s01 g768693 ( .a(n_12181), .b(n_12273), .o(n_12331) );
na02s01 g768694 ( .a(n_12108), .b(n_11852), .o(n_12154) );
oa12s01 g768695 ( .a(n_11571), .b(n_44451), .c(n_11890), .o(n_12199) );
no02s01 g768696 ( .a(n_12108), .b(n_12071), .o(n_12072) );
ao12s01 g768697 ( .a(n_11728), .b(n_44450), .c(n_11632), .o(n_12140) );
oa12s01 g768698 ( .a(n_11935), .b(n_44451), .c(n_12003), .o(n_12202) );
in01s01 g768699 ( .a(n_12292), .o(n_12225) );
in01s02 g768701 ( .a(n_12238), .o(n_12239) );
ao12m06 g768702 ( .a(n_12148), .b(FE_OCP_RBN2394_n_45697), .c(delay_xor_ln21_unr9_stage4_stallmux_q_14_), .o(n_12238) );
oa12m06 g768703 ( .a(n_12019), .b(n_12173), .c(n_12091), .o(n_12260) );
ao12s06 g768704 ( .a(n_12136), .b(FE_OCPN1606_n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_14_), .o(n_12416) );
in01s01 g768705 ( .a(n_13054), .o(n_12245) );
oa12s01 g768706 ( .a(n_12123), .b(n_12122), .c(n_12121), .o(n_13054) );
oa12s01 g768707 ( .a(n_12175), .b(n_12174), .c(n_12173), .o(n_13095) );
in01m02 g768709 ( .a(n_12145), .o(n_12102) );
oa22s01 g768711 ( .a(n_44450), .b(n_12049), .c(n_44451), .d(n_12048), .o(n_12720) );
in01s01 g768712 ( .a(n_12134), .o(n_12135) );
ao12s01 g768713 ( .a(n_12031), .b(n_12030), .c(n_12029), .o(n_12134) );
in01s02 g768714 ( .a(n_12068), .o(n_12064) );
in01s02 g768716 ( .a(n_12158), .o(n_12133) );
ao12s02 g768720 ( .a(n_11617), .b(n_12024), .c(n_11752), .o(n_12025) );
oa12s02 g768721 ( .a(n_11580), .b(n_11989), .c(n_11712), .o(n_11990) );
oa12m04 g768722 ( .a(n_11613), .b(n_12024), .c(n_11656), .o(n_12023) );
ao12s04 g768723 ( .a(n_11578), .b(n_11989), .c(n_11716), .o(n_11988) );
in01m02 g768724 ( .a(n_12162), .o(n_12132) );
in01s01 g768726 ( .a(n_12247), .o(n_12942) );
oa12s01 g768727 ( .a(n_12126), .b(n_12125), .c(n_12124), .o(n_12247) );
in01s01 g768728 ( .a(n_12283), .o(n_12284) );
oa12s01 g768729 ( .a(n_12178), .b(n_12177), .c(n_12176), .o(n_12283) );
in01s01 g768733 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_24_), .o(n_12834) );
in01s06 g768735 ( .a(n_12148), .o(n_12149) );
no02s20 g768736 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_14_), .b(FE_OCP_RBN2394_n_45697), .o(n_12148) );
in01s01 g768737 ( .a(n_12204), .o(n_12205) );
na02s01 g768738 ( .a(n_12130), .b(n_12042), .o(n_12204) );
na02s06 g768739 ( .a(n_12129), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_4_), .o(n_12248) );
na02s10 g768740 ( .a(n_11998), .b(FE_OCPN4935_n_11993), .o(n_12039) );
na02s08 g768742 ( .a(n_12128), .b(n_12127), .o(n_12273) );
in01s01 g768745 ( .a(n_12182), .o(n_12183) );
no02s06 g768746 ( .a(n_12129), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_4_), .o(n_12182) );
no02m06 g768747 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_14_), .b(FE_OCPN1606_n_45697), .o(n_12136) );
in01s01 g768748 ( .a(n_12180), .o(n_12181) );
no02s08 g768749 ( .a(n_12128), .b(n_12127), .o(n_12180) );
na02s06 g768750 ( .a(n_11998), .b(n_11997), .o(n_11999) );
na02s01 g768751 ( .a(n_12125), .b(n_12124), .o(n_12126) );
na02s01 g768752 ( .a(n_12093), .b(n_12179), .o(n_12249) );
na02s01 g768753 ( .a(n_12122), .b(n_12121), .o(n_12123) );
no02s01 g768754 ( .a(n_12030), .b(n_12029), .o(n_12031) );
na02s01 g768755 ( .a(n_12177), .b(n_12176), .o(n_12178) );
na02s01 g768756 ( .a(n_12174), .b(n_12173), .o(n_12175) );
na02f10 g768757 ( .a(n_12065), .b(n_11758), .o(n_12108) );
in01s01 g768759 ( .a(n_12144), .o(n_12112) );
ao12s02 g768761 ( .a(n_12035), .b(n_12034), .c(n_12033), .o(n_12789) );
in01s01 g768762 ( .a(n_12223), .o(n_12224) );
ao12s01 g768763 ( .a(n_12096), .b(n_12095), .c(n_12094), .o(n_12223) );
in01m02 g768764 ( .a(n_12027), .o(n_12028) );
na02f02 TIMEBOOST_cell_5582 ( .a(n_11063), .b(n_11197), .o(TIMEBOOST_net_1739) );
oa12s02 g768768 ( .a(n_11698), .b(n_11958), .c(n_11924), .o(n_11964) );
no02s04 g768769 ( .a(n_11925), .b(n_11654), .o(n_11987) );
in01s02 g768771 ( .a(n_12098), .o(n_12099) );
na02s01 TIMEBOOST_cell_7899 ( .a(TIMEBOOST_net_2580), .b(n_35956), .o(TIMEBOOST_net_1304) );
oa12s02 g768773 ( .a(n_11598), .b(n_11914), .c(n_11520), .o(n_11986) );
ao12s02 g768774 ( .a(n_11478), .b(n_45748), .c(n_11518), .o(n_12022) );
in01s02 g768775 ( .a(n_12037), .o(n_12114) );
ao22m02 g768776 ( .a(n_11958), .b(FE_OCP_RBN3425_n_11754), .c(n_11754), .d(n_11874), .o(n_12037) );
ao12s02 g768777 ( .a(n_11677), .b(n_11459), .c(n_11958), .o(n_11959) );
oa12s04 g768778 ( .a(n_11715), .b(n_11874), .c(n_11514), .o(n_11985) );
in01s01 g768780 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_24_), .o(n_12254) );
na02s06 g768783 ( .a(n_12026), .b(n_11983), .o(n_11984) );
na02s03 g768784 ( .a(n_11956), .b(n_11766), .o(n_11957) );
na02f06 TIMEBOOST_cell_6766 ( .a(TIMEBOOST_net_2140), .b(n_16442), .o(n_16466) );
no02s01 g768786 ( .a(n_12097), .b(n_12069), .o(n_12177) );
no02m06 TIMEBOOST_cell_1598 ( .a(TIMEBOOST_net_413), .b(n_35196), .o(n_35262) );
no02s01 g768788 ( .a(n_12095), .b(n_12094), .o(n_12096) );
in01s01 g768789 ( .a(n_12041), .o(n_12042) );
no02s06 g768790 ( .a(n_12021), .b(delay_add_ln22_unr8_stage4_stallmux_q_3_), .o(n_12041) );
na02s08 g768792 ( .a(n_11956), .b(n_11955), .o(n_11994) );
na02m10 g768793 ( .a(n_11956), .b(n_11955), .o(n_11962) );
na02s06 g768794 ( .a(n_12062), .b(n_12061), .o(n_12179) );
in01s01 g768795 ( .a(n_12092), .o(n_12093) );
no02s06 g768796 ( .a(n_12062), .b(n_12061), .o(n_12092) );
no02s01 g768797 ( .a(n_12020), .b(n_12091), .o(n_12174) );
na02s06 g768798 ( .a(n_12021), .b(delay_add_ln22_unr8_stage4_stallmux_q_3_), .o(n_12130) );
no02s01 g768799 ( .a(n_12034), .b(n_12033), .o(n_12035) );
no02s02 g768800 ( .a(n_11958), .b(n_11924), .o(n_11925) );
ao12m08 g768801 ( .a(n_12147), .b(n_45685), .c(delay_xor_ln21_unr9_stage4_stallmux_q_13_), .o(n_12477) );
in01s01 g768802 ( .a(n_12207), .o(n_12208) );
ao12s02 g768803 ( .a(n_12402), .b(FE_OCPN1606_n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_13_), .o(n_12207) );
na02s06 g768804 ( .a(n_11853), .b(n_11776), .o(n_11989) );
no02m08 g768805 ( .a(FE_OCP_RBN6237_n_11853), .b(n_11847), .o(n_12024) );
oa12f10 g768807 ( .a(n_11687), .b(n_11929), .c(n_11635), .o(n_12065) );
oa12s02 g768808 ( .a(FE_OCP_RBN3407_n_11560), .b(n_11915), .c(n_11870), .o(n_11954) );
na02s01 TIMEBOOST_cell_4185 ( .a(n_27462), .b(FE_RN_345_0), .o(TIMEBOOST_net_1183) );
in01s02 g768810 ( .a(n_11922), .o(n_11923) );
oa12s04 g768811 ( .a(n_11753), .b(n_11823), .c(n_11676), .o(n_11922) );
oa12s01 g768812 ( .a(n_11648), .b(n_11929), .c(n_11631), .o(n_12030) );
in01m02 g768813 ( .a(n_12060), .o(n_12131) );
in01m02 g768815 ( .a(n_11952), .o(n_11953) );
ao12s06 g768816 ( .a(n_11685), .b(n_11850), .c(n_11597), .o(n_11952) );
no02s01 TIMEBOOST_cell_5581 ( .a(FE_OCP_RBN3342_n_39942), .b(TIMEBOOST_net_1738), .o(n_40271) );
ao12s01 g768818 ( .a(n_11966), .b(n_12005), .c(delay_add_ln22_unr8_stage4_stallmux_q_1_), .o(n_12125) );
ao12m08 g768819 ( .a(n_11872), .b(n_12005), .c(n_11875), .o(n_12176) );
na02m04 g768821 ( .a(n_11822), .b(n_11883), .o(n_11980) );
ao12m06 g768822 ( .a(n_11880), .b(n_11884), .c(n_12036), .o(n_12173) );
ao12s01 g768823 ( .a(n_11996), .b(n_12036), .c(delay_sub_ln21_0_unr8_stage4_stallmux_q_1_), .o(n_12122) );
na02m04 TIMEBOOST_cell_7089 ( .a(n_36565), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_2303) );
no02s01 g768827 ( .a(n_11876), .b(n_11686), .o(n_12034) );
na03f04 TIMEBOOST_cell_7339 ( .a(n_37717), .b(n_37760), .c(FE_OCP_RBN4033_n_37690), .o(n_37761) );
na02m08 TIMEBOOST_cell_6672 ( .a(TIMEBOOST_net_2093), .b(n_24522), .o(n_24683) );
no02s01 g768830 ( .a(n_12005), .b(delay_add_ln22_unr8_stage4_stallmux_q_1_), .o(n_11966) );
no02m06 g768831 ( .a(n_11941), .b(delay_add_ln22_unr8_stage4_stallmux_q_2_), .o(n_12069) );
in01s02 g768833 ( .a(n_11956), .o(n_11917) );
in01s01 g768835 ( .a(n_12019), .o(n_12020) );
na02m06 g768836 ( .a(n_11978), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_2_), .o(n_12019) );
no02m06 g768837 ( .a(n_11978), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_2_), .o(n_12091) );
no02s01 g768839 ( .a(n_12036), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_1_), .o(n_11996) );
in01s01 g768840 ( .a(n_12402), .o(n_12059) );
no02m03 g768841 ( .a(FE_OCPN1606_n_45697), .b(delay_xor_ln22_unr9_stage4_stallmux_q_13_), .o(n_12402) );
no02m06 g768842 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_13_), .b(n_45685), .o(n_12147) );
ao12s04 g768843 ( .a(n_12056), .b(n_45685), .c(delay_xor_ln21_unr9_stage4_stallmux_q_12_), .o(n_12456) );
oa12s01 g768844 ( .a(n_11933), .b(n_12088), .c(n_12011), .o(n_12095) );
no02m04 TIMEBOOST_cell_4184 ( .a(n_22476), .b(TIMEBOOST_net_1182), .o(FE_RN_1327_0) );
ao12m02 g768846 ( .a(n_11821), .b(n_11699), .c(FE_OCP_RBN4480_n_11439), .o(n_11822) );
ao12s02 g768849 ( .a(n_11836), .b(n_11835), .c(n_11834), .o(n_12699) );
in01s01 g768850 ( .a(n_12221), .o(n_12222) );
oa12s01 g768851 ( .a(n_12089), .b(n_12088), .c(n_12087), .o(n_12221) );
in01s02 g768854 ( .a(n_12058), .o(n_12150) );
na02f04 TIMEBOOST_cell_6784 ( .a(TIMEBOOST_net_2149), .b(n_9971), .o(n_10198) );
oa12s01 g768860 ( .a(n_11657), .b(n_44356), .c(n_11647), .o(n_11913) );
ao12s02 g768861 ( .a(n_11458), .b(n_44355), .c(n_11658), .o(n_11947) );
in01s03 g768864 ( .a(n_11958), .o(n_11874) );
no02s06 g768867 ( .a(n_11736), .b(n_11821), .o(n_11958) );
in01s01 g768869 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_23_), .o(n_11886) );
na02m08 g768874 ( .a(n_12124), .b(n_11871), .o(n_11875) );
in01s06 g768875 ( .a(n_11909), .o(n_11910) );
no02s10 g768876 ( .a(n_11927), .b(n_11919), .o(n_11909) );
no02m08 g768877 ( .a(n_12124), .b(n_11871), .o(n_11872) );
no02s03 g768880 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_12_), .b(n_45685), .o(n_12056) );
no02s06 g768881 ( .a(n_12121), .b(n_11879), .o(n_11880) );
na02s06 g768882 ( .a(n_12121), .b(n_11879), .o(n_11884) );
in01s01 g768884 ( .a(n_11929), .o(n_11876) );
na02f10 g768885 ( .a(n_11787), .b(n_11543), .o(n_11929) );
no02s01 g768886 ( .a(n_11835), .b(n_11834), .o(n_11836) );
no02m06 g768887 ( .a(n_11847), .b(n_11723), .o(n_11848) );
na02s01 g768888 ( .a(n_12088), .b(n_12087), .o(n_12089) );
na02s06 TIMEBOOST_cell_4216 ( .a(TIMEBOOST_net_1198), .b(n_12427), .o(n_12530) );
no02s04 g768890 ( .a(n_11726), .b(n_11661), .o(n_11736) );
in01s03 g768891 ( .a(n_11945), .o(n_11946) );
ao12s06 g768892 ( .a(n_11888), .b(FE_OCPN7085_n_45697), .c(delay_xor_ln21_unr9_stage4_stallmux_q_10_), .o(n_11945) );
ao12s01 g768893 ( .a(n_12055), .b(n_45685), .c(delay_xor_ln22_unr9_stage4_stallmux_q_12_), .o(n_12393) );
in01s01 g768894 ( .a(n_11944), .o(n_12724) );
ao12s01 g768895 ( .a(n_11846), .b(n_11845), .c(delay_add_ln22_unr8_stage4_stallmux_q_0_), .o(n_11944) );
in01s04 g768899 ( .a(n_11850), .o(n_11870) );
in01s06 g768901 ( .a(n_11823), .o(n_11850) );
in01s06 g768902 ( .a(n_11777), .o(n_11823) );
na02m02 g768906 ( .a(n_44356), .b(n_11662), .o(n_11883) );
in01s01 g768907 ( .a(n_12747), .o(n_11943) );
oa12s01 g768908 ( .a(n_11843), .b(n_11842), .c(delay_sub_ln21_0_unr8_stage4_stallmux_q_0_), .o(n_12747) );
in01s06 g768913 ( .a(n_11927), .o(n_11833) );
no02s01 g768915 ( .a(n_11845), .b(delay_add_ln22_unr8_stage4_stallmux_q_0_), .o(n_11846) );
no02s06 g768916 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_12_), .b(FE_OCPN1606_n_45697), .o(n_12055) );
no02s01 g768917 ( .a(n_12053), .b(n_11895), .o(n_12054) );
na02m10 g768918 ( .a(n_11760), .b(delay_add_ln22_unr8_stage4_stallmux_q_0_), .o(n_12124) );
no02s10 g768920 ( .a(n_11881), .b(n_11844), .o(n_11907) );
no02m08 g768921 ( .a(n_11761), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_0_), .o(n_12121) );
no02s10 g768922 ( .a(n_45697), .b(delay_xor_ln21_unr9_stage4_stallmux_q_10_), .o(n_11888) );
na02s01 g768923 ( .a(n_11842), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_0_), .o(n_11843) );
na02s01 g768924 ( .a(n_12213), .b(n_11968), .o(n_12220) );
na02s01 g768925 ( .a(n_12213), .b(n_12168), .o(n_12214) );
na02s06 g768927 ( .a(n_11600), .b(n_11664), .o(n_11821) );
in01m06 g768928 ( .a(n_11776), .o(n_11847) );
na02m08 TIMEBOOST_cell_7438 ( .a(n_40455), .b(n_40809), .o(TIMEBOOST_net_2350) );
in01s01 g768930 ( .a(n_12110), .o(n_12111) );
ao12s02 g768931 ( .a(n_12043), .b(FE_OCPN1606_n_45697), .c(delay_xor_ln21_unr9_stage4_stallmux_q_11_), .o(n_12110) );
in01s02 g768932 ( .a(n_11938), .o(n_11939) );
ao12s06 g768933 ( .a(n_12311), .b(FE_OCPN1606_n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_10_), .o(n_11938) );
na02s03 g768942 ( .a(n_11698), .b(FE_OCPN1218_n_11012), .o(n_11699) );
oa12s01 g768943 ( .a(n_11525), .b(n_11775), .c(n_11607), .o(n_11835) );
in01s01 g768945 ( .a(n_11787), .o(n_12088) );
oa12f10 g768946 ( .a(n_11637), .b(n_11775), .c(n_11636), .o(n_11787) );
ao22f01 g768949 ( .a(n_11775), .b(n_11680), .c(n_11665), .d(n_11681), .o(n_12692) );
in01s02 g768950 ( .a(n_11873), .o(n_11841) );
no02s02 g768952 ( .a(n_11661), .b(n_11555), .o(n_11662) );
in01s02 g768953 ( .a(n_11778), .o(n_11725) );
in01s01 g768955 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_22_), .o(n_13024) );
in01s01 g768959 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_22_), .o(n_11868) );
na02s20 g768963 ( .a(FE_OCP_RBN5508_FE_RN_1997_0), .b(n_11762), .o(n_11881) );
no02m08 g768964 ( .a(n_11730), .b(FE_OCP_RBN5510_FE_RN_1997_0), .o(n_11819) );
no02s06 g768965 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_10_), .b(FE_OCPN1606_n_45697), .o(n_12311) );
na02s01 g768967 ( .a(n_11852), .b(n_11798), .o(n_11825) );
no02m03 g768968 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_11_), .b(FE_OCPN1606_n_45697), .o(n_12043) );
na02s01 g768969 ( .a(n_12085), .b(n_12084), .o(n_12086) );
oa12m01 g768970 ( .a(n_11976), .b(n_11866), .c(FE_OCP_RBN5445_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_12053) );
in01s08 g768971 ( .a(n_12193), .o(n_11867) );
na02s10 g768972 ( .a(n_11852), .b(n_11751), .o(n_12193) );
in01s06 g768974 ( .a(n_11772), .o(n_11773) );
in01s01 g768976 ( .a(n_12281), .o(n_12213) );
na02s04 g768977 ( .a(n_12085), .b(n_12013), .o(n_12281) );
ao12s01 g768978 ( .a(n_12278), .b(FE_OCP_RBN2394_n_45697), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_29_), .o(n_12706) );
in01s06 g768979 ( .a(n_11734), .o(n_11735) );
in01m08 g768981 ( .a(n_11817), .o(n_11818) );
ao12s06 g768984 ( .a(n_11975), .b(n_45685), .c(delay_xor_ln22_unr9_stage4_stallmux_q_11_), .o(n_12017) );
in01s01 g768985 ( .a(n_11900), .o(n_11901) );
ao12s02 g768986 ( .a(n_11860), .b(FE_OCPN7085_n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_9_), .o(n_11900) );
no02s06 g768987 ( .a(n_11656), .b(n_47279), .o(n_11729) );
in01s01 g768989 ( .a(n_11770), .o(n_11771) );
oa12s06 g768991 ( .a(n_11769), .b(n_11659), .c(FE_OCP_RBN6314_n_45224), .o(n_11983) );
ao12s02 g768992 ( .a(n_11885), .b(FE_OCPN7085_n_45697), .c(delay_xor_ln21_unr9_stage4_stallmux_q_9_), .o(n_12295) );
in01s01 g768993 ( .a(n_11877), .o(n_11878) );
ao12s01 g768994 ( .a(n_11756), .b(n_45697), .c(delay_xor_ln21_unr9_stage4_stallmux_q_8_), .o(n_11877) );
in01s04 g768995 ( .a(n_11815), .o(n_11816) );
ao12s06 g768996 ( .a(n_11780), .b(n_45697), .c(delay_xor_ln21_unr9_stage4_stallmux_q_7_), .o(n_11815) );
ao22s10 g768998 ( .a(n_11595), .b(FE_OCP_RBN3975_n_45224), .c(FE_OCP_RBN6523_n_45224), .d(delay_xor_ln21_unr9_stage4_stallmux_q_6_), .o(n_11767) );
in01s02 g768999 ( .a(n_11765), .o(n_11766) );
ao12s10 g769000 ( .a(n_11693), .b(n_45697), .c(delay_xor_ln21_unr9_stage4_stallmux_q_5_), .o(n_11765) );
in01s06 g769001 ( .a(n_11763), .o(n_11764) );
in01m04 g769005 ( .a(n_11813), .o(n_11814) );
ao12s02 g769008 ( .a(n_11840), .b(n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_8_), .o(n_12105) );
oa12s06 g769009 ( .a(n_11993), .b(n_11689), .c(FE_OCP_RBN6310_n_45224), .o(n_11997) );
no02m04 TIMEBOOST_cell_1403 ( .a(n_24359), .b(FE_OCP_RBN5670_n_24288), .o(TIMEBOOST_net_316) );
oa22s01 g769012 ( .a(n_12219), .b(FE_OCP_RBN5395_cordic_combinational_sub_ln23_0_unr12_z_0_), .c(n_12218), .d(FE_OCP_RBN5392_cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n_12671) );
oa12m06 g769013 ( .a(n_11538), .b(n_11477), .c(n_11473), .o(n_11603) );
no02s01 TIMEBOOST_cell_1420 ( .a(n_13698), .b(TIMEBOOST_net_324), .o(n_13798) );
na02s04 g769015 ( .a(n_11604), .b(n_11498), .o(n_11661) );
in01s01 g769016 ( .a(n_11761), .o(n_11842) );
ao12m04 g769018 ( .a(n_11420), .b(n_11454), .c(n_11434), .o(n_11535) );
in01s01 g769019 ( .a(n_11698), .o(n_11654) );
no02s02 TIMEBOOST_cell_7030 ( .a(TIMEBOOST_net_2273), .b(n_3714), .o(n_3899) );
no04f02 TIMEBOOST_cell_8339 ( .a(n_9686), .b(n_9615), .c(n_9639), .d(n_9616), .o(n_10029) );
in01s01 g769022 ( .a(n_11760), .o(n_11845) );
no02s03 g769027 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_9_), .b(n_45697), .o(n_11860) );
no02s10 g769028 ( .a(n_11633), .b(n_11738), .o(n_11758) );
no02s10 g769029 ( .a(n_11728), .b(n_11727), .o(n_11852) );
no02s01 g769030 ( .a(FE_OCP_RBN2394_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_29_), .o(n_12278) );
in01s08 g769031 ( .a(n_11786), .o(n_11704) );
in01s02 g769033 ( .a(n_11975), .o(n_11899) );
no02m03 g769034 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_11_), .b(FE_OCPN1606_n_45697), .o(n_11975) );
no02s03 g769035 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_8_), .b(n_45697), .o(n_11840) );
no02s40 g769036 ( .a(FE_OCP_RBN6315_n_45224), .b(delay_xor_ln22_unr9_stage4_stallmux_q_4_), .o(n_11918) );
no02s10 g769037 ( .a(FE_OCP_RBN6523_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_7_), .o(n_11780) );
no02s01 TIMEBOOST_cell_5013 ( .a(TIMEBOOST_net_1454), .b(n_29046), .o(n_29130) );
no02s03 g769040 ( .a(n_45697), .b(delay_xor_ln22_unr9_stage4_stallmux_q_7_), .o(n_11694) );
no02s10 g769042 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_9_), .b(n_45697), .o(n_11885) );
no02m06 g769043 ( .a(n_45697), .b(delay_xor_ln21_unr9_stage4_stallmux_q_6_), .o(n_11643) );
in01s03 g769044 ( .a(n_11693), .o(n_11955) );
no02m06 g769045 ( .a(FE_OCP_RBN6311_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_5_), .o(n_11693) );
no02s20 g769046 ( .a(FE_OCP_RBN6308_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_2_), .o(n_11844) );
in01s02 g769047 ( .a(n_11762), .o(n_11730) );
na02s20 g769048 ( .a(n_45224), .b(FE_OCP_RBN6444_delay_xor_ln21_unr9_stage4_stallmux_q_1_), .o(n_11762) );
no02s20 g769053 ( .a(FE_OCP_RBN6307_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_3_), .o(n_11882) );
no02s10 g769054 ( .a(FE_OCP_RBN6312_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_4_), .o(n_11737) );
in01s01 g769055 ( .a(n_11756), .o(n_11757) );
no02s06 g769056 ( .a(n_45697), .b(delay_xor_ln21_unr9_stage4_stallmux_q_8_), .o(n_11756) );
no02s40 g769060 ( .a(FE_OCP_RBN6316_n_45224), .b(delay_xor_ln22_unr9_stage4_stallmux_q_3_), .o(n_11919) );
na02s03 g769061 ( .a(FE_OCP_RBN6314_n_45224), .b(n_11689), .o(n_11993) );
in01s02 g769063 ( .a(n_11769), .o(n_11718) );
na02s06 g769064 ( .a(n_45224), .b(n_11659), .o(n_11769) );
in01s01 g769066 ( .a(n_11656), .o(n_11716) );
na02s06 g769067 ( .a(n_11552), .b(n_11580), .o(n_11656) );
no02m04 g769068 ( .a(n_11497), .b(FE_OCP_RBN3243_n_10676), .o(n_11530) );
no02s01 TIMEBOOST_cell_1419 ( .a(n_13700), .b(n_13271), .o(TIMEBOOST_net_324) );
ao12s02 g769071 ( .a(n_11972), .b(n_12016), .c(n_11794), .o(n_12051) );
in01s01 g769072 ( .a(n_11775), .o(n_11665) );
no02f10 g769073 ( .a(n_11537), .b(n_11640), .o(n_11775) );
no02s10 g769074 ( .a(n_11602), .b(n_11686), .o(n_11687) );
na02s02 g769075 ( .a(n_12157), .b(n_12081), .o(n_12279) );
no03s20 TIMEBOOST_cell_3440 ( .a(n_32595), .b(n_32522), .c(n_32599), .o(n_32596) );
no02s01 TIMEBOOST_cell_6987 ( .a(n_14439), .b(n_15142), .o(TIMEBOOST_net_2252) );
na02s01 TIMEBOOST_cell_1379 ( .a(n_33498), .b(n_33513), .o(TIMEBOOST_net_304) );
na02s01 g769080 ( .a(n_11715), .b(n_11459), .o(n_11754) );
na02m04 g769081 ( .a(n_11568), .b(n_11357), .o(n_11569) );
na02s02 g769083 ( .a(n_11753), .b(n_11675), .o(n_11810) );
in01s01 g769084 ( .a(n_11700), .o(n_11701) );
no02s01 g769085 ( .a(n_11497), .b(n_11517), .o(n_11700) );
in01s01 g769086 ( .a(n_11808), .o(n_11809) );
na02s01 g769087 ( .a(n_11580), .b(n_11752), .o(n_11808) );
no03s02 TIMEBOOST_cell_7740 ( .a(n_9335), .b(n_9268), .c(n_9389), .o(TIMEBOOST_net_2501) );
na02m04 g769089 ( .a(n_11568), .b(n_11358), .o(n_11599) );
na02s02 g769090 ( .a(FE_OCP_RBN3407_n_11560), .b(n_11532), .o(n_11685) );
na02s01 g769091 ( .a(n_11509), .b(n_11485), .o(n_11555) );
in01s02 g769092 ( .a(n_11638), .o(n_11639) );
na02s06 g769093 ( .a(n_11518), .b(n_11598), .o(n_11638) );
no02s01 TIMEBOOST_cell_7029 ( .a(n_3705), .b(n_3323), .o(TIMEBOOST_net_2273) );
na02s02 g769096 ( .a(n_11658), .b(n_11657), .o(n_11713) );
no02m04 g769097 ( .a(n_11482), .b(n_11313), .o(n_11484) );
in01s01 g769098 ( .a(n_11596), .o(n_11597) );
na02s04 g769099 ( .a(n_11510), .b(n_11516), .o(n_11596) );
oa12s06 g769100 ( .a(FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n_11611), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_12_), .o(n_11751) );
oa12s02 g769102 ( .a(n_45685), .b(n_12014), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_24_), .o(n_12085) );
oa12s02 g769103 ( .a(FE_OCPN1606_n_45697), .b(n_11889), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_26_), .o(n_12013) );
oa12s02 g769104 ( .a(n_45685), .b(n_12076), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_28_), .o(n_12168) );
in01s01 g769105 ( .a(n_11806), .o(n_11807) );
na02s02 g769106 ( .a(n_11673), .b(n_11649), .o(n_11806) );
in01s01 g769109 ( .a(n_11749), .o(n_11750) );
in01s02 g769111 ( .a(n_11856), .o(n_11805) );
no02s01 TIMEBOOST_cell_1406 ( .a(TIMEBOOST_net_317), .b(n_13636), .o(n_13696) );
in01s01 g769113 ( .a(n_11803), .o(n_11804) );
na02s01 g769114 ( .a(n_11626), .b(n_11671), .o(n_11803) );
in01s01 g769115 ( .a(n_11801), .o(n_11802) );
no02s02 g769116 ( .a(n_47279), .b(n_11622), .o(n_11801) );
oa12s02 g769117 ( .a(FE_OCP_RBN3383_n_11405), .b(n_11582), .c(n_11581), .o(n_11652) );
na02s01 TIMEBOOST_cell_1408 ( .a(n_13638), .b(TIMEBOOST_net_318), .o(n_13675) );
in01s01 g769119 ( .a(n_11747), .o(n_11748) );
no02s01 g769120 ( .a(n_11623), .b(n_11608), .o(n_11747) );
in01s01 g769121 ( .a(n_11745), .o(n_11746) );
no03s40 TIMEBOOST_cell_4589 ( .a(n_27970), .b(n_27937), .c(n_27936), .o(n_28037) );
in01s02 g769123 ( .a(n_11731), .o(n_11682) );
na03f02 TIMEBOOST_cell_8244 ( .a(FE_RN_854_0), .b(FE_RN_855_0), .c(FE_RN_856_0), .o(FE_RN_857_0) );
ao12s01 g769125 ( .a(n_11372), .b(n_11480), .c(n_11479), .o(n_11523) );
na02s02 g769126 ( .a(n_11481), .b(n_11392), .o(n_11553) );
in01s01 g769127 ( .a(n_11743), .o(n_11744) );
na03m10 TIMEBOOST_cell_8377 ( .a(n_25855), .b(FE_RN_93_0), .c(FE_RN_94_0), .o(n_46962) );
in01s01 g769129 ( .a(n_11741), .o(n_11742) );
no02f06 TIMEBOOST_cell_1394 ( .a(TIMEBOOST_net_311), .b(FE_RN_2041_0), .o(n_14503) );
in01s01 g769131 ( .a(n_11799), .o(n_11800) );
na02s02 g769132 ( .a(n_11678), .b(n_11624), .o(n_11799) );
in01s01 g769133 ( .a(n_11739), .o(n_11740) );
no04s02 TIMEBOOST_cell_4591 ( .a(FE_RN_2539_0), .b(FE_RN_2541_0), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_16_), .d(FE_RN_2537_0), .o(FE_RN_2542_0) );
in01s01 g769135 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_21_), .o(n_11663) );
in01s40 g769145 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_2_), .o(n_11696) );
in01s06 g769147 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_5_), .o(n_11659) );
in01s01 g769150 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_19_), .o(n_11492) );
in01s03 g769155 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_6_), .o(n_11595) );
in01s06 g769162 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_0_), .o(n_11593) );
in01m01 g769169 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_6_), .o(n_11689) );
na02s01 g769173 ( .a(n_11971), .b(n_11893), .o(n_12170) );
no02m10 g769175 ( .a(n_11606), .b(n_11549), .o(n_11637) );
na02m20 g769176 ( .a(n_11547), .b(n_11590), .o(n_11636) );
na02s10 g769177 ( .a(n_11546), .b(n_11634), .o(n_11635) );
na02s10 g769178 ( .a(n_11601), .b(n_11544), .o(n_11602) );
na02m03 g769179 ( .a(n_11797), .b(n_11710), .o(n_12071) );
na02s10 g769180 ( .a(n_11571), .b(n_11570), .o(n_11728) );
no02s02 g769182 ( .a(n_12083), .b(n_12082), .o(n_12157) );
no02s02 g769183 ( .a(n_12080), .b(n_12079), .o(n_12081) );
no02s02 g769185 ( .a(n_12077), .b(n_12078), .o(n_12119) );
na02s01 g769186 ( .a(n_11976), .b(n_11897), .o(n_11898) );
no02s01 g769187 ( .a(n_11686), .b(n_11630), .o(n_11648) );
no02s01 g769188 ( .a(n_11838), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_18_), .o(n_11866) );
no02s01 g769189 ( .a(n_12083), .b(n_12014), .o(n_12610) );
ao12f08 g769190 ( .a(FE_OCP_RBN5393_cordic_combinational_sub_ln23_0_unr12_z_0_), .b(FE_OCP_RBN5438_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .c(n_45224), .o(n_11537) );
no02s01 g769191 ( .a(n_11974), .b(n_11973), .o(n_12567) );
na02s01 g769192 ( .a(n_12016), .b(n_12050), .o(n_12544) );
in01s01 g769193 ( .a(n_12218), .o(n_12219) );
ao12s01 g769194 ( .a(n_11640), .b(FE_OCP_RBN5439_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .c(FE_OCP_RBN2398_n_45697), .o(n_12218) );
no02s01 g769195 ( .a(n_12077), .b(n_12076), .o(n_12678) );
na02s01 g769196 ( .a(n_12084), .b(n_12047), .o(n_12702) );
in01s06 g769197 ( .a(n_11632), .o(n_11633) );
no02s01 g769199 ( .a(n_11896), .b(n_11895), .o(n_12513) );
in01s01 g769200 ( .a(n_12165), .o(n_12166) );
na02s01 g769201 ( .a(n_12115), .b(n_12008), .o(n_12165) );
na02s01 g769202 ( .a(n_11897), .b(n_11960), .o(n_12470) );
in01s01 g769203 ( .a(n_12048), .o(n_12049) );
no02s01 g769204 ( .a(n_12003), .b(n_11936), .o(n_12048) );
na02s01 g769205 ( .a(n_11798), .b(n_11797), .o(n_12153) );
no02s01 g769206 ( .a(n_11796), .b(n_11795), .o(n_12264) );
na02s01 g769207 ( .a(n_11601), .b(n_11634), .o(n_12029) );
no02s01 g769208 ( .a(n_11631), .b(n_11630), .o(n_12033) );
in01s01 g769209 ( .a(n_11680), .o(n_11681) );
no02s01 g769210 ( .a(n_11607), .b(n_11606), .o(n_11680) );
na02s01 g769211 ( .a(n_11548), .b(n_11590), .o(n_11834) );
no02s01 g769212 ( .a(n_12011), .b(n_11934), .o(n_12087) );
no02s01 g769213 ( .a(n_11738), .b(n_11727), .o(n_12139) );
in01s02 g769214 ( .a(n_11520), .o(n_11518) );
in01s01 g769216 ( .a(n_11451), .o(n_11520) );
na02s02 g769217 ( .a(n_11439), .b(FE_OCP_RBN3229_n_10644), .o(n_11451) );
no02s02 TIMEBOOST_cell_7050 ( .a(TIMEBOOST_net_2283), .b(n_10618), .o(TIMEBOOST_net_1145) );
no02s02 TIMEBOOST_cell_1367 ( .a(n_37794), .b(n_37838), .o(TIMEBOOST_net_298) );
no02s01 g769222 ( .a(FE_OCP_RBN3386_n_11439), .b(n_45300), .o(n_11589) );
no02s02 g769223 ( .a(n_11486), .b(FE_OCP_RBN3243_n_10676), .o(n_11608) );
in01s01 g769224 ( .a(n_11587), .o(n_11588) );
na02s02 g769225 ( .a(n_11474), .b(n_11538), .o(n_11587) );
no02s04 TIMEBOOST_cell_1393 ( .a(n_13418), .b(n_14466), .o(TIMEBOOST_net_311) );
na02s02 g769227 ( .a(FE_OCP_RBN6882_n_11486), .b(n_10543), .o(n_11678) );
na02s06 g769228 ( .a(FE_OCP_RBN6209_n_11486), .b(n_10935), .o(n_11552) );
na02s01 g769229 ( .a(FE_OCP_RBN6209_n_11486), .b(n_10935), .o(n_11626) );
in01s01 g769230 ( .a(n_11715), .o(n_11677) );
na02s06 g769231 ( .a(FE_OCP_RBN4483_n_11439), .b(FE_OCPN6933_FE_OCP_RBN6087_n_10852), .o(n_11715) );
in01s01 g769232 ( .a(n_11675), .o(n_11676) );
na02s02 g769233 ( .a(FE_OCP_RBN3398_n_11486), .b(FE_OCPN4859_n_10369), .o(n_11675) );
na02s06 g769234 ( .a(FE_OCP_RBN6882_n_11486), .b(FE_OCP_RBN3147_n_10369), .o(n_11753) );
in01s01 g769235 ( .a(n_12493), .o(n_12494) );
ao12s01 g769236 ( .a(n_11970), .b(FE_OCP_RBN2394_n_45697), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_22_), .o(n_12493) );
in01s01 g769237 ( .a(n_12429), .o(n_12430) );
ao12s01 g769238 ( .a(n_12082), .b(FE_OCP_RBN2394_n_45697), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_24_), .o(n_12429) );
na03f06 TIMEBOOST_cell_8346 ( .a(n_25976), .b(n_25937), .c(n_23317), .o(n_26087) );
ao12s01 g769240 ( .a(n_11863), .b(n_11707), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_18_), .o(n_12485) );
oa12s01 g769241 ( .a(n_11570), .b(n_11707), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_9_), .o(n_12198) );
ao12s01 g769242 ( .a(n_11709), .b(n_11707), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_12_), .o(n_12241) );
in01s01 g769243 ( .a(n_11658), .o(n_11647) );
na02s02 g769244 ( .a(FE_OCP_RBN4482_n_11439), .b(n_11435), .o(n_11658) );
no02s01 TIMEBOOST_cell_1405 ( .a(n_13255), .b(n_13346), .o(TIMEBOOST_net_317) );
na02s01 g769246 ( .a(FE_OCP_RBN3398_n_11486), .b(n_10480), .o(n_11624) );
in01s01 g769248 ( .a(n_11497), .o(n_11532) );
no02m02 g769249 ( .a(n_11475), .b(FE_OCP_RBN3214_n_10568), .o(n_11497) );
in01s01 g769250 ( .a(n_11516), .o(n_11517) );
na02s02 g769251 ( .a(n_11475), .b(FE_OCP_RBN3214_n_10568), .o(n_11516) );
no02s01 g769252 ( .a(n_10676), .b(FE_OCP_RBN3398_n_11486), .o(n_11623) );
na02s02 g769253 ( .a(FE_OCP_RBN6883_n_11486), .b(n_11031), .o(n_11673) );
na02s01 g769254 ( .a(FE_OCP_RBN6209_n_11486), .b(FE_OCP_RBN6117_n_11004), .o(n_11649) );
ao12s01 g769255 ( .a(n_12080), .b(FE_OCP_RBN2394_n_45697), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_26_), .o(n_12740) );
na02s01 g769256 ( .a(FE_OCP_RBN3386_n_11439), .b(n_10962), .o(n_11586) );
no02s01 g769257 ( .a(FE_OCP_RBN6209_n_11486), .b(n_10915), .o(n_11622) );
na02s01 g769258 ( .a(n_11480), .b(n_11479), .o(n_11481) );
no02s06 TIMEBOOST_cell_5484 ( .a(n_35256), .b(FE_OCP_RBN5944_n_35207), .o(TIMEBOOST_net_1690) );
na02s01 g769261 ( .a(FE_OCP_RBN3384_n_11439), .b(n_11012), .o(n_11485) );
na02s04 TIMEBOOST_cell_8618 ( .a(n_10856), .b(n_10456), .o(TIMEBOOST_net_2796) );
na02s01 g769263 ( .a(FE_OCP_RBN6882_n_11486), .b(n_10910), .o(n_11671) );
na03s04 TIMEBOOST_cell_4590 ( .a(n_1608), .b(n_1633), .c(n_1662), .o(n_1671) );
in01s01 g769265 ( .a(n_11500), .o(n_11501) );
na02s01 g769266 ( .a(n_11454), .b(n_11407), .o(n_11500) );
in01s01 g769267 ( .a(n_11752), .o(n_11712) );
na02s03 g769268 ( .a(FE_OCP_RBN6883_n_11486), .b(n_10802), .o(n_11752) );
in01s01 g769270 ( .a(n_11458), .o(n_11657) );
no02s04 g769271 ( .a(n_11439), .b(n_11435), .o(n_11458) );
in01s01 g769274 ( .a(n_11459), .o(n_11514) );
na02s03 g769275 ( .a(n_11439), .b(FE_OCP_RBN3265_n_10852), .o(n_11459) );
no02s01 g769276 ( .a(FE_OCP_RBN4483_n_11439), .b(FE_OCP_RBN4385_n_10570), .o(n_11620) );
no02s06 TIMEBOOST_cell_7543 ( .a(TIMEBOOST_net_2402), .b(FE_OCP_RBN6634_n_9304), .o(n_8229) );
na02s01 TIMEBOOST_cell_1407 ( .a(n_13077), .b(n_13621), .o(TIMEBOOST_net_318) );
in01s01 g769281 ( .a(n_11580), .o(n_11617) );
na02s04 g769282 ( .a(FE_OCP_RBN6208_n_11486), .b(n_10797), .o(n_11580) );
ao12s01 g769283 ( .a(n_12078), .b(FE_OCP_RBN2394_n_45697), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_28_), .o(n_12710) );
na02s01 g769284 ( .a(FE_OCP_RBN3386_n_11439), .b(FE_OCPN1217_n_11012), .o(n_11557) );
na02s01 g769285 ( .a(FE_OCP_RBN3386_n_11439), .b(n_11112), .o(n_11579) );
in01s01 g769287 ( .a(n_11478), .o(n_11598) );
no02s04 g769288 ( .a(n_11439), .b(FE_OCP_RBN3229_n_10644), .o(n_11478) );
na02m04 g769289 ( .a(n_11456), .b(n_11398), .o(n_11511) );
ao12m04 g769290 ( .a(n_11337), .b(n_11410), .c(n_11392), .o(n_11434) );
no02s06 g769293 ( .a(FE_OCP_RBN3398_n_11486), .b(FE_OCPN4551_n_10545), .o(n_11560) );
in01s01 g769295 ( .a(n_11578), .o(n_11613) );
no02s06 g769296 ( .a(FE_OCP_RBN6207_n_11486), .b(n_10936), .o(n_11578) );
na02m06 g769299 ( .a(n_11407), .b(n_11379), .o(n_11482) );
na02s02 TIMEBOOST_cell_8164 ( .a(n_44454), .b(n_11078), .o(TIMEBOOST_net_2713) );
oa12m04 g769301 ( .a(n_11425), .b(n_11476), .c(n_11405), .o(n_11477) );
in01s01 g769302 ( .a(n_11510), .o(n_11915) );
na02s02 g769303 ( .a(n_11475), .b(n_10544), .o(n_11510) );
in01m02 g769304 ( .a(n_11669), .o(n_11759) );
ao22m04 g769305 ( .a(n_11504), .b(n_11427), .c(n_11503), .d(n_11426), .o(n_11669) );
in01s01 g769306 ( .a(n_11509), .o(n_11924) );
na02s01 g769307 ( .a(FE_OCP_RBN3384_n_11439), .b(n_10977), .o(n_11509) );
oa22s01 g769309 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_), .c(n_10812), .d(FE_OCP_RBN5445_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_12442) );
oa22s01 g769310 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_), .c(n_10387), .d(FE_OCP_RBN5445_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_12201) );
ao22s01 g769311 ( .a(n_12164), .b(FE_OCP_RBN5445_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .c(n_11707), .d(delay_sub_ln23_0_unr8_stage4_stallmux_q_14_), .o(n_12356) );
oa22s01 g769312 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_4_), .c(n_11542), .d(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_12094) );
in01s01 g769313 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_20_), .o(n_12693) );
in01s01 g769315 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_19_), .o(n_11528) );
in01s01 g769317 ( .a(n_11972), .o(n_12050) );
no02s01 g769318 ( .a(FE_OCPN1606_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_20_), .o(n_11972) );
na02s01 g769319 ( .a(FE_OCPN1606_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_20_), .o(n_12016) );
in01s01 g769320 ( .a(n_11794), .o(n_11895) );
na02s01 g769321 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_19_), .o(n_11794) );
in01s01 g769322 ( .a(n_11894), .o(n_11973) );
na02s01 g769323 ( .a(FE_OCPN1606_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_21_), .o(n_11894) );
in01s01 g769324 ( .a(n_11970), .o(n_11971) );
no02s01 g769325 ( .a(FE_OCPN1606_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_22_), .o(n_11970) );
in01s01 g769326 ( .a(n_11974), .o(n_11893) );
no02s01 g769327 ( .a(FE_OCPN1606_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_21_), .o(n_11974) );
no02s01 g769329 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_18_), .o(n_11863) );
na02s01 g769330 ( .a(FE_OCP_RBN5445_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n_11784), .o(n_11960) );
no02s02 g769331 ( .a(FE_OCP_RBN5445_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n_10708), .o(n_11795) );
in01s06 g769332 ( .a(n_11548), .o(n_11549) );
na02m10 g769333 ( .a(FE_OCP_RBN6442_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_2_), .o(n_11548) );
in01m08 g769334 ( .a(n_11525), .o(n_11606) );
na02s10 g769335 ( .a(FE_OCP_RBN6442_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_1_), .o(n_11525) );
no02m06 g769336 ( .a(n_45224), .b(FE_OCP_RBN5439_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .o(n_11640) );
na02s20 g769337 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(FE_OCP_RBN5441_delay_sub_ln23_0_unr8_stage4_stallmux_q_2_), .o(n_11590) );
in01m10 g769338 ( .a(n_11607), .o(n_11547) );
no02s20 g769339 ( .a(FE_OCP_RBN6442_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_1_), .o(n_11607) );
in01s03 g769340 ( .a(n_11631), .o(n_11546) );
no02s06 g769341 ( .a(FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_5_), .o(n_11631) );
na02s06 g769342 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n_10035), .o(n_11634) );
in01s01 g769343 ( .a(n_11544), .o(n_11630) );
na02s10 g769344 ( .a(FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_5_), .o(n_11544) );
na02s10 g769345 ( .a(FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_6_), .o(n_11601) );
no02s06 g769346 ( .a(FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_10_), .o(n_11738) );
no02s10 g769347 ( .a(FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_), .o(n_12003) );
in01m01 g769348 ( .a(n_11711), .o(n_11797) );
no02s03 g769349 ( .a(FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_11_), .o(n_11711) );
in01m01 g769350 ( .a(n_11709), .o(n_11710) );
no02s03 g769351 ( .a(FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_12_), .o(n_11709) );
no02s03 g769352 ( .a(FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_13_), .o(n_11796) );
in01s06 g769353 ( .a(n_11798), .o(n_11611) );
na02s03 g769354 ( .a(FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_11_), .o(n_11798) );
no02s03 g769355 ( .a(FE_OCP_RBN5445_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n_10419), .o(n_11727) );
na02s06 g769356 ( .a(n_11507), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_9_), .o(n_11570) );
in01s01 g769357 ( .a(n_11838), .o(n_11897) );
no02s01 g769358 ( .a(FE_OCP_RBN5445_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n_11784), .o(n_11838) );
no02s01 g769360 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_19_), .o(n_11896) );
in01s02 g769361 ( .a(n_11892), .o(n_12014) );
na02s02 g769362 ( .a(FE_OCPN1606_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_23_), .o(n_11892) );
in01s01 g769363 ( .a(n_12084), .o(n_11889) );
na02s02 g769364 ( .a(FE_OCPN1606_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_25_), .o(n_12084) );
in01s01 g769365 ( .a(n_11968), .o(n_12076) );
na02s02 g769366 ( .a(FE_OCPN1606_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_27_), .o(n_11968) );
no02s02 g769367 ( .a(FE_OCPN1606_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_23_), .o(n_12083) );
no02s01 g769368 ( .a(FE_OCPN1606_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_24_), .o(n_12082) );
no02s02 g769369 ( .a(n_45685), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_26_), .o(n_12080) );
in01s01 g769370 ( .a(n_12079), .o(n_12047) );
no02s02 g769371 ( .a(n_45685), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_25_), .o(n_12079) );
in01s01 g769372 ( .a(n_12077), .o(n_12046) );
no02s02 g769373 ( .a(FE_OCP_RBN2394_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_27_), .o(n_12077) );
no02s01 g769374 ( .a(FE_OCP_RBN2394_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_28_), .o(n_12078) );
na02s01 g769375 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_), .o(n_12115) );
in01s01 g769376 ( .a(n_12007), .o(n_12008) );
no02s01 g769377 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_), .o(n_12007) );
in01s01 g769378 ( .a(n_11935), .o(n_11936) );
na02s01 g769379 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_), .o(n_11935) );
in01s01 g769380 ( .a(n_11933), .o(n_11934) );
na02s01 g769381 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_), .o(n_11933) );
no02s01 g769382 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_), .o(n_12011) );
na02s04 g769383 ( .a(n_11378), .b(n_10451), .o(n_11454) );
oa12s06 g769385 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n_11542), .c(n_9777), .o(n_11543) );
no02s06 TIMEBOOST_cell_4894 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_5_), .b(FE_OCP_RBN6517_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(TIMEBOOST_net_1395) );
na02s06 TIMEBOOST_cell_3843 ( .a(n_32699), .b(FE_RN_2200_0), .o(TIMEBOOST_net_1012) );
in01s01 g769389 ( .a(n_11407), .o(n_11420) );
na02m06 g769390 ( .a(n_11377), .b(FE_OCP_RBN3161_n_10399), .o(n_11407) );
oa12s01 g769391 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_), .o(n_11976) );
ao12s01 g769392 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_), .o(n_11890) );
in01s01 g769393 ( .a(n_11473), .o(n_11474) );
no02s06 g769394 ( .a(FE_OCP_RBN6188_n_11403), .b(n_10293), .o(n_11473) );
no02s06 TIMEBOOST_cell_4873 ( .a(n_32525), .b(TIMEBOOST_net_1384), .o(FE_RN_445_0) );
na02s06 g769396 ( .a(FE_OCP_RBN6189_n_11403), .b(n_10293), .o(n_11538) );
oa22s02 g769397 ( .a(n_11384), .b(n_10383), .c(n_11385), .d(n_10384), .o(n_11433) );
in01s02 g769416 ( .a(n_11453), .o(n_11422) );
na02s01 TIMEBOOST_cell_1374 ( .a(TIMEBOOST_net_301), .b(n_19404), .o(n_19524) );
in01s01 g769419 ( .a(n_11582), .o(n_11575) );
na02s04 g769420 ( .a(n_11430), .b(n_11476), .o(n_11582) );
no02m10 g769431 ( .a(n_11355), .b(n_11336), .o(n_11439) );
in01s08 g769444 ( .a(n_11475), .o(n_11486) );
in01m02 g769446 ( .a(n_11527), .o(n_11655) );
ao22m04 g769447 ( .a(n_11413), .b(n_11388), .c(n_11414), .d(n_11389), .o(n_11527) );
in01s02 g769452 ( .a(n_11480), .o(n_11456) );
na02s02 TIMEBOOST_cell_2828 ( .a(FE_RN_2542_0), .b(FE_RN_2536_0), .o(TIMEBOOST_net_705) );
in01m02 g769478 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11707) );
in01s20 g769486 ( .a(FE_OCP_RBN5445_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11507) );
in01s01 g769488 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_20_), .o(n_11524) );
no02m08 g769557 ( .a(n_11328), .b(n_11280), .o(n_11355) );
na02s01 TIMEBOOST_cell_1373 ( .a(n_19402), .b(n_18808), .o(TIMEBOOST_net_301) );
no02m08 TIMEBOOST_cell_8535 ( .a(TIMEBOOST_net_2754), .b(TIMEBOOST_net_1888), .o(n_24748) );
in01s04 g769560 ( .a(n_11503), .o(n_11504) );
na02m08 g769561 ( .a(n_11416), .b(n_11374), .o(n_11503) );
na02s02 g769562 ( .a(n_11415), .b(n_11419), .o(n_11430) );
in01s01 g769563 ( .a(n_11464), .o(n_11465) );
na02s02 g769564 ( .a(n_11425), .b(FE_OCP_RBN3383_n_11405), .o(n_11464) );
in01s02 g769565 ( .a(n_11398), .o(n_11399) );
na02s03 g769566 ( .a(n_11392), .b(n_11479), .o(n_11398) );
no02s06 g769567 ( .a(n_11327), .b(FE_OCP_RBN3358_n_11275), .o(n_11336) );
na02m06 g769568 ( .a(FE_OCP_RBN3382_n_11405), .b(n_11395), .o(n_11429) );
in01m02 g769572 ( .a(n_11495), .o(n_11605) );
ao22f02 g769573 ( .a(n_11383), .b(n_11360), .c(n_11400), .d(n_11359), .o(n_11495) );
na02m06 g769574 ( .a(n_11376), .b(n_47185), .o(n_11476) );
no02m04 g769575 ( .a(n_11335), .b(n_11353), .o(n_11379) );
no02m06 g769576 ( .a(n_11352), .b(n_11386), .o(n_11410) );
in01s02 g769577 ( .a(n_11377), .o(n_11378) );
in01s02 g769579 ( .a(n_11494), .o(n_11463) );
no02f04 TIMEBOOST_cell_1498 ( .a(TIMEBOOST_net_363), .b(n_30105), .o(n_30168) );
no02s04 g769585 ( .a(n_47182), .b(n_11394), .o(n_11395) );
no02m08 g769589 ( .a(n_11381), .b(n_11380), .o(n_11405) );
no02s02 TIMEBOOST_cell_1497 ( .a(n_30104), .b(n_29818), .o(TIMEBOOST_net_363) );
na02m04 g769591 ( .a(n_11375), .b(n_11374), .o(n_11376) );
in01s01 g769592 ( .a(n_11425), .o(n_11581) );
na02s02 g769593 ( .a(n_11381), .b(n_11380), .o(n_11425) );
in01s02 g769594 ( .a(n_11388), .o(n_11389) );
no02m02 g769595 ( .a(n_11386), .b(n_11351), .o(n_11388) );
in01s02 g769596 ( .a(n_11337), .o(n_11479) );
no02s04 g769597 ( .a(n_11320), .b(FE_OCP_RBN3137_n_10326), .o(n_11337) );
in01m02 g769598 ( .a(n_11318), .o(n_11335) );
in01s01 g769600 ( .a(n_11392), .o(n_11372) );
na02m02 g769601 ( .a(FE_OCP_RBN3137_n_10326), .b(n_11320), .o(n_11318) );
na02s03 g769602 ( .a(n_11320), .b(FE_OCP_RBN3137_n_10326), .o(n_11392) );
na02m02 g769603 ( .a(n_11345), .b(n_11325), .o(n_11353) );
in01s04 g769604 ( .a(n_11415), .o(n_11416) );
no02m06 g769605 ( .a(n_11383), .b(n_11394), .o(n_11415) );
in01m02 g769606 ( .a(n_11413), .o(n_11414) );
no02m06 g769607 ( .a(n_11367), .b(n_11269), .o(n_11413) );
no02m04 g769608 ( .a(n_11269), .b(n_11351), .o(n_11352) );
in01s02 g769609 ( .a(n_11426), .o(n_11427) );
na02s02 g769610 ( .a(n_11375), .b(n_11419), .o(n_11426) );
no02f04 TIMEBOOST_cell_5559 ( .a(TIMEBOOST_net_1727), .b(n_25922), .o(n_26021) );
no02m06 TIMEBOOST_cell_3977 ( .a(FE_OCP_RBN2842_n_9044), .b(FE_OFN4770_n_8309), .o(TIMEBOOST_net_1079) );
in01s01 g769615 ( .a(n_11384), .o(n_11385) );
oa12s01 g769616 ( .a(n_10250), .b(n_11333), .c(n_10341), .o(n_11384) );
in01m04 g769617 ( .a(n_11327), .o(n_11328) );
na03m04 TIMEBOOST_cell_7169 ( .a(n_29475), .b(n_29477), .c(n_29454), .o(n_29574) );
in01m04 g769619 ( .a(n_11370), .o(n_11371) );
no02f04 TIMEBOOST_cell_1358 ( .a(TIMEBOOST_net_293), .b(FE_RN_1015_0), .o(n_13703) );
oa22s01 g769621 ( .a(n_11342), .b(n_10343), .c(n_11333), .d(n_10344), .o(n_11402) );
in01s02 g769622 ( .a(n_11411), .o(n_11396) );
na02s01 TIMEBOOST_cell_1376 ( .a(n_19369), .b(TIMEBOOST_net_302), .o(n_19521) );
in01s01 g769624 ( .a(n_11349), .o(n_11350) );
oa12s02 g769625 ( .a(n_11249), .b(n_11294), .c(n_11131), .o(n_11349) );
in01s02 g769626 ( .a(n_11409), .o(n_11490) );
ao22m02 g769627 ( .a(n_11340), .b(n_11332), .c(n_11317), .d(n_11331), .o(n_11409) );
in01s01 g769628 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_17_), .o(n_12672) );
no02m04 g769630 ( .a(n_11183), .b(FE_OCP_RBN3348_n_47269), .o(n_11251) );
in01s04 g769635 ( .a(FE_OCP_RBN3358_n_11275), .o(n_11280) );
na02f04 TIMEBOOST_cell_8733 ( .a(TIMEBOOST_net_2853), .b(n_13731), .o(TIMEBOOST_net_2409) );
na02s01 TIMEBOOST_cell_1375 ( .a(n_18582), .b(n_19400), .o(TIMEBOOST_net_302) );
no02m02 g769640 ( .a(n_11301), .b(FE_OCP_RBN3116_n_10198), .o(n_11351) );
na02s02 g769641 ( .a(n_11310), .b(n_11259), .o(n_11326) );
in01s02 g769643 ( .a(n_11383), .o(n_11400) );
no02m08 g769644 ( .a(n_11358), .b(n_11357), .o(n_11383) );
in01s01 g769645 ( .a(n_47182), .o(n_11419) );
in01s04 g769648 ( .a(n_11366), .o(n_11367) );
na02m08 g769649 ( .a(n_11317), .b(n_11345), .o(n_11366) );
na02m04 g769650 ( .a(n_11308), .b(FE_OCP_RBN3095_n_10023), .o(n_11375) );
in01s04 g769651 ( .a(n_11325), .o(n_11386) );
na02m04 g769652 ( .a(n_11301), .b(FE_OCP_RBN3116_n_10198), .o(n_11325) );
in01m02 g769653 ( .a(n_11323), .o(n_11324) );
no02m06 g769654 ( .a(n_11258), .b(n_11194), .o(n_11323) );
na02m06 g769656 ( .a(n_11333), .b(n_10285), .o(n_11364) );
no02f02 TIMEBOOST_cell_1357 ( .a(FE_OCP_RBN2540_n_12880), .b(n_13536), .o(TIMEBOOST_net_293) );
no02f08 TIMEBOOST_cell_5990 ( .a(TIMEBOOST_net_1846), .b(TIMEBOOST_net_217), .o(n_23513) );
oa12s04 g769659 ( .a(FE_OCP_RBN6130_n_46424), .b(n_11247), .c(FE_OCP_RBN3347_n_47269), .o(n_11274) );
na02f08 TIMEBOOST_cell_7913 ( .a(TIMEBOOST_net_2587), .b(n_26032), .o(n_26188) );
na02m06 g769661 ( .a(n_11299), .b(n_11231), .o(n_11315) );
oa22s01 g769662 ( .a(n_11288), .b(n_10381), .c(n_11287), .d(n_10382), .o(n_11344) );
na02m06 g769663 ( .a(n_11314), .b(n_11281), .o(n_11381) );
in01f02 g769664 ( .a(n_11356), .o(n_11334) );
no02m10 TIMEBOOST_cell_5957 ( .a(n_22927), .b(n_22748), .o(TIMEBOOST_net_1830) );
in01f02 g769666 ( .a(n_46986), .o(n_11412) );
in01s01 g769668 ( .a(n_11362), .o(n_11363) );
ao12s01 g769669 ( .a(n_11104), .b(n_11316), .c(n_47199), .o(n_11362) );
na02m06 g769670 ( .a(n_11245), .b(n_11210), .o(n_11320) );
in01s01 g769671 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_16_), .o(n_12537) );
no02s04 g769675 ( .a(n_11229), .b(n_11230), .o(n_11258) );
na02m04 g769676 ( .a(n_11272), .b(n_11264), .o(n_11314) );
na02s03 g769677 ( .a(n_11271), .b(n_11263), .o(n_11281) );
na02m08 g769678 ( .a(n_11256), .b(n_44511), .o(n_11299) );
no03m03 TIMEBOOST_cell_3429 ( .a(n_12003), .b(FE_RN_1558_0), .c(FE_OCP_RBN5444_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11632) );
no02s06 g769680 ( .a(n_44855), .b(n_44516), .o(n_11205) );
no02m04 g769681 ( .a(n_44855), .b(n_44498), .o(n_11183) );
no02s02 g769682 ( .a(n_11209), .b(n_46424), .o(n_11227) );
na02s02 TIMEBOOST_cell_4913 ( .a(TIMEBOOST_net_1404), .b(n_41208), .o(n_40935) );
na03f04 TIMEBOOST_cell_8361 ( .a(FE_OCP_RBN1839_n_20273), .b(n_45065), .c(n_20297), .o(n_20417) );
no02s04 g769686 ( .a(n_11256), .b(n_44511), .o(n_11257) );
in01s01 g769688 ( .a(n_11333), .o(n_11342) );
no02m06 g769689 ( .a(n_11268), .b(n_10246), .o(n_11333) );
in01s01 g769691 ( .a(n_11317), .o(n_11340) );
na02m08 g769692 ( .a(n_11313), .b(n_11312), .o(n_11317) );
na02f04 g769693 ( .a(n_11316), .b(n_11187), .o(n_11361) );
na02m04 g769694 ( .a(n_11247), .b(n_11168), .o(n_11245) );
na03s02 TIMEBOOST_cell_4795 ( .a(n_4525), .b(n_4255), .c(n_4539), .o(n_4762) );
na02m04 g769696 ( .a(n_11243), .b(n_11157), .o(n_11295) );
in01s01 g769698 ( .a(n_11294), .o(n_11310) );
no02s06 g769699 ( .a(n_11226), .b(n_11179), .o(n_11294) );
no02m06 g769700 ( .a(n_11285), .b(n_11284), .o(n_11357) );
in01s01 g769701 ( .a(n_11331), .o(n_11332) );
na02s02 g769702 ( .a(n_11345), .b(n_11289), .o(n_11331) );
in01s02 g769703 ( .a(n_11359), .o(n_11360) );
na02s04 g769704 ( .a(n_11374), .b(n_11306), .o(n_11359) );
na02m02 g769705 ( .a(n_11209), .b(n_11167), .o(n_11210) );
in01f02 g769707 ( .a(n_11369), .o(n_11338) );
no02f06 TIMEBOOST_cell_2996 ( .a(FE_RN_2584_0), .b(FE_OCPN1709_FE_OFN739_n_17093), .o(TIMEBOOST_net_789) );
no02s06 g769709 ( .a(n_11225), .b(n_11262), .o(n_11358) );
no02f04 TIMEBOOST_cell_7816 ( .a(n_38534), .b(TIMEBOOST_net_1255), .o(TIMEBOOST_net_2539) );
in01m02 g769715 ( .a(n_11271), .o(n_11272) );
in01m04 g769716 ( .a(n_11229), .o(n_11271) );
na02m06 g769717 ( .a(n_11198), .b(n_11200), .o(n_11229) );
no02s04 g769718 ( .a(n_11201), .b(n_11230), .o(n_11231) );
na02m04 g769719 ( .a(n_11199), .b(n_11218), .o(n_11244) );
in01f02 g769720 ( .a(n_11242), .o(n_11243) );
na02f04 g769721 ( .a(n_11173), .b(n_11106), .o(n_11242) );
in01s02 g769722 ( .a(n_11225), .o(n_11226) );
na02s06 g769723 ( .a(n_11172), .b(n_11159), .o(n_11225) );
na02s06 g769724 ( .a(n_11293), .b(n_11292), .o(n_11374) );
no02s06 TIMEBOOST_cell_8523 ( .a(TIMEBOOST_net_2748), .b(n_682), .o(n_686) );
in01s02 g769726 ( .a(n_11394), .o(n_11306) );
no02s06 g769727 ( .a(n_11293), .b(n_11292), .o(n_11394) );
na02s06 g769728 ( .a(n_11254), .b(FE_OCPN4549_FE_OCP_RBN3086_n_10015), .o(n_11345) );
na02f08 TIMEBOOST_cell_2995 ( .a(n_13697), .b(TIMEBOOST_net_788), .o(n_13765) );
na02f04 g769730 ( .a(n_11239), .b(n_11043), .o(n_11291) );
na02s08 g769733 ( .a(n_11241), .b(n_11073), .o(n_11316) );
no03s03 TIMEBOOST_cell_3428 ( .a(FE_RN_118_0), .b(FE_RN_117_0), .c(n_6708), .o(n_6612) );
in01s02 g769736 ( .a(n_11269), .o(n_11289) );
no02s06 g769737 ( .a(n_11254), .b(FE_OCPN4549_FE_OCP_RBN3086_n_10015), .o(n_11269) );
in01s01 g769738 ( .a(n_11287), .o(n_11288) );
oa12s01 g769739 ( .a(n_11266), .b(n_11267), .c(n_10124), .o(n_11287) );
ao12m04 g769740 ( .a(n_10211), .b(n_11267), .c(n_11266), .o(n_11268) );
oa22s01 g769741 ( .a(n_11213), .b(n_10248), .c(n_11214), .d(n_10249), .o(n_11286) );
oa22s01 g769742 ( .a(n_11267), .b(n_10296), .c(n_11233), .d(n_10297), .o(n_11305) );
in01m04 g769743 ( .a(n_11223), .o(n_11256) );
no02s02 TIMEBOOST_cell_1274 ( .a(TIMEBOOST_net_251), .b(n_38003), .o(n_38004) );
in01s04 g769745 ( .a(n_11209), .o(n_11247) );
no02s04 TIMEBOOST_cell_5136 ( .a(n_9012), .b(n_8983), .o(TIMEBOOST_net_1516) );
in01f02 g769748 ( .a(n_11297), .o(n_11265) );
no02s01 TIMEBOOST_cell_2976 ( .a(n_18594), .b(n_18548), .o(TIMEBOOST_net_779) );
na02m06 g769750 ( .a(n_11240), .b(n_11175), .o(n_11313) );
no02f04 TIMEBOOST_cell_7680 ( .a(n_44871), .b(n_37414), .o(TIMEBOOST_net_2471) );
na02m08 g769754 ( .a(n_11196), .b(n_11228), .o(n_11312) );
in01s01 g769756 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_15_), .o(n_11298) );
in01s02 g769758 ( .a(n_11200), .o(n_11201) );
no02s06 g769759 ( .a(n_46423), .b(n_44453), .o(n_11200) );
na02m06 g769760 ( .a(n_11122), .b(n_11123), .o(n_11124) );
no02m04 TIMEBOOST_cell_5135 ( .a(TIMEBOOST_net_1515), .b(n_38627), .o(n_38676) );
no02s08 TIMEBOOST_cell_3255 ( .a(TIMEBOOST_net_918), .b(n_10702), .o(n_10797) );
no02s02 TIMEBOOST_cell_1273 ( .a(n_44867), .b(n_38269), .o(TIMEBOOST_net_251) );
no02s01 TIMEBOOST_cell_4329 ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .b(n_38778), .o(TIMEBOOST_net_1255) );
no02s04 g769767 ( .a(n_46423), .b(n_11145), .o(n_11221) );
in01m02 g769768 ( .a(n_11263), .o(n_11264) );
no02m04 g769769 ( .a(n_11193), .b(n_11194), .o(n_11263) );
no02m04 g769770 ( .a(FE_OCP_RBN3331_n_11087), .b(n_44516), .o(n_11148) );
na02m02 g769771 ( .a(n_47269), .b(FE_OCP_RBN4443_n_46424), .o(n_11168) );
no02s02 g769772 ( .a(FE_OCP_RBN3346_n_47269), .b(n_46424), .o(n_11167) );
in01s02 g769773 ( .a(n_11198), .o(n_11199) );
na02m06 g769774 ( .a(n_11144), .b(n_11134), .o(n_11198) );
no02s02 TIMEBOOST_cell_4899 ( .a(TIMEBOOST_net_1397), .b(n_6776), .o(n_6918) );
na02s02 g769776 ( .a(n_11235), .b(n_11152), .o(n_11262) );
in01s02 g769777 ( .a(n_11303), .o(n_11304) );
no02m04 g769778 ( .a(n_11284), .b(n_11283), .o(n_11303) );
in01f02 g769779 ( .a(n_11172), .o(n_11173) );
no02f08 g769780 ( .a(n_11113), .b(n_10984), .o(n_11172) );
na02f02 g769781 ( .a(n_11113), .b(n_11064), .o(n_11197) );
in01s03 g769782 ( .a(n_11240), .o(n_11241) );
no02s06 g769783 ( .a(n_11208), .b(n_11047), .o(n_11240) );
in01m02 g769784 ( .a(n_11238), .o(n_11239) );
na02m04 g769785 ( .a(n_11208), .b(n_10982), .o(n_11238) );
na02s04 TIMEBOOST_cell_2975 ( .a(TIMEBOOST_net_778), .b(n_13954), .o(n_14144) );
no02s04 g769788 ( .a(n_11166), .b(n_47200), .o(n_11175) );
in01s01 g769789 ( .a(n_11236), .o(n_11237) );
na02s02 g769790 ( .a(n_11195), .b(n_11228), .o(n_11236) );
na02m06 g769791 ( .a(n_11137), .b(n_11138), .o(n_11254) );
in01m02 g769792 ( .a(n_11252), .o(n_11220) );
na02f08 TIMEBOOST_cell_1346 ( .a(TIMEBOOST_net_287), .b(n_19381), .o(n_19528) );
na02m06 g769794 ( .a(n_11191), .b(n_11190), .o(n_11293) );
in01m02 g769795 ( .a(n_11307), .o(n_11282) );
na02s01 TIMEBOOST_cell_4175 ( .a(FE_OFN5083_n_36750), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_1178) );
in01s01 g769797 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_14_), .o(n_12468) );
in01s02 g769800 ( .a(n_11144), .o(n_11145) );
na02s06 g769801 ( .a(n_11118), .b(FE_OFN756_n_44464), .o(n_11144) );
in01m02 g769808 ( .a(n_11194), .o(n_11218) );
no02s06 g769809 ( .a(n_11132), .b(n_44511), .o(n_11194) );
na02m06 g769810 ( .a(n_11052), .b(FE_OCPN4845_FE_OFN4779_n_44490), .o(n_11123) );
no02m04 g769811 ( .a(n_11192), .b(FE_OFN4799_n_44498), .o(n_11193) );
no02s06 g769812 ( .a(n_11192), .b(FE_OFN4799_n_44498), .o(n_11230) );
na02s02 g769817 ( .a(n_11164), .b(n_44454), .o(n_11181) );
no02s04 g769818 ( .a(n_11165), .b(n_44453), .o(n_11217) );
no02s02 g769821 ( .a(n_11052), .b(FE_OCP_RBN5955_FE_OFN4772_n_44463), .o(n_11053) );
na02m06 TIMEBOOST_cell_3259 ( .a(TIMEBOOST_net_920), .b(FE_OCP_RBN6116_n_11004), .o(n_11146) );
no02s02 g769823 ( .a(n_11083), .b(FE_OCP_RBN6128_n_11026), .o(n_11114) );
na03f20 TIMEBOOST_cell_3427 ( .a(n_40653), .b(n_40654), .c(n_40641), .o(n_40660) );
no02f06 TIMEBOOST_cell_4174 ( .a(TIMEBOOST_net_1177), .b(n_36581), .o(n_36646) );
in01s04 g769826 ( .a(n_11235), .o(n_11284) );
na02s04 g769827 ( .a(n_46987), .b(FE_OCP_RBN5980_n_9682), .o(n_11235) );
na02m04 g769828 ( .a(n_11082), .b(n_10986), .o(n_11130) );
in01s01 g769830 ( .a(n_11113), .o(n_11139) );
oa12f08 g769831 ( .a(n_10953), .b(n_10971), .c(n_10941), .o(n_11113) );
na02s04 g769832 ( .a(n_11086), .b(n_11024), .o(n_11138) );
na02s04 TIMEBOOST_cell_3262 ( .a(n_11029), .b(FE_OFN4800_n_44498), .o(TIMEBOOST_net_922) );
na02m04 TIMEBOOST_cell_1345 ( .a(n_19430), .b(n_17881), .o(TIMEBOOST_net_287) );
in01s03 g769835 ( .a(n_11166), .o(n_11228) );
no02s06 g769836 ( .a(FE_OCP_RBN3064_n_9892), .b(n_11128), .o(n_11166) );
no02s03 g769837 ( .a(n_46987), .b(FE_OCP_RBN5980_n_9682), .o(n_11283) );
na02m08 g769838 ( .a(n_11129), .b(n_10983), .o(n_11208) );
na02s02 TIMEBOOST_cell_6632 ( .a(TIMEBOOST_net_2073), .b(n_18440), .o(n_18509) );
na02s04 g769840 ( .a(n_11136), .b(n_11103), .o(n_11190) );
na02f02 g769841 ( .a(n_11162), .b(n_11016), .o(n_11189) );
no02s02 g769842 ( .a(n_11178), .b(n_11131), .o(n_11215) );
na02m04 g769843 ( .a(n_11128), .b(FE_OCP_RBN3064_n_9892), .o(n_11195) );
in01s01 g769844 ( .a(n_11213), .o(n_11214) );
oa12s01 g769845 ( .a(n_10208), .b(n_11180), .c(n_10119), .o(n_11213) );
in01s01 g769847 ( .a(n_11267), .o(n_11233) );
oa12m06 g769848 ( .a(n_10161), .b(n_11180), .c(n_10160), .o(n_11267) );
no02s02 TIMEBOOST_cell_3839 ( .a(n_27959), .b(n_27991), .o(TIMEBOOST_net_1010) );
in01m02 g769850 ( .a(n_11278), .o(n_11232) );
no02s06 TIMEBOOST_cell_1468 ( .a(TIMEBOOST_net_348), .b(n_7713), .o(n_7756) );
in01s01 g769852 ( .a(FE_OCP_RBN6117_n_11004), .o(n_11031) );
in01s01 g769856 ( .a(FE_OCP_RBN3330_n_11087), .o(n_11112) );
no02f06 TIMEBOOST_cell_5064 ( .a(FE_RN_1623_0), .b(n_13599), .o(TIMEBOOST_net_1480) );
na02s01 g769862 ( .a(n_11180), .b(n_10240), .o(n_11211) );
no04m04 TIMEBOOST_cell_4637 ( .a(n_41912), .b(n_41828), .c(n_41531), .d(n_41532), .o(FE_RN_856_0) );
no02s02 g769864 ( .a(n_11048), .b(n_44453), .o(n_11136) );
no02f06 TIMEBOOST_cell_3261 ( .a(n_6266), .b(TIMEBOOST_net_921), .o(n_46195) );
no02s04 g769866 ( .a(FE_OCP_RBN6127_n_11026), .b(n_11027), .o(n_11086) );
in01s02 g769867 ( .a(n_11164), .o(n_11165) );
in01s02 g769868 ( .a(n_11134), .o(n_11164) );
no02m06 g769869 ( .a(n_11074), .b(n_11048), .o(n_11134) );
in01s02 g769870 ( .a(n_11083), .o(n_11084) );
in01s04 g769871 ( .a(n_11056), .o(n_11083) );
na02m08 g769872 ( .a(n_10998), .b(n_11000), .o(n_11056) );
na02s02 g769873 ( .a(n_11072), .b(n_11035), .o(n_11110) );
in01f01 g769875 ( .a(n_11129), .o(n_11162) );
ao12f06 g769876 ( .a(n_10903), .b(n_11032), .c(n_10872), .o(n_11129) );
no02s01 TIMEBOOST_cell_1467 ( .a(n_7634), .b(n_7683), .o(TIMEBOOST_net_348) );
na02m04 g769878 ( .a(n_11097), .b(n_10920), .o(n_11161) );
na02m04 g769880 ( .a(n_47199), .b(n_11076), .o(n_11187) );
in01s02 g769881 ( .a(n_11259), .o(n_11260) );
na02s04 g769882 ( .a(n_11249), .b(n_11152), .o(n_11259) );
oa22s01 g769883 ( .a(n_11069), .b(n_10206), .c(n_11070), .d(n_10207), .o(n_11153) );
in01s02 g769884 ( .a(n_11177), .o(n_11151) );
na02s01 TIMEBOOST_cell_4053 ( .a(n_24429), .b(FE_OCP_RBN5926_n_25211), .o(TIMEBOOST_net_1117) );
na03s03 TIMEBOOST_cell_8380 ( .a(n_20536), .b(n_20456), .c(n_20533), .o(n_20634) );
in01s02 g769887 ( .a(n_11081), .o(n_11082) );
oa12m04 g769888 ( .a(n_10979), .b(n_11003), .c(n_10923), .o(n_11081) );
in01s01 g769889 ( .a(n_11178), .o(n_11179) );
na03s08 TIMEBOOST_cell_3478 ( .a(n_6596), .b(n_6890), .c(n_6845), .o(n_6990) );
in01m04 g769891 ( .a(n_11132), .o(n_11192) );
na03s06 TIMEBOOST_cell_8407 ( .a(FE_OCP_RBN4354_n_4585), .b(FE_OCP_RBN4342_n_4198), .c(n_4641), .o(n_4809) );
in01s02 g769894 ( .a(n_11052), .o(n_11029) );
no02s02 TIMEBOOST_cell_4463 ( .a(n_21730), .b(n_21539), .o(TIMEBOOST_net_1322) );
no02f06 TIMEBOOST_cell_1316 ( .a(TIMEBOOST_net_272), .b(n_12800), .o(n_12879) );
no02s02 TIMEBOOST_cell_3376 ( .a(n_31518), .b(n_31599), .o(TIMEBOOST_net_979) );
no02s03 g769900 ( .a(n_10965), .b(n_10918), .o(n_10970) );
no02m04 g769901 ( .a(n_11045), .b(n_10989), .o(n_11080) );
no02f06 TIMEBOOST_cell_1315 ( .a(FE_OCP_RBN6564_n_12753), .b(n_12865), .o(TIMEBOOST_net_272) );
na02s02 TIMEBOOST_cell_8878 ( .a(FE_OCP_RBN6204_n_31819), .b(n_31034), .o(TIMEBOOST_net_2926) );
na02s06 g769906 ( .a(n_10915), .b(n_44498), .o(n_10939) );
in01s01 g769911 ( .a(n_11048), .o(n_11078) );
no02s06 g769912 ( .a(n_10992), .b(FE_OCP_RBN5955_FE_OFN4772_n_44463), .o(n_11048) );
na02s03 g769913 ( .a(n_10991), .b(FE_OCP_RBN5955_FE_OFN4772_n_44463), .o(n_11033) );
na04s02 TIMEBOOST_cell_8399 ( .a(n_25542), .b(n_24794), .c(n_25589), .d(n_25624), .o(n_25697) );
no02m06 TIMEBOOST_cell_7546 ( .a(TIMEBOOST_net_2082), .b(n_13751), .o(TIMEBOOST_net_2404) );
no02s04 g769916 ( .a(n_10945), .b(FE_OCPN4844_FE_OFN4779_n_44490), .o(n_11001) );
in01s01 g769918 ( .a(n_11000), .o(n_11027) );
na02s06 g769919 ( .a(n_10919), .b(FE_OFN756_n_44464), .o(n_11000) );
na02s06 g769920 ( .a(n_10878), .b(FE_OFN756_n_44464), .o(n_10912) );
na02s08 g769922 ( .a(n_10974), .b(FE_OCPN4845_FE_OFN4779_n_44490), .o(n_11122) );
na02s06 g769923 ( .a(n_10974), .b(FE_OCP_RBN5955_FE_OFN4772_n_44463), .o(n_11026) );
no02s01 g769924 ( .a(n_10910), .b(n_10802), .o(n_10936) );
no03s02 TIMEBOOST_cell_8690 ( .a(n_28025), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_15_), .c(n_27923), .o(TIMEBOOST_net_2832) );
na02m04 g769928 ( .a(n_11005), .b(FE_OCP_RBN6805_n_9742), .o(n_11035) );
in01s01 g769930 ( .a(n_11076), .o(n_11104) );
na02s03 g769931 ( .a(n_9742), .b(n_11006), .o(n_11076) );
na02m02 g769932 ( .a(n_11022), .b(n_11014), .o(n_11075) );
no02f08 g769933 ( .a(n_10948), .b(n_10891), .o(n_10971) );
in01s02 g769936 ( .a(n_11131), .o(n_11152) );
no02s06 g769937 ( .a(n_11058), .b(FE_OCP_RBN3029_n_9584), .o(n_11131) );
na02f10 TIMEBOOST_cell_5155 ( .a(TIMEBOOST_net_1525), .b(FE_RN_295_0), .o(n_25178) );
in01s02 g769939 ( .a(n_11158), .o(n_11249) );
no02m04 g769940 ( .a(n_11059), .b(n_9620), .o(n_11158) );
in01m01 g769941 ( .a(n_11156), .o(n_11157) );
na02m02 g769942 ( .a(n_11107), .b(n_11159), .o(n_11156) );
na02s01 g769943 ( .a(n_10962), .b(FE_OCP_RBN3265_n_10852), .o(n_10977) );
in01s01 g769945 ( .a(n_11180), .o(n_11154) );
na02m06 g769946 ( .a(n_11042), .b(n_10154), .o(n_11180) );
in01s02 g769947 ( .a(n_11102), .o(n_11103) );
in01m01 g769948 ( .a(n_11074), .o(n_11102) );
in01m02 g769950 ( .a(n_10880), .o(n_10881) );
oa12s04 g769951 ( .a(n_10734), .b(n_10278), .c(n_10767), .o(n_10880) );
in01m02 g769952 ( .a(n_11212), .o(n_11184) );
na02s02 TIMEBOOST_cell_1458 ( .a(TIMEBOOST_net_343), .b(n_2342), .o(n_2457) );
in01m02 g769954 ( .a(n_11096), .o(n_11097) );
ao12m02 g769955 ( .a(n_10836), .b(n_11019), .c(n_10899), .o(n_11096) );
oa12m04 g769957 ( .a(n_10825), .b(n_10857), .c(FE_OCP_RBN4359_n_10100), .o(n_10946) );
in01s02 g769958 ( .a(n_11072), .o(n_11073) );
na02s06 TIMEBOOST_cell_8601 ( .a(TIMEBOOST_net_2787), .b(n_39131), .o(n_39278) );
in01s01 g769960 ( .a(n_11024), .o(n_11025) );
in01s02 g769961 ( .a(n_10998), .o(n_11024) );
no02m06 TIMEBOOST_cell_7022 ( .a(TIMEBOOST_net_2269), .b(n_9937), .o(n_10146) );
in01s01 g769963 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_13_), .o(n_11101) );
no02m04 TIMEBOOST_cell_7021 ( .a(FE_OCP_RBN3065_n_9892), .b(FE_OCP_RBN5931_n_44563), .o(TIMEBOOST_net_2269) );
na02f08 TIMEBOOST_cell_1068 ( .a(TIMEBOOST_net_148), .b(n_23237), .o(n_23253) );
na02s03 g769970 ( .a(n_10956), .b(n_10995), .o(n_11045) );
in01m02 g769971 ( .a(n_10965), .o(n_10966) );
no02f06 TIMEBOOST_cell_3246 ( .a(n_15862), .b(n_14650), .o(TIMEBOOST_net_914) );
na02m06 g769973 ( .a(n_11018), .b(n_9494), .o(n_11159) );
na02s02 g769974 ( .a(n_11017), .b(FE_OCP_RBN3039_n_9494), .o(n_11107) );
na02s06 g769975 ( .a(n_11008), .b(n_10801), .o(n_11032) );
in01m02 g769976 ( .a(n_11043), .o(n_11044) );
no02f02 g769977 ( .a(n_11047), .b(n_10993), .o(n_11043) );
na03s10 TIMEBOOST_cell_3421 ( .a(n_37006), .b(n_36465), .c(n_46254), .o(n_37128) );
na02s02 g769979 ( .a(n_11037), .b(n_10925), .o(n_11071) );
no02f06 TIMEBOOST_cell_8566 ( .a(n_14317), .b(n_14614), .o(TIMEBOOST_net_2770) );
in01s01 g769981 ( .a(n_11069), .o(n_11070) );
ao12s01 g769982 ( .a(n_11041), .b(n_11057), .c(n_10036), .o(n_11069) );
oa12m04 g769983 ( .a(n_10082), .b(n_11057), .c(n_11041), .o(n_11042) );
in01s03 g769984 ( .a(n_10992), .o(n_11049) );
no02f08 TIMEBOOST_cell_3378 ( .a(n_31667), .b(n_31523), .o(TIMEBOOST_net_980) );
oa22s01 g769986 ( .a(n_10972), .b(n_10157), .c(n_11057), .d(n_10156), .o(n_11068) );
in01m02 g769987 ( .a(n_11058), .o(n_11059) );
no02f08 TIMEBOOST_cell_5991 ( .a(n_28011), .b(n_28012), .o(TIMEBOOST_net_1847) );
in01s06 g769989 ( .a(n_10919), .o(n_10974) );
na03f04 TIMEBOOST_cell_5880 ( .a(FE_OCP_RBN1171_n_25817), .b(n_25829), .c(n_25856), .o(n_25931) );
in01s01 g769992 ( .a(n_11003), .o(n_11022) );
in01s02 g769993 ( .a(n_10948), .o(n_11003) );
oa12f08 g769994 ( .a(n_10811), .b(n_10874), .c(n_10748), .o(n_10948) );
in01s02 g769995 ( .a(n_11055), .o(n_11098) );
no02m06 TIMEBOOST_cell_1338 ( .a(TIMEBOOST_net_283), .b(n_7869), .o(n_8269) );
in01s01 g770001 ( .a(n_10991), .o(n_11012) );
in01s02 g770002 ( .a(n_10991), .o(n_10978) );
na02m06 TIMEBOOST_cell_1268 ( .a(n_28894), .b(TIMEBOOST_net_248), .o(n_28952) );
na02s01 TIMEBOOST_cell_4267 ( .a(n_7472), .b(FE_RN_186_0), .o(TIMEBOOST_net_1224) );
in01s02 g770009 ( .a(n_11005), .o(n_11006) );
na02f08 TIMEBOOST_cell_1310 ( .a(n_13729), .b(TIMEBOOST_net_269), .o(n_13815) );
in01s01 g770013 ( .a(n_10962), .o(n_11007) );
in01s01 g770014 ( .a(n_10944), .o(n_10962) );
in01s02 g770015 ( .a(n_10944), .o(n_10945) );
in01s01 g770019 ( .a(n_10910), .o(n_10935) );
in01s01 g770020 ( .a(n_10878), .o(n_10910) );
in01s02 g770021 ( .a(n_10878), .o(n_10879) );
in01s01 g770024 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_12_), .o(n_12462) );
in01s01 g770026 ( .a(n_10917), .o(n_10918) );
no02s02 g770027 ( .a(n_10884), .b(n_10883), .o(n_10917) );
na02s03 g770029 ( .a(n_10958), .b(n_10957), .o(n_10989) );
na02s06 g770030 ( .a(n_10833), .b(FE_OFN4800_n_44498), .o(n_10894) );
no02s08 g770031 ( .a(n_10797), .b(FE_OFN756_n_44464), .o(n_10826) );
na02s02 g770032 ( .a(n_10852), .b(FE_OFN756_n_44464), .o(n_10877) );
na02s06 g770033 ( .a(n_10922), .b(FE_OCPN4845_FE_OFN4779_n_44490), .o(n_10995) );
na02m08 TIMEBOOST_cell_5474 ( .a(n_21489), .b(n_21611), .o(TIMEBOOST_net_1685) );
na02f08 TIMEBOOST_cell_1067 ( .a(FE_RN_59_0), .b(n_23113), .o(TIMEBOOST_net_148) );
no03s04 TIMEBOOST_cell_5404 ( .a(n_26453), .b(n_26416), .c(n_26514), .o(TIMEBOOST_net_1650) );
in01s02 g770037 ( .a(n_10955), .o(n_10956) );
no02s06 g770038 ( .a(n_10922), .b(FE_OCPN4845_FE_OFN4779_n_44490), .o(n_10955) );
no02s08 TIMEBOOST_cell_3377 ( .a(n_31554), .b(TIMEBOOST_net_979), .o(n_31685) );
no02s04 g770040 ( .a(n_10827), .b(FE_OCPN1932_n_9114), .o(n_10857) );
na02s02 g770041 ( .a(n_10933), .b(n_10930), .o(n_10988) );
in01m02 g770042 ( .a(n_11063), .o(n_11064) );
na02m04 g770043 ( .a(n_11106), .b(n_10985), .o(n_11063) );
no02s02 TIMEBOOST_cell_4972 ( .a(FE_RN_2080_0), .b(FE_RN_2079_0), .o(TIMEBOOST_net_1434) );
no02s06 g770045 ( .a(n_10766), .b(n_10469), .o(n_10800) );
no02s04 g770046 ( .a(n_10732), .b(n_10733), .o(n_10767) );
no02m02 g770047 ( .a(n_10906), .b(FE_OCP_RBN3034_n_9629), .o(n_10993) );
na02f06 TIMEBOOST_cell_7857 ( .a(TIMEBOOST_net_2559), .b(n_35455), .o(n_35512) );
no02s02 g770049 ( .a(n_10889), .b(n_10835), .o(n_10934) );
no02s04 TIMEBOOST_cell_7679 ( .a(TIMEBOOST_net_2470), .b(n_2889), .o(n_3040) );
no02f04 TIMEBOOST_cell_7921 ( .a(TIMEBOOST_net_2591), .b(n_5605), .o(n_5717) );
no02m04 TIMEBOOST_cell_1337 ( .a(FE_OCP_RBN6621_n_7821), .b(n_7379), .o(TIMEBOOST_net_283) );
no02f06 g770053 ( .a(n_10907), .b(n_9629), .o(n_11047) );
na02s02 TIMEBOOST_cell_1309 ( .a(n_12900), .b(n_12864), .o(TIMEBOOST_net_269) );
na02m04 g770055 ( .a(n_10832), .b(n_10851), .o(n_10908) );
in01s01 g770057 ( .a(n_11019), .o(n_11037) );
in01f01 g770058 ( .a(n_11008), .o(n_11019) );
in01f02 g770060 ( .a(n_11017), .o(n_11018) );
oa22f02 g770061 ( .a(FE_OCP_RBN6122_n_10904), .b(n_10845), .c(n_10904), .d(n_10846), .o(n_11017) );
in01s02 g770062 ( .a(n_11061), .o(n_11036) );
no02m04 TIMEBOOST_cell_6050 ( .a(TIMEBOOST_net_1876), .b(n_19177), .o(TIMEBOOST_net_1478) );
na02s06 g770065 ( .a(n_10898), .b(n_10897), .o(n_10958) );
no02s06 g770066 ( .a(n_10762), .b(n_10809), .o(n_10884) );
in01s01 g770067 ( .a(n_10932), .o(n_10933) );
no02s02 g770068 ( .a(n_10898), .b(n_10875), .o(n_10932) );
no02m06 g770069 ( .a(n_10823), .b(n_10875), .o(n_10957) );
na02s06 g770070 ( .a(n_10791), .b(n_10792), .o(n_10883) );
in01m02 g770071 ( .a(n_10831), .o(n_10832) );
na02f04 g770072 ( .a(n_10792), .b(n_10763), .o(n_10831) );
in01s02 g770073 ( .a(n_10930), .o(n_10931) );
na02s04 g770074 ( .a(n_10897), .b(n_10849), .o(n_10930) );
na02s04 g770075 ( .a(n_10950), .b(FE_OCP_RBN4316_n_9292), .o(n_11106) );
na02m06 g770076 ( .a(n_10940), .b(n_10914), .o(n_10941) );
na02s03 g770077 ( .a(n_10673), .b(n_10733), .o(n_10734) );
in01s02 g770078 ( .a(n_10986), .o(n_10987) );
na02m02 g770079 ( .a(n_10940), .b(n_10953), .o(n_10986) );
in01m02 g770080 ( .a(n_10984), .o(n_10985) );
no02f04 g770081 ( .a(n_10950), .b(FE_OCP_RBN4316_n_9292), .o(n_10984) );
in01s02 g770082 ( .a(n_10855), .o(n_10856) );
in01s02 g770083 ( .a(n_10827), .o(n_10855) );
na02s02 g770085 ( .a(n_10761), .b(FE_OCPN1932_n_9114), .o(n_10825) );
in01s04 g770086 ( .a(n_10765), .o(n_10766) );
in01s03 g770087 ( .a(n_10732), .o(n_10765) );
na02f08 TIMEBOOST_cell_6752 ( .a(TIMEBOOST_net_2133), .b(n_15743), .o(n_15915) );
na02s02 g770090 ( .a(n_10893), .b(n_10746), .o(n_10952) );
in01m01 g770091 ( .a(n_11015), .o(n_11016) );
na02m02 g770092 ( .a(n_10983), .b(n_10982), .o(n_11015) );
in01s01 g770093 ( .a(n_11057), .o(n_10972) );
oa12m06 g770094 ( .a(n_10077), .b(n_10951), .c(n_9951), .o(n_11057) );
in01s01 g770095 ( .a(n_10959), .o(n_10928) );
na02m06 TIMEBOOST_cell_1334 ( .a(TIMEBOOST_net_281), .b(FE_OCP_RBN4181_n_19599), .o(n_19747) );
oa12s01 g770097 ( .a(n_10943), .b(n_10951), .c(n_10942), .o(n_10981) );
in01s01 g770100 ( .a(n_10797), .o(n_10802) );
in01s03 g770101 ( .a(n_10797), .o(n_10778) );
na03f02 TIMEBOOST_cell_7256 ( .a(n_38703), .b(n_38697), .c(n_38728), .o(n_38765) );
in01s01 g770103 ( .a(n_10889), .o(n_10890) );
in01s01 g770104 ( .a(n_10874), .o(n_10889) );
oa12f08 g770105 ( .a(n_10634), .b(n_10821), .c(n_10678), .o(n_10874) );
na02s02 TIMEBOOST_cell_5552 ( .a(n_6179), .b(n_6116), .o(TIMEBOOST_net_1724) );
no02m08 TIMEBOOST_cell_4031 ( .a(n_46958), .b(FE_OCPN5300_n_27130), .o(TIMEBOOST_net_1106) );
oa12s04 g770111 ( .a(n_10347), .b(n_10770), .c(n_10768), .o(n_10798) );
na02m08 TIMEBOOST_cell_8614 ( .a(FE_OCPN1382_n_45026), .b(FE_OCP_RBN1868_n_21358), .o(TIMEBOOST_net_2794) );
ao12s04 g770113 ( .a(n_10360), .b(n_44852), .c(n_10699), .o(n_10731) );
na02m06 g770114 ( .a(n_10700), .b(n_10280), .o(n_10764) );
in01f02 g770115 ( .a(n_10906), .o(n_10907) );
in01s02 g770117 ( .a(n_10833), .o(n_10806) );
no02s06 g770118 ( .a(n_10704), .b(n_10729), .o(n_10833) );
na02s01 g770122 ( .a(n_10951), .b(n_10942), .o(n_10943) );
no02m04 g770124 ( .a(n_10804), .b(n_10691), .o(n_10904) );
no02s06 g770125 ( .a(n_10803), .b(n_10755), .o(n_10898) );
in01s02 g770126 ( .a(n_10850), .o(n_10851) );
na02s04 g770127 ( .a(n_10809), .b(n_10791), .o(n_10850) );
na02s06 g770128 ( .a(n_10730), .b(FE_OCP_RBN5938_n_44563), .o(n_10792) );
na02s06 g770129 ( .a(n_10810), .b(n_44492), .o(n_10897) );
na02s02 g770130 ( .a(n_10742), .b(FE_OCPN1067_n_44461), .o(n_10782) );
no02m04 g770131 ( .a(n_10810), .b(FE_OFN756_n_44464), .o(n_10823) );
na02m02 g770132 ( .a(n_10787), .b(FE_OCP_RBN6740_n_44563), .o(n_10849) );
no02s02 g770133 ( .a(n_10676), .b(n_44492), .o(n_10704) );
no03f20 TIMEBOOST_cell_4603 ( .a(n_23195), .b(FE_RN_748_0), .c(n_23077), .o(n_23328) );
no02s06 g770135 ( .a(FE_OCP_RBN3242_n_10676), .b(FE_OCP_RBN5953_FE_OFN4772_n_44463), .o(n_10729) );
in01f02 g770136 ( .a(n_10762), .o(n_10763) );
no02m06 g770137 ( .a(n_10730), .b(FE_OCPN4847_FE_OFN4778_n_44490), .o(n_10762) );
na02m04 g770138 ( .a(n_10828), .b(FE_OCP_RBN2924_n_9198), .o(n_10940) );
no02s01 TIMEBOOST_cell_1255 ( .a(n_37733), .b(n_37716), .o(TIMEBOOST_net_242) );
na02s04 g770140 ( .a(n_10902), .b(n_44821), .o(n_10983) );
na02f04 TIMEBOOST_cell_7824 ( .a(n_26055), .b(FE_OCPN1390_n_26054), .o(TIMEBOOST_net_2543) );
no02s04 g770142 ( .a(n_44852), .b(n_10412), .o(n_10702) );
na02s04 TIMEBOOST_cell_8706 ( .a(n_40720), .b(FE_RN_902_0), .o(TIMEBOOST_net_2840) );
in01s01 g770144 ( .a(n_10672), .o(n_10673) );
na02s06 g770145 ( .a(n_10599), .b(n_10329), .o(n_10672) );
no02m06 g770146 ( .a(n_10871), .b(n_10805), .o(n_10872) );
na02m06 g770147 ( .a(n_10829), .b(FE_OCP_RBN6750_n_9198), .o(n_10953) );
na02m04 g770148 ( .a(n_44852), .b(n_10699), .o(n_10700) );
no02f06 g770149 ( .a(n_10862), .b(n_10864), .o(n_10865) );
na02s02 g770150 ( .a(n_10788), .b(n_10714), .o(n_10861) );
no03f04 TIMEBOOST_cell_4786 ( .a(FE_OCP_RBN4319_n_14768), .b(n_16535), .c(n_16474), .o(n_16536) );
in01s02 g770152 ( .a(n_10760), .o(n_10761) );
na02s02 TIMEBOOST_cell_7507 ( .a(TIMEBOOST_net_2384), .b(n_12686), .o(n_12743) );
in01s02 g770155 ( .a(n_10920), .o(n_10921) );
no02m02 g770156 ( .a(n_10903), .b(n_10871), .o(n_10920) );
in01m02 g770157 ( .a(n_10927), .o(n_10982) );
no02m04 g770158 ( .a(n_10902), .b(n_44821), .o(n_10927) );
in01s01 g770159 ( .a(n_10892), .o(n_10893) );
oa12s02 g770160 ( .a(n_10653), .b(n_10813), .c(n_10864), .o(n_10892) );
na03m20 TIMEBOOST_cell_6400 ( .a(n_22708), .b(delay_xor_ln21_unr15_stage6_stallmux_q_1_), .c(FE_OCP_RBN6463_n_44061), .o(n_22746) );
in01s02 g770162 ( .a(n_46988), .o(n_10980) );
no02f06 g770164 ( .a(n_10862), .b(n_10608), .o(n_10863) );
in01s01 g770166 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_17_), .o(n_11784) );
in01s01 g770168 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_11_), .o(n_12452) );
in01s02 g770170 ( .a(n_10803), .o(n_10804) );
na02s06 g770171 ( .a(n_10754), .b(n_10724), .o(n_10803) );
in01m02 g770172 ( .a(n_10789), .o(n_10790) );
no02m04 g770173 ( .a(n_10759), .b(n_10601), .o(n_10789) );
na02s06 g770174 ( .a(n_10759), .b(n_10735), .o(n_10809) );
na02m04 g770175 ( .a(n_10796), .b(n_10772), .o(n_10847) );
na02s06 g770176 ( .a(n_10727), .b(n_10664), .o(n_10875) );
na03m10 TIMEBOOST_cell_6399 ( .a(n_22634), .b(n_45204), .c(FE_OCP_RBN5459_n_44061), .o(n_22672) );
no02s06 g770178 ( .a(n_10669), .b(n_10601), .o(n_10791) );
in01s02 g770179 ( .a(n_10845), .o(n_10846) );
na02m04 g770180 ( .a(n_10710), .b(n_10756), .o(n_10845) );
in01s02 g770181 ( .a(n_10757), .o(n_10758) );
na02m04 g770182 ( .a(n_10670), .b(n_10735), .o(n_10757) );
na02s01 g770183 ( .a(n_10813), .b(n_10684), .o(n_10900) );
in01s01 g770184 ( .a(n_11013), .o(n_11014) );
na02s02 g770185 ( .a(n_10914), .b(n_10979), .o(n_11013) );
no02f08 g770186 ( .a(n_10779), .b(n_10584), .o(n_10862) );
no02m04 g770187 ( .a(n_10784), .b(FE_OCP_RBN2984_n_9247), .o(n_10871) );
no02m04 g770188 ( .a(n_10785), .b(n_9247), .o(n_10903) );
oa12m06 g770190 ( .a(n_9953), .b(n_10869), .c(n_10039), .o(n_10951) );
oa12s01 g770191 ( .a(n_10818), .b(n_10817), .c(n_10816), .o(n_10868) );
oa12s01 g770192 ( .a(n_10842), .b(n_10869), .c(n_10841), .o(n_10913) );
in01s01 g770193 ( .a(n_10821), .o(n_10788) );
ao12f08 g770194 ( .a(n_10556), .b(n_10745), .c(n_10603), .o(n_10821) );
in01s01 g770195 ( .a(n_10799), .o(n_10885) );
ao12s01 g770196 ( .a(n_10726), .b(n_10745), .c(n_10725), .o(n_10799) );
no02m04 TIMEBOOST_cell_1036 ( .a(TIMEBOOST_net_132), .b(n_23126), .o(n_23228) );
na02m06 TIMEBOOST_cell_4504 ( .a(TIMEBOOST_net_1342), .b(n_5718), .o(n_5881) );
in01s02 g770202 ( .a(n_10828), .o(n_10829) );
oa22f02 g770203 ( .a(n_10722), .b(n_10692), .c(n_10723), .d(n_10693), .o(n_10828) );
in01s04 g770204 ( .a(n_10711), .o(n_10770) );
na02m04 TIMEBOOST_cell_1232 ( .a(n_18703), .b(TIMEBOOST_net_230), .o(n_18702) );
in01m01 g770211 ( .a(n_10810), .o(n_10787) );
na02s01 TIMEBOOST_cell_5555 ( .a(TIMEBOOST_net_1725), .b(n_16977), .o(n_17321) );
no02s01 TIMEBOOST_cell_1242 ( .a(TIMEBOOST_net_235), .b(n_7413), .o(n_45864) );
na02s02 TIMEBOOST_cell_8861 ( .a(TIMEBOOST_net_2917), .b(n_6269), .o(TIMEBOOST_net_1733) );
na02s01 g770222 ( .a(n_10869), .b(n_10841), .o(n_10842) );
no02s06 g770223 ( .a(n_10667), .b(n_10696), .o(n_10759) );
no02f04 TIMEBOOST_cell_6981 ( .a(FE_OCP_RBN4923_n_34980), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(TIMEBOOST_net_2249) );
no02s01 TIMEBOOST_cell_6083 ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .b(n_38778), .o(TIMEBOOST_net_1893) );
in01s02 g770226 ( .a(n_10755), .o(n_10756) );
no02m06 g770227 ( .a(n_10709), .b(FE_OCPN4847_FE_OFN4778_n_44490), .o(n_10755) );
na02s03 g770228 ( .a(n_10568), .b(FE_OCP_RBN5949_FE_OFN4772_n_44463), .o(n_10594) );
na02s02 g770229 ( .a(n_10709), .b(FE_OCP_RBN6740_n_44563), .o(n_10727) );
na02s02 g770230 ( .a(n_10709), .b(FE_OCP_RBN5937_n_44563), .o(n_10710) );
na02s01 TIMEBOOST_cell_5554 ( .a(FE_OCP_RBN3111_n_15817), .b(n_17032), .o(TIMEBOOST_net_1725) );
no02s02 g770232 ( .a(n_10644), .b(n_44492), .o(n_10671) );
na02s08 TIMEBOOST_cell_3199 ( .a(n_26013), .b(TIMEBOOST_net_890), .o(n_26146) );
na02s06 g770234 ( .a(n_10629), .b(FE_OCPN1063_n_44461), .o(n_10735) );
in01m02 g770235 ( .a(n_10669), .o(n_10670) );
no02m06 g770236 ( .a(n_10629), .b(FE_OCPN1063_n_44461), .o(n_10669) );
na02s01 g770237 ( .a(n_10817), .b(n_10816), .o(n_10818) );
no02s01 TIMEBOOST_cell_4536 ( .a(TIMEBOOST_net_1358), .b(TIMEBOOST_net_982), .o(n_31858) );
no02s01 TIMEBOOST_cell_1241 ( .a(n_45858), .b(n_6862), .o(TIMEBOOST_net_235) );
na03s02 TIMEBOOST_cell_8263 ( .a(FE_OCP_RBN5769_n_3338), .b(n_2913), .c(n_3339), .o(n_3428) );
in01s02 g770241 ( .a(n_10925), .o(n_10926) );
na02s02 g770242 ( .a(n_10801), .b(n_10899), .o(n_10925) );
in01s01 g770244 ( .a(n_10914), .o(n_10923) );
na02m04 g770245 ( .a(n_46989), .b(FE_OCP_RBN2934_n_9075), .o(n_10914) );
na02s06 g770246 ( .a(n_10569), .b(n_10592), .o(n_10620) );
no02s02 TIMEBOOST_cell_2135 ( .a(n_21075), .b(n_44277), .o(TIMEBOOST_net_682) );
no02s01 g770248 ( .a(n_10745), .b(n_10725), .o(n_10726) );
in01s02 g770249 ( .a(n_10891), .o(n_10979) );
no02s06 g770250 ( .a(n_46989), .b(FE_OCP_RBN2933_n_9075), .o(n_10891) );
in01m02 g770251 ( .a(n_10795), .o(n_10796) );
in01f02 g770252 ( .a(n_10754), .o(n_10795) );
na02f08 g770253 ( .a(n_10666), .b(n_10647), .o(n_10754) );
oa12s01 g770254 ( .a(n_10753), .b(n_10752), .c(n_10751), .o(n_10815) );
oa12s01 g770255 ( .a(n_10777), .b(n_10776), .c(n_10775), .o(n_10840) );
in01s01 g770256 ( .a(n_10848), .o(n_10814) );
oa22s01 g770257 ( .a(n_10740), .b(n_10554), .c(n_10681), .d(n_10555), .o(n_10848) );
in01s01 g770260 ( .a(n_10779), .o(n_10813) );
in01m02 g770262 ( .a(n_10784), .o(n_10785) );
oa22m04 g770263 ( .a(FE_OCP_RBN6093_n_10660), .b(n_10615), .c(n_10660), .d(n_10616), .o(n_10784) );
in01s01 g770264 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_), .o(n_10812) );
na02s01 g770268 ( .a(n_10776), .b(n_10775), .o(n_10777) );
na02s01 g770269 ( .a(n_10752), .b(n_10751), .o(n_10753) );
in01s02 g770270 ( .a(n_10772), .o(n_10773) );
na02m04 g770271 ( .a(n_10690), .b(n_10724), .o(n_10772) );
in01s02 g770272 ( .a(n_10736), .o(n_10737) );
no02m02 g770273 ( .a(n_10601), .b(n_10696), .o(n_10736) );
na02s01 TIMEBOOST_cell_6263 ( .a(FE_OCPN1663_n_4556), .b(n_4675), .o(TIMEBOOST_net_1983) );
in01s01 g770276 ( .a(n_10801), .o(n_10836) );
na02m04 g770277 ( .a(n_10781), .b(FE_OCP_RBN2989_n_9182), .o(n_10801) );
in01s01 g770278 ( .a(n_10618), .o(n_10619) );
na02s02 g770279 ( .a(n_10573), .b(n_10592), .o(n_10618) );
na02s02 TIMEBOOST_cell_1231 ( .a(n_18701), .b(n_18449), .o(TIMEBOOST_net_230) );
in01s01 g770281 ( .a(n_10834), .o(n_10835) );
na02s02 g770282 ( .a(n_10749), .b(n_10811), .o(n_10834) );
in01s02 g770283 ( .a(n_10517), .o(n_10518) );
na02s04 g770284 ( .a(n_10485), .b(n_47263), .o(n_10517) );
in01m01 g770285 ( .a(n_10805), .o(n_10899) );
no02m04 g770286 ( .a(n_10781), .b(FE_OCP_RBN2989_n_9182), .o(n_10805) );
na02m08 TIMEBOOST_cell_5063 ( .a(TIMEBOOST_net_1479), .b(n_14477), .o(n_14645) );
in01s02 g770288 ( .a(n_10722), .o(n_10723) );
ao12f02 g770289 ( .a(n_10604), .b(n_10626), .c(n_10677), .o(n_10722) );
in01m01 g770291 ( .a(n_10667), .o(n_10694) );
ao12f06 g770292 ( .a(n_10571), .b(n_10478), .c(n_10548), .o(n_10667) );
oa12s01 g770294 ( .a(n_9915), .b(n_10720), .c(n_9824), .o(n_10817) );
in01s01 g770295 ( .a(n_10739), .o(n_10721) );
oa12s01 g770296 ( .a(n_10641), .b(n_10650), .c(n_10640), .o(n_10739) );
oa12f08 g770297 ( .a(n_10454), .b(n_10650), .c(n_10523), .o(n_10745) );
no02m02 TIMEBOOST_cell_8792 ( .a(TIMEBOOST_net_1242), .b(n_24621), .o(TIMEBOOST_net_2883) );
ao12s06 g770300 ( .a(n_10148), .b(n_10406), .c(n_10484), .o(n_10507) );
oa12s04 g770301 ( .a(FE_OCP_RBN4357_n_10100), .b(n_10541), .c(n_8908), .o(n_10569) );
na03m06 TIMEBOOST_cell_7315 ( .a(n_16918), .b(n_16834), .c(n_16954), .o(n_17199) );
na02s01 g770310 ( .a(n_10720), .b(n_9955), .o(n_10776) );
na02s02 g770312 ( .a(n_10654), .b(n_10682), .o(n_10719) );
no02f08 TIMEBOOST_cell_3193 ( .a(TIMEBOOST_net_887), .b(n_39110), .o(n_39145) );
na02m06 g770314 ( .a(n_10612), .b(n_44492), .o(n_10724) );
no02m06 g770318 ( .a(n_10538), .b(FE_OFN756_n_44464), .o(n_10601) );
in01s02 g770319 ( .a(n_10692), .o(n_10693) );
na02m02 g770320 ( .a(n_10614), .b(n_10665), .o(n_10692) );
in01s01 g770321 ( .a(n_10690), .o(n_10691) );
na02s02 g770322 ( .a(FE_OCP_RBN3241_n_10612), .b(FE_OCPN4847_FE_OFN4778_n_44490), .o(n_10664) );
na02m04 g770323 ( .a(FE_OCP_RBN3240_n_10612), .b(FE_OCP_RBN5938_n_44563), .o(n_10690) );
na02s04 g770324 ( .a(n_10570), .b(FE_OCP_RBN5952_FE_OFN4772_n_44463), .o(n_10591) );
no02s10 TIMEBOOST_cell_3355 ( .a(n_32026), .b(TIMEBOOST_net_968), .o(n_32107) );
no02s04 g770326 ( .a(n_10537), .b(FE_OFN4775_n_44463), .o(n_10696) );
na02s06 TIMEBOOST_cell_4444 ( .a(TIMEBOOST_net_1312), .b(FE_OCP_RBN6056_n_46957), .o(n_30960) );
no02s01 g770328 ( .a(n_10543), .b(FE_OCP_RBN3147_n_10369), .o(n_10545) );
na02s01 g770329 ( .a(n_10650), .b(n_10640), .o(n_10641) );
na02s01 g770330 ( .a(n_10543), .b(FE_OCP_RBN3147_n_10369), .o(n_10544) );
na02s06 g770331 ( .a(n_10541), .b(n_10241), .o(n_10573) );
na02s06 g770332 ( .a(n_10405), .b(n_10324), .o(n_10485) );
na02m06 g770333 ( .a(n_10707), .b(FE_OCP_RBN4262_n_9009), .o(n_10811) );
in01s01 g770334 ( .a(n_10748), .o(n_10749) );
no02m06 g770335 ( .a(n_10707), .b(FE_OCP_RBN4262_n_9009), .o(n_10748) );
ao12s01 g770337 ( .a(n_9775), .b(n_10689), .c(n_9870), .o(n_10752) );
na02s02 TIMEBOOST_cell_4277 ( .a(n_33557), .b(n_33817), .o(TIMEBOOST_net_1229) );
no02f04 g770340 ( .a(n_10597), .b(n_10508), .o(n_10660) );
no02s01 TIMEBOOST_cell_1184 ( .a(TIMEBOOST_net_206), .b(n_37826), .o(n_37854) );
oa12s01 g770342 ( .a(n_10688), .b(n_10687), .c(n_10686), .o(n_10744) );
oa12s01 g770343 ( .a(n_10658), .b(n_10689), .c(n_10657), .o(n_10717) );
in01s02 g770344 ( .a(n_10746), .o(n_10747) );
oa22s01 g770345 ( .a(n_10712), .b(FE_OCP_RBN2936_n_8981), .c(n_10630), .d(n_8981), .o(n_10746) );
na02m04 g770346 ( .a(n_10639), .b(n_10656), .o(n_10781) );
in01s01 g770347 ( .a(n_10740), .o(n_10681) );
oa12f06 g770348 ( .a(n_10393), .b(n_10659), .c(n_10380), .o(n_10740) );
in01s01 g770349 ( .a(n_10716), .o(n_10783) );
ao12s01 g770350 ( .a(n_10638), .b(n_10659), .c(n_10637), .o(n_10716) );
in01s01 g770351 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_13_), .o(n_10708) );
in01s01 g770353 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_14_), .o(n_12164) );
na02s01 g770357 ( .a(n_10687), .b(n_10686), .o(n_10688) );
na02s01 g770358 ( .a(n_10689), .b(n_10657), .o(n_10658) );
no02m04 g770359 ( .a(n_10567), .b(n_10586), .o(n_10597) );
na02m02 g770360 ( .a(n_10567), .b(n_10610), .o(n_10656) );
in01s02 g770362 ( .a(n_10626), .o(n_10654) );
no02f02 g770363 ( .a(n_10624), .b(n_44053), .o(n_10626) );
no02m06 g770364 ( .a(n_10547), .b(n_10508), .o(n_10548) );
na02s02 g770365 ( .a(n_10588), .b(n_10609), .o(n_10639) );
na02m04 g770366 ( .a(n_10582), .b(FE_OFN757_n_44464), .o(n_10665) );
in01m02 g770367 ( .a(n_10615), .o(n_10616) );
no02m02 g770368 ( .a(n_10536), .b(n_10547), .o(n_10615) );
no02s01 TIMEBOOST_cell_1183 ( .a(n_37751), .b(n_37784), .o(TIMEBOOST_net_206) );
na02s02 g770370 ( .a(n_10564), .b(FE_OCPN4847_FE_OFN4778_n_44490), .o(n_10614) );
in01s01 g770371 ( .a(n_10713), .o(n_10714) );
no02s02 g770372 ( .a(n_10635), .b(n_10678), .o(n_10713) );
no02s01 g770373 ( .a(n_10659), .b(n_10637), .o(n_10638) );
na02m06 g770374 ( .a(n_10689), .b(n_9829), .o(n_10720) );
na02s04 g770375 ( .a(n_10535), .b(n_10506), .o(n_10571) );
in01s01 g770377 ( .a(n_10541), .o(n_10511) );
oa12s08 g770378 ( .a(n_10145), .b(n_10404), .c(n_10116), .o(n_10541) );
in01m03 g770381 ( .a(n_10480), .o(n_10543) );
oa12f06 g770384 ( .a(n_10489), .b(n_10575), .c(n_10417), .o(n_10650) );
na02f06 TIMEBOOST_cell_1306 ( .a(TIMEBOOST_net_267), .b(n_29233), .o(n_29380) );
in01s01 g770388 ( .a(FE_OCP_RBN4385_n_10570), .o(n_10613) );
no02f06 TIMEBOOST_cell_4511 ( .a(n_39645), .b(n_39674), .o(TIMEBOOST_net_1346) );
in01s01 g770394 ( .a(n_10636), .o(n_10705) );
ao12s01 g770395 ( .a(n_10566), .b(n_10575), .c(n_10565), .o(n_10636) );
in01s02 g770397 ( .a(n_10405), .o(n_10445) );
in01s02 g770398 ( .a(n_10405), .o(n_10406) );
oa12s08 g770399 ( .a(n_10153), .b(n_10243), .c(n_10197), .o(n_10405) );
in01f02 g770400 ( .a(n_10537), .o(n_10538) );
na02f08 TIMEBOOST_cell_7004 ( .a(TIMEBOOST_net_2260), .b(n_10594), .o(n_10730) );
in01s01 g770402 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_8_), .o(n_10611) );
in01s01 g770405 ( .a(n_10567), .o(n_10588) );
na02m08 g770406 ( .a(FE_OCP_RBN6058_n_10478), .b(n_10331), .o(n_10567) );
na02f02 g770407 ( .a(n_44054), .b(n_10514), .o(n_10587) );
na02s20 TIMEBOOST_cell_914 ( .a(TIMEBOOST_net_71), .b(FE_OCP_RBN5542_n_23044), .o(n_23195) );
no02s04 g770409 ( .a(n_10483), .b(FE_OFN4775_n_44463), .o(n_10547) );
na02s02 g770411 ( .a(n_10677), .b(n_10598), .o(n_10682) );
in01m01 g770412 ( .a(n_10535), .o(n_10536) );
na02m04 g770413 ( .a(n_10483), .b(FE_OFN4778_n_44490), .o(n_10535) );
no02f04 g770414 ( .a(n_10477), .b(FE_OCP_RBN5949_FE_OFN4772_n_44463), .o(n_10505) );
in01m02 g770415 ( .a(n_10609), .o(n_10610) );
no02m02 g770416 ( .a(n_10586), .b(n_10508), .o(n_10609) );
no02s06 TIMEBOOST_cell_4510 ( .a(TIMEBOOST_net_1345), .b(n_16518), .o(n_16570) );
in01s01 TIMEBOOST_cell_7380 ( .a(n_36750), .o(TIMEBOOST_net_2316) );
no02f08 TIMEBOOST_cell_4436 ( .a(TIMEBOOST_net_1308), .b(n_16094), .o(n_16230) );
na02m04 g770420 ( .a(n_10579), .b(FE_OCP_RBN2936_n_8981), .o(n_10608) );
no02s06 g770421 ( .a(n_10607), .b(FE_OCP_RBN4247_n_8904), .o(n_10678) );
no02s01 g770422 ( .a(n_10575), .b(n_10565), .o(n_10566) );
na02s01 g770424 ( .a(n_10653), .b(n_10579), .o(n_10684) );
na02f06 TIMEBOOST_cell_1305 ( .a(n_29143), .b(FE_OFN774_n_25834), .o(TIMEBOOST_net_267) );
no02m04 g770426 ( .a(n_10526), .b(n_10562), .o(n_10585) );
in01s01 g770427 ( .a(n_10634), .o(n_10635) );
na02m04 g770428 ( .a(n_10607), .b(FE_OCP_RBN4247_n_8904), .o(n_10634) );
oa12m06 g770429 ( .a(n_9773), .b(n_10551), .c(n_9776), .o(n_10689) );
oa12s01 g770430 ( .a(n_9811), .b(n_10633), .c(n_9772), .o(n_10687) );
oa12s01 g770432 ( .a(n_10578), .b(n_10577), .c(n_10576), .o(n_10632) );
oa22s01 g770433 ( .a(n_10633), .b(n_9813), .c(n_10551), .d(n_9814), .o(n_10652) );
in01s01 g770434 ( .a(n_10582), .o(n_10564) );
ao12f06 g770436 ( .a(n_10349), .b(n_10572), .c(n_10423), .o(n_10659) );
in01s01 g770437 ( .a(n_10631), .o(n_10680) );
ao12s01 g770438 ( .a(n_10561), .b(n_10572), .c(n_10560), .o(n_10631) );
in01s01 g770439 ( .a(n_10712), .o(n_10630) );
na02m04 g770440 ( .a(n_10531), .b(n_10550), .o(n_10712) );
na02s01 g770444 ( .a(n_10577), .b(n_10576), .o(n_10578) );
in01s01 g770449 ( .a(n_10598), .o(n_10604) );
na03s40 TIMEBOOST_cell_913 ( .a(FE_OCP_RBN2422_n_23023), .b(FE_OCP_RBN3979_n_22972), .c(FE_OCP_RBN5522_n_23078), .o(TIMEBOOST_net_71) );
no02s02 g770453 ( .a(n_10401), .b(FE_OFN757_n_44464), .o(n_10586) );
in01s02 g770455 ( .a(n_10562), .o(n_10563) );
na02s02 g770456 ( .a(n_10473), .b(n_10503), .o(n_10562) );
na02s02 g770457 ( .a(n_10513), .b(FE_OCP_RBN6741_n_44563), .o(n_10514) );
na02s02 g770458 ( .a(n_10513), .b(FE_OCPN4847_FE_OFN4778_n_44490), .o(n_10677) );
no02m06 g770462 ( .a(n_10437), .b(FE_OFN4778_n_44490), .o(n_10508) );
no02s01 g770463 ( .a(n_10572), .b(n_10560), .o(n_10561) );
na02s01 g770464 ( .a(n_10557), .b(n_10603), .o(n_10725) );
in01m02 g770466 ( .a(n_10579), .o(n_10864) );
na02m04 g770467 ( .a(n_10559), .b(FE_OCP_RBN2903_n_8902), .o(n_10579) );
na02s02 g770468 ( .a(n_10499), .b(n_10402), .o(n_10531) );
in01s01 g770469 ( .a(n_10584), .o(n_10653) );
no02m06 g770470 ( .a(n_10559), .b(FE_OCP_RBN2903_n_8902), .o(n_10584) );
na02s04 g770471 ( .a(n_10500), .b(n_10403), .o(n_10550) );
no02f06 g770473 ( .a(n_10328), .b(n_10368), .o(n_10478) );
in01s02 g770474 ( .a(n_10440), .o(n_10441) );
in01s02 g770475 ( .a(n_10404), .o(n_10440) );
oa12m08 g770476 ( .a(n_9942), .b(n_10277), .c(n_9978), .o(n_10404) );
oa12f06 g770477 ( .a(n_10251), .b(n_10481), .c(n_10342), .o(n_10575) );
na02s01 TIMEBOOST_cell_6363 ( .a(FE_OCP_RBN6175_n_16923), .b(n_15901), .o(TIMEBOOST_net_2033) );
ao22f02 g770483 ( .a(n_10195), .b(n_10150), .c(FE_OCP_RBN3113_n_10195), .d(n_10149), .o(n_10369) );
oa12s01 g770484 ( .a(n_10472), .b(n_10481), .c(n_10471), .o(n_10530) );
no02s02 TIMEBOOST_cell_3176 ( .a(n_4104), .b(n_4006), .o(TIMEBOOST_net_879) );
in01s01 g770486 ( .a(FE_OCP_RBN3181_n_10477), .o(n_11435) );
in01s01 g770490 ( .a(n_10320), .o(n_10321) );
in01s02 g770491 ( .a(n_10243), .o(n_10320) );
oa12s08 g770492 ( .a(n_10022), .b(n_10101), .c(n_10020), .o(n_10243) );
na02s04 g770494 ( .a(n_10474), .b(n_10433), .o(n_10475) );
in01s01 g770495 ( .a(n_10330), .o(n_10331) );
na02s02 g770496 ( .a(n_10319), .b(n_10096), .o(n_10330) );
no02m04 TIMEBOOST_cell_5503 ( .a(TIMEBOOST_net_1699), .b(n_11047), .o(n_11072) );
na02m04 g770498 ( .a(n_10332), .b(n_10104), .o(n_10368) );
na02s02 g770500 ( .a(n_10394), .b(FE_OCPN4847_FE_OFN4778_n_44490), .o(n_10473) );
na02f04 g770501 ( .a(n_10411), .b(FE_OFN757_n_44464), .o(n_10503) );
in01s01 g770502 ( .a(n_10402), .o(n_10403) );
na02s01 g770503 ( .a(n_10319), .b(n_10332), .o(n_10402) );
na02s02 g770504 ( .a(n_10274), .b(FE_OFN756_n_44464), .o(n_10325) );
na02s04 TIMEBOOST_cell_3175 ( .a(TIMEBOOST_net_878), .b(n_34754), .o(n_34878) );
in01s01 g770506 ( .a(n_10365), .o(n_10366) );
na02s02 g770507 ( .a(n_10324), .b(n_47263), .o(n_10365) );
na02s01 g770508 ( .a(n_10481), .b(n_10471), .o(n_10472) );
na02s06 g770509 ( .a(n_10529), .b(FE_OCP_RBN4238_n_8781), .o(n_10603) );
in01s01 g770510 ( .a(n_10556), .o(n_10557) );
no02s06 g770511 ( .a(n_10529), .b(FE_OCP_RBN4238_n_8781), .o(n_10556) );
in01s01 g770512 ( .a(n_10412), .o(n_10413) );
na02s01 g770513 ( .a(n_10280), .b(n_10282), .o(n_10412) );
na02s02 g770514 ( .a(n_10153), .b(n_10230), .o(n_10318) );
no02s02 g770515 ( .a(n_10197), .b(n_10228), .o(n_10317) );
ao12s01 g770516 ( .a(n_9651), .b(n_10527), .c(n_9730), .o(n_10577) );
in01s01 g770518 ( .a(n_10551), .o(n_10633) );
na02s04 TIMEBOOST_cell_8624 ( .a(n_10884), .b(n_10894), .o(TIMEBOOST_net_2799) );
in01s02 g770520 ( .a(n_10525), .o(n_10526) );
oa12m04 g770521 ( .a(n_10398), .b(n_10474), .c(n_10286), .o(n_10525) );
in01m02 g770522 ( .a(n_10499), .o(n_10500) );
ao12m02 g770523 ( .a(n_10265), .b(n_10435), .c(n_10313), .o(n_10499) );
oa12s01 g770524 ( .a(n_10492), .b(n_10527), .c(n_10491), .o(n_10549) );
oa12f06 g770525 ( .a(n_10174), .b(n_10498), .c(n_10257), .o(n_10572) );
in01m02 g770527 ( .a(n_10401), .o(n_10437) );
na02f04 g770530 ( .a(n_10362), .b(n_10397), .o(n_10513) );
in01s01 g770531 ( .a(FE_OCP_RBN3161_n_10399), .o(n_10451) );
oa12s01 g770535 ( .a(n_10432), .b(n_10431), .c(n_10430), .o(n_10496) );
oa12s01 g770536 ( .a(n_10462), .b(n_10498), .c(n_10461), .o(n_10524) );
in01s01 g770537 ( .a(n_10554), .o(n_10555) );
oa12s01 g770538 ( .a(n_46420), .b(n_10465), .c(n_10464), .o(n_10554) );
na02m08 TIMEBOOST_cell_6660 ( .a(TIMEBOOST_net_2087), .b(TIMEBOOST_net_1471), .o(n_19609) );
in01s01 g770540 ( .a(n_10494), .o(n_10495) );
na02s01 g770541 ( .a(n_10396), .b(n_10359), .o(n_10494) );
in01s01 g770542 ( .a(n_10469), .o(n_10470) );
oa22s01 g770543 ( .a(n_10148), .b(n_10733), .c(n_10278), .d(n_9200), .o(n_10469) );
in01s01 g770544 ( .a(n_10363), .o(n_10364) );
oa22s01 g770545 ( .a(n_10148), .b(n_10484), .c(n_10194), .d(n_8937), .o(n_10363) );
in01s01 g770546 ( .a(n_10467), .o(n_10468) );
na02s02 g770547 ( .a(n_10337), .b(n_10279), .o(n_10467) );
na02s01 g770551 ( .a(n_10527), .b(n_10491), .o(n_10492) );
no02m04 TIMEBOOST_cell_8584 ( .a(n_35053), .b(n_30612), .o(TIMEBOOST_net_2779) );
na02m02 TIMEBOOST_cell_8022 ( .a(n_16388), .b(n_16389), .o(TIMEBOOST_net_2642) );
in01s02 g770554 ( .a(n_10433), .o(n_10434) );
na02s06 g770555 ( .a(n_10287), .b(n_10398), .o(n_10433) );
na02m04 g770556 ( .a(FE_OCP_RBN3138_n_10326), .b(FE_OCPN1067_n_44461), .o(n_10397) );
na02f02 g770557 ( .a(n_10326), .b(FE_OCP_RBN5949_FE_OFN4772_n_44463), .o(n_10362) );
na02m04 g770558 ( .a(n_10193), .b(FE_OCP_RBN5906_n_44563), .o(n_10332) );
na02s02 g770559 ( .a(n_10192), .b(FE_OCP_RBN5934_n_44563), .o(n_10319) );
oa12f06 g770560 ( .a(n_10162), .b(n_10261), .c(n_10170), .o(n_10481) );
na02s01 g770561 ( .a(n_10278), .b(n_9121), .o(n_10279) );
no02s01 g770562 ( .a(FE_OCP_RBN3255_n_10454), .b(n_10523), .o(n_10640) );
na02s01 g770563 ( .a(n_10148), .b(FE_OCP_RBN2841_n_9044), .o(n_10337) );
na02s01 g770564 ( .a(n_10278), .b(n_9188), .o(n_10396) );
na02s01 g770565 ( .a(n_10194), .b(n_9041), .o(n_10282) );
na02s02 g770566 ( .a(n_10278), .b(n_9041), .o(n_10699) );
na02m08 g770570 ( .a(n_10102), .b(n_10016), .o(n_10277) );
in01f01 g770572 ( .a(n_10101), .o(n_10195) );
na02f06 g770573 ( .a(n_10021), .b(n_9974), .o(n_10101) );
in01s01 g770575 ( .a(n_10197), .o(n_10230) );
na02s01 g770577 ( .a(n_10431), .b(n_10430), .o(n_10432) );
in01s01 g770580 ( .a(n_10153), .o(n_10228) );
na02s03 g770581 ( .a(FE_OCP_DRV_N7077_n_10105), .b(n_10106), .o(n_10153) );
in01s01 g770584 ( .a(n_10280), .o(n_10360) );
na02m01 g770585 ( .a(FE_OCP_DRV_N7079_n_8992), .b(n_10148), .o(n_10280) );
na02s01 g770586 ( .a(n_10498), .b(n_10461), .o(n_10462) );
na02s01 g770587 ( .a(n_10148), .b(FE_OCP_RBN2869_n_9188), .o(n_10359) );
in01s01 g770588 ( .a(n_47263), .o(n_10276) );
na02m04 TIMEBOOST_cell_6708 ( .a(TIMEBOOST_net_2111), .b(n_47253), .o(n_13582) );
na02s01 g770593 ( .a(n_10194), .b(n_9146), .o(n_10329) );
no02f04 TIMEBOOST_cell_4057 ( .a(n_20446), .b(FE_OCP_RBN1840_n_20439), .o(TIMEBOOST_net_1119) );
in01s01 g770595 ( .a(FE_OCP_RBN3135_n_10274), .o(n_10293) );
oa12s01 g770600 ( .a(n_10426), .b(n_10425), .c(n_10424), .o(n_10490) );
ao12s01 g770601 ( .a(n_10429), .b(n_10428), .c(FE_OCP_RBN4252_n_8687), .o(n_10637) );
in01s01 g770602 ( .a(n_10411), .o(n_10394) );
no02f04 g770603 ( .a(n_10267), .b(n_10201), .o(n_10411) );
na02s01 g770604 ( .a(n_10148), .b(n_9204), .o(n_10357) );
na02s06 g770606 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_9_), .o(n_10458) );
in01m02 g770607 ( .a(n_10286), .o(n_10287) );
no02s04 g770609 ( .a(n_10270), .b(FE_OFN757_n_44464), .o(n_10286) );
na02s03 g770611 ( .a(n_10270), .b(n_44492), .o(n_10398) );
no02m04 g770612 ( .a(FE_OCP_RBN3114_n_10198), .b(FE_OCPN1064_n_44461), .o(n_10267) );
in01m02 g770613 ( .a(n_10338), .o(n_10339) );
na02m06 g770614 ( .a(n_10313), .b(n_10264), .o(n_10338) );
no02s02 g770615 ( .a(n_10198), .b(FE_OCP_RBN5936_n_44563), .o(n_10201) );
na02s06 g770616 ( .a(FE_OCP_RBN4253_n_8687), .b(n_10379), .o(n_10393) );
no02s01 g770617 ( .a(n_10428), .b(FE_OCP_RBN4252_n_8687), .o(n_10429) );
na02m06 g770619 ( .a(n_10410), .b(FE_OCP_RBN4222_n_8732), .o(n_10454) );
no02m02 g770620 ( .a(n_10355), .b(n_10310), .o(n_10356) );
na02s01 g770621 ( .a(n_10418), .b(n_10489), .o(n_10565) );
na02s02 g770622 ( .a(n_10022), .b(n_10065), .o(n_10150) );
no02s02 g770623 ( .a(n_10063), .b(n_10020), .o(n_10149) );
no02m06 g770624 ( .a(n_10410), .b(FE_OCP_RBN4222_n_8732), .o(n_10523) );
no02m02 TIMEBOOST_cell_6260 ( .a(TIMEBOOST_net_1981), .b(n_4941), .o(n_5110) );
na02s01 g770626 ( .a(n_10425), .b(n_10424), .o(n_10426) );
oa12f06 g770627 ( .a(n_10165), .b(n_10169), .c(n_10256), .o(n_10498) );
na02s01 g770628 ( .a(n_10423), .b(n_10350), .o(n_10560) );
no02s06 g770629 ( .a(n_10379), .b(FE_OCP_RBN4253_n_8687), .o(n_10380) );
in01s01 g770630 ( .a(n_10422), .o(n_10527) );
oa12m04 g770631 ( .a(n_9735), .b(n_10373), .c(n_9649), .o(n_10422) );
in01s02 g770632 ( .a(n_10474), .o(n_10421) );
in01s04 g770633 ( .a(n_10377), .o(n_10474) );
oa12m06 g770634 ( .a(n_10242), .b(n_10355), .c(n_10190), .o(n_10377) );
in01m04 g770635 ( .a(n_10354), .o(n_10435) );
in01f04 g770636 ( .a(n_10328), .o(n_10354) );
oa12f06 g770637 ( .a(n_10094), .b(n_10181), .c(n_10025), .o(n_10328) );
oa12s01 g770638 ( .a(n_10352), .b(n_10373), .c(n_10351), .o(n_10420) );
in01s01 g770644 ( .a(n_10148), .o(n_10278) );
in01s06 g770649 ( .a(n_10148), .o(n_10194) );
in01s08 g770650 ( .a(n_10106), .o(n_10148) );
no02m08 g770651 ( .a(n_9946), .b(n_9936), .o(n_10106) );
oa12f04 g770652 ( .a(n_9935), .b(n_9898), .c(FE_OCP_RBN5974_FE_RN_2033_0), .o(n_10021) );
na02m04 g770653 ( .a(n_10307), .b(n_10260), .o(n_10465) );
oa12f02 g770657 ( .a(FE_OCP_RBN5989_FE_RN_1865_0), .b(n_10068), .c(FE_OCP_RBN4349_n_9975), .o(n_10200) );
ao12f04 g770658 ( .a(FE_OCP_RBN5990_FE_RN_1865_0), .b(n_9975), .c(FE_OCP_RBN6003_n_10068), .o(n_10203) );
oa12s01 g770659 ( .a(n_10164), .b(n_10353), .c(n_10083), .o(n_10431) );
oa12s01 g770660 ( .a(n_10289), .b(n_10353), .c(n_10288), .o(n_10392) );
oa12f06 g770661 ( .a(n_9947), .b(n_10030), .c(FE_OCP_RBN5988_FE_RN_1865_0), .o(n_10102) );
in01s01 g770662 ( .a(n_10225), .o(n_11380) );
in01m02 g770665 ( .a(n_10192), .o(n_10193) );
in01s01 g770667 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_10_), .o(n_10419) );
na02s01 g770671 ( .a(n_10373), .b(n_10351), .o(n_10352) );
na02s02 g770672 ( .a(n_10057), .b(FE_OCP_RBN5934_n_44563), .o(n_10096) );
na02s08 g770673 ( .a(n_10109), .b(FE_OFN4775_n_44463), .o(n_10313) );
in01s02 g770674 ( .a(n_10310), .o(n_10311) );
na02s04 g770675 ( .a(n_10191), .b(n_10242), .o(n_10310) );
in01s01 g770676 ( .a(n_10264), .o(n_10265) );
na02s02 g770677 ( .a(n_10072), .b(FE_OFN757_n_44464), .o(n_10104) );
na02s04 g770678 ( .a(n_10072), .b(FE_OFN757_n_44464), .o(n_10264) );
in01s01 g770679 ( .a(n_10349), .o(n_10350) );
no02m04 g770680 ( .a(n_10309), .b(FE_OCP_RBN4218_n_8597), .o(n_10349) );
na02s02 g770681 ( .a(n_10145), .b(n_10186), .o(n_10263) );
no02s02 g770682 ( .a(n_10188), .b(n_10116), .o(n_10262) );
in01m02 g770683 ( .a(n_9982), .o(n_9983) );
na02m02 g770684 ( .a(n_9897), .b(n_9974), .o(n_9982) );
in01s01 g770686 ( .a(n_10020), .o(n_10065) );
no02m04 g770687 ( .a(n_9941), .b(FE_OCPN6283_FE_OCP_RBN2783_n_8664), .o(n_10020) );
no02f04 g770688 ( .a(n_9896), .b(n_9862), .o(n_9935) );
na02s01 g770689 ( .a(n_10353), .b(n_10288), .o(n_10289) );
in01s01 g770690 ( .a(n_10322), .o(n_10323) );
na02s01 g770691 ( .a(n_10241), .b(n_10185), .o(n_10322) );
na02s02 g770692 ( .a(n_10181), .b(n_10112), .o(n_10307) );
na02m04 g770693 ( .a(n_10375), .b(n_10374), .o(n_10489) );
in01s01 g770694 ( .a(n_10417), .o(n_10418) );
no02m06 g770695 ( .a(n_10375), .b(n_10374), .o(n_10417) );
na02m04 g770696 ( .a(n_10309), .b(FE_OCP_RBN4218_n_8597), .o(n_10423) );
no02m06 g770697 ( .a(n_9861), .b(n_9111), .o(n_9946) );
in01s01 g770699 ( .a(n_10022), .o(n_10063) );
na02m04 g770700 ( .a(n_9941), .b(FE_OCPN6283_FE_OCP_RBN2783_n_8664), .o(n_10022) );
no02f06 g770701 ( .a(n_10223), .b(n_10031), .o(n_10261) );
no02s04 g770702 ( .a(n_9860), .b(n_9173), .o(n_9936) );
na02m04 g770703 ( .a(n_10220), .b(n_10113), .o(n_10260) );
in01s01 g770704 ( .a(n_10390), .o(n_10391) );
no02s01 g770705 ( .a(n_10290), .b(n_10768), .o(n_10390) );
ao12f04 g770706 ( .a(FE_OCP_RBN5976_FE_RN_2033_0), .b(n_10017), .c(FE_OCP_RBN3068_n_9910), .o(n_10062) );
oa12m02 g770707 ( .a(FE_OCP_RBN5975_FE_RN_2033_0), .b(n_9910), .c(FE_OCP_RBN4347_n_10017), .o(n_10095) );
no02m06 g770708 ( .a(n_10098), .b(n_10061), .o(n_10270) );
no02s06 TIMEBOOST_cell_956 ( .a(TIMEBOOST_net_92), .b(n_23211), .o(n_23313) );
in01s01 g770712 ( .a(n_10379), .o(n_10428) );
na02s01 TIMEBOOST_cell_1278 ( .a(n_28926), .b(TIMEBOOST_net_253), .o(n_28992) );
oa12s01 g770714 ( .a(n_10204), .b(n_10334), .c(n_10125), .o(n_10425) );
oa12s01 g770715 ( .a(n_10303), .b(n_10334), .c(n_10302), .o(n_10389) );
na02m06 g770716 ( .a(n_10258), .b(n_10259), .o(n_10410) );
in01s01 g770717 ( .a(n_10415), .o(n_10416) );
na02s01 g770718 ( .a(n_10245), .b(n_10304), .o(n_10415) );
in01s01 g770719 ( .a(n_10305), .o(n_10306) );
oa22s01 g770720 ( .a(FE_OCP_RBN3052_n_10100), .b(n_8865), .c(FE_OCP_RBN4357_n_10100), .d(n_8908), .o(n_10305) );
in01s01 g770721 ( .a(n_10456), .o(n_10457) );
oa22s01 g770722 ( .a(FE_OCP_RBN4359_n_10100), .b(n_9197), .c(FE_OCP_RBN3052_n_10100), .d(n_9114), .o(n_10456) );
in01s01 g770723 ( .a(n_10521), .o(n_10522) );
no02s06 TIMEBOOST_cell_3296 ( .a(n_10573), .b(n_8865), .o(TIMEBOOST_net_939) );
in01s01 g770725 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_5_), .o(n_10371) );
no02f10 TIMEBOOST_cell_3842 ( .a(n_244), .b(TIMEBOOST_net_1011), .o(n_258) );
na02m04 g770728 ( .a(n_10179), .b(n_10177), .o(n_10259) );
na02s04 g770729 ( .a(n_10180), .b(n_10176), .o(n_10258) );
no02s06 g770730 ( .a(n_10142), .b(n_9965), .o(n_10236) );
na02s01 TIMEBOOST_cell_1277 ( .a(n_28991), .b(n_28925), .o(TIMEBOOST_net_253) );
no02m02 g770732 ( .a(n_10015), .b(FE_OCP_RBN5931_n_44563), .o(n_10061) );
na02s06 g770733 ( .a(n_10146), .b(FE_OCP_RBN5906_n_44563), .o(n_10242) );
in01s02 g770734 ( .a(n_10112), .o(n_10113) );
na02s04 g770735 ( .a(FE_OCP_RBN3112_n_10025), .b(n_10094), .o(n_10112) );
in01s02 g770736 ( .a(n_10190), .o(n_10191) );
no02s06 g770737 ( .a(n_10146), .b(FE_OCP_RBN5912_n_44563), .o(n_10190) );
no02m04 g770738 ( .a(FE_OCP_RBN6002_n_10015), .b(FE_OCPN1064_n_44461), .o(n_10098) );
na02s02 g770739 ( .a(FE_OCP_RBN5975_FE_RN_2033_0), .b(n_10017), .o(n_10019) );
no02s02 g770740 ( .a(FE_OCP_RBN5974_FE_RN_2033_0), .b(FE_OCP_RBN4347_n_10017), .o(n_10060) );
in01s01 g770742 ( .a(n_10145), .o(n_10188) );
na02m03 g770743 ( .a(n_10100), .b(FE_OCP_RBN2776_n_8637), .o(n_10145) );
na02m02 g770744 ( .a(n_9819), .b(FE_OCP_RBN2779_n_8599), .o(n_9974) );
in01s01 g770746 ( .a(n_10116), .o(n_10186) );
no02s04 g770747 ( .a(n_10100), .b(FE_OCP_RBN2776_n_8637), .o(n_10116) );
no02s01 g770748 ( .a(FE_OCP_RBN3052_n_10100), .b(FE_OCPN1092_n_9014), .o(n_10768) );
na02s01 g770749 ( .a(FE_OCP_RBN3052_n_10100), .b(FE_OCP_RBN2790_n_8767), .o(n_10241) );
na02s01 g770750 ( .a(FE_OCP_RBN4357_n_10100), .b(n_10183), .o(n_10185) );
na02s01 g770751 ( .a(FE_OCP_RBN4357_n_10100), .b(n_10183), .o(n_10592) );
no02s04 TIMEBOOST_cell_955 ( .a(FE_RN_65_0), .b(n_23390), .o(TIMEBOOST_net_92) );
in01s01 g770753 ( .a(n_9896), .o(n_9897) );
no02f04 g770754 ( .a(n_9819), .b(FE_OCP_RBN2779_n_8599), .o(n_9896) );
no03f08 TIMEBOOST_cell_8401 ( .a(TIMEBOOST_net_1285), .b(n_30497), .c(n_30142), .o(n_30598) );
na02s01 g770756 ( .a(FE_OCP_RBN3057_n_10100), .b(n_9148), .o(n_10304) );
na02s01 g770757 ( .a(FE_OCP_RBN4356_n_10100), .b(n_9162), .o(n_10245) );
no02s01 g770758 ( .a(n_10175), .b(n_10257), .o(n_10461) );
no02f06 g770759 ( .a(n_10212), .b(n_10067), .o(n_10256) );
no02m08 TIMEBOOST_cell_7044 ( .a(TIMEBOOST_net_2280), .b(TIMEBOOST_net_894), .o(n_39635) );
no02s01 g770761 ( .a(n_10252), .b(n_10342), .o(n_10471) );
no02s01 TIMEBOOST_cell_4523 ( .a(FE_OCP_RBN6173_n_16923), .b(n_17139), .o(TIMEBOOST_net_1352) );
in01s01 g770764 ( .a(n_10290), .o(n_10347) );
no02s01 g770765 ( .a(FE_OCP_RBN4356_n_10100), .b(FE_OCP_RBN5813_n_9014), .o(n_10290) );
na02s01 g770766 ( .a(n_10334), .b(n_10302), .o(n_10303) );
oa12m06 g770767 ( .a(n_9601), .b(n_10255), .c(n_9695), .o(n_10373) );
in01s01 g770768 ( .a(n_10355), .o(n_10254) );
oa12s01 g770770 ( .a(n_10238), .b(n_10255), .c(n_10237), .o(n_10301) );
oa12s01 g770771 ( .a(n_10219), .b(n_10218), .c(n_10217), .o(n_10295) );
na02s04 TIMEBOOST_cell_1222 ( .a(TIMEBOOST_net_225), .b(n_33852), .o(n_33903) );
in01f02 g770776 ( .a(n_10030), .o(n_10068) );
no02f04 TIMEBOOST_cell_8653 ( .a(TIMEBOOST_net_2813), .b(n_16567), .o(TIMEBOOST_net_1737) );
in01m04 g770780 ( .a(n_10072), .o(n_10109) );
in01m04 g770781 ( .a(n_10057), .o(n_10072) );
oa22m04 g770782 ( .a(FE_OCP_RBN5931_n_44563), .b(n_9859), .c(FE_OCP_RBN3062_n_9859), .d(FE_OCP_RBN5910_n_44563), .o(n_10057) );
in01s01 g770784 ( .a(n_10223), .o(n_10353) );
oa12f04 g770785 ( .a(n_10034), .b(n_10182), .c(n_9959), .o(n_10223) );
in01m02 g770786 ( .a(n_9860), .o(n_9861) );
oa12m04 g770787 ( .a(n_9422), .b(n_9855), .c(n_9420), .o(n_9860) );
oa12s01 g770788 ( .a(n_10140), .b(n_10182), .c(n_10139), .o(n_10222) );
no02s04 TIMEBOOST_cell_7007 ( .a(n_10518), .b(n_10363), .o(TIMEBOOST_net_2262) );
no02s02 TIMEBOOST_cell_8067 ( .a(TIMEBOOST_net_2664), .b(n_6373), .o(n_6418) );
na02s01 g770794 ( .a(FE_OCP_RBN3052_n_10100), .b(n_9260), .o(n_10300) );
in01s01 g770796 ( .a(n_10181), .o(n_10220) );
oa12m06 g770797 ( .a(n_9869), .b(n_10071), .c(n_9909), .o(n_10181) );
in01s06 g770798 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_), .o(n_10387) );
in01s01 g770800 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_4_), .o(n_12127) );
na02s01 g770802 ( .a(n_10218), .b(n_10217), .o(n_10219) );
na02s01 g770803 ( .a(n_10255), .b(n_10237), .o(n_10238) );
in01s02 g770804 ( .a(n_10179), .o(n_10180) );
no02m02 g770805 ( .a(n_10111), .b(n_10092), .o(n_10179) );
na02s01 TIMEBOOST_cell_1221 ( .a(n_33851), .b(n_33366), .o(TIMEBOOST_net_225) );
no02m06 g770809 ( .a(FE_OCP_RBN3172_n_10134), .b(n_10053), .o(n_10216) );
in01m02 g770810 ( .a(n_10141), .o(n_10142) );
na02s03 g770811 ( .a(n_10071), .b(n_9854), .o(n_10141) );
in01s02 g770812 ( .a(n_10176), .o(n_10177) );
na02s04 g770813 ( .a(n_10051), .b(n_10107), .o(n_10176) );
no02m04 g770815 ( .a(n_9944), .b(FE_OFN757_n_44464), .o(n_10025) );
na02m04 g770816 ( .a(n_9944), .b(FE_OCP_RBN5905_n_44563), .o(n_10094) );
no02m04 g770817 ( .a(n_9908), .b(n_9928), .o(n_9934) );
na02f04 TIMEBOOST_cell_5471 ( .a(TIMEBOOST_net_1683), .b(n_39616), .o(n_39643) );
in01s01 g770819 ( .a(n_10251), .o(n_10252) );
na02m04 g770820 ( .a(n_10215), .b(FE_OCP_RBN4216_FE_OCPN3565_n_10214), .o(n_10251) );
no02m06 g770821 ( .a(n_10215), .b(FE_OCP_RBN4216_FE_OCPN3565_n_10214), .o(n_10342) );
in01m02 g770823 ( .a(n_9862), .o(n_10017) );
no02f02 g770824 ( .a(n_9809), .b(FE_OCP_RBN6684_FE_OCPN4529_FE_OCP_RBN2748_n_8474), .o(n_9862) );
in01s01 g770825 ( .a(n_10174), .o(n_10175) );
na02m03 g770826 ( .a(n_10138), .b(n_10137), .o(n_10174) );
in01s02 g770827 ( .a(n_10032), .o(n_10033) );
na02s02 g770828 ( .a(n_9931), .b(n_10016), .o(n_10032) );
no02m04 g770829 ( .a(n_9808), .b(n_9749), .o(n_9867) );
na02s02 g770834 ( .a(n_10010), .b(n_9942), .o(n_10090) );
no02s02 g770835 ( .a(n_9978), .b(n_10008), .o(n_10089) );
na02s01 g770836 ( .a(n_10182), .b(n_10139), .o(n_10140) );
no02s06 g770837 ( .a(n_9930), .b(n_47260), .o(n_9947) );
no02m04 g770838 ( .a(n_10138), .b(n_10137), .o(n_10257) );
no02s02 TIMEBOOST_cell_4954 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .b(n_33242), .o(TIMEBOOST_net_1425) );
in01f01 g770840 ( .a(n_9970), .o(n_9971) );
na02f01 g770841 ( .a(n_9908), .b(n_9741), .o(n_9970) );
na02s02 TIMEBOOST_cell_3346 ( .a(n_36271), .b(n_36307), .o(TIMEBOOST_net_964) );
oa12s01 g770843 ( .a(n_10133), .b(n_10132), .c(n_10171), .o(n_10213) );
na02m10 g770862 ( .a(n_9932), .b(n_9866), .o(n_10100) );
in01m02 g770868 ( .a(n_9898), .o(n_9910) );
no02s06 g770869 ( .a(n_9755), .b(n_9727), .o(n_9898) );
in01s01 g770870 ( .a(n_10212), .o(n_10334) );
ao12f04 g770871 ( .a(n_9919), .b(n_10171), .c(n_9999), .o(n_10212) );
no02f02 TIMEBOOST_cell_6385 ( .a(n_26327), .b(n_26208), .o(TIMEBOOST_net_2044) );
na02s06 g770874 ( .a(n_9851), .b(n_9676), .o(n_9866) );
na02m08 g770875 ( .a(n_9852), .b(FE_OCP_RBN2971_n_9676), .o(n_9932) );
no02m06 g770877 ( .a(n_10007), .b(n_9744), .o(n_10134) );
na02m04 g770878 ( .a(n_9968), .b(n_9716), .o(n_10092) );
no02f04 g770879 ( .a(n_10006), .b(n_9899), .o(n_10111) );
no02m06 g770880 ( .a(n_9853), .b(n_9868), .o(n_9869) );
in01m02 g770881 ( .a(n_10053), .o(n_10054) );
na02m04 g770882 ( .a(n_9968), .b(n_9900), .o(n_10053) );
no02s02 g770883 ( .a(n_10013), .b(FE_OCP_RBN3030_n_9624), .o(n_10014) );
na02s01 TIMEBOOST_cell_3345 ( .a(TIMEBOOST_net_963), .b(n_26978), .o(n_27033) );
no02m02 g770885 ( .a(n_9892), .b(FE_OCP_RBN5906_n_44563), .o(n_9937) );
na02m04 TIMEBOOST_cell_3279 ( .a(TIMEBOOST_net_930), .b(FE_RN_1234_0), .o(n_21118) );
na02f06 g770887 ( .a(n_10013), .b(n_9820), .o(n_10071) );
in01s02 g770888 ( .a(n_10050), .o(n_10051) );
no02m04 g770889 ( .a(n_9992), .b(FE_OCP_RBN5913_n_44563), .o(n_10050) );
na02m04 g770890 ( .a(n_9992), .b(FE_OCP_RBN5913_n_44563), .o(n_10107) );
in01s02 g770891 ( .a(n_9965), .o(n_9966) );
no02s04 g770892 ( .a(n_9868), .b(n_9909), .o(n_9965) );
no02s01 g770893 ( .a(n_10128), .b(n_10163), .o(n_10430) );
na02m02 g770894 ( .a(FE_OCPN1086_n_8499), .b(n_9864), .o(n_10016) );
na02m06 g770895 ( .a(n_10127), .b(n_10027), .o(n_10170) );
na02f04 g770896 ( .a(n_9762), .b(n_9740), .o(n_9908) );
in01s01 g770898 ( .a(n_9978), .o(n_10010) );
no02s03 g770899 ( .a(n_9904), .b(n_8562), .o(n_9978) );
in01f02 g770900 ( .a(n_9807), .o(n_9808) );
na02f02 g770901 ( .a(n_9723), .b(n_9674), .o(n_9807) );
no02s06 g770902 ( .a(n_9723), .b(n_9726), .o(n_9755) );
in01s01 g770904 ( .a(n_9942), .o(n_10008) );
na02m03 g770905 ( .a(n_9904), .b(n_8562), .o(n_9942) );
na02s01 g770906 ( .a(n_10132), .b(n_10171), .o(n_10133) );
in01s01 g770907 ( .a(n_9930), .o(n_9931) );
no02m04 g770908 ( .a(n_9864), .b(FE_OCPN1086_n_8499), .o(n_9930) );
na02f04 g770909 ( .a(n_10129), .b(n_10070), .o(n_10169) );
no02s01 g770910 ( .a(n_10166), .b(n_10130), .o(n_10424) );
in01s01 g770911 ( .a(n_9855), .o(n_9754) );
ao12m06 g770913 ( .a(n_9481), .b(n_10131), .c(n_9548), .o(n_10255) );
ao12s01 g770914 ( .a(n_9434), .b(n_10131), .c(n_9505), .o(n_10218) );
oa12s01 g770915 ( .a(n_10087), .b(n_10131), .c(n_10086), .o(n_10168) );
ao22f02 g770916 ( .a(n_9890), .b(n_9745), .c(n_9901), .d(n_9746), .o(n_10138) );
na02m06 g770917 ( .a(n_9991), .b(n_10048), .o(n_10215) );
oa12s01 g770918 ( .a(n_10005), .b(n_10049), .c(n_10004), .o(n_10088) );
no02f02 g770920 ( .a(n_9675), .b(n_9671), .o(n_9809) );
oa12f04 g770921 ( .a(n_9838), .b(n_10049), .c(n_9918), .o(n_10182) );
in01s01 g770922 ( .a(FE_OCP_RBN3063_n_9859), .o(n_11292) );
no02s08 TIMEBOOST_cell_3148 ( .a(FE_OCP_RBN3102_n_15768), .b(n_15524), .o(TIMEBOOST_net_865) );
in01s06 g770926 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_), .o(n_10167) );
na02s01 TIMEBOOST_cell_4177 ( .a(n_35782), .b(n_35587), .o(TIMEBOOST_net_1179) );
no02s02 g770930 ( .a(n_9580), .b(n_9456), .o(n_9671) );
na02s01 g770931 ( .a(n_10131), .b(n_10086), .o(n_10087) );
in01s02 g770932 ( .a(n_9853), .o(n_9854) );
na02m06 g770933 ( .a(n_9806), .b(n_9624), .o(n_9853) );
na02m04 g770934 ( .a(n_9979), .b(n_9850), .o(n_9991) );
na02m04 g770935 ( .a(n_9980), .b(n_9849), .o(n_10048) );
in01m02 g770936 ( .a(n_10006), .o(n_10007) );
na02f06 g770937 ( .a(n_9926), .b(n_9804), .o(n_10006) );
in01s01 g770938 ( .a(n_10013), .o(n_9964) );
no02f06 g770939 ( .a(n_9890), .b(n_9685), .o(n_10013) );
na02m04 g770940 ( .a(n_9895), .b(FE_OCP_RBN5930_n_44563), .o(n_9968) );
no02m04 g770941 ( .a(n_9747), .b(FE_OCP_RBN5905_n_44563), .o(n_9868) );
in01s02 g770942 ( .a(n_9899), .o(n_9900) );
no02m04 g770943 ( .a(FE_OCP_RBN6731_n_44579), .b(n_9895), .o(n_9899) );
no02f04 TIMEBOOST_cell_4406 ( .a(TIMEBOOST_net_1293), .b(n_25997), .o(TIMEBOOST_net_1107) );
na02s04 g770946 ( .a(n_9806), .b(n_9820), .o(n_9893) );
no02m06 g770947 ( .a(FE_OCP_RBN5930_n_44563), .b(n_9748), .o(n_9909) );
na02s08 TIMEBOOST_cell_3147 ( .a(TIMEBOOST_net_864), .b(n_15768), .o(n_15908) );
na02s01 g770949 ( .a(n_10049), .b(n_10004), .o(n_10005) );
in01s01 g770950 ( .a(n_10165), .o(n_10166) );
na02s06 g770951 ( .a(n_10043), .b(n_8427), .o(n_10165) );
na02s01 g770952 ( .a(n_10027), .b(n_10164), .o(n_10288) );
in01s01 g770953 ( .a(n_10162), .o(n_10163) );
na02m06 g770954 ( .a(n_10041), .b(n_8429), .o(n_10162) );
na02s02 g770955 ( .a(FE_OCP_RBN5989_FE_RN_1865_0), .b(n_9975), .o(n_9987) );
no02s02 g770956 ( .a(FE_OCP_RBN4350_n_9975), .b(FE_OCP_RBN5988_FE_RN_1865_0), .o(n_10047) );
in01s01 g770957 ( .a(n_10129), .o(n_10130) );
na02f02 g770958 ( .a(n_10042), .b(n_8426), .o(n_10129) );
in01s01 g770959 ( .a(n_10127), .o(n_10128) );
na02m04 g770960 ( .a(n_10040), .b(n_8428), .o(n_10127) );
na02f06 g770961 ( .a(n_9625), .b(n_9670), .o(n_9723) );
in01m04 g770963 ( .a(n_9851), .o(n_9852) );
oa12m06 g770964 ( .a(n_9594), .b(n_9571), .c(n_9764), .o(n_9851) );
na02m04 g770966 ( .a(n_9541), .b(n_9579), .o(n_9626) );
no02m02 g770967 ( .a(n_9463), .b(n_9582), .o(n_9583) );
no02f08 TIMEBOOST_cell_5989 ( .a(FE_OCP_RBN2479_n_47245), .b(FE_OCPN1687_n_23097), .o(TIMEBOOST_net_1846) );
no02s01 TIMEBOOST_cell_4479 ( .a(n_23259), .b(FE_OFN748_n_22641), .o(TIMEBOOST_net_1330) );
oa12s01 g770971 ( .a(n_10003), .b(n_10045), .c(n_10002), .o(n_10085) );
oa12f04 g770973 ( .a(n_9836), .b(n_10045), .c(n_9905), .o(n_10171) );
in01f01 g770975 ( .a(n_9762), .o(n_9856) );
ao12m04 g770976 ( .a(n_9555), .b(n_9637), .c(n_9659), .o(n_9762) );
no02s06 TIMEBOOST_cell_5980 ( .a(TIMEBOOST_net_1841), .b(n_18069), .o(n_18160) );
in01s01 g770981 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_3_), .o(n_12061) );
na02m04 g770983 ( .a(n_9503), .b(n_9363), .o(n_9507) );
na02f06 TIMEBOOST_cell_4176 ( .a(n_36632), .b(TIMEBOOST_net_1178), .o(TIMEBOOST_net_996) );
na02s02 g770985 ( .a(n_9579), .b(n_9465), .o(n_9580) );
na02s04 g770986 ( .a(FE_OCP_RBN5920_n_9456), .b(n_9465), .o(n_9541) );
no02s02 g770987 ( .a(n_9461), .b(n_9456), .o(n_9463) );
in01s02 g770988 ( .a(n_9550), .o(n_9551) );
na02m02 g770989 ( .a(n_9503), .b(n_9504), .o(n_9550) );
in01s02 g770990 ( .a(n_9849), .o(n_9850) );
na02m04 g770991 ( .a(n_9804), .b(n_9743), .o(n_9849) );
no03s01 TIMEBOOST_cell_7508 ( .a(n_1940), .b(n_2343), .c(n_1687), .o(TIMEBOOST_net_2385) );
na02m06 g770993 ( .a(n_9666), .b(FE_OCP_RBN5930_n_44563), .o(n_9806) );
na02m08 g770994 ( .a(FE_OCP_RBN5907_n_44563), .b(n_9667), .o(n_9820) );
na02s04 TIMEBOOST_cell_5425 ( .a(TIMEBOOST_net_1660), .b(n_5045), .o(n_5215) );
in01s01 g770996 ( .a(n_10031), .o(n_10164) );
no02s04 g770997 ( .a(n_9989), .b(n_9988), .o(n_10031) );
na02m02 g770998 ( .a(n_9888), .b(n_9845), .o(n_9927) );
no02s02 g770999 ( .a(n_9928), .b(n_9763), .o(n_9963) );
no02f08 TIMEBOOST_cell_6702 ( .a(TIMEBOOST_net_2108), .b(n_14864), .o(n_14988) );
na02s01 g771004 ( .a(n_10045), .b(n_10002), .o(n_10003) );
na02s01 g771005 ( .a(n_9960), .b(n_10034), .o(n_10139) );
na02s01 g771006 ( .a(n_10070), .b(n_10204), .o(n_10302) );
na02s01 TIMEBOOST_cell_3269 ( .a(TIMEBOOST_net_925), .b(n_31815), .o(n_31939) );
in01s02 g771008 ( .a(n_47260), .o(n_9975) );
in01s02 g771014 ( .a(n_9749), .o(n_9750) );
no02m02 g771015 ( .a(n_9726), .b(n_9672), .o(n_9749) );
in01s01 g771017 ( .a(n_10027), .o(n_10083) );
na02m04 g771018 ( .a(n_9989), .b(n_9988), .o(n_10027) );
in01s01 g771020 ( .a(n_9890), .o(n_9901) );
oa12f04 g771021 ( .a(n_9593), .b(n_9703), .c(n_9542), .o(n_9890) );
ao12m06 g771022 ( .a(n_9596), .b(n_10001), .c(n_9516), .o(n_10131) );
in01s02 g771023 ( .a(n_9979), .o(n_9980) );
in01m02 g771024 ( .a(n_9926), .o(n_9979) );
oa12s01 g771026 ( .a(n_9962), .b(n_10001), .c(n_9961), .o(n_10044) );
oa12s01 g771027 ( .a(n_9925), .b(n_9924), .c(n_9923), .o(n_10000) );
in01s02 g771028 ( .a(n_10042), .o(n_10043) );
ao22f02 g771029 ( .a(n_9883), .b(n_9665), .c(n_9831), .d(n_9664), .o(n_10042) );
na02m06 g771030 ( .a(n_9644), .b(n_9717), .o(n_9895) );
in01s02 g771031 ( .a(n_10040), .o(n_10041) );
no02s02 TIMEBOOST_cell_8866 ( .a(n_25753), .b(FE_OCP_RBN2977_n_25509), .o(TIMEBOOST_net_2920) );
ao12f04 g771033 ( .a(n_9787), .b(n_9822), .c(n_9698), .o(n_10049) );
ao22m02 g771036 ( .a(FE_OCP_RBN6792_n_9510), .b(n_9413), .c(n_9510), .d(FE_OCP_RBN2992_n_9413), .o(n_9682) );
in01m01 g771038 ( .a(n_9625), .o(n_9668) );
ao12f06 g771039 ( .a(n_9366), .b(n_9496), .c(n_9213), .o(n_9625) );
in01s02 g771040 ( .a(n_9747), .o(n_9748) );
in01s02 g771043 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_6_), .o(n_10035) );
na02m06 g771050 ( .a(n_9362), .b(FE_OCP_RBN5880_FE_RN_314_0), .o(n_9456) );
no02s02 g771051 ( .a(n_9419), .b(n_8362), .o(n_9420) );
na02s04 g771052 ( .a(n_9360), .b(n_8362), .o(n_9504) );
no02s06 g771054 ( .a(n_9417), .b(n_8362), .o(n_9582) );
na02s02 g771055 ( .a(n_9359), .b(n_8232), .o(n_9579) );
in01m06 g771058 ( .a(n_9461), .o(n_9465) );
no02m08 g771060 ( .a(n_9359), .b(n_8232), .o(n_9461) );
na02s02 g771061 ( .a(n_9419), .b(n_8362), .o(n_9422) );
na02s01 g771062 ( .a(n_10001), .b(n_9961), .o(n_9962) );
na02s04 g771063 ( .a(n_9621), .b(FE_OCP_RBN6738_n_44563), .o(n_9804) );
na02m04 g771064 ( .a(FE_OCP_RBN3033_n_9629), .b(FE_OCP_RBN6738_n_44563), .o(n_9717) );
na02s03 g771065 ( .a(n_9629), .b(FE_OCP_RBN6731_n_44579), .o(n_9644) );
in01m02 g771066 ( .a(n_9745), .o(n_9746) );
no02m04 g771067 ( .a(FE_OCP_RBN3031_n_9624), .b(n_9685), .o(n_9745) );
in01s02 g771068 ( .a(n_9743), .o(n_9744) );
na02s02 g771069 ( .a(FE_OCP_RBN3045_n_9621), .b(FE_OCP_RBN6731_n_44579), .o(n_9716) );
na02s04 g771070 ( .a(FE_OCP_RBN3045_n_9621), .b(FE_OCP_RBN5930_n_44563), .o(n_9743) );
in01s02 g771071 ( .a(n_9800), .o(n_9801) );
na02s02 g771072 ( .a(n_9741), .b(n_9740), .o(n_9800) );
in01s01 g771074 ( .a(n_9928), .o(n_9888) );
in01s01 g771076 ( .a(n_10067), .o(n_10204) );
no02f02 g771077 ( .a(n_10029), .b(n_10028), .o(n_10067) );
na02s02 TIMEBOOST_cell_4125 ( .a(n_10855), .b(n_10457), .o(TIMEBOOST_net_1153) );
na02m02 g771079 ( .a(n_9907), .b(n_9906), .o(n_10034) );
in01s01 g771080 ( .a(n_9959), .o(n_9960) );
no02m02 g771081 ( .a(n_9907), .b(n_9906), .o(n_9959) );
in01s01 g771083 ( .a(n_9763), .o(n_9845) );
no02s02 g771084 ( .a(n_9704), .b(FE_OCP_RBN6679_n_8288), .o(n_9763) );
in01s01 g771086 ( .a(n_10070), .o(n_10125) );
na02f02 g771087 ( .a(n_10029), .b(n_10028), .o(n_10070) );
na02s01 g771088 ( .a(n_9924), .b(n_9923), .o(n_9925) );
in01s02 g771089 ( .a(n_9718), .o(n_9719) );
na02s02 g771090 ( .a(n_9674), .b(n_9670), .o(n_9718) );
no02m08 TIMEBOOST_cell_7547 ( .a(TIMEBOOST_net_2404), .b(n_13750), .o(n_13918) );
no02m06 g771092 ( .a(n_9515), .b(FE_OCP_RBN5738_n_8402), .o(n_9726) );
no02m02 g771093 ( .a(n_9514), .b(FE_OCP_RBN2737_n_8402), .o(n_9672) );
na02s01 g771094 ( .a(n_9843), .b(n_9999), .o(n_10132) );
oa12s02 g771095 ( .a(n_9492), .b(n_9553), .c(n_9552), .o(n_9628) );
no02m04 g771096 ( .a(n_9554), .b(FE_OCP_RBN2888_n_9492), .o(n_9638) );
ao12f04 g771097 ( .a(n_9721), .b(n_9921), .c(n_9786), .o(n_10045) );
in01m04 g771098 ( .a(n_9666), .o(n_9667) );
in01s02 g771100 ( .a(n_9713), .o(n_9714) );
in01m01 g771101 ( .a(n_9637), .o(n_9713) );
ao12m06 g771102 ( .a(n_9402), .b(n_9502), .c(n_9486), .o(n_9637) );
in01m01 g771103 ( .a(n_9764), .o(n_9712) );
oa12s01 g771105 ( .a(n_9886), .b(n_9885), .c(n_9921), .o(n_9958) );
na02m04 g771110 ( .a(n_9844), .b(n_9795), .o(n_9989) );
in01s06 g771114 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_1_), .o(n_11871) );
in01m01 g771117 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_1_), .o(n_11879) );
na02s04 TIMEBOOST_cell_5684 ( .a(FE_OCPN1950_delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n_36566), .o(TIMEBOOST_net_1790) );
no02m02 g771120 ( .a(n_9553), .b(n_9552), .o(n_9554) );
na02s06 g771124 ( .a(n_9570), .b(n_9594), .o(n_9676) );
na02f04 g771125 ( .a(n_47259), .b(n_9447), .o(n_9542) );
na02m02 g771126 ( .a(n_9618), .b(n_9757), .o(n_9795) );
na02m02 g771127 ( .a(n_9758), .b(n_9617), .o(n_9844) );
no02m04 g771128 ( .a(n_9546), .b(FE_OCP_RBN5930_n_44563), .o(n_9685) );
na02m06 g771132 ( .a(n_9546), .b(FE_OCP_RBN6731_n_44579), .o(n_9624) );
in01m01 g771133 ( .a(n_9706), .o(n_9707) );
na02m02 g771134 ( .a(n_9635), .b(FE_RN_319_0), .o(n_9706) );
in01m02 g771135 ( .a(n_9664), .o(n_9665) );
na02m02 g771136 ( .a(n_47259), .b(n_9593), .o(n_9664) );
na02s02 g771137 ( .a(n_9509), .b(FE_OCPN3568_n_8348), .o(n_9670) );
in01s01 g771138 ( .a(n_9663), .o(n_9741) );
no02m04 g771139 ( .a(n_9623), .b(FE_OCP_RBN2692_n_8221), .o(n_9663) );
na02m04 g771140 ( .a(n_9789), .b(n_8240), .o(n_9999) );
na02s02 g771141 ( .a(n_9623), .b(FE_OCP_RBN2692_n_8221), .o(n_9740) );
in01m01 g771142 ( .a(n_9578), .o(n_9674) );
no02m04 g771143 ( .a(FE_OCPN3568_n_8348), .b(n_9509), .o(n_9578) );
na02s01 g771144 ( .a(n_9885), .b(n_9921), .o(n_9886) );
in01s02 g771146 ( .a(n_9843), .o(n_9919) );
na02s02 g771147 ( .a(n_9788), .b(n_8239), .o(n_9843) );
no02s01 g771148 ( .a(n_9839), .b(n_9918), .o(n_10004) );
in01s02 g771152 ( .a(n_9362), .o(n_9363) );
ao12m06 g771154 ( .a(n_9385), .b(n_9884), .c(n_9475), .o(n_10001) );
ao12s02 g771155 ( .a(n_9446), .b(n_9639), .c(n_9447), .o(n_9831) );
no02f02 TIMEBOOST_cell_6991 ( .a(n_15041), .b(n_15098), .o(TIMEBOOST_net_2254) );
oa12s01 g771157 ( .a(n_9738), .b(n_9794), .c(n_9737), .o(n_9842) );
oa12s01 g771158 ( .a(n_9882), .b(n_9881), .c(n_9880), .o(n_9957) );
oa12s01 g771159 ( .a(n_9816), .b(n_9884), .c(n_9815), .o(n_9917) );
na02s02 TIMEBOOST_cell_5399 ( .a(TIMEBOOST_net_1647), .b(n_3948), .o(n_4126) );
na02m02 TIMEBOOST_cell_5108 ( .a(FE_RN_2021_0), .b(n_8870), .o(TIMEBOOST_net_1502) );
no02s04 TIMEBOOST_cell_4473 ( .a(FE_OCPN1942_n_20723), .b(n_22028), .o(TIMEBOOST_net_1327) );
in01s01 g771164 ( .a(FE_OCP_RBN3029_n_9584), .o(n_9620) );
ao22m04 g771167 ( .a(n_9374), .b(n_9291), .c(FE_OCP_RBN5941_n_9374), .d(n_9290), .o(n_9584) );
in01s01 g771168 ( .a(n_9840), .o(n_9841) );
in01f02 g771169 ( .a(n_9761), .o(n_9840) );
ao12f04 g771170 ( .a(n_9532), .b(n_9720), .c(n_9586), .o(n_9761) );
in01m02 g771175 ( .a(n_9514), .o(n_9515) );
no02m02 TIMEBOOST_cell_4381 ( .a(n_26162), .b(n_26163), .o(TIMEBOOST_net_1281) );
na02m02 g771178 ( .a(n_9572), .b(n_9538), .o(n_9704) );
in01s01 g771179 ( .a(n_9822), .o(n_9924) );
oa12m04 g771180 ( .a(n_9560), .b(n_9656), .c(n_9794), .o(n_9822) );
in01s01 g771182 ( .a(n_9496), .o(n_9510) );
ao12m06 g771183 ( .a(n_9135), .b(n_9212), .c(n_9354), .o(n_9496) );
na02m04 g771185 ( .a(n_9144), .b(n_9161), .o(n_9360) );
in01s02 g771187 ( .a(n_9359), .o(n_9417) );
no02m08 g771188 ( .a(n_9195), .b(n_9145), .o(n_9359) );
na02m08 TIMEBOOST_cell_2820 ( .a(FE_RN_633_0), .b(FE_RN_635_0), .o(TIMEBOOST_net_701) );
in01s06 g771190 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_4_), .o(n_11542) );
in01m04 g771192 ( .a(n_9573), .o(n_9574) );
in01m04 g771193 ( .a(n_9553), .o(n_9573) );
na02f06 g771194 ( .a(n_9495), .b(n_9351), .o(n_9553) );
na02m02 g771195 ( .a(n_9489), .b(n_9409), .o(n_9572) );
na02m02 g771197 ( .a(n_9452), .b(n_9408), .o(n_9538) );
no02m06 TIMEBOOST_cell_5217 ( .a(TIMEBOOST_net_1556), .b(n_24267), .o(n_24369) );
no02s03 g771199 ( .a(n_9091), .b(FE_OCP_DRV_N3506_n_8189), .o(n_9145) );
in01s02 g771200 ( .a(n_9570), .o(n_9571) );
na02s02 g771202 ( .a(n_9057), .b(n_8232), .o(n_9144) );
na02s06 g771203 ( .a(n_9450), .b(n_8362), .o(n_9594) );
na02s02 g771204 ( .a(n_9424), .b(FE_OCP_RBN5882_FE_RN_2220_0), .o(n_9543) );
no02s02 g771205 ( .a(n_9468), .b(FE_RN_2220_0), .o(n_9569) );
no02s02 g771206 ( .a(n_9552), .b(FE_OCP_RBN2889_n_9492), .o(n_9476) );
na02s02 g771207 ( .a(n_9492), .b(n_9415), .o(n_9493) );
na02s04 g771208 ( .a(n_9058), .b(FE_OCP_RBN4146_n_7743), .o(n_9161) );
no03m08 TIMEBOOST_cell_674 ( .a(n_6090), .b(n_6089), .c(n_6028), .o(n_6130) );
no02f04 TIMEBOOST_cell_8555 ( .a(TIMEBOOST_net_2764), .b(n_8285), .o(n_8454) );
no02m06 g771211 ( .a(n_9092), .b(FE_OFN4768_n_8309), .o(n_9195) );
na02m08 TIMEBOOST_cell_3962 ( .a(TIMEBOOST_net_1071), .b(FE_RN_1071_0), .o(n_24436) );
na02s01 g771213 ( .a(n_9881), .b(n_9880), .o(n_9882) );
na02s01 g771214 ( .a(n_9884), .b(n_9815), .o(n_9816) );
in01s02 g771215 ( .a(n_9757), .o(n_9758) );
no02s02 g771216 ( .a(n_9720), .b(n_9407), .o(n_9757) );
no02f02 g771218 ( .a(FE_OCP_RBN5835_n_44563), .b(n_9535), .o(n_9556) );
no02f04 g771219 ( .a(n_9639), .b(n_9446), .o(n_9703) );
no02s01 TIMEBOOST_cell_5448 ( .a(n_4875), .b(n_4759), .o(TIMEBOOST_net_1672) );
no02s02 g771221 ( .a(FE_OCP_RBN5842_n_44563), .b(n_9411), .o(n_9462) );
na02f02 g771224 ( .a(n_9535), .b(FE_OCP_RBN6730_n_44579), .o(n_9635) );
na02s01 TIMEBOOST_cell_6316 ( .a(TIMEBOOST_net_2009), .b(n_36385), .o(n_46953) );
na02s06 g771226 ( .a(FE_OCP_RBN6786_n_9410), .b(FE_OCP_RBN6733_n_44579), .o(n_9593) );
no02m06 TIMEBOOST_cell_6949 ( .a(FE_OCP_RBN2611_n_29298), .b(FE_RN_1099_0), .o(TIMEBOOST_net_2233) );
no02m04 g771228 ( .a(n_9791), .b(n_9790), .o(n_9918) );
no02s01 g771229 ( .a(n_9837), .b(n_9905), .o(n_10002) );
no02s02 TIMEBOOST_cell_8701 ( .a(TIMEBOOST_net_2837), .b(n_6759), .o(FE_RN_2132_0) );
na02s01 g771231 ( .a(n_9794), .b(n_9737), .o(n_9738) );
in01s01 g771232 ( .a(n_9838), .o(n_9839) );
na02s03 g771233 ( .a(n_9791), .b(n_9790), .o(n_9838) );
na02s01 g771234 ( .a(n_9162), .b(FE_OCP_RBN5813_n_9014), .o(n_9260) );
na02f04 TIMEBOOST_cell_8570 ( .a(n_186), .b(n_29854), .o(TIMEBOOST_net_2772) );
no02s04 TIMEBOOST_cell_5394 ( .a(FE_OCPN3573_n_30345), .b(FE_RN_1279_0), .o(TIMEBOOST_net_1645) );
na02s01 g771238 ( .a(n_9613), .b(n_9659), .o(n_9660) );
no02s01 g771239 ( .a(n_9568), .b(n_9555), .o(n_9701) );
in01s01 g771241 ( .a(n_9502), .o(n_9565) );
na02m08 g771242 ( .a(n_9356), .b(n_9397), .o(n_9502) );
oa12s01 g771243 ( .a(n_9835), .b(n_9834), .c(n_9833), .o(n_9916) );
in01m02 g771248 ( .a(n_9788), .o(n_9789) );
oa12s01 g771251 ( .a(n_9783), .b(n_9782), .c(n_9781), .o(n_9878) );
no02m04 g771252 ( .a(n_9314), .b(n_9298), .o(n_9509) );
no03m08 TIMEBOOST_cell_5883 ( .a(n_26725), .b(n_26332), .c(TIMEBOOST_net_1736), .o(n_26874) );
oa12s01 g771254 ( .a(n_9689), .b(n_9688), .c(n_9687), .o(n_9760) );
na02m06 g771255 ( .a(n_9371), .b(n_9302), .o(n_9546) );
na02m04 g771256 ( .a(n_9350), .b(n_9288), .o(n_9457) );
no02s01 TIMEBOOST_cell_4466 ( .a(n_43664), .b(TIMEBOOST_net_1323), .o(n_43744) );
no02s02 g771258 ( .a(n_9353), .b(n_9347), .o(n_9489) );
na02s02 g771259 ( .a(FE_OCP_RBN2866_n_9347), .b(n_9372), .o(n_9452) );
na02f06 g771260 ( .a(n_9353), .b(n_9318), .o(n_9495) );
in01s01 g771261 ( .a(n_9552), .o(n_9415) );
no02m06 g771262 ( .a(n_9313), .b(n_8232), .o(n_9552) );
na02s06 g771267 ( .a(n_9313), .b(n_8232), .o(n_9492) );
no02f04 TIMEBOOST_cell_8116 ( .a(n_20722), .b(FE_OCP_RBN5386_n_20638), .o(TIMEBOOST_net_2689) );
in01s01 g771270 ( .a(n_9424), .o(n_9468) );
na02m04 g771271 ( .a(n_9342), .b(FE_OFN4771_n_8309), .o(n_9424) );
na02s04 g771272 ( .a(n_9194), .b(FE_OCP_RBN4235_n_9089), .o(n_9299) );
na02f04 TIMEBOOST_cell_8168 ( .a(n_21116), .b(n_21063), .o(TIMEBOOST_net_2715) );
no02m02 g771274 ( .a(n_9150), .b(n_9050), .o(n_9298) );
na02f02 g771275 ( .a(n_9531), .b(n_9406), .o(n_9532) );
in01s02 g771276 ( .a(n_9657), .o(n_9658) );
na02m02 g771277 ( .a(n_9588), .b(n_9379), .o(n_9657) );
na02m02 g771278 ( .a(n_9292), .b(FE_OCPN880_n_44593), .o(n_9302) );
no02m04 g771279 ( .a(n_9588), .b(n_9341), .o(n_9720) );
in01s02 g771280 ( .a(n_9617), .o(n_9618) );
na02s02 g771281 ( .a(n_9531), .b(n_9586), .o(n_9617) );
in01m02 g771282 ( .a(n_9615), .o(n_9616) );
na02m04 g771283 ( .a(n_9447), .b(n_9464), .o(n_9615) );
na02m04 g771284 ( .a(FE_OCP_RBN4317_n_9292), .b(n_44594), .o(n_9371) );
no02s01 g771285 ( .a(n_9787), .b(n_9699), .o(n_9923) );
na02s01 g771286 ( .a(n_9688), .b(n_9687), .o(n_9689) );
na02s01 g771287 ( .a(n_9786), .b(n_9722), .o(n_9885) );
in01s01 g771288 ( .a(n_9836), .o(n_9837) );
na02s03 g771289 ( .a(n_9785), .b(n_9784), .o(n_9836) );
na02s01 g771290 ( .a(n_9834), .b(n_9833), .o(n_9835) );
in01s01 g771291 ( .a(n_9659), .o(n_9568) );
na02m04 g771292 ( .a(FE_OCPN1208_n_8185), .b(n_9513), .o(n_9659) );
in01s01 g771294 ( .a(n_9555), .o(n_9613) );
no02m04 g771295 ( .a(n_9513), .b(FE_OCPN1208_n_8185), .o(n_9555) );
no02s02 g771297 ( .a(n_9214), .b(n_9366), .o(n_9413) );
na02s02 g771298 ( .a(n_9266), .b(n_9108), .o(n_9297) );
no02s04 g771299 ( .a(n_9267), .b(n_9051), .o(n_9357) );
no02m04 g771301 ( .a(n_9785), .b(n_9784), .o(n_9905) );
na02m06 g771302 ( .a(n_9152), .b(n_9355), .o(n_9356) );
na02s01 g771303 ( .a(n_9782), .b(n_9781), .o(n_9783) );
oa12m06 g771304 ( .a(n_9310), .b(n_9654), .c(n_9311), .o(n_9884) );
ao12s01 g771305 ( .a(n_9308), .b(n_9780), .c(n_9380), .o(n_9881) );
in01s01 g771310 ( .a(n_9639), .o(n_9686) );
ao12f04 g771311 ( .a(n_9346), .b(n_9567), .c(n_9376), .o(n_9639) );
oa22s01 g771312 ( .a(n_9780), .b(n_9435), .c(n_9654), .d(n_9436), .o(n_9832) );
oa22m02 g771315 ( .a(n_9137), .b(n_9178), .c(n_9138), .d(n_9177), .o(n_9411) );
in01s01 g771318 ( .a(n_9148), .o(n_9162) );
in01s01 g771319 ( .a(n_9091), .o(n_9148) );
in01m02 g771320 ( .a(n_9091), .o(n_9092) );
in01s01 g771329 ( .a(n_9111), .o(n_9173) );
in01s02 g771330 ( .a(n_9090), .o(n_9111) );
no02s04 TIMEBOOST_cell_8613 ( .a(TIMEBOOST_net_2793), .b(FE_OCP_RBN3238_n_5307), .o(n_5484) );
no02f04 g771334 ( .a(n_9564), .b(n_9609), .o(n_9794) );
in01f01 g771336 ( .a(n_9354), .o(n_9374) );
na02f06 g771337 ( .a(n_9205), .b(n_9202), .o(n_9354) );
in01s01 g771339 ( .a(n_9114), .o(n_9197) );
in01s01 g771340 ( .a(n_9057), .o(n_9114) );
in01s02 g771341 ( .a(n_9057), .o(n_9058) );
na02f02 g771346 ( .a(n_9344), .b(n_9294), .o(n_9535) );
na02f04 TIMEBOOST_cell_8659 ( .a(TIMEBOOST_net_2816), .b(n_16763), .o(n_16916) );
no02m04 TIMEBOOST_cell_2960 ( .a(n_23872), .b(n_24092), .o(TIMEBOOST_net_771) );
in01s02 g771349 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_), .o(n_9777) );
in01s02 g771352 ( .a(n_9353), .o(n_9372) );
no02f06 g771353 ( .a(n_9208), .b(n_9163), .o(n_9353) );
no02s06 g771355 ( .a(n_9347), .b(n_9191), .o(n_9351) );
na02m04 TIMEBOOST_cell_5661 ( .a(TIMEBOOST_net_1778), .b(n_17049), .o(n_17294) );
no02f08 TIMEBOOST_cell_4274 ( .a(TIMEBOOST_net_1227), .b(n_2318), .o(FE_RN_780_0) );
no02s02 TIMEBOOST_cell_8875 ( .a(TIMEBOOST_net_2924), .b(n_31400), .o(n_31465) );
in01s02 g771359 ( .a(n_9408), .o(n_9409) );
na02s04 g771360 ( .a(n_9318), .b(n_9253), .o(n_9408) );
na02s04 g771361 ( .a(FE_OCP_RBN2867_n_9347), .b(n_9210), .o(n_9350) );
no02s02 g771362 ( .a(n_9163), .b(n_9347), .o(n_9348) );
na02m02 g771363 ( .a(FE_OCP_RBN4235_n_9089), .b(n_9047), .o(n_9150) );
no02f04 TIMEBOOST_cell_8774 ( .a(FE_OCP_RBN4229_n_13962), .b(n_14932), .o(TIMEBOOST_net_2874) );
na02s02 g771365 ( .a(n_9188), .b(n_8232), .o(n_9254) );
in01s02 g771366 ( .a(n_9261), .o(n_9194) );
no02m06 g771367 ( .a(n_9113), .b(n_9112), .o(n_9261) );
na02f02 g771368 ( .a(n_9345), .b(n_9243), .o(n_9346) );
no02s02 g771370 ( .a(n_9567), .b(FE_OCP_RBN4282_n_9243), .o(n_9611) );
na02m04 g771371 ( .a(n_9485), .b(n_9378), .o(n_9588) );
na02s02 g771373 ( .a(n_9345), .b(n_9376), .o(n_9425) );
na02s06 g771377 ( .a(n_9370), .b(FE_OCP_RBN6731_n_44579), .o(n_9447) );
na02f02 g771378 ( .a(n_9400), .b(n_44594), .o(n_9531) );
na02s02 g771379 ( .a(n_9247), .b(n_44576), .o(n_9294) );
na02f02 g771380 ( .a(FE_OCP_RBN6734_n_44579), .b(FE_OCP_RBN2985_n_9247), .o(n_9344) );
na02m06 g771381 ( .a(n_9401), .b(FE_OCPN880_n_44593), .o(n_9586) );
in01m04 g771384 ( .a(n_9446), .o(n_9464) );
no02m06 g771385 ( .a(n_9370), .b(FE_OCP_RBN5833_n_44563), .o(n_9446) );
in01s02 g771386 ( .a(n_9266), .o(n_9267) );
in01f01 g771387 ( .a(n_9152), .o(n_9266) );
no02m06 g771388 ( .a(n_9093), .b(n_9099), .o(n_9152) );
in01s01 g771389 ( .a(n_9698), .o(n_9699) );
na02m02 g771390 ( .a(n_9643), .b(n_9642), .o(n_9698) );
in01s02 g771393 ( .a(n_9527), .o(n_9528) );
na02s02 g771394 ( .a(n_9486), .b(n_9403), .o(n_9527) );
in01s01 g771395 ( .a(n_9213), .o(n_9214) );
na02m06 g771396 ( .a(n_9088), .b(FE_OCP_RBN2752_FE_RN_1223_0), .o(n_9213) );
no02s02 g771397 ( .a(n_9643), .b(n_9642), .o(n_9787) );
in01s01 g771398 ( .a(n_9721), .o(n_9722) );
no02m02 g771399 ( .a(n_9641), .b(n_9640), .o(n_9721) );
na02f04 g771400 ( .a(n_9116), .b(n_9201), .o(n_9205) );
no02s02 TIMEBOOST_cell_5363 ( .a(TIMEBOOST_net_1629), .b(n_31349), .o(n_31350) );
no02f02 g771402 ( .a(n_9563), .b(n_9687), .o(n_9564) );
na02f02 g771403 ( .a(n_9166), .b(n_8927), .o(n_9215) );
no02f04 g771404 ( .a(n_9167), .b(n_8905), .o(n_9293) );
no02s01 g771405 ( .a(n_9609), .b(n_9563), .o(n_9688) );
no02s01 g771406 ( .a(n_9561), .b(n_9656), .o(n_9737) );
na02f02 g771407 ( .a(n_9641), .b(n_9640), .o(n_9786) );
na02s04 g771408 ( .a(n_9523), .b(n_9440), .o(n_9549) );
no02s01 g771409 ( .a(n_9634), .b(n_9604), .o(n_9834) );
oa12s01 g771410 ( .a(n_9607), .b(n_9606), .c(n_9605), .o(n_9782) );
na02s01 TIMEBOOST_cell_3236 ( .a(n_20675), .b(n_20519), .o(TIMEBOOST_net_909) );
in01s01 g771415 ( .a(n_9655), .o(n_9833) );
no02m04 g771417 ( .a(n_9340), .b(n_9274), .o(n_9513) );
na02s01 TIMEBOOST_cell_6923 ( .a(n_2175), .b(FE_RN_824_0), .o(TIMEBOOST_net_2220) );
na03f08 TIMEBOOST_cell_8288 ( .a(n_29635), .b(n_29613), .c(n_29591), .o(n_29716) );
no02s01 TIMEBOOST_cell_4039 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n_45840), .o(TIMEBOOST_net_1110) );
no02s03 g771424 ( .a(n_9044), .b(FE_OCPN4535_n_9012), .o(n_9095) );
no02s04 g771428 ( .a(n_9190), .b(FE_OCPN4535_n_9012), .o(n_9191) );
na02s04 g771429 ( .a(n_9134), .b(n_8309), .o(n_9253) );
no02m06 g771433 ( .a(FE_OCP_RBN2839_n_8974), .b(FE_OCP_DRV_N3506_n_8189), .o(n_9089) );
in01s01 g771434 ( .a(n_9112), .o(n_9047) );
no02s04 g771435 ( .a(n_8974), .b(FE_OCP_RBN4146_n_7743), .o(n_9112) );
na02s04 g771436 ( .a(n_9190), .b(FE_OCPN4535_n_9012), .o(n_9318) );
na02s02 g771437 ( .a(n_9082), .b(FE_OFN4770_n_8309), .o(n_9140) );
in01s01 g771439 ( .a(n_9163), .o(n_9210) );
no02s04 g771440 ( .a(n_9080), .b(n_8309), .o(n_9163) );
no02m02 g771441 ( .a(n_9521), .b(n_9398), .o(n_9562) );
in01s01 g771442 ( .a(n_9406), .o(n_9407) );
no02m02 g771443 ( .a(n_9317), .b(n_9269), .o(n_9406) );
no02m06 g771444 ( .a(n_9377), .b(n_9337), .o(n_9567) );
no02f08 TIMEBOOST_cell_3235 ( .a(TIMEBOOST_net_908), .b(n_5944), .o(n_6062) );
na02f02 g771446 ( .a(n_9185), .b(FE_OCP_RBN5837_n_44563), .o(n_9345) );
in01m02 g771447 ( .a(n_9404), .o(n_9405) );
no02s02 g771448 ( .a(n_9317), .b(n_9341), .o(n_9404) );
na02s06 g771449 ( .a(FE_OCP_RBN6751_n_9185), .b(FE_OCPN880_n_44593), .o(n_9376) );
na02s01 g771450 ( .a(FE_OCP_RBN2841_n_9044), .b(FE_OCP_DRV_N7079_n_8992), .o(n_9146) );
no02f02 g771451 ( .a(n_9441), .b(n_7978), .o(n_9563) );
no02m04 g771452 ( .a(n_9246), .b(n_9132), .o(n_9340) );
in01m01 g771453 ( .a(n_9113), .o(n_9050) );
in01s01 g771455 ( .a(n_9560), .o(n_9561) );
na02s03 g771456 ( .a(n_9526), .b(n_9525), .o(n_9560) );
in01s01 g771457 ( .a(n_9633), .o(n_9634) );
na02s04 g771458 ( .a(n_9520), .b(n_8025), .o(n_9633) );
na02s04 g771459 ( .a(n_9305), .b(FE_OCP_RBN2661_n_9304), .o(n_9486) );
no02s02 g771460 ( .a(n_9245), .b(n_9074), .o(n_9274) );
na02s01 g771461 ( .a(n_9606), .b(n_9605), .o(n_9607) );
in01s02 g771462 ( .a(n_9290), .o(n_9291) );
na02m02 g771463 ( .a(n_9212), .b(n_9136), .o(n_9290) );
oa12s04 g771464 ( .a(n_7678), .b(FE_OCP_RBN2798_n_8817), .c(FE_OCPN1210_n_8846), .o(n_8914) );
no02s02 TIMEBOOST_cell_8859 ( .a(TIMEBOOST_net_2916), .b(n_32223), .o(FE_RN_374_0) );
no02m04 g771466 ( .a(n_9442), .b(n_7979), .o(n_9609) );
no02s04 g771467 ( .a(n_9526), .b(n_9525), .o(n_9656) );
in01f02 g771468 ( .a(n_9166), .o(n_9167) );
in01f01 g771469 ( .a(n_9116), .o(n_9166) );
no02f04 g771470 ( .a(n_9046), .b(n_8936), .o(n_9116) );
in01s01 g771471 ( .a(n_9603), .o(n_9604) );
na02m02 g771472 ( .a(n_9519), .b(n_8024), .o(n_9603) );
na02s01 g771473 ( .a(n_9121), .b(n_9041), .o(n_9204) );
in01s01 g771474 ( .a(n_9402), .o(n_9403) );
no02m04 g771475 ( .a(n_9305), .b(FE_OCP_RBN2661_n_9304), .o(n_9402) );
in01m02 g771476 ( .a(n_8943), .o(n_8944) );
ao12m06 g771477 ( .a(n_7622), .b(FE_OCP_RBN2799_n_8817), .c(n_7633), .o(n_8943) );
in01s02 g771478 ( .a(n_8941), .o(n_8942) );
ao12s02 g771479 ( .a(n_7744), .b(FE_OCP_RBN2798_n_8817), .c(n_7738), .o(n_8941) );
in01s02 g771480 ( .a(n_9288), .o(n_9289) );
in01s02 g771481 ( .a(n_9208), .o(n_9288) );
oa12f06 g771482 ( .a(n_9189), .b(n_9074), .c(n_9077), .o(n_9208) );
in01s01 g771484 ( .a(n_9654), .o(n_9780) );
ao12m06 g771485 ( .a(n_9225), .b(n_9595), .c(n_9323), .o(n_9654) );
in01s01 g771486 ( .a(n_9523), .o(n_9524) );
in01s02 g771487 ( .a(n_9485), .o(n_9523) );
na02s03 TIMEBOOST_cell_7619 ( .a(TIMEBOOST_net_2440), .b(n_2726), .o(n_2864) );
in01m02 g771489 ( .a(n_9400), .o(n_9401) );
oa22f02 g771490 ( .a(n_9182), .b(n_44594), .c(FE_OCP_RBN2988_n_9182), .d(FE_OCP_RBN6710_n_44570), .o(n_9400) );
in01s02 g771491 ( .a(n_9137), .o(n_9138) );
in01m01 g771492 ( .a(n_9093), .o(n_9137) );
ao12m04 g771493 ( .a(n_47244), .b(n_8922), .c(n_47243), .o(n_9093) );
ao22f02 g771497 ( .a(n_9017), .b(n_8930), .c(FE_OCP_RBN2886_n_9017), .d(n_8929), .o(n_9198) );
in01s02 g771498 ( .a(n_9087), .o(n_9088) );
oa12s01 g771500 ( .a(n_9559), .b(n_9595), .c(n_9558), .o(n_9653) );
no02s02 TIMEBOOST_cell_4331 ( .a(n_38213), .b(n_38200), .o(TIMEBOOST_net_1256) );
in01s01 g771510 ( .a(n_8951), .o(n_9014) );
in01s02 g771511 ( .a(n_8951), .o(n_8952) );
na02s02 TIMEBOOST_cell_5574 ( .a(n_6172), .b(n_6311), .o(TIMEBOOST_net_1735) );
na02m06 g771517 ( .a(n_9153), .b(n_9101), .o(n_9370) );
na02s01 TIMEBOOST_cell_2051 ( .a(n_24013), .b(n_24041), .o(TIMEBOOST_net_640) );
no02s02 g771521 ( .a(n_8985), .b(FE_OCP_RBN2786_n_8767), .o(n_8986) );
in01m02 g771522 ( .a(n_9245), .o(n_9246) );
na02m04 g771523 ( .a(n_9078), .b(n_9189), .o(n_9245) );
na02s01 g771524 ( .a(n_9595), .b(n_9558), .o(n_9559) );
na02m04 g771529 ( .a(FE_OCP_RBN4314_n_9396), .b(n_9327), .o(n_9521) );
no02m04 TIMEBOOST_cell_6908 ( .a(n_24068), .b(TIMEBOOST_net_2212), .o(TIMEBOOST_net_1458) );
no02s08 TIMEBOOST_cell_6873 ( .a(n_11770), .b(n_11910), .o(TIMEBOOST_net_2195) );
no02m02 g771532 ( .a(n_9102), .b(n_44579), .o(n_9317) );
na03f06 TIMEBOOST_cell_8371 ( .a(n_4316), .b(FE_OCP_RBN6111_n_5444), .c(n_5495), .o(n_5644) );
na02m04 g771534 ( .a(FE_OCP_RBN6760_n_9075), .b(n_44594), .o(n_9153) );
no02s04 g771535 ( .a(FE_OCP_RBN4330_n_9102), .b(FE_OCP_RBN5838_n_44563), .o(n_9341) );
in01s02 g771536 ( .a(n_9398), .o(n_9399) );
no02m04 g771537 ( .a(FE_OCP_RBN4283_n_9243), .b(n_9337), .o(n_9398) );
na02f02 g771538 ( .a(n_9075), .b(FE_OCP_RBN6733_n_44579), .o(n_9101) );
in01s01 g771540 ( .a(n_9135), .o(n_9136) );
no02m06 g771541 ( .a(n_9086), .b(FE_OCP_RBN2701_n_8187), .o(n_9135) );
na02f02 TIMEBOOST_cell_5207 ( .a(TIMEBOOST_net_1551), .b(n_8584), .o(n_8729) );
na03f10 TIMEBOOST_cell_2212 ( .a(n_27920), .b(FE_RN_361_0), .c(FE_RN_360_0), .o(n_46961) );
na02s06 g771544 ( .a(n_9086), .b(FE_OCP_RBN2701_n_8187), .o(n_9212) );
in01s01 g771546 ( .a(n_9083), .o(n_9084) );
in01s01 g771547 ( .a(n_9046), .o(n_9083) );
oa12f04 g771548 ( .a(n_8887), .b(n_8911), .c(n_8861), .o(n_9046) );
oa22f02 g771552 ( .a(n_9009), .b(n_44576), .c(FE_OCP_RBN4263_n_9009), .d(FE_OCP_RBN6710_n_44570), .o(n_9185) );
na02s03 g771553 ( .a(n_9276), .b(n_9355), .o(n_9397) );
oa12s01 g771554 ( .a(n_9393), .b(n_9392), .c(FE_OFN381_n_9391), .o(n_9474) );
in01s01 g771555 ( .a(n_9506), .o(n_9606) );
no02f04 TIMEBOOST_cell_7571 ( .a(TIMEBOOST_net_2416), .b(n_29210), .o(n_29318) );
in01m01 g771558 ( .a(n_9441), .o(n_9442) );
oa22m02 g771559 ( .a(n_9234), .b(n_9128), .c(n_9235), .d(n_9127), .o(n_9441) );
in01s01 g771560 ( .a(n_10733), .o(n_9200) );
in01s01 g771561 ( .a(FE_OCP_RBN2859_n_9082), .o(n_10733) );
na02f04 g771564 ( .a(n_9076), .b(n_9201), .o(n_9202) );
in01s02 g771565 ( .a(n_9519), .o(n_9520) );
na02m04 g771567 ( .a(n_9079), .b(n_9115), .o(n_9305) );
oa12s01 g771568 ( .a(n_9781), .b(n_9332), .c(n_9331), .o(n_9428) );
in01s02 g771573 ( .a(n_9190), .o(n_9134) );
no02f08 TIMEBOOST_cell_4233 ( .a(n_40806), .b(n_41084), .o(TIMEBOOST_net_1207) );
in01s01 g771577 ( .a(FE_OCP_RBN2841_n_9044), .o(n_9121) );
na02m02 g771582 ( .a(n_8881), .b(n_8880), .o(n_8985) );
na02s02 g771583 ( .a(n_9025), .b(n_9007), .o(n_9079) );
na02m02 g771584 ( .a(n_9026), .b(n_9006), .o(n_9115) );
na02s04 TIMEBOOST_cell_4232 ( .a(TIMEBOOST_net_1206), .b(n_33397), .o(n_33446) );
in01m02 g771587 ( .a(n_9077), .o(n_9078) );
in01s03 g771589 ( .a(n_8989), .o(n_9189) );
no02m02 g771590 ( .a(n_8953), .b(n_8309), .o(n_8989) );
no02s02 g771592 ( .a(n_8923), .b(FE_OFN4770_n_8309), .o(n_8973) );
in01s01 g771594 ( .a(n_10385), .o(n_10386) );
no02s01 g771595 ( .a(n_10340), .b(n_10341), .o(n_10385) );
no02s01 g771596 ( .a(n_10283), .b(n_10284), .o(n_10285) );
in01s01 g771598 ( .a(n_9268), .o(n_9335) );
no02m04 g771599 ( .a(n_9168), .b(n_9203), .o(n_9268) );
na02m04 TIMEBOOST_cell_5331 ( .a(TIMEBOOST_net_1613), .b(n_15809), .o(n_15992) );
in01m02 g771602 ( .a(n_9333), .o(n_9396) );
no02m04 g771603 ( .a(n_9236), .b(FE_OCP_RBN6723_n_44055), .o(n_9333) );
na02m02 g771605 ( .a(n_9238), .b(n_9265), .o(n_9365) );
na02s01 g771607 ( .a(n_10210), .b(n_10209), .o(n_10211) );
in01s01 g771608 ( .a(n_10296), .o(n_10297) );
na02s01 g771609 ( .a(n_10210), .b(n_11266), .o(n_10296) );
no02m04 g771610 ( .a(n_9165), .b(n_44576), .o(n_9337) );
in01s01 g771611 ( .a(n_10383), .o(n_10384) );
no02s01 g771612 ( .a(n_10340), .b(n_10283), .o(n_10383) );
na02m04 g771614 ( .a(n_9165), .b(FE_OCP_RBN5837_n_44563), .o(n_9243) );
in01s02 g771615 ( .a(n_9439), .o(n_9440) );
na02m04 g771616 ( .a(n_9379), .b(n_9378), .o(n_9439) );
in01s01 g771617 ( .a(n_10343), .o(n_10344) );
no02s01 g771618 ( .a(n_10341), .b(n_10284), .o(n_10343) );
no02s02 g771619 ( .a(n_9130), .b(n_9070), .o(n_9170) );
na02m02 g771620 ( .a(n_9201), .b(FE_OCP_RBN2923_n_9070), .o(n_9242) );
na02s02 g771621 ( .a(n_9275), .b(FE_OFN381_n_9391), .o(n_9687) );
na02s01 g771622 ( .a(n_9392), .b(FE_OFN381_n_9391), .o(n_9393) );
no02s01 g771623 ( .a(n_9328), .b(n_9286), .o(n_9368) );
na02s01 g771624 ( .a(n_9355), .b(n_9237), .o(n_9438) );
na02s02 g771625 ( .a(n_9237), .b(n_9036), .o(n_9276) );
na02s04 g771626 ( .a(n_9332), .b(n_9331), .o(n_9781) );
na02f02 g771627 ( .a(n_9027), .b(n_8862), .o(n_9076) );
no02s02 TIMEBOOST_cell_2049 ( .a(n_3331), .b(n_2641), .o(TIMEBOOST_net_639) );
oa12m06 g771632 ( .a(n_9206), .b(n_9482), .c(n_9322), .o(n_9595) );
oa12f02 g771634 ( .a(n_8858), .b(n_8891), .c(n_8813), .o(n_9017) );
oa12s01 g771635 ( .a(n_9430), .b(n_9482), .c(n_9429), .o(n_9518) );
oa12m04 g771642 ( .a(FE_OCP_RBN5846_FE_RN_987_0), .b(n_8872), .c(FE_OCP_RBN5848_FE_RN_2187_0), .o(n_8922) );
ao12f04 g771644 ( .a(FE_OCP_RBN5850_FE_RN_2187_0), .b(FE_OCP_RBN4269_n_8872), .c(FE_OCP_RBN5847_FE_RN_987_0), .o(n_9042) );
in01m01 g771646 ( .a(n_9074), .o(n_9132) );
na02f06 g771647 ( .a(n_8972), .b(n_8970), .o(n_9074) );
in01s02 g771648 ( .a(n_9010), .o(n_9011) );
na02s02 TIMEBOOST_cell_5526 ( .a(n_6025), .b(n_5791), .o(TIMEBOOST_net_1711) );
no02s01 TIMEBOOST_cell_7509 ( .a(TIMEBOOST_net_2385), .b(n_2445), .o(TIMEBOOST_net_1247) );
no02s10 TIMEBOOST_cell_8824 ( .a(TIMEBOOST_net_1632), .b(n_16086), .o(TIMEBOOST_net_2899) );
no02s06 g771655 ( .a(n_8885), .b(n_7571), .o(n_8939) );
no02s06 TIMEBOOST_cell_8691 ( .a(TIMEBOOST_net_2832), .b(FE_RN_728_0), .o(FE_RN_731_0) );
na02f04 g771658 ( .a(n_8969), .b(n_8971), .o(n_8972) );
no02m04 g771659 ( .a(n_8968), .b(n_8919), .o(n_8970) );
in01m02 g771660 ( .a(n_9025), .o(n_9026) );
na02m02 g771661 ( .a(n_8920), .b(n_8971), .o(n_9025) );
no02f04 TIMEBOOST_cell_5043 ( .a(TIMEBOOST_net_1469), .b(n_37883), .o(n_37943) );
na02s01 g771666 ( .a(n_9482), .b(n_9429), .o(n_9430) );
in01s02 g771667 ( .a(n_9264), .o(n_9265) );
in01s02 g771668 ( .a(n_9203), .o(n_9264) );
na02m04 g771669 ( .a(n_9097), .b(n_9005), .o(n_9203) );
no02s01 g771670 ( .a(n_9065), .b(n_44511), .o(n_10283) );
na02s01 g771671 ( .a(n_10073), .b(n_44516), .o(n_11266) );
in01s01 g771672 ( .a(n_10284), .o(n_10250) );
no02s01 g771673 ( .a(n_44511), .b(n_9029), .o(n_10284) );
no02s01 g771674 ( .a(n_9066), .b(n_44516), .o(n_10340) );
in01m02 g771675 ( .a(n_9269), .o(n_9379) );
no02m02 g771676 ( .a(n_9240), .b(n_44579), .o(n_9269) );
in01s01 g771677 ( .a(n_9389), .o(n_9390) );
na02m02 g771678 ( .a(n_9232), .b(n_9330), .o(n_9389) );
no02s01 g771679 ( .a(FE_OFN810_n_9028), .b(n_44516), .o(n_10341) );
in01s01 g771680 ( .a(n_10124), .o(n_10210) );
no02s01 g771681 ( .a(n_44516), .b(n_10073), .o(n_10124) );
na02s04 g771682 ( .a(n_9240), .b(n_44575), .o(n_9378) );
in01m01 g771683 ( .a(n_9238), .o(n_9239) );
no02m02 g771684 ( .a(n_9169), .b(n_9168), .o(n_9238) );
in01s01 g771686 ( .a(n_9237), .o(n_9286) );
na02f02 g771687 ( .a(n_9125), .b(FE_OCP_RBN6630_n_8269), .o(n_9237) );
in01s01 g771689 ( .a(n_9201), .o(n_9130) );
na02m06 g771690 ( .a(n_8965), .b(FE_OCP_RBN5697_n_8342), .o(n_9201) );
in01s01 g771692 ( .a(n_9355), .o(n_9328) );
in01m01 g771695 ( .a(n_9027), .o(n_9070) );
na02f02 g771696 ( .a(FE_OCP_RBN6645_n_8342), .b(n_8964), .o(n_9027) );
no02f04 g771697 ( .a(n_8848), .b(n_8794), .o(n_8911) );
oa12s02 g771698 ( .a(n_7554), .b(n_8863), .c(n_8840), .o(n_8864) );
no02s01 TIMEBOOST_cell_6718 ( .a(TIMEBOOST_net_2116), .b(n_2987), .o(n_3035) );
ao12m06 g771700 ( .a(n_7584), .b(n_44057), .c(n_8699), .o(n_8746) );
na02f04 g771701 ( .a(n_8786), .b(n_8795), .o(n_8881) );
no02m04 g771702 ( .a(n_8791), .b(n_8784), .o(n_8880) );
no02m02 g771704 ( .a(n_9236), .b(n_9105), .o(n_9284) );
in01s02 g771705 ( .a(n_9234), .o(n_9235) );
no02s01 TIMEBOOST_cell_8536 ( .a(TIMEBOOST_net_2095), .b(n_14044), .o(TIMEBOOST_net_2755) );
na02s04 g771708 ( .a(n_9180), .b(n_9119), .o(n_9306) );
na02m04 g771710 ( .a(n_9327), .b(n_9228), .o(n_9387) );
in01s01 g771711 ( .a(n_9275), .o(n_9392) );
ao22s02 g771712 ( .a(n_8995), .b(FE_OCP_RBN4244_n_44594), .c(n_9032), .d(FE_OCP_RBN4240_n_44594), .o(n_9275) );
in01s01 g771717 ( .a(n_8865), .o(n_8908) );
in01s01 g771718 ( .a(n_8842), .o(n_8865) );
in01m02 g771719 ( .a(n_8842), .o(n_8828) );
in01s01 g771723 ( .a(FE_OCP_DRV_N7079_n_8992), .o(n_9041) );
in01s01 g771724 ( .a(n_8983), .o(n_8992) );
in01m02 g771725 ( .a(n_8923), .o(n_8983) );
oa22m04 g771730 ( .a(n_44576), .b(FE_OCP_RBN4246_n_8904), .c(FE_OCP_RBN4239_n_44594), .d(FE_OFN5066_n_8904), .o(n_9165) );
oa12s01 g771731 ( .a(n_9326), .b(n_9325), .c(n_9324), .o(n_9437) );
in01s01 g771732 ( .a(n_10484), .o(n_8937) );
in01m01 g771733 ( .a(FE_OCPN1079_n_8915), .o(n_10484) );
ao22s02 g771736 ( .a(n_9035), .b(FE_OCP_RBN4244_n_44594), .c(FE_OCP_RBN4241_n_44594), .d(FE_OCP_RBN5843_n_9035), .o(n_9332) );
na02s01 TIMEBOOST_cell_6315 ( .a(n_35795), .b(n_35717), .o(TIMEBOOST_net_2009) );
in01s02 g771740 ( .a(n_9006), .o(n_9007) );
no02m02 g771741 ( .a(n_8969), .b(n_8968), .o(n_9006) );
na02f04 g771743 ( .a(n_8787), .b(FE_OCP_RBN4223_n_8784), .o(n_8850) );
na02m02 g771744 ( .a(n_8790), .b(FE_OCP_DRV_N3506_n_8189), .o(n_8795) );
in01s01 g771745 ( .a(n_8919), .o(n_8920) );
no02f02 g771746 ( .a(n_8879), .b(FE_OCP_DRV_N3506_n_8189), .o(n_8919) );
na02s02 g771747 ( .a(n_8879), .b(n_8189), .o(n_8971) );
no02f02 g771748 ( .a(n_8790), .b(FE_OCP_DRV_N3506_n_8189), .o(n_8791) );
no02s01 g771749 ( .a(n_9830), .b(n_9876), .o(n_9915) );
no02s01 g771750 ( .a(n_10120), .b(n_10123), .o(n_10161) );
na02s01 g771751 ( .a(n_10158), .b(n_10159), .o(n_10160) );
in01s01 g771752 ( .a(n_10239), .o(n_10240) );
na02s01 g771753 ( .a(n_10159), .b(n_10208), .o(n_10239) );
in01s01 g771754 ( .a(n_10248), .o(n_10249) );
na02s01 g771755 ( .a(n_10158), .b(n_10121), .o(n_10248) );
na02m02 g771756 ( .a(n_9110), .b(n_44575), .o(n_9330) );
in01s01 g771757 ( .a(n_10381), .o(n_10382) );
na02s01 g771758 ( .a(n_10247), .b(n_10209), .o(n_10381) );
no02m02 g771759 ( .a(n_9002), .b(FE_OCP_RBN6711_n_44570), .o(n_9169) );
no02s02 g771760 ( .a(n_44594), .b(n_9001), .o(n_9168) );
na02s02 g771761 ( .a(n_8980), .b(n_44575), .o(n_9005) );
na02m02 g771762 ( .a(n_8980), .b(FE_OCP_RBN4240_n_44594), .o(n_9053) );
na02s40 TIMEBOOST_cell_7405 ( .a(n_16972), .b(TIMEBOOST_net_2333), .o(n_17192) );
na02s02 g771764 ( .a(n_9061), .b(n_44594), .o(n_9232) );
na02m04 TIMEBOOST_cell_7743 ( .a(TIMEBOOST_net_2502), .b(FE_OCP_RBN5915_n_3750), .o(n_4023) );
na02s02 g771767 ( .a(n_9034), .b(FE_OCP_RBN4241_n_44594), .o(n_9180) );
in01s02 g771768 ( .a(n_9127), .o(n_9128) );
in01s02 g771769 ( .a(n_9097), .o(n_9127) );
na02m04 g771770 ( .a(n_8995), .b(n_44575), .o(n_9097) );
na02s02 g771771 ( .a(FE_OCP_RBN6722_n_9034), .b(FE_OCP_RBN4244_n_44594), .o(n_9119) );
in01s01 g771772 ( .a(n_9229), .o(n_9230) );
na02s02 g771774 ( .a(n_9035), .b(n_44579), .o(n_9229) );
no02s04 g771775 ( .a(n_9020), .b(FE_OCP_RBN4244_n_44594), .o(n_9236) );
no02s02 TIMEBOOST_cell_3059 ( .a(TIMEBOOST_net_820), .b(n_38523), .o(n_38570) );
na02s04 g771777 ( .a(n_9157), .b(FE_OCP_RBN4241_n_44594), .o(n_9327) );
no02m02 g771778 ( .a(n_9021), .b(n_44579), .o(n_9105) );
na02s04 g771779 ( .a(n_9124), .b(FE_OCP_RBN4244_n_44594), .o(n_9228) );
na02s01 g771780 ( .a(n_9325), .b(n_9324), .o(n_9326) );
in01s02 g771781 ( .a(n_9177), .o(n_9178) );
no02s02 g771782 ( .a(n_9099), .b(n_9051), .o(n_9177) );
no02m06 g771783 ( .a(n_8863), .b(n_7592), .o(n_8885) );
in01s01 g771784 ( .a(n_8966), .o(n_8967) );
no02s02 g771785 ( .a(n_8905), .b(n_8936), .o(n_8966) );
in01m01 g771787 ( .a(n_8891), .o(n_8934) );
in01m01 g771788 ( .a(n_8848), .o(n_8891) );
oa12f04 g771789 ( .a(n_8682), .b(n_8751), .c(n_8661), .o(n_8848) );
na02s01 g771790 ( .a(n_9877), .b(n_9955), .o(n_9956) );
no02m06 g771791 ( .a(n_9263), .b(n_9218), .o(n_9482) );
in01s01 g771792 ( .a(FE_OFN810_n_9028), .o(n_9029) );
ao12s01 g771793 ( .a(n_8933), .b(n_8932), .c(n_8931), .o(n_9028) );
no03f06 TIMEBOOST_cell_5358 ( .a(n_15109), .b(n_15038), .c(n_15108), .o(TIMEBOOST_net_1627) );
ao12f04 g771800 ( .a(n_8714), .b(n_8766), .c(n_8771), .o(n_8872) );
in01m02 g771807 ( .a(n_8964), .o(n_8965) );
na02f04 g771808 ( .a(n_8849), .b(n_8839), .o(n_8964) );
ao12s01 g771809 ( .a(n_8869), .b(n_8868), .c(n_8867), .o(n_10073) );
in01s01 g771810 ( .a(n_9065), .o(n_9066) );
oa12s01 g771811 ( .a(n_8963), .b(n_8962), .c(n_8961), .o(n_9065) );
na02f04 g771812 ( .a(FE_OCP_RBN6713_n_8800), .b(n_8562), .o(n_8849) );
na02m02 g771813 ( .a(n_8800), .b(n_8610), .o(n_8839) );
na02s01 g771814 ( .a(n_8962), .b(n_8961), .o(n_8963) );
no02s01 g771815 ( .a(n_8932), .b(n_8931), .o(n_8933) );
no02s01 g771816 ( .a(n_8867), .b(n_8868), .o(n_8869) );
no02s03 g771817 ( .a(n_9309), .b(n_9308), .o(n_9310) );
no02s01 g771818 ( .a(n_9825), .b(n_9876), .o(n_9877) );
na02s02 g771819 ( .a(n_9480), .b(n_9431), .o(n_9481) );
no02s01 g771820 ( .a(n_9433), .b(n_9547), .o(n_9548) );
na02s01 g771821 ( .a(n_9592), .b(n_9730), .o(n_9696) );
na02s02 g771822 ( .a(n_9281), .b(n_9380), .o(n_9311) );
na02s01 g771823 ( .a(n_9811), .b(n_9733), .o(n_9776) );
na02s01 g771824 ( .a(n_9693), .b(n_9728), .o(n_9729) );
in01s01 g771825 ( .a(n_9955), .o(n_9830) );
no02s01 g771826 ( .a(n_9775), .b(n_9774), .o(n_9955) );
no02s01 g771827 ( .a(n_9770), .b(n_9828), .o(n_9829) );
no02s01 g771828 ( .a(n_10037), .b(n_10081), .o(n_10082) );
no02s01 g771829 ( .a(n_9772), .b(n_9771), .o(n_9773) );
na02s01 g771830 ( .a(n_9874), .b(n_9873), .o(n_9875) );
na02s01 g771831 ( .a(n_9728), .b(n_9730), .o(n_10491) );
no02s01 g771832 ( .a(n_9517), .b(n_9596), .o(n_9961) );
na02s01 g771833 ( .a(n_9323), .b(n_9226), .o(n_9558) );
na02s01 g771834 ( .a(n_9386), .b(n_9475), .o(n_9815) );
no02m04 g771835 ( .a(n_9219), .b(n_9324), .o(n_9263) );
no02s01 g771836 ( .a(n_9602), .b(n_9695), .o(n_10237) );
na02s01 g771837 ( .a(n_9650), .b(n_9735), .o(n_10351) );
in01s01 g771838 ( .a(n_9813), .o(n_9814) );
na02s01 g771839 ( .a(n_9648), .b(n_9811), .o(n_9813) );
no02s01 g771840 ( .a(n_9771), .b(n_9734), .o(n_10686) );
na02s01 g771841 ( .a(n_9826), .b(n_9873), .o(n_10816) );
in01s01 g771842 ( .a(n_10156), .o(n_10157) );
no02s01 g771843 ( .a(n_11041), .b(n_10081), .o(n_10156) );
in01s01 g771844 ( .a(n_10123), .o(n_10208) );
no02s01 g771845 ( .a(n_44516), .b(n_10079), .o(n_10123) );
na02s01 g771846 ( .a(n_44511), .b(n_10122), .o(n_10209) );
no02m04 TIMEBOOST_cell_6294 ( .a(TIMEBOOST_net_1998), .b(n_35404), .o(n_35470) );
no02s01 g771848 ( .a(n_9694), .b(n_9591), .o(n_10576) );
na02s01 g771849 ( .a(n_44516), .b(n_10078), .o(n_10158) );
in01s01 g771850 ( .a(n_10120), .o(n_10121) );
no02s01 g771851 ( .a(n_44516), .b(n_10078), .o(n_10120) );
in01s01 g771852 ( .a(n_9435), .o(n_9436) );
na02s01 g771853 ( .a(n_9283), .b(n_9380), .o(n_9435) );
in01s01 g771854 ( .a(n_10159), .o(n_10119) );
na02s01 g771855 ( .a(n_10079), .b(n_44516), .o(n_10159) );
no02s01 g771856 ( .a(n_9219), .b(n_9218), .o(n_9325) );
in01s01 g771857 ( .a(n_10206), .o(n_10207) );
na02s01 g771858 ( .a(n_10154), .b(n_10038), .o(n_10206) );
no02s01 g771859 ( .a(n_9954), .b(n_10039), .o(n_10841) );
na02s01 g771860 ( .a(n_9692), .b(n_9870), .o(n_10657) );
no02s01 g771861 ( .a(n_9774), .b(n_9828), .o(n_10751) );
in01s01 g771862 ( .a(n_10246), .o(n_10247) );
no02s01 g771863 ( .a(n_10122), .b(n_44511), .o(n_10246) );
no02s01 g771864 ( .a(n_9432), .b(n_9547), .o(n_10217) );
na02s01 g771865 ( .a(n_10077), .b(n_9952), .o(n_10942) );
no02s01 g771866 ( .a(n_9309), .b(n_9282), .o(n_9880) );
na02s01 g771867 ( .a(n_9827), .b(n_9874), .o(n_10775) );
na02s01 g771868 ( .a(n_9480), .b(n_9505), .o(n_10086) );
no02s01 g771869 ( .a(n_9207), .b(n_9322), .o(n_9429) );
no02s02 g771870 ( .a(n_44575), .b(n_8902), .o(n_8988) );
in01s01 g771872 ( .a(n_9051), .o(n_9108) );
in01s01 g771873 ( .a(n_9036), .o(n_9051) );
na02m02 g771874 ( .a(FE_OCP_RBN2633_n_9003), .b(n_9004), .o(n_9036) );
no02s02 g771875 ( .a(n_9004), .b(FE_OCP_RBN2633_n_9003), .o(n_9099) );
in01s02 g771876 ( .a(n_8863), .o(n_8819) );
no02f08 g771877 ( .a(n_8748), .b(n_7570), .o(n_8863) );
in01s01 g771878 ( .a(n_8929), .o(n_8930) );
na02s02 g771879 ( .a(n_8860), .b(n_8887), .o(n_8929) );
in01s01 g771881 ( .a(n_8905), .o(n_8927) );
in01s02 g771882 ( .a(n_8862), .o(n_8905) );
na02s02 g771883 ( .a(n_8838), .b(n_46991), .o(n_8862) );
oa12m02 g771884 ( .a(n_7569), .b(n_8747), .c(n_8742), .o(n_8769) );
no02s06 TIMEBOOST_cell_6073 ( .a(n_24438), .b(n_24547), .o(TIMEBOOST_net_1888) );
no02s02 g771886 ( .a(n_46991), .b(n_8838), .o(n_8936) );
na02f04 g771887 ( .a(n_8860), .b(n_8770), .o(n_8861) );
in01m02 g771888 ( .a(n_8703), .o(n_8704) );
oa12f04 g771890 ( .a(n_8635), .b(n_45503), .c(n_8634), .o(n_8703) );
in01f02 g771891 ( .a(n_8786), .o(n_8787) );
no02m10 TIMEBOOST_cell_3223 ( .a(TIMEBOOST_net_902), .b(FE_RN_1112_0), .o(n_25458) );
no02m04 g771893 ( .a(n_8805), .b(n_8857), .o(n_8969) );
na02f02 g771895 ( .a(n_8698), .b(n_8678), .o(n_8784) );
in01s02 g771897 ( .a(n_9157), .o(n_9124) );
na02s06 TIMEBOOST_cell_6605 ( .a(n_17582), .b(n_17581), .o(TIMEBOOST_net_2060) );
ao12s02 g771899 ( .a(n_8560), .b(FE_OCP_RBN6704_n_8762), .c(n_8561), .o(n_8836) );
na02f02 g771900 ( .a(n_8508), .b(n_8798), .o(n_8859) );
ao22f02 g771903 ( .a(FE_OCP_RBN6705_n_8762), .b(n_8671), .c(n_8762), .d(n_8670), .o(n_8904) );
in01s01 g771905 ( .a(FE_OCP_RBN2790_n_8767), .o(n_10183) );
in01m02 g771909 ( .a(n_9020), .o(n_9021) );
in01m01 g771913 ( .a(n_8980), .o(n_8990) );
ao22f02 g771914 ( .a(n_8875), .b(FE_OCP_RBN4217_n_8597), .c(n_44570), .d(n_8597), .o(n_8980) );
ao22m06 g771917 ( .a(n_44575), .b(n_8514), .c(FE_OCP_RBN6708_n_44570), .d(FE_OCP_RBN4214_FE_OCPN3565_n_10214), .o(n_9035) );
ao22m04 g771920 ( .a(n_44575), .b(n_10374), .c(FE_OCP_RBN6708_n_44570), .d(FE_OCPN1206_n_46990), .o(n_9034) );
in01s01 g771922 ( .a(n_8995), .o(n_9032) );
no02m04 g771923 ( .a(n_8876), .b(n_8916), .o(n_8995) );
no02m02 TIMEBOOST_cell_4272 ( .a(TIMEBOOST_net_1226), .b(n_37976), .o(n_38041) );
in01s02 g771929 ( .a(n_9110), .o(n_9061) );
no02m04 g771930 ( .a(n_8925), .b(n_8955), .o(n_9110) );
in01m02 g771931 ( .a(n_9001), .o(n_9002) );
no02s02 TIMEBOOST_cell_2076 ( .a(TIMEBOOST_net_652), .b(n_39154), .o(n_39249) );
no02m06 g771934 ( .a(n_8747), .b(n_7537), .o(n_8748) );
no02s02 g771935 ( .a(n_8747), .b(n_7600), .o(n_8741) );
na02s02 TIMEBOOST_cell_2077 ( .a(n_42296), .b(n_42363), .o(TIMEBOOST_net_653) );
no03m10 TIMEBOOST_cell_5819 ( .a(TIMEBOOST_net_1106), .b(FE_OCPN1404_n_30823), .c(n_30814), .o(n_30958) );
no02s02 g771942 ( .a(n_8803), .b(FE_OCPN931_n_7817), .o(n_8805) );
na02m02 g771943 ( .a(n_8696), .b(FE_OCP_RBN4138_n_7743), .o(n_8698) );
na02s02 TIMEBOOST_cell_2099 ( .a(n_20850), .b(n_20495), .o(TIMEBOOST_net_664) );
in01s01 g771946 ( .a(n_9693), .o(n_9694) );
na02s01 g771947 ( .a(FE_OCP_RBN5907_n_44563), .b(n_9544), .o(n_9693) );
na02s01 g771948 ( .a(FE_OFN4778_n_44490), .b(n_9598), .o(n_9811) );
no02s02 g771949 ( .a(FE_OFN757_n_44464), .b(n_9913), .o(n_10039) );
no02s01 g771950 ( .a(FE_OFN4775_n_44463), .b(n_9681), .o(n_9771) );
in01s01 g771951 ( .a(n_9206), .o(n_9207) );
na02s06 g771952 ( .a(FE_OCP_RBN4240_n_44594), .b(n_9151), .o(n_9206) );
in01s01 g771953 ( .a(n_9480), .o(n_9434) );
na02s01 g771954 ( .a(FE_OCP_RBN5907_n_44563), .b(n_9367), .o(n_9480) );
no02s01 g771955 ( .a(FE_OCP_RBN5907_n_44563), .b(n_9381), .o(n_9547) );
in01s01 g771956 ( .a(n_9308), .o(n_9283) );
no02s01 g771957 ( .a(FE_OCP_RBN5838_n_44563), .b(n_9223), .o(n_9308) );
na02s02 g771958 ( .a(FE_OCP_RBN6737_n_44563), .b(n_9172), .o(n_9323) );
na02s01 g771959 ( .a(FE_OFN4775_n_44463), .b(n_9587), .o(n_9735) );
na02s01 g771960 ( .a(FE_OFN4775_n_44463), .b(n_9631), .o(n_9730) );
in01s01 g771961 ( .a(n_9651), .o(n_9728) );
no02s01 g771962 ( .a(FE_OFN4775_n_44463), .b(n_9631), .o(n_9651) );
in01s01 g771963 ( .a(n_9591), .o(n_9592) );
no02s01 g771964 ( .a(FE_OFN757_n_44464), .b(n_9544), .o(n_9591) );
in01s01 g771965 ( .a(n_9770), .o(n_9870) );
no02s01 g771966 ( .a(n_44492), .b(n_9647), .o(n_9770) );
no02s01 g771967 ( .a(n_44492), .b(n_8689), .o(n_9828) );
no02s01 g771968 ( .a(FE_OFN4778_n_44490), .b(n_8688), .o(n_9774) );
in01s01 g771969 ( .a(n_9876), .o(n_9827) );
no02s01 g771970 ( .a(FE_OCPN1061_n_44460), .b(n_9768), .o(n_9876) );
in01s01 g771971 ( .a(n_9953), .o(n_9954) );
na02s02 g771972 ( .a(FE_OFN4802_n_44498), .b(n_9913), .o(n_9953) );
in01s01 g771973 ( .a(n_9951), .o(n_9952) );
no02s02 g771974 ( .a(FE_OFN4802_n_44498), .b(FE_OFN809_n_9939), .o(n_9951) );
in01s01 g771975 ( .a(n_10037), .o(n_10038) );
no02s01 g771976 ( .a(FE_OFN4802_n_44498), .b(n_9994), .o(n_10037) );
na02s01 g771977 ( .a(n_44516), .b(n_9994), .o(n_10154) );
no02m02 g771978 ( .a(n_44575), .b(FE_OCP_RBN4237_n_8781), .o(n_9019) );
na02s01 g771979 ( .a(n_9767), .b(FE_OFN4778_n_44490), .o(n_9873) );
in01s01 g771980 ( .a(n_9516), .o(n_9517) );
na02s02 g771981 ( .a(FE_OCP_RBN5907_n_44563), .b(n_9369), .o(n_9516) );
in01s01 g771982 ( .a(n_9649), .o(n_9650) );
no02s01 g771983 ( .a(FE_OFN4778_n_44490), .b(n_9587), .o(n_9649) );
no02s01 TIMEBOOST_cell_5012 ( .a(n_29129), .b(n_29071), .o(TIMEBOOST_net_1454) );
no02s02 g771985 ( .a(FE_OCP_RBN5907_n_44563), .b(n_9369), .o(n_9596) );
in01s01 g771986 ( .a(n_9601), .o(n_9602) );
na02s02 g771987 ( .a(FE_OFN757_n_44464), .b(n_9478), .o(n_9601) );
no02s02 g771988 ( .a(n_44592), .b(n_8809), .o(n_8955) );
in01s01 g771989 ( .a(n_9225), .o(n_9226) );
no02s02 g771990 ( .a(n_44579), .b(n_9172), .o(n_9225) );
no02s02 g771991 ( .a(n_44570), .b(n_10137), .o(n_8916) );
na02s02 g771992 ( .a(FE_OCP_RBN5828_n_44579), .b(n_9223), .o(n_9380) );
no02s02 g771993 ( .a(n_44575), .b(n_7862), .o(n_9218) );
na02s02 g771994 ( .a(FE_OFN809_n_9939), .b(FE_OFN4802_n_44498), .o(n_10077) );
in01s01 g771995 ( .a(n_10081), .o(n_10036) );
no02s01 g771996 ( .a(FE_OFN4802_n_44498), .b(n_8810), .o(n_10081) );
no02s06 g771997 ( .a(FE_OCP_RBN6737_n_44563), .b(n_9151), .o(n_9322) );
in01s01 g771998 ( .a(n_9772), .o(n_9648) );
no02s01 g771999 ( .a(FE_OFN4778_n_44490), .b(n_9598), .o(n_9772) );
in01s01 g772000 ( .a(n_9825), .o(n_9826) );
no02s01 g772001 ( .a(FE_OCPN1061_n_44460), .b(n_9767), .o(n_9825) );
no02s06 g772002 ( .a(n_44576), .b(n_7861), .o(n_9219) );
no02s02 g772003 ( .a(n_8875), .b(n_8539), .o(n_8876) );
no02s04 g772004 ( .a(FE_OCP_RBN5779_n_44570), .b(n_10464), .o(n_8925) );
no02s02 g772005 ( .a(FE_OFN757_n_44464), .b(n_9478), .o(n_9695) );
no02s01 g772006 ( .a(n_8811), .b(n_44511), .o(n_11041) );
in01s01 g772007 ( .a(n_9281), .o(n_9282) );
na02s02 g772008 ( .a(FE_OCP_RBN5827_n_44579), .b(n_9220), .o(n_9281) );
in01s01 g772009 ( .a(n_9385), .o(n_9386) );
no02s02 g772010 ( .a(FE_OCP_RBN6730_n_44579), .b(n_9321), .o(n_9385) );
in01s01 g772011 ( .a(n_9431), .o(n_9432) );
na02s01 g772012 ( .a(FE_OCP_RBN5907_n_44563), .b(n_9381), .o(n_9431) );
in01s01 g772013 ( .a(n_9433), .o(n_9505) );
no02s01 g772014 ( .a(FE_OCP_RBN5907_n_44563), .b(n_9367), .o(n_9433) );
in01s01 g772015 ( .a(n_9874), .o(n_9824) );
na02s01 g772016 ( .a(FE_OFN4778_n_44490), .b(n_9768), .o(n_9874) );
in01s01 g772017 ( .a(n_9692), .o(n_9775) );
na02s01 g772018 ( .a(n_44492), .b(n_9647), .o(n_9692) );
in01s01 g772019 ( .a(n_9733), .o(n_9734) );
na02s01 g772020 ( .a(FE_OFN4775_n_44463), .b(n_9681), .o(n_9733) );
na02s02 g772021 ( .a(FE_OCPN1061_n_44460), .b(n_9321), .o(n_9475) );
no02s02 g772022 ( .a(FE_OCP_RBN5827_n_44579), .b(n_9220), .o(n_9309) );
na02m02 g772023 ( .a(FE_OCP_RBN6704_n_8762), .b(n_8561), .o(n_8798) );
na02m06 g772024 ( .a(n_8783), .b(FE_OCP_RBN2655_FE_OCPN914_n_8091), .o(n_8887) );
no02f04 g772025 ( .a(n_8711), .b(n_8560), .o(n_8751) );
na02s02 g772027 ( .a(n_8950), .b(n_47243), .o(n_9030) );
na02f04 g772028 ( .a(n_8782), .b(FE_OCP_RBN2656_FE_OCPN914_n_8091), .o(n_8860) );
ao12s01 g772029 ( .a(n_8081), .b(n_8852), .c(n_8110), .o(n_8932) );
ao12s01 g772030 ( .a(n_8085), .b(n_8824), .c(n_8031), .o(n_8868) );
ao12s01 g772031 ( .a(n_8151), .b(n_8900), .c(n_8172), .o(n_8962) );
ao12s01 g772032 ( .a(n_8773), .b(n_8824), .c(n_8772), .o(n_10078) );
ao12s02 g772033 ( .a(n_8651), .b(FE_OCP_RBN5825_n_8692), .c(FE_OCP_RBN4220_n_8594), .o(n_8815) );
na02s04 g772034 ( .a(FE_OCP_RBN5819_n_8651), .b(n_8793), .o(n_8825) );
oa12m04 g772035 ( .a(FE_OCP_RBN4219_n_8594), .b(n_8692), .c(n_8651), .o(n_8766) );
ao12s01 g772036 ( .a(n_8822), .b(n_8821), .c(n_8820), .o(n_10079) );
ao22m02 g772039 ( .a(FE_OCP_RBN5826_n_8692), .b(n_8775), .c(FE_OCP_RBN2854_n_8692), .d(n_8774), .o(n_8902) );
oa22s01 g772041 ( .a(n_8900), .b(n_8166), .c(n_8852), .d(n_8167), .o(n_10122) );
ao22m02 g772042 ( .a(n_8831), .b(FE_OCP_RBN5750_n_8599), .c(n_8599), .d(n_8832), .o(n_9004) );
no02s01 g772043 ( .a(n_8821), .b(n_8820), .o(n_8822) );
na02s02 g772045 ( .a(FE_OCP_RBN4220_n_8594), .b(FE_OCP_RBN5826_n_8692), .o(n_8793) );
in01s02 g772046 ( .a(n_8898), .o(n_8899) );
na02m02 g772047 ( .a(n_8770), .b(n_8858), .o(n_8898) );
no02s01 g772048 ( .a(n_8824), .b(n_8772), .o(n_8773) );
in01s02 g772049 ( .a(n_8998), .o(n_8999) );
na02s02 g772050 ( .a(FE_OCP_RBN5849_FE_RN_2187_0), .b(FE_OCP_RBN5847_FE_RN_987_0), .o(n_8998) );
in01s01 g772051 ( .a(n_47244), .o(n_8950) );
in01s03 g772053 ( .a(n_45503), .o(n_8700) );
ao12m04 g772054 ( .a(n_8531), .b(n_8471), .c(n_7594), .o(n_8532) );
in01s02 g772056 ( .a(n_8747), .o(n_8694) );
ao12f08 g772057 ( .a(n_7568), .b(n_8621), .c(n_7581), .o(n_8747) );
na02s01 TIMEBOOST_cell_2816 ( .a(FE_OCPN6913_n_1715), .b(n_1714), .o(TIMEBOOST_net_699) );
in01f02 g772203 ( .a(n_8857), .o(n_8895) );
na02f04 g772204 ( .a(n_8812), .b(n_8761), .o(n_8857) );
na02f04 g772206 ( .a(n_8641), .b(n_8633), .o(n_8739) );
in01m02 g772207 ( .a(n_8782), .o(n_8783) );
in01s01 g772217 ( .a(n_8765), .o(n_10105) );
in01m02 g772218 ( .a(n_8765), .o(n_8764) );
na02m04 g772219 ( .a(n_8622), .b(n_8668), .o(n_8765) );
in01m02 g772224 ( .a(n_8711), .o(n_8762) );
ao12f04 g772225 ( .a(n_8487), .b(n_8632), .c(n_8535), .o(n_8711) );
na02s02 g772229 ( .a(n_8621), .b(n_7609), .o(n_8622) );
na02s04 g772230 ( .a(FE_OCP_RBN4187_n_8621), .b(n_7610), .o(n_8668) );
in01s01 g772231 ( .a(n_8852), .o(n_8900) );
no02s01 g772232 ( .a(n_8144), .b(n_8734), .o(n_8852) );
na02f04 g772234 ( .a(n_8609), .b(FE_OCP_RBN4138_n_7743), .o(n_8678) );
na02s02 g772235 ( .a(n_8727), .b(n_8104), .o(n_8761) );
na02s04 g772236 ( .a(n_8608), .b(n_8104), .o(n_8633) );
na02m06 g772239 ( .a(n_8728), .b(FE_OCPN931_n_7817), .o(n_8799) );
in01f01 g772248 ( .a(n_8794), .o(n_8858) );
no02f04 g772249 ( .a(FE_OCPN917_n_8753), .b(FE_OCP_RBN6627_n_7832), .o(n_8794) );
in01s01 g772251 ( .a(n_8770), .o(n_8813) );
na02s06 g772252 ( .a(FE_OCPN917_n_8753), .b(FE_OCP_RBN6627_n_7832), .o(n_8770) );
oa12s01 g772253 ( .a(n_8045), .b(n_8760), .c(n_8038), .o(n_8821) );
no02f10 TIMEBOOST_cell_2815 ( .a(n_222), .b(TIMEBOOST_net_698), .o(n_244) );
in01s02 g772255 ( .a(n_8680), .o(n_8681) );
in01m01 g772256 ( .a(n_8641), .o(n_8680) );
na02m02 TIMEBOOST_cell_4064 ( .a(TIMEBOOST_net_1122), .b(n_4386), .o(n_4548) );
in01s02 g772258 ( .a(n_8831), .o(n_8832) );
in01f01 g772259 ( .a(n_8812), .o(n_8831) );
na02f04 g772260 ( .a(n_8729), .b(n_8730), .o(n_8812) );
oa12f06 g772266 ( .a(n_8590), .b(n_8585), .c(n_8642), .o(n_8692) );
ao12s01 g772268 ( .a(n_8113), .b(n_8684), .c(n_8048), .o(n_8824) );
ao22s01 g772269 ( .a(n_8760), .b(n_8087), .c(n_8690), .d(n_8086), .o(n_9994) );
in01s01 g772270 ( .a(n_8810), .o(n_8811) );
ao12s01 g772271 ( .a(n_8737), .b(n_8736), .c(n_8735), .o(n_8810) );
in01m02 g772272 ( .a(n_8809), .o(n_10464) );
oa22m02 g772274 ( .a(FE_OCP_RBN6691_n_8629), .b(n_8685), .c(n_8629), .d(n_8647), .o(n_8809) );
no02s01 g772275 ( .a(n_8736), .b(n_8735), .o(n_8737) );
in01s02 g772278 ( .a(n_8471), .o(n_8523) );
ao12f08 g772279 ( .a(n_7531), .b(n_8409), .c(n_7559), .o(n_8471) );
oa12f08 g772281 ( .a(n_7530), .b(n_8504), .c(n_7511), .o(n_8621) );
in01s01 g772282 ( .a(n_8733), .o(n_8734) );
in01f02 g772284 ( .a(n_8666), .o(n_8667) );
no02f04 g772285 ( .a(n_8576), .b(n_8545), .o(n_8666) );
oa12s01 g772286 ( .a(n_8723), .b(n_8722), .c(n_8721), .o(n_9913) );
ao12s01 g772288 ( .a(n_8708), .b(n_8707), .c(n_8706), .o(n_9939) );
no02m04 TIMEBOOST_cell_5576 ( .a(n_26724), .b(n_26333), .o(TIMEBOOST_net_1736) );
ao12f02 g772297 ( .a(n_8604), .b(n_8620), .c(FE_OCP_RBN4139_n_7743), .o(n_8730) );
ao12f04 g772301 ( .a(n_8478), .b(n_8492), .c(FE_OCPN931_n_7817), .o(n_8578) );
in01s01 g772303 ( .a(n_8562), .o(n_8610) );
in01s01 g772304 ( .a(n_8548), .o(n_8562) );
ao12s01 g772307 ( .a(n_8726), .b(n_8725), .c(n_8724), .o(n_9768) );
in01s02 g772308 ( .a(n_8653), .o(n_8654) );
in01m01 g772309 ( .a(n_8632), .o(n_8653) );
oa12m04 g772310 ( .a(n_8484), .b(n_8553), .c(n_8423), .o(n_8632) );
in01f02 g772312 ( .a(n_8727), .o(n_8728) );
in01m02 g772314 ( .a(n_8608), .o(n_8609) );
in01s01 g772316 ( .a(n_8760), .o(n_8690) );
in01s01 g772317 ( .a(n_8684), .o(n_8760) );
no02s01 g772319 ( .a(n_8725), .b(n_8724), .o(n_8726) );
na02s01 g772320 ( .a(n_8722), .b(n_8721), .o(n_8723) );
no02s01 g772321 ( .a(n_8706), .b(n_8707), .o(n_8708) );
no02s01 TIMEBOOST_cell_8771 ( .a(TIMEBOOST_net_2872), .b(n_14050), .o(n_16111) );
na02s02 g772323 ( .a(n_8491), .b(FE_OCP_RBN5634_n_7708), .o(n_8528) );
no02f02 g772324 ( .a(n_8332), .b(n_8507), .o(n_8576) );
na02s06 TIMEBOOST_cell_6644 ( .a(TIMEBOOST_net_2079), .b(FE_OCP_RBN4113_n_33533), .o(n_33627) );
no02s02 g772326 ( .a(n_8511), .b(n_8574), .o(n_8587) );
na02s02 g772328 ( .a(n_8660), .b(n_8682), .o(n_8719) );
na02s02 g772330 ( .a(n_8771), .b(FE_OCP_RBN2864_n_8714), .o(n_8806) );
na02f04 g772331 ( .a(n_8660), .b(n_8561), .o(n_8661) );
no02f04 g772333 ( .a(n_8659), .b(n_8628), .o(n_8755) );
oa12s01 g772334 ( .a(n_8718), .b(n_8717), .c(n_8716), .o(n_9647) );
ao12s01 g772335 ( .a(n_8082), .b(n_8656), .c(n_7916), .o(n_8736) );
in01s01 g772336 ( .a(n_8688), .o(n_8689) );
ao12s01 g772337 ( .a(n_8607), .b(n_8606), .c(n_8605), .o(n_8688) );
ao12s01 g772342 ( .a(n_8589), .b(n_8613), .c(n_8588), .o(n_9767) );
in01s01 g772344 ( .a(n_8585), .o(n_8629) );
oa12m06 g772345 ( .a(n_8555), .b(n_44058), .c(n_8482), .o(n_8585) );
in01m02 g772346 ( .a(n_8434), .o(n_8435) );
in01s02 g772347 ( .a(n_8409), .o(n_8434) );
oa12f08 g772348 ( .a(n_7536), .b(n_8304), .c(n_7502), .o(n_8409) );
in01s02 g772349 ( .a(n_8546), .o(n_8547) );
in01m02 g772350 ( .a(n_8504), .o(n_8546) );
ao12m08 g772351 ( .a(n_7466), .b(n_8407), .c(n_7501), .o(n_8504) );
no02s01 g772352 ( .a(n_8606), .b(n_8605), .o(n_8607) );
no02s01 g772353 ( .a(n_8613), .b(n_8588), .o(n_8589) );
na02s01 g772354 ( .a(n_8717), .b(n_8716), .o(n_8718) );
no02f02 g772355 ( .a(n_8627), .b(n_8596), .o(n_8659) );
na02f04 g772356 ( .a(n_8477), .b(n_8413), .o(n_8478) );
na02m02 g772357 ( .a(n_8603), .b(n_8626), .o(n_8628) );
na02m02 g772358 ( .a(n_8603), .b(n_8515), .o(n_8604) );
na02s02 g772359 ( .a(n_8521), .b(n_8477), .o(n_8545) );
no02s04 g772361 ( .a(n_8677), .b(FE_OCP_RBN6580_n_8676), .o(n_8714) );
na02m04 g772363 ( .a(n_8627), .b(n_8626), .o(n_8657) );
na02f02 g772364 ( .a(n_8571), .b(n_7957), .o(n_8660) );
na02s04 g772365 ( .a(n_8677), .b(FE_OCP_RBN6580_n_8676), .o(n_8771) );
na02s06 g772366 ( .a(n_8572), .b(n_7941), .o(n_8682) );
oa12s01 g772367 ( .a(n_8105), .b(n_8573), .c(n_7996), .o(n_8722) );
no02s02 TIMEBOOST_cell_1904 ( .a(TIMEBOOST_net_566), .b(n_27119), .o(n_27234) );
oa12s01 g772369 ( .a(n_7955), .b(n_8519), .c(n_7997), .o(n_8725) );
in01f02 g772370 ( .a(n_8506), .o(n_8507) );
ao12m04 g772371 ( .a(n_8440), .b(n_8411), .c(FE_OCPN935_n_7802), .o(n_8506) );
in01m02 g772372 ( .a(n_8601), .o(n_8602) );
no02f04 g772373 ( .a(n_8441), .b(n_8522), .o(n_8601) );
in01s02 g772374 ( .a(n_8574), .o(n_8575) );
in01s01 g772375 ( .a(n_8553), .o(n_8574) );
oa12m06 g772376 ( .a(n_8340), .b(n_8392), .c(n_8460), .o(n_8553) );
in01s03 g772377 ( .a(n_46990), .o(n_10374) );
in01s01 g772386 ( .a(n_8499), .o(n_8554) );
in01s01 g772387 ( .a(n_8498), .o(n_8499) );
in01m02 g772388 ( .a(n_8498), .o(n_8465) );
in01f02 g772393 ( .a(n_8491), .o(n_8492) );
ao22f02 g772394 ( .a(n_8380), .b(FE_OCP_RBN5634_n_7708), .c(n_8379), .d(FE_OCPN931_n_7817), .o(n_8491) );
in01s02 g772395 ( .a(n_8619), .o(n_8620) );
in01s01 TIMEBOOST_cell_5908 ( .a(TIMEBOOST_net_1796), .o(TIMEBOOST_net_1797) );
no02s01 g772397 ( .a(n_8518), .b(n_8027), .o(n_8606) );
no02f08 g772398 ( .a(n_8517), .b(n_8550), .o(n_8613) );
no02s01 g772399 ( .a(n_8015), .b(n_8573), .o(n_8656) );
na02m02 g772400 ( .a(n_8525), .b(FE_OCP_RBN4139_n_7743), .o(n_8603) );
no02f04 TIMEBOOST_cell_7840 ( .a(n_38662), .b(n_45192), .o(TIMEBOOST_net_2551) );
no04s04 TIMEBOOST_cell_8192 ( .a(n_12281), .b(FE_RN_796_0), .c(FE_RN_797_0), .d(delay_sub_ln23_0_unr8_stage4_stallmux_q_29_), .o(FE_RN_800_0) );
in01s01 g772403 ( .a(n_8595), .o(n_8596) );
na02m04 g772404 ( .a(n_8526), .b(FE_OCPN935_n_7802), .o(n_8595) );
na02f04 g772405 ( .a(n_8410), .b(FE_OCP_RBN4139_n_7743), .o(n_8477) );
in01m02 g772406 ( .a(n_8521), .o(n_8522) );
no02m04 g772407 ( .a(n_8414), .b(FE_OCP_RBN6663_n_8355), .o(n_8521) );
na02f04 g772408 ( .a(n_8420), .b(n_8540), .o(n_8627) );
na02s02 g772409 ( .a(n_8421), .b(n_8466), .o(n_8520) );
no02s02 g772410 ( .a(n_8440), .b(n_8332), .o(n_8441) );
in01s02 g772411 ( .a(n_8670), .o(n_8671) );
na02s02 g772412 ( .a(n_8508), .b(n_8561), .o(n_8670) );
no02f02 g772415 ( .a(n_8530), .b(FE_OCP_RBN5742_n_8540), .o(n_8584) );
in01s01 g772416 ( .a(n_8774), .o(n_8775) );
na02s02 g772417 ( .a(FE_OCP_RBN5819_n_8651), .b(FE_OCP_RBN4220_n_8594), .o(n_8774) );
oa12s01 g772418 ( .a(n_7889), .b(n_8503), .c(n_7922), .o(n_8717) );
ao12s01 g772419 ( .a(n_8495), .b(n_8503), .c(n_8494), .o(n_9681) );
in01s01 g772422 ( .a(n_44058), .o(n_8542) );
in01s02 g772424 ( .a(n_8571), .o(n_8572) );
oa22f02 g772425 ( .a(FE_OCP_RBN6680_n_8448), .b(n_8221), .c(FE_OCP_RBN2690_n_8221), .d(n_8448), .o(n_8571) );
ao12s01 g772426 ( .a(n_8640), .b(n_8639), .c(n_8638), .o(n_9598) );
in01s01 g772427 ( .a(n_8518), .o(n_8519) );
no02s01 g772428 ( .a(n_8503), .b(n_7952), .o(n_8518) );
no02s01 g772429 ( .a(n_8639), .b(n_8638), .o(n_8640) );
no02s01 g772430 ( .a(n_8503), .b(n_8494), .o(n_8495) );
no02s02 g772435 ( .a(n_8580), .b(n_7900), .o(n_8594) );
in01s04 g772439 ( .a(n_8508), .o(n_8560) );
na02f04 g772440 ( .a(n_8489), .b(FE_OCP_RBN6604_n_7881), .o(n_8508) );
in01s01 g772441 ( .a(n_8496), .o(n_8497) );
no02s01 g772442 ( .a(n_8443), .b(FE_OCP_RBN5700_n_45828), .o(n_8496) );
na02m06 g772450 ( .a(n_8490), .b(FE_OCP_RBN6605_n_7881), .o(n_8561) );
oa12m06 g772451 ( .a(n_8406), .b(n_8354), .c(n_45212), .o(n_8407) );
ao12f06 g772452 ( .a(n_8303), .b(n_8231), .c(n_8302), .o(n_8304) );
oa12m06 g772453 ( .a(n_45213), .b(n_8387), .c(n_7464), .o(n_8476) );
ao12s04 g772454 ( .a(n_45212), .b(n_8386), .c(n_8406), .o(n_8461) );
in01m02 g772455 ( .a(n_8381), .o(n_8382) );
oa12m04 g772456 ( .a(n_8302), .b(FE_OCP_RBN6657_n_44352), .c(n_8303), .o(n_8381) );
in01s01 g772457 ( .a(n_8517), .o(n_8573) );
no02f08 g772458 ( .a(n_8503), .b(n_8061), .o(n_8517) );
ao12f02 g772460 ( .a(n_8398), .b(n_8462), .c(FE_OCP_RBN4139_n_7743), .o(n_8515) );
oa12m04 g772461 ( .a(n_8326), .b(n_8385), .c(FE_OCP_RBN2597_n_7743), .o(n_8440) );
no02f02 TIMEBOOST_cell_3228 ( .a(n_20282), .b(n_20321), .o(TIMEBOOST_net_905) );
in01m02 g772464 ( .a(n_8413), .o(n_8414) );
ao12m04 g772465 ( .a(n_8306), .b(n_8385), .c(FE_OCPN931_n_7817), .o(n_8413) );
in01m01 g772467 ( .a(n_8460), .o(n_8466) );
oa12m06 g772468 ( .a(n_8263), .b(n_8403), .c(n_8313), .o(n_8460) );
oa12s01 g772469 ( .a(n_8470), .b(n_8469), .c(n_8468), .o(n_9544) );
in01s01 g772470 ( .a(n_10214), .o(n_8514) );
no03s08 TIMEBOOST_cell_7165 ( .a(n_7785), .b(n_7676), .c(TIMEBOOST_net_2086), .o(n_7974) );
in01s01 g772474 ( .a(FE_OCPN1084_n_8388), .o(n_8750) );
in01s01 g772475 ( .a(n_8380), .o(n_8388) );
in01m02 g772476 ( .a(n_8380), .o(n_8379) );
in01s02 g772478 ( .a(n_10137), .o(n_8539) );
na02s06 g772479 ( .a(n_8415), .b(n_8464), .o(n_10137) );
ao12s01 g772486 ( .a(n_8650), .b(n_8649), .c(n_8648), .o(n_9631) );
in01s02 g772487 ( .a(n_8525), .o(n_8526) );
in01m02 g772489 ( .a(n_8410), .o(n_8411) );
na02s01 g772491 ( .a(n_8469), .b(n_8468), .o(n_8470) );
no02s01 g772492 ( .a(n_8649), .b(n_8648), .o(n_8650) );
no02s02 TIMEBOOST_cell_2075 ( .a(n_39089), .b(FE_OCP_RBN4180_n_38592), .o(TIMEBOOST_net_652) );
no02s01 g772494 ( .a(n_8617), .b(n_8642), .o(n_8647) );
na02s01 g772495 ( .a(n_8591), .b(n_8590), .o(n_8685) );
na02s01 g772496 ( .a(n_8400), .b(n_8292), .o(n_8415) );
na02s02 g772497 ( .a(n_8401), .b(n_8291), .o(n_8464) );
na02s02 g772498 ( .a(n_8509), .b(n_8535), .o(n_8536) );
no02s02 g772499 ( .a(n_8487), .b(n_8488), .o(n_8570) );
no02m06 g772500 ( .a(n_8374), .b(n_45827), .o(n_8443) );
na02s01 g772501 ( .a(n_8344), .b(n_8403), .o(n_8404) );
no02m06 TIMEBOOST_cell_5004 ( .a(n_37707), .b(n_37709), .o(TIMEBOOST_net_1450) );
ao12f08 g772503 ( .a(n_8010), .b(n_8369), .c(n_7989), .o(n_8503) );
in01m02 g772504 ( .a(n_8533), .o(n_8534) );
no02m04 g772505 ( .a(n_8456), .b(n_8457), .o(n_8533) );
no02f04 g772507 ( .a(n_8378), .b(n_8365), .o(n_8448) );
ao12s01 g772508 ( .a(n_8432), .b(n_8431), .c(n_8430), .o(n_9587) );
oa12s01 g772509 ( .a(n_8028), .b(n_8433), .c(n_7988), .o(n_8639) );
in01f02 g772510 ( .a(n_8489), .o(n_8490) );
oa12s01 g772512 ( .a(n_8646), .b(n_8645), .c(n_8644), .o(n_9478) );
na02s01 g772515 ( .a(n_8433), .b(n_8009), .o(n_8469) );
no02s01 g772516 ( .a(n_8431), .b(n_8430), .o(n_8432) );
na02s01 g772517 ( .a(n_8645), .b(n_8644), .o(n_8646) );
na02m04 g772518 ( .a(n_8307), .b(n_8355), .o(n_8365) );
no02m04 g772519 ( .a(n_8332), .b(n_8327), .o(n_8378) );
na02s04 g772520 ( .a(n_8395), .b(FE_OCP_RBN2740_n_8398), .o(n_8457) );
no02s02 g772521 ( .a(n_8419), .b(n_8455), .o(n_8456) );
in01s01 g772522 ( .a(n_8535), .o(n_8488) );
na02m04 g772523 ( .a(n_8454), .b(n_8453), .o(n_8535) );
in01s01 g772525 ( .a(n_8487), .o(n_8509) );
no02s04 g772526 ( .a(n_8454), .b(n_8453), .o(n_8487) );
in01s01 g772528 ( .a(n_8590), .o(n_8617) );
na02m03 g772529 ( .a(n_8569), .b(n_8568), .o(n_8590) );
in01s01 g772530 ( .a(n_8642), .o(n_8591) );
no02m04 g772531 ( .a(n_8569), .b(n_8568), .o(n_8642) );
oa12f08 g772535 ( .a(n_7492), .b(n_8186), .c(n_7460), .o(n_8231) );
in01s04 g772537 ( .a(n_8386), .o(n_8387) );
in01m04 g772538 ( .a(n_8376), .o(n_8386) );
in01m02 g772539 ( .a(n_8354), .o(n_8376) );
ao12f08 g772540 ( .a(n_7411), .b(n_8261), .c(n_7444), .o(n_8354) );
oa12s01 g772541 ( .a(n_7928), .b(n_8337), .c(n_7914), .o(n_8649) );
oa12s01 g772548 ( .a(n_8558), .b(n_8557), .c(n_8556), .o(n_9367) );
oa12s01 g772549 ( .a(n_8373), .b(n_8372), .c(n_8371), .o(n_9381) );
in01s01 g772556 ( .a(n_8403), .o(n_8375) );
in01s01 g772558 ( .a(n_8428), .o(n_8429) );
oa12s01 g772559 ( .a(n_8353), .b(n_8352), .c(n_8351), .o(n_8428) );
in01s01 g772560 ( .a(n_8400), .o(n_8401) );
in01s01 g772561 ( .a(n_8374), .o(n_8400) );
ao12m04 g772562 ( .a(n_8216), .b(n_8256), .c(n_8182), .o(n_8374) );
in01s01 g772563 ( .a(n_8426), .o(n_8427) );
oa12s01 g772564 ( .a(n_8360), .b(n_8359), .c(n_8358), .o(n_8426) );
oa22f02 g772565 ( .a(n_8321), .b(FE_OCP_RBN4141_n_7743), .c(n_8322), .d(FE_OCP_RBN4159_FE_OCPN857_n_7802), .o(n_8462) );
na02m06 g772566 ( .a(n_8248), .b(n_8277), .o(n_8385) );
na02s01 g772567 ( .a(n_8372), .b(n_8371), .o(n_8373) );
na02s01 g772568 ( .a(n_8557), .b(n_8556), .o(n_8558) );
no02s01 g772569 ( .a(n_8324), .b(n_7927), .o(n_8431) );
in01s01 g772570 ( .a(n_8326), .o(n_8327) );
na02s04 g772571 ( .a(n_8296), .b(FE_OCP_RBN2616_FE_OCPN857_n_7802), .o(n_8326) );
na02m06 g772572 ( .a(FE_OCP_RBN2690_n_8221), .b(FE_OCPN861_n_7743), .o(n_8277) );
na02s02 g772573 ( .a(n_8221), .b(FE_OCP_RBN5609_n_7730), .o(n_8248) );
no02m02 g772575 ( .a(n_8335), .b(FE_OCP_RBN5632_n_7708), .o(n_8398) );
in01s01 g772576 ( .a(n_8306), .o(n_8307) );
no02s04 g772577 ( .a(n_8296), .b(FE_OCP_RBN2616_FE_OCPN857_n_7802), .o(n_8306) );
no02f04 g772578 ( .a(n_8336), .b(FE_OCP_RBN4141_n_7743), .o(n_8455) );
na02s01 g772579 ( .a(n_8359), .b(n_8358), .o(n_8360) );
na02s01 g772580 ( .a(n_8352), .b(n_8351), .o(n_8353) );
in01s01 g772581 ( .a(n_8566), .o(n_8567) );
na02s02 g772582 ( .a(n_8483), .b(n_8555), .o(n_8566) );
no02f06 g772584 ( .a(n_8437), .b(n_8396), .o(n_8530) );
in01m02 g772585 ( .a(n_8439), .o(n_8370) );
na02m06 g772586 ( .a(n_8332), .b(n_8355), .o(n_8439) );
in01m02 g772587 ( .a(n_8511), .o(n_8512) );
na02m02 g772588 ( .a(n_8484), .b(n_8424), .o(n_8511) );
in01s01 g772589 ( .a(n_8369), .o(n_8433) );
oa12s01 g772591 ( .a(n_7831), .b(n_8305), .c(n_7858), .o(n_8645) );
na02m04 TIMEBOOST_cell_2936 ( .a(n_41447), .b(n_41382), .o(TIMEBOOST_net_759) );
na02m04 g772593 ( .a(n_8425), .b(n_8450), .o(n_8569) );
na02s01 g772594 ( .a(n_8305), .b(n_7860), .o(n_8372) );
na02s04 g772595 ( .a(FE_OCP_RBN2701_n_8187), .b(n_8394), .o(n_8450) );
no02m06 TIMEBOOST_cell_4266 ( .a(n_33849), .b(TIMEBOOST_net_1223), .o(n_33873) );
na02s01 TIMEBOOST_cell_4936 ( .a(n_7077), .b(n_7150), .o(TIMEBOOST_net_1416) );
na02s02 g772598 ( .a(n_8393), .b(FE_OCP_RBN6656_n_8187), .o(n_8425) );
in01m01 g772599 ( .a(n_8482), .o(n_8483) );
no02m06 g772600 ( .a(n_8445), .b(FE_OCPN1618_n_8444), .o(n_8482) );
in01m01 g772601 ( .a(n_8423), .o(n_8424) );
no02f02 g772602 ( .a(n_8390), .b(n_8389), .o(n_8423) );
na02s06 g772603 ( .a(n_8445), .b(FE_OCPN1618_n_8444), .o(n_8555) );
na02s02 g772604 ( .a(n_8390), .b(n_8389), .o(n_8484) );
no02m01 g772606 ( .a(n_8392), .b(n_8293), .o(n_8421) );
in01s02 g772607 ( .a(n_8294), .o(n_8295) );
in01s02 g772608 ( .a(n_8261), .o(n_8294) );
oa12m08 g772609 ( .a(n_7423), .b(n_8191), .c(n_7384), .o(n_8261) );
in01s02 g772610 ( .a(n_8206), .o(n_8207) );
in01s02 g772611 ( .a(n_8186), .o(n_8206) );
ao12s01 g772613 ( .a(n_7697), .b(n_8289), .c(n_7827), .o(n_8557) );
in01s01 g772614 ( .a(n_8337), .o(n_8324) );
na02f08 g772615 ( .a(n_8283), .b(n_7859), .o(n_8337) );
in01s01 g772616 ( .a(n_8419), .o(n_8420) );
in01s02 g772617 ( .a(n_8396), .o(n_8419) );
no02f08 g772618 ( .a(n_8320), .b(n_8368), .o(n_8396) );
no02s06 g772620 ( .a(n_8230), .b(n_8219), .o(n_8355) );
na02m08 g772624 ( .a(FE_OCP_RBN2722_n_8243), .b(n_8250), .o(n_8332) );
in01s01 g772625 ( .a(n_8437), .o(n_8395) );
na02m06 g772626 ( .a(n_8319), .b(n_8364), .o(n_8437) );
na02s01 g772628 ( .a(n_8252), .b(n_8170), .o(n_8352) );
oa12m04 g772629 ( .a(n_8224), .b(n_8255), .c(n_8123), .o(n_8256) );
oa12s01 g772630 ( .a(n_8274), .b(n_8275), .c(n_8273), .o(n_9988) );
na02s01 g772631 ( .a(n_8225), .b(n_8145), .o(n_8359) );
oa12s01 g772637 ( .a(n_8282), .b(n_8289), .c(n_8281), .o(n_9369) );
in01s01 g772639 ( .a(n_8348), .o(n_8366) );
in01s01 g772640 ( .a(n_8321), .o(n_8348) );
in01m02 g772641 ( .a(n_8321), .o(n_8322) );
oa12s01 g772643 ( .a(n_8246), .b(n_8255), .c(n_8245), .o(n_10028) );
no02s01 TIMEBOOST_cell_6649 ( .a(FE_OCP_RBN4103_n_12880), .b(FE_OCP_RBN4097_n_12880), .o(TIMEBOOST_net_2082) );
in01m02 g772645 ( .a(n_8335), .o(n_8336) );
na02s01 g772647 ( .a(n_8289), .b(n_8281), .o(n_8282) );
in01m02 g772648 ( .a(n_8393), .o(n_8394) );
na02m04 g772649 ( .a(n_8368), .b(n_8364), .o(n_8393) );
in01s02 g772650 ( .a(n_8284), .o(n_8285) );
na02f02 g772651 ( .a(n_8243), .b(n_8220), .o(n_8284) );
na02s02 g772652 ( .a(n_8229), .b(FE_OCP_RBN4161_FE_OCPN857_n_7802), .o(n_8250) );
no02m04 g772653 ( .a(n_8318), .b(FE_OCP_RBN4141_n_7743), .o(n_8320) );
na02m04 g772654 ( .a(n_8318), .b(FE_OCP_RBN4141_n_7743), .o(n_8319) );
no02s02 g772655 ( .a(n_8229), .b(FE_OCP_RBN4162_FE_OCPN857_n_7802), .o(n_8230) );
na02s03 TIMEBOOST_cell_4076 ( .a(n_31314), .b(TIMEBOOST_net_1128), .o(n_31456) );
na02f04 TIMEBOOST_cell_8787 ( .a(TIMEBOOST_net_2880), .b(n_15022), .o(n_15198) );
na02s01 g772658 ( .a(n_8275), .b(n_8273), .o(n_8274) );
in01s02 g772660 ( .a(n_8293), .o(n_8340) );
no02s02 g772661 ( .a(n_8271), .b(FE_OCPN6919_n_7726), .o(n_8293) );
in01s01 g772662 ( .a(n_46418), .o(n_8367) );
na02m06 g772666 ( .a(n_8346), .b(n_45828), .o(n_8316) );
na02s01 g772667 ( .a(n_8255), .b(n_8245), .o(n_8246) );
na02s01 g772668 ( .a(n_8275), .b(n_8251), .o(n_8252) );
na02s01 g772669 ( .a(n_8255), .b(n_8224), .o(n_8225) );
in01s01 g772670 ( .a(n_8283), .o(n_8305) );
no02s01 TIMEBOOST_cell_4263 ( .a(n_18032), .b(n_18010), .o(TIMEBOOST_net_1222) );
na02s01 TIMEBOOST_cell_5248 ( .a(n_26605), .b(FE_OCP_RBN6858_n_26160), .o(TIMEBOOST_net_1572) );
ao12s01 g772674 ( .a(n_8481), .b(n_8480), .c(n_8479), .o(n_9321) );
no02s01 g772675 ( .a(n_8480), .b(n_8479), .o(n_8481) );
in01s01 g772676 ( .a(n_8215), .o(n_8289) );
in01s01 g772678 ( .a(n_8344), .o(n_8345) );
no02s01 g772679 ( .a(n_8264), .b(n_8313), .o(n_8344) );
no02s01 TIMEBOOST_cell_5122 ( .a(n_4093), .b(FE_OFN4765_n_3029), .o(TIMEBOOST_net_1509) );
no02s02 g772681 ( .a(n_8300), .b(FE_OCP_RBN6644_n_8342), .o(n_8315) );
na02s06 g772682 ( .a(n_8236), .b(FE_OFN4701_n_7702), .o(n_8493) );
na02m04 g772683 ( .a(n_8235), .b(n_7728), .o(n_8346) );
na03m06 TIMEBOOST_cell_8353 ( .a(n_15395), .b(n_15266), .c(TIMEBOOST_net_1272), .o(n_15595) );
na02s02 g772685 ( .a(n_8237), .b(n_8269), .o(n_8270) );
in01s02 g772687 ( .a(n_8101), .o(n_8111) );
oa12m06 g772688 ( .a(n_7432), .b(n_7986), .c(n_7395), .o(n_8101) );
in01s01 g772689 ( .a(n_8211), .o(n_8212) );
in01s02 g772690 ( .a(n_8191), .o(n_8211) );
ao12m08 g772691 ( .a(n_7349), .b(n_8106), .c(n_7382), .o(n_8191) );
no02s06 TIMEBOOST_cell_2898 ( .a(n_13412), .b(n_12634), .o(TIMEBOOST_net_740) );
in01s02 g772694 ( .a(n_8219), .o(n_8220) );
na02s03 g772695 ( .a(n_8162), .b(FE_OCP_RBN2702_FE_RN_299_0), .o(n_8219) );
na02m08 g772696 ( .a(n_8268), .b(n_8259), .o(n_8368) );
no02s02 TIMEBOOST_cell_5927 ( .a(n_36151), .b(n_35989), .o(TIMEBOOST_net_1815) );
ao12m06 g772698 ( .a(n_8052), .b(n_8197), .c(n_8122), .o(n_8255) );
ao12m04 g772699 ( .a(n_8102), .b(n_8204), .c(n_8158), .o(n_8275) );
in01s01 g772711 ( .a(n_8239), .o(n_8240) );
oa12s01 g772712 ( .a(n_8181), .b(n_8180), .c(n_8197), .o(n_8239) );
ao12s01 g772715 ( .a(n_8193), .b(n_8192), .c(n_8204), .o(n_9906) );
na02s02 TIMEBOOST_cell_2844 ( .a(n_7146), .b(n_7147), .o(TIMEBOOST_net_713) );
na02s02 TIMEBOOST_cell_4075 ( .a(n_31393), .b(n_31394), .o(TIMEBOOST_net_1128) );
na02m02 g772718 ( .a(n_8195), .b(FE_OCP_RBN2634_n_9003), .o(n_8196) );
na02s08 TIMEBOOST_cell_4074 ( .a(TIMEBOOST_net_1127), .b(n_30564), .o(n_46959) );
na02s02 g772720 ( .a(n_8107), .b(FE_OCP_RBN5609_n_7730), .o(n_8162) );
na02s06 TIMEBOOST_cell_2843 ( .a(n_7507), .b(TIMEBOOST_net_712), .o(n_7560) );
na02m06 g772722 ( .a(n_8266), .b(FE_OCP_RBN4137_n_7743), .o(n_8268) );
no02m06 TIMEBOOST_cell_2897 ( .a(TIMEBOOST_net_739), .b(n_29145), .o(n_29262) );
na02s02 TIMEBOOST_cell_4182 ( .a(TIMEBOOST_net_1181), .b(n_22601), .o(n_22682) );
no02s03 TIMEBOOST_cell_6619 ( .a(n_32857), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_15_), .o(TIMEBOOST_net_2067) );
no03f08 TIMEBOOST_cell_8237 ( .a(n_18564), .b(n_18437), .c(n_17661), .o(n_18681) );
na02s01 g772727 ( .a(n_8180), .b(n_8197), .o(n_8181) );
no02s03 g772728 ( .a(n_8227), .b(n_8226), .o(n_8313) );
no02m04 g772730 ( .a(n_8259), .b(n_8258), .o(n_8300) );
in01s01 g772731 ( .a(n_8263), .o(n_8264) );
na02s04 g772732 ( .a(n_8227), .b(n_8226), .o(n_8263) );
in01s01 g772733 ( .a(n_8291), .o(n_8292) );
no02s01 g772734 ( .a(FE_OCP_RBN5700_n_45828), .b(n_45827), .o(n_8291) );
in01m01 g772735 ( .a(n_8237), .o(n_8238) );
no02m02 g772736 ( .a(FE_RN_299_0), .b(n_8213), .o(n_8237) );
no02s01 g772737 ( .a(n_8204), .b(n_8192), .o(n_8193) );
oa12s01 g772738 ( .a(n_7830), .b(n_8169), .c(n_7740), .o(n_8480) );
ao12s01 g772739 ( .a(n_8161), .b(n_8169), .c(n_8160), .o(n_9220) );
in01m02 g772740 ( .a(n_8235), .o(n_8236) );
in01s01 TIMEBOOST_cell_7374 ( .a(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_2310) );
no02m02 g772742 ( .a(n_8133), .b(n_47240), .o(n_8195) );
na02s01 TIMEBOOST_cell_8845 ( .a(TIMEBOOST_net_2909), .b(n_42970), .o(TIMEBOOST_net_2610) );
no02m06 TIMEBOOST_cell_5257 ( .a(n_20238), .b(TIMEBOOST_net_1576), .o(n_20325) );
no02s01 g772746 ( .a(n_8169), .b(n_8160), .o(n_8161) );
no02s01 g772750 ( .a(n_8234), .b(FE_RN_976_0), .o(n_8351) );
no02s01 g772751 ( .a(n_8216), .b(n_8183), .o(n_8358) );
in01s01 g772753 ( .a(n_8106), .o(n_8138) );
oa12m08 g772754 ( .a(FE_OCPN4524_n_7360), .b(n_8042), .c(n_7307), .o(n_8106) );
in01s02 g772755 ( .a(n_8043), .o(n_8044) );
in01s01 g772756 ( .a(n_7986), .o(n_8043) );
ao12m06 g772757 ( .a(n_7368), .b(n_7905), .c(n_7403), .o(n_7986) );
no02s04 g772758 ( .a(n_8134), .b(n_8078), .o(n_8213) );
oa12m06 g772759 ( .a(n_8094), .b(n_8155), .c(FE_OCP_RBN5614_n_7730), .o(n_8258) );
no02s06 g772760 ( .a(n_8095), .b(n_8177), .o(n_8259) );
na02m04 g772763 ( .a(n_8109), .b(n_47242), .o(n_8227) );
oa12m04 g772764 ( .a(n_8039), .b(n_8140), .c(n_8084), .o(n_8204) );
ao12s01 g772765 ( .a(n_8098), .b(n_8097), .c(n_8096), .o(n_9223) );
oa12s01 g772766 ( .a(n_8142), .b(n_8141), .c(n_8140), .o(n_9790) );
na03m08 TIMEBOOST_cell_5738 ( .a(n_19154), .b(n_18427), .c(FE_OCP_RBN3711_n_19116), .o(n_19270) );
oa12s01 g772769 ( .a(n_8126), .b(n_8125), .c(n_8124), .o(n_9784) );
oa12m06 g772775 ( .a(n_8054), .b(n_8057), .c(n_8006), .o(n_8197) );
no02f08 TIMEBOOST_cell_2070 ( .a(TIMEBOOST_net_649), .b(n_42098), .o(n_42128) );
in01m02 g772777 ( .a(n_8107), .o(n_8108) );
no02s02 g772779 ( .a(FE_OCP_RBN6622_n_7943), .b(n_7414), .o(n_7990) );
no02s01 TIMEBOOST_cell_8502 ( .a(n_7608), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_), .o(TIMEBOOST_net_2738) );
no02s01 g772781 ( .a(n_8097), .b(n_8096), .o(n_8098) );
in01s02 g772782 ( .a(n_8127), .o(n_8128) );
na02s04 g772783 ( .a(n_8095), .b(n_8094), .o(n_8127) );
no02s02 g772784 ( .a(n_8154), .b(FE_OCP_RBN6601_n_7708), .o(n_8177) );
no02s06 g772785 ( .a(FE_OCP_RBN6643_n_8342), .b(FE_OCPN849_n_7712), .o(n_8176) );
in01s01 g772786 ( .a(n_8093), .o(n_8169) );
oa12f06 g772787 ( .a(n_7760), .b(n_8041), .c(n_7757), .o(n_8093) );
no02s02 g772788 ( .a(n_8077), .b(FE_OCP_RBN6601_n_7708), .o(n_8078) );
no03m04 TIMEBOOST_cell_8214 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_), .b(n_23606), .c(n_23629), .o(n_23775) );
na02s02 g772791 ( .a(n_8175), .b(n_8174), .o(n_8208) );
no02s01 g772793 ( .a(FE_RN_974_0), .b(n_8159), .o(n_8273) );
in01s01 g772794 ( .a(n_8182), .o(n_8183) );
na02s04 g772795 ( .a(n_8136), .b(n_8135), .o(n_8182) );
no02s02 g772796 ( .a(n_8175), .b(n_8174), .o(n_8234) );
no02s03 g772797 ( .a(n_8136), .b(n_8135), .o(n_8216) );
na02s01 g772798 ( .a(n_8125), .b(n_8124), .o(n_8126) );
no02s01 g772799 ( .a(n_8123), .b(n_8121), .o(n_8245) );
na02m02 g772800 ( .a(FE_OCP_RBN2649_n_8073), .b(FE_OCP_RBN2609_n_47235), .o(n_8109) );
na02s01 g772801 ( .a(n_8141), .b(n_8140), .o(n_8142) );
in01s01 g772802 ( .a(n_8133), .o(n_8134) );
no02m04 g772803 ( .a(n_8073), .b(n_47241), .o(n_8133) );
na02s02 TIMEBOOST_cell_5254 ( .a(n_3506), .b(FE_OCP_RBN5770_n_3338), .o(TIMEBOOST_net_1575) );
no02s01 g772805 ( .a(n_8041), .b(n_7782), .o(n_8097) );
in01s01 g772807 ( .a(n_8159), .o(n_8170) );
no02s02 g772808 ( .a(n_8115), .b(n_8114), .o(n_8159) );
in01s01 g772809 ( .a(n_8224), .o(n_8121) );
na02s03 g772810 ( .a(n_8100), .b(FE_OCPN4526_n_8099), .o(n_8224) );
na02s01 g772811 ( .a(n_8103), .b(n_8158), .o(n_8192) );
in01s01 g772813 ( .a(n_8123), .o(n_8145) );
no02s04 g772814 ( .a(n_8100), .b(n_8099), .o(n_8123) );
na02m02 g772817 ( .a(n_8115), .b(n_8114), .o(n_8251) );
na02s01 g772818 ( .a(n_8122), .b(n_8053), .o(n_8180) );
no02s06 TIMEBOOST_cell_5253 ( .a(TIMEBOOST_net_1574), .b(n_3437), .o(n_3598) );
in01s02 g772820 ( .a(n_8074), .o(n_8075) );
in01s02 g772821 ( .a(n_8042), .o(n_8074) );
ao12m08 g772822 ( .a(n_7301), .b(n_7949), .c(n_7326), .o(n_8042) );
in01s01 g772824 ( .a(n_7905), .o(n_7943) );
oa12m08 g772825 ( .a(n_7371), .b(n_7798), .c(n_7341), .o(n_7905) );
ao12m06 g772828 ( .a(FE_OCP_RBN4075_n_7708), .b(n_7959), .c(FE_OCP_RBN6582_n_8021), .o(n_8073) );
ao12s01 g772830 ( .a(n_8065), .b(n_8064), .c(n_8063), .o(n_9642) );
na02s10 TIMEBOOST_cell_4211 ( .a(n_32732), .b(n_32665), .o(TIMEBOOST_net_1196) );
na02m06 TIMEBOOST_cell_4253 ( .a(n_13388), .b(FE_OCP_RBN4112_n_12880), .o(TIMEBOOST_net_1217) );
ao12m04 g772833 ( .a(n_7987), .b(n_7966), .c(n_7931), .o(n_8140) );
na02s02 TIMEBOOST_cell_1967 ( .a(n_37056), .b(n_37561), .o(TIMEBOOST_net_598) );
in01s01 TIMEBOOST_cell_5917 ( .a(FE_OFN1_n_43918), .o(TIMEBOOST_net_1806) );
in01s01 g772838 ( .a(n_8057), .o(n_8124) );
ao12m06 g772839 ( .a(n_7936), .b(n_8066), .c(n_7984), .o(n_8057) );
ao12s01 g772840 ( .a(n_7977), .b(n_7976), .c(n_7975), .o(n_9172) );
ao12s01 g772841 ( .a(n_8068), .b(n_8067), .c(n_8066), .o(n_9640) );
in01m02 g772843 ( .a(n_8154), .o(n_8155) );
no02s02 g772845 ( .a(n_7821), .b(n_7378), .o(n_7869) );
na02s06 TIMEBOOST_cell_4170 ( .a(n_32279), .b(TIMEBOOST_net_1175), .o(n_32360) );
no02m02 TIMEBOOST_cell_4948 ( .a(n_18096), .b(n_18024), .o(TIMEBOOST_net_1422) );
na02s04 g772848 ( .a(n_7969), .b(n_7331), .o(n_8011) );
no02f06 g772849 ( .a(n_7976), .b(n_7783), .o(n_8041) );
no02s01 g772850 ( .a(n_7976), .b(n_7975), .o(n_7977) );
na02s01 g772852 ( .a(n_7967), .b(FE_OCP_RBN6627_n_7832), .o(n_8008) );
na02m08 TIMEBOOST_cell_4210 ( .a(TIMEBOOST_net_1195), .b(n_12378), .o(n_12450) );
no02s02 g772854 ( .a(n_8001), .b(FE_OCP_RBN6582_n_8021), .o(n_8022) );
no02s06 TIMEBOOST_cell_5128 ( .a(n_34180), .b(n_34206), .o(TIMEBOOST_net_1512) );
no02s01 g772857 ( .a(n_8067), .b(n_8066), .o(n_8068) );
na02s04 g772858 ( .a(n_8051), .b(n_8050), .o(n_8158) );
in01s01 g772859 ( .a(n_8052), .o(n_8053) );
no02s02 g772860 ( .a(n_8017), .b(n_8016), .o(n_8052) );
in01s01 g772861 ( .a(n_8102), .o(n_8103) );
no02s03 g772862 ( .a(n_8051), .b(n_8050), .o(n_8102) );
no02s01 g772863 ( .a(n_8040), .b(n_8084), .o(n_8141) );
na02s03 g772864 ( .a(n_8017), .b(n_8016), .o(n_8122) );
no02s01 g772865 ( .a(n_8064), .b(n_8063), .o(n_8065) );
na02s01 g772866 ( .a(n_8007), .b(n_8054), .o(n_8125) );
in01s01 g772868 ( .a(n_7985), .o(n_8019) );
in01s01 g772870 ( .a(n_8024), .o(n_8025) );
ao12s01 g772871 ( .a(n_7940), .b(n_7939), .c(n_7938), .o(n_8024) );
na02s04 TIMEBOOST_cell_2100 ( .a(TIMEBOOST_net_664), .b(n_20822), .o(n_20935) );
oa12s01 g772874 ( .a(n_8005), .b(n_8004), .c(n_8003), .o(n_9525) );
na02s02 g772875 ( .a(n_8153), .b(n_8143), .o(n_8200) );
in01s01 g772877 ( .a(n_8006), .o(n_8007) );
no02s03 g772878 ( .a(n_7974), .b(n_7973), .o(n_8006) );
in01s01 g772879 ( .a(n_8039), .o(n_8040) );
na02s03 g772880 ( .a(n_7992), .b(n_7991), .o(n_8039) );
no02s04 TIMEBOOST_cell_4015 ( .a(n_8850), .b(FE_OCP_RBN5747_n_8637), .o(TIMEBOOST_net_1098) );
no02m04 g772883 ( .a(n_7992), .b(n_7991), .o(n_8084) );
na02s02 g772884 ( .a(n_7974), .b(n_7973), .o(n_8054) );
na02s01 g772886 ( .a(n_8004), .b(n_8003), .o(n_8005) );
no02s01 g772887 ( .a(n_7939), .b(n_7938), .o(n_7940) );
no02s01 g772888 ( .a(n_7987), .b(n_7932), .o(n_8064) );
na02s01 g772889 ( .a(n_7984), .b(n_7937), .o(n_8067) );
in01s01 g772891 ( .a(n_7798), .o(n_7821) );
ao12m08 g772892 ( .a(n_7338), .b(n_7731), .c(n_7355), .o(n_7798) );
in01s02 g772893 ( .a(n_7969), .o(n_7970) );
in01m01 g772894 ( .a(n_7949), .o(n_7969) );
oa12m08 g772895 ( .a(n_7268), .b(n_45875), .c(n_7291), .o(n_7949) );
ao12f06 g772896 ( .a(n_7698), .b(n_7902), .c(n_7751), .o(n_7976) );
in01s01 g772897 ( .a(n_8001), .o(n_8002) );
in01s02 g772898 ( .a(n_7959), .o(n_8001) );
no02m06 g772899 ( .a(n_7887), .b(n_7722), .o(n_7959) );
in01s01 g772900 ( .a(n_7967), .o(n_7968) );
in01s02 g772901 ( .a(n_7948), .o(n_7967) );
na02s06 g772902 ( .a(n_7843), .b(n_7720), .o(n_7948) );
no02s02 TIMEBOOST_cell_1983 ( .a(n_33020), .b(FE_OCP_RBN2483_FE_RN_657_0), .o(TIMEBOOST_net_606) );
na02s01 TIMEBOOST_cell_3833 ( .a(n_1393), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_), .o(TIMEBOOST_net_1007) );
oa12s02 g772906 ( .a(n_7871), .b(n_7902), .c(n_7870), .o(n_9151) );
oa12s01 g772907 ( .a(n_7935), .b(n_7934), .c(n_7933), .o(n_9605) );
in01s01 g772908 ( .a(n_7978), .o(n_7979) );
oa12s01 g772909 ( .a(n_7898), .b(n_7897), .c(n_7896), .o(n_7978) );
in01s01 g772910 ( .a(n_7966), .o(n_8063) );
oa12m04 g772911 ( .a(n_7912), .b(n_7865), .c(n_7810), .o(n_7966) );
no02s08 TIMEBOOST_cell_2008 ( .a(TIMEBOOST_net_618), .b(n_33871), .o(n_33942) );
na02s02 g772916 ( .a(n_7750), .b(n_7365), .o(n_7804) );
na02s02 g772917 ( .a(n_45875), .b(n_7318), .o(n_7868) );
na03m06 TIMEBOOST_cell_5761 ( .a(TIMEBOOST_net_1244), .b(FE_OCP_RBN4136_n_7743), .c(FE_OCP_RBN6654_n_8187), .o(n_8318) );
na02s01 g772920 ( .a(n_7902), .b(n_7870), .o(n_7871) );
no02s01 g772921 ( .a(n_7953), .b(n_7849), .o(n_8028) );
na02s03 g772923 ( .a(n_7835), .b(FE_OCP_RBN6602_n_7881), .o(n_7852) );
no02s04 TIMEBOOST_cell_6729 ( .a(FE_OCPN5128_n_22280), .b(n_24688), .o(TIMEBOOST_net_2122) );
na03s20 TIMEBOOST_cell_8173 ( .a(n_10167), .b(n_10387), .c(n_11507), .o(n_11571) );
na02s02 g772928 ( .a(FE_OCP_RBN2654_FE_OCPN914_n_8091), .b(n_7730), .o(n_8094) );
no02f06 TIMEBOOST_cell_4921 ( .a(TIMEBOOST_net_1408), .b(n_23176), .o(n_23250) );
in01s01 g772930 ( .a(n_7936), .o(n_7937) );
no02s02 g772931 ( .a(n_7875), .b(n_7874), .o(n_7936) );
na02s02 g772932 ( .a(n_7875), .b(n_7874), .o(n_7984) );
na02s01 g772933 ( .a(n_7897), .b(n_7896), .o(n_7898) );
na02s01 g772934 ( .a(n_7934), .b(n_7933), .o(n_7935) );
na02s04 g772935 ( .a(n_8009), .b(n_7850), .o(n_8010) );
in01s01 g772937 ( .a(n_7931), .o(n_7932) );
na02s04 g772938 ( .a(n_7884), .b(n_7883), .o(n_7931) );
no02s03 g772939 ( .a(n_7884), .b(n_7883), .o(n_7987) );
na02s01 g772940 ( .a(n_7912), .b(n_7866), .o(n_8004) );
na02s01 g772941 ( .a(n_7847), .b(n_7844), .o(n_7939) );
oa12s01 g772943 ( .a(FE_OCP_RBN4139_n_7743), .b(n_8151), .c(n_8150), .o(n_8153) );
in01s02 g772944 ( .a(n_7894), .o(n_7895) );
in01s02 g772945 ( .a(n_7843), .o(n_7894) );
no02s06 g772946 ( .a(n_7799), .b(n_7689), .o(n_7843) );
in01m02 g772948 ( .a(n_7887), .o(n_7929) );
na02m06 g772949 ( .a(n_7834), .b(n_7701), .o(n_7887) );
na02m04 g772950 ( .a(n_7846), .b(n_7825), .o(n_7992) );
na02s01 TIMEBOOST_cell_3344 ( .a(n_26863), .b(n_26862), .o(TIMEBOOST_net_963) );
no02s01 g772955 ( .a(n_8550), .b(n_7995), .o(n_8105) );
no02s01 g772956 ( .a(n_7927), .b(n_7913), .o(n_7928) );
na02s01 g772957 ( .a(n_8046), .b(n_7999), .o(n_8082) );
na02m02 g772958 ( .a(n_7814), .b(n_8568), .o(n_7846) );
na03m02 TIMEBOOST_cell_7297 ( .a(FE_RN_1936_0), .b(FE_RN_1937_0), .c(n_5279), .o(n_47002) );
na02s02 g772960 ( .a(n_7813), .b(n_7509), .o(n_7825) );
na02s06 g772961 ( .a(n_7748), .b(n_7027), .o(n_7847) );
in01s01 g772962 ( .a(n_7865), .o(n_7866) );
no02s04 g772963 ( .a(n_7820), .b(n_7819), .o(n_7865) );
in01s01 g772964 ( .a(n_8009), .o(n_7953) );
no02s02 g772965 ( .a(n_7927), .b(n_7818), .o(n_8009) );
na02s02 g772966 ( .a(n_7747), .b(n_7026), .o(n_7844) );
na02s03 g772967 ( .a(n_7820), .b(n_7819), .o(n_7912) );
no03m10 TIMEBOOST_cell_6581 ( .a(n_21350), .b(FE_OCP_RBN3250_n_21312), .c(FE_OCPN1382_n_45026), .o(n_21537) );
in01s01 g772971 ( .a(n_7749), .o(n_7750) );
in01s01 g772972 ( .a(n_7731), .o(n_7749) );
oa12m08 g772973 ( .a(n_7305), .b(n_7662), .c(n_7262), .o(n_7731) );
oa12f06 g772974 ( .a(n_7681), .b(n_7803), .c(n_7727), .o(n_7902) );
in01s02 g772975 ( .a(n_7835), .o(n_7836) );
in01s02 g772976 ( .a(n_7799), .o(n_7835) );
na02s06 g772977 ( .a(n_7677), .b(n_7756), .o(n_7799) );
in01s02 g772978 ( .a(n_7863), .o(n_7864) );
in01s02 g772979 ( .a(n_7834), .o(n_7863) );
no02m06 g772980 ( .a(n_7766), .b(n_7680), .o(n_7834) );
in01s01 g772981 ( .a(n_7861), .o(n_7862) );
oa12s01 g772982 ( .a(n_7787), .b(n_7803), .c(n_7786), .o(n_7861) );
in01s01 TIMEBOOST_cell_8895 ( .a(TIMEBOOST_net_2938), .o(TIMEBOOST_net_2939) );
oa12s01 g772984 ( .a(n_7797), .b(n_7796), .c(n_7795), .o(n_7934) );
oa12s01 g772985 ( .a(n_7790), .b(n_7789), .c(n_7788), .o(n_7897) );
oa12m04 g772986 ( .a(n_7407), .b(n_7754), .c(n_7388), .o(n_7938) );
oa12m01 g772988 ( .a(n_7773), .b(n_45846), .c(n_45871), .o(n_8091) );
in01s01 g772989 ( .a(n_7810), .o(n_8003) );
na02m08 TIMEBOOST_cell_5194 ( .a(TIMEBOOST_net_646), .b(FE_RN_2248_0), .o(TIMEBOOST_net_1545) );
na02m01 g772994 ( .a(n_45846), .b(n_45871), .o(n_7773) );
na02s01 g772995 ( .a(n_7803), .b(n_7786), .o(n_7787) );
na02s01 g772996 ( .a(n_8172), .b(n_8119), .o(n_8173) );
no02s02 TIMEBOOST_cell_5193 ( .a(TIMEBOOST_net_1544), .b(n_3421), .o(TIMEBOOST_net_1259) );
na02m08 TIMEBOOST_cell_8811 ( .a(TIMEBOOST_net_2892), .b(n_10912), .o(n_11052) );
no02s01 g773001 ( .a(n_7965), .b(n_7964), .o(n_7999) );
na02s02 g773002 ( .a(n_7713), .b(n_7683), .o(n_7777) );
no02s01 g773003 ( .a(n_8027), .b(n_7954), .o(n_7955) );
no02s02 g773004 ( .a(n_7752), .b(n_8444), .o(n_7753) );
no02s01 g773005 ( .a(n_7775), .b(n_7807), .o(n_7831) );
na02s01 g773006 ( .a(n_7796), .b(n_7795), .o(n_7797) );
in01s02 g773007 ( .a(n_8046), .o(n_8550) );
ao12s02 g773008 ( .a(n_8027), .b(n_7924), .c(FE_OCP_RBN2587_n_7743), .o(n_8046) );
na02s01 g773009 ( .a(n_7789), .b(n_7788), .o(n_7790) );
na02s02 g773010 ( .a(n_7860), .b(n_7809), .o(n_7927) );
in01s01 g773011 ( .a(n_8143), .o(n_8144) );
ao12s02 g773012 ( .a(n_8113), .b(n_8032), .c(FE_OCP_RBN4139_n_7743), .o(n_8143) );
in01s02 g773013 ( .a(n_7784), .o(n_7785) );
in01s03 g773014 ( .a(n_7756), .o(n_7784) );
na03f08 TIMEBOOST_cell_5729 ( .a(n_12863), .b(n_12718), .c(n_12860), .o(n_12861) );
ao12s01 g773016 ( .a(FE_OCP_RBN2587_n_7743), .b(n_8110), .c(n_8062), .o(n_8151) );
in01s02 g773017 ( .a(n_7813), .o(n_7814) );
in01s02 g773018 ( .a(n_7766), .o(n_7813) );
na02m06 g773019 ( .a(n_7752), .b(n_7672), .o(n_7766) );
ao12s01 g773020 ( .a(n_7762), .b(n_7761), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_0_), .o(n_9324) );
no02s01 TIMEBOOST_cell_5467 ( .a(TIMEBOOST_net_1681), .b(n_47278), .o(n_22336) );
in01s01 g773022 ( .a(n_7747), .o(n_7748) );
no02s01 g773024 ( .a(n_7761), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_0_), .o(n_7762) );
no02s01 g773025 ( .a(n_8037), .b(n_8081), .o(n_8172) );
in01s01 g773026 ( .a(n_8166), .o(n_8167) );
na02s01 g773027 ( .a(n_8110), .b(n_8047), .o(n_8166) );
na02m02 g773028 ( .a(n_7703), .b(n_7702), .o(n_7704) );
na02s02 TIMEBOOST_cell_4092 ( .a(TIMEBOOST_net_1136), .b(FE_OCP_RBN6834_n_31073), .o(n_31236) );
in01s01 g773031 ( .a(n_7686), .o(n_7687) );
in01s01 g773032 ( .a(n_7662), .o(n_7686) );
ao12m08 g773033 ( .a(n_7235), .b(n_7636), .c(n_7252), .o(n_7662) );
no02f08 g773034 ( .a(n_7679), .b(FE_OCP_RBN2558_n_7665), .o(n_7803) );
na02s02 g773035 ( .a(n_7951), .b(n_7998), .o(n_8061) );
ao12s01 g773037 ( .a(n_8118), .b(n_8362), .c(n_8150), .o(n_8961) );
ao12s01 g773040 ( .a(FE_OCP_RBN5610_n_7730), .b(n_7889), .c(n_7888), .o(n_8027) );
oa12s01 g773041 ( .a(FE_OCPN858_n_7802), .b(n_7849), .c(n_7848), .o(n_7850) );
ao12s01 g773042 ( .a(FE_OCP_RBN4080_n_7708), .b(n_7824), .c(n_7908), .o(n_7965) );
ao12s01 g773043 ( .a(FE_OCP_RBN2587_n_7743), .b(n_8045), .c(n_7982), .o(n_8113) );
ao12s01 g773044 ( .a(n_7730), .b(n_7763), .c(n_7828), .o(n_7818) );
in01s01 g773046 ( .a(n_7713), .o(n_7718) );
na02s06 g773047 ( .a(n_7626), .b(n_7693), .o(n_7713) );
oa12s01 g773048 ( .a(FE_OCPN850_n_7712), .b(n_7807), .c(n_7801), .o(n_7809) );
in01s01 g773049 ( .a(n_7860), .o(n_7775) );
na02s02 g773050 ( .a(n_7717), .b(FE_OCP_RBN6598_n_7708), .o(n_7860) );
in01s01 g773051 ( .a(n_7752), .o(n_7724) );
in01s01 g773053 ( .a(FE_OCP_RBN6583_n_8021), .o(n_8069) );
ao12s01 g773054 ( .a(n_7629), .b(n_7636), .c(n_7628), .o(n_8021) );
no02s01 g773056 ( .a(n_7706), .b(n_7742), .o(n_7832) );
in01s01 g773057 ( .a(n_7754), .o(n_7796) );
na02s02 g773058 ( .a(n_7656), .b(n_7685), .o(n_7754) );
in01s01 g773059 ( .a(n_7745), .o(n_7789) );
na02s03 g773060 ( .a(n_45826), .b(n_7647), .o(n_7745) );
no02s01 g773061 ( .a(n_7636), .b(n_7628), .o(n_7629) );
no02m06 g773062 ( .a(n_7667), .b(n_167), .o(n_7679) );
no02s01 g773063 ( .a(n_7696), .b(n_7227), .o(n_7742) );
no02s01 g773064 ( .a(n_45887), .b(n_7228), .o(n_7706) );
in01s01 g773066 ( .a(n_7951), .o(n_7952) );
no02s01 g773067 ( .a(n_7855), .b(n_7922), .o(n_7951) );
in01s01 g773068 ( .a(n_8014), .o(n_8015) );
no02s01 g773069 ( .a(n_7920), .b(n_7996), .o(n_8014) );
no02s02 g773070 ( .a(n_7839), .b(n_7858), .o(n_7859) );
no02s01 g773071 ( .a(n_7997), .b(n_7918), .o(n_7998) );
no02s01 g773074 ( .a(n_7961), .b(n_8038), .o(n_8048) );
no02s02 g773075 ( .a(n_7909), .b(n_7988), .o(n_7989) );
no02s01 g773077 ( .a(n_8058), .b(n_8012), .o(n_8735) );
no02s01 g773078 ( .a(n_7914), .b(n_7913), .o(n_8430) );
na02s01 g773079 ( .a(n_7716), .b(n_7827), .o(n_8281) );
na02s01 g773080 ( .a(n_7716), .b(n_7715), .o(n_7717) );
in01s01 g773081 ( .a(n_8118), .o(n_8119) );
no02s01 g773082 ( .a(FE_OCP_RBN4139_n_7743), .b(n_8150), .o(n_8118) );
na02s01 g773083 ( .a(n_7768), .b(n_7830), .o(n_8160) );
na02s01 g773084 ( .a(n_7665), .b(n_7668), .o(n_7761) );
in01s01 g773086 ( .a(n_8086), .o(n_8087) );
na02s01 g773087 ( .a(n_7993), .b(n_8045), .o(n_8086) );
in01s01 g773088 ( .a(n_8081), .o(n_8047) );
no02s01 g773089 ( .a(FE_OCP_RBN2595_n_7743), .b(n_7950), .o(n_8081) );
no02s01 g773090 ( .a(n_7962), .b(n_8085), .o(n_8772) );
na02s01 g773092 ( .a(n_7811), .b(n_7921), .o(n_8468) );
na02s01 g773093 ( .a(n_7712), .b(n_7957), .o(n_7720) );
na02s01 g773094 ( .a(n_7641), .b(n_8226), .o(n_7656) );
no02s02 g773095 ( .a(FE_OCP_RBN4075_n_7708), .b(n_8676), .o(n_7722) );
na02s02 g773096 ( .a(n_7646), .b(n_45821), .o(n_7647) );
na02s01 g773097 ( .a(n_7627), .b(n_7611), .o(n_7685) );
na02s01 g773098 ( .a(n_7739), .b(n_7841), .o(n_8371) );
no02s01 g773099 ( .a(n_7996), .b(n_7995), .o(n_8588) );
no02s01 g773100 ( .a(n_7759), .b(n_7711), .o(n_8096) );
no02s01 g773101 ( .a(n_7783), .b(n_7782), .o(n_7975) );
na02s02 g773102 ( .a(FE_OCP_RBN2605_FE_OCPN855_n_7721), .b(n_7950), .o(n_8110) );
na02s01 g773103 ( .a(n_7699), .b(n_7751), .o(n_7870) );
na02s01 g773104 ( .a(n_7880), .b(n_7923), .o(n_7924) );
no02s01 g773105 ( .a(n_7980), .b(n_7964), .o(n_8706) );
na02s01 g773106 ( .a(n_8031), .b(n_8030), .o(n_8032) );
no02s01 g773107 ( .a(n_7997), .b(n_7954), .o(n_8605) );
no02s01 g773108 ( .a(n_7922), .b(n_7829), .o(n_8494) );
no02s01 g773109 ( .a(n_7682), .b(n_7727), .o(n_7786) );
na02s02 g773110 ( .a(n_7741), .b(n_7710), .o(n_7757) );
oa12s01 g773111 ( .a(n_7854), .b(n_8362), .c(n_7888), .o(n_8716) );
ao12s01 g773112 ( .a(n_7806), .b(n_8232), .c(n_7215), .o(n_8556) );
ao12s01 g773113 ( .a(n_7816), .b(FE_OFN4767_n_8309), .c(n_7105), .o(n_8479) );
oa12s01 g773114 ( .a(n_8059), .b(n_8232), .c(n_8030), .o(n_8867) );
oa12s01 g773115 ( .a(n_7960), .b(n_8232), .c(n_7982), .o(n_8820) );
oa12s01 g773116 ( .a(n_8036), .b(n_8232), .c(n_8062), .o(n_8931) );
oa12s01 g773117 ( .a(n_7891), .b(n_8362), .c(n_7828), .o(n_8648) );
oa12s01 g773118 ( .a(n_7919), .b(n_8362), .c(n_7908), .o(n_8721) );
oa12s01 g773119 ( .a(n_7917), .b(n_8362), .c(n_7923), .o(n_8724) );
oa12s01 g773120 ( .a(n_7840), .b(n_8362), .c(n_7296), .o(n_8644) );
oa12s01 g773121 ( .a(n_7910), .b(n_8362), .c(n_7356), .o(n_8638) );
in01s01 g773122 ( .a(n_7693), .o(n_7675) );
na02m06 g773124 ( .a(n_7654), .b(n_45825), .o(n_7703) );
no02m02 g773125 ( .a(n_7646), .b(n_7644), .o(n_7692) );
in01s01 g773126 ( .a(n_7741), .o(n_7782) );
na02s01 g773127 ( .a(n_7708), .b(n_7707), .o(n_7741) );
in01s01 g773128 ( .a(n_7698), .o(n_7699) );
no02s02 g773129 ( .a(n_7674), .b(n_7663), .o(n_7698) );
no02s02 g773130 ( .a(n_7712), .b(n_7707), .o(n_7783) );
no02s01 g773131 ( .a(FE_OCP_RBN2587_n_7743), .b(n_7915), .o(n_8058) );
in01s01 g773132 ( .a(n_7710), .o(n_7711) );
na02s01 g773133 ( .a(n_7617), .b(n_7690), .o(n_7710) );
na02s01 g773134 ( .a(FE_OCP_RBN2612_FE_OCPN857_n_7802), .b(n_8030), .o(n_8059) );
in01s01 g773135 ( .a(n_7857), .o(n_7914) );
na02s01 g773136 ( .a(FE_OCP_RBN5610_n_7730), .b(n_7723), .o(n_7857) );
in01s01 g773137 ( .a(n_8018), .o(n_8085) );
na02s01 g773138 ( .a(FE_OCP_RBN2587_n_7743), .b(n_7945), .o(n_8018) );
na02s02 g773139 ( .a(n_7712), .b(FE_OCPN1204_n_7663), .o(n_7751) );
no02s01 g773140 ( .a(n_7617), .b(n_7881), .o(n_7689) );
in01s01 g773141 ( .a(n_7667), .o(n_7668) );
no02f04 g773142 ( .a(n_7634), .b(FE_OCPN1614_n_7630), .o(n_7667) );
in01s01 g773143 ( .a(n_7768), .o(n_7740) );
na02s01 g773144 ( .a(n_7708), .b(n_7714), .o(n_7768) );
no02s01 g773145 ( .a(FE_OCP_RBN6597_n_7708), .b(n_7794), .o(n_7922) );
na02s01 g773146 ( .a(n_7599), .b(n_7676), .o(n_7677) );
in01s01 g773147 ( .a(n_7716), .o(n_7697) );
na02s01 g773148 ( .a(n_7674), .b(n_7163), .o(n_7716) );
in01s01 g773149 ( .a(n_7909), .o(n_7910) );
no02s01 g773150 ( .a(FE_OCPN858_n_7802), .b(n_7848), .o(n_7909) );
in01s01 g773151 ( .a(n_7824), .o(n_7995) );
na02s01 g773152 ( .a(FE_OCPN849_n_7712), .b(n_7812), .o(n_7824) );
no02s01 g773153 ( .a(FE_OCP_RBN2593_n_7743), .b(n_7877), .o(n_7964) );
in01s01 g773154 ( .a(n_7767), .o(n_7830) );
no02s02 g773155 ( .a(FE_OCPN850_n_7712), .b(n_7714), .o(n_7767) );
no02s01 g773157 ( .a(n_7612), .b(n_8135), .o(n_7646) );
no02s01 g773159 ( .a(FE_OCPN861_n_7743), .b(n_7812), .o(n_7996) );
in01s01 g773160 ( .a(n_7849), .o(n_7811) );
no02s01 g773161 ( .a(n_7730), .b(n_7771), .o(n_7849) );
na02s01 g773162 ( .a(FE_OCP_RBN5609_n_7730), .b(n_7885), .o(n_8045) );
in01s01 g773163 ( .a(n_7889), .o(n_7829) );
na02s01 g773164 ( .a(FE_OCP_RBN2612_FE_OCPN857_n_7802), .b(n_7794), .o(n_7889) );
in01s01 g773165 ( .a(n_7880), .o(n_7954) );
na02s01 g773166 ( .a(FE_OCP_RBN2612_FE_OCPN857_n_7802), .b(n_7853), .o(n_7880) );
in01s01 g773167 ( .a(n_7921), .o(n_7988) );
na02s01 g773168 ( .a(FE_OCP_RBN4075_n_7708), .b(n_7771), .o(n_7921) );
na02s01 g773169 ( .a(n_7730), .b(n_7164), .o(n_7827) );
in01s01 g773170 ( .a(n_7839), .o(n_7840) );
no02s01 g773171 ( .a(FE_OCPN858_n_7802), .b(n_7801), .o(n_7839) );
in01s01 g773172 ( .a(n_7858), .o(n_7841) );
no02s01 g773173 ( .a(FE_OCPN850_n_7712), .b(n_7700), .o(n_7858) );
in01s01 g773174 ( .a(n_7919), .o(n_7920) );
na02s01 g773175 ( .a(FE_OCP_RBN5610_n_7730), .b(n_7908), .o(n_7919) );
in01s01 g773176 ( .a(n_7963), .o(n_8012) );
na02s01 g773177 ( .a(FE_OCP_RBN2612_FE_OCPN857_n_7802), .b(n_7915), .o(n_7963) );
no02m20 TIMEBOOST_cell_8505 ( .a(FE_OCPN3550_n_28381), .b(TIMEBOOST_net_2739), .o(n_28437) );
no02s01 TIMEBOOST_cell_1927 ( .a(n_11915), .b(n_11560), .o(TIMEBOOST_net_578) );
na02f04 g773181 ( .a(n_7615), .b(n_7630), .o(n_7665) );
na02s02 g773182 ( .a(n_7708), .b(n_7925), .o(n_7701) );
no02s01 g773183 ( .a(n_7634), .b(n_8568), .o(n_7680) );
in01s01 g773184 ( .a(n_45825), .o(n_7644) );
in01s01 g773186 ( .a(n_7854), .o(n_7855) );
na02s01 g773187 ( .a(FE_OCP_RBN5610_n_7730), .b(n_7888), .o(n_7854) );
in01s01 g773189 ( .a(n_7627), .o(n_7641) );
no02s06 g773190 ( .a(n_7612), .b(n_8174), .o(n_7627) );
in01s01 g773191 ( .a(n_8036), .o(n_8037) );
na02s01 g773192 ( .a(FE_OCP_RBN4162_FE_OCPN857_n_7802), .b(n_8062), .o(n_8036) );
na02s02 g773193 ( .a(n_7650), .b(n_8444), .o(n_7672) );
in01s01 g773194 ( .a(n_7917), .o(n_7918) );
na02s01 g773195 ( .a(FE_OCP_RBN4075_n_7708), .b(n_7923), .o(n_7917) );
in01s01 g773196 ( .a(n_7739), .o(n_7807) );
na02s01 g773197 ( .a(n_7650), .b(n_7700), .o(n_7739) );
in01s01 g773198 ( .a(n_7805), .o(n_7806) );
na02s01 g773199 ( .a(n_7730), .b(n_7715), .o(n_7805) );
in01s01 g773200 ( .a(n_7916), .o(n_7980) );
na02s01 g773201 ( .a(FE_OCP_RBN5610_n_7730), .b(n_7877), .o(n_7916) );
na02m01 g773202 ( .a(n_7599), .b(n_7726), .o(n_7626) );
in01s01 g773203 ( .a(n_7681), .o(n_7682) );
na02s06 g773204 ( .a(n_7674), .b(n_7673), .o(n_7681) );
in01s01 g773205 ( .a(n_7913), .o(n_7763) );
no02s01 g773206 ( .a(FE_OCP_RBN4075_n_7708), .b(n_7723), .o(n_7913) );
na02s01 g773207 ( .a(FE_OCP_RBN5610_n_7730), .b(n_7828), .o(n_7891) );
in01s01 g773208 ( .a(n_7815), .o(n_7816) );
na02s01 g773209 ( .a(FE_OCP_RBN6598_n_7708), .b(n_7769), .o(n_7815) );
no02s01 g773210 ( .a(FE_OCP_RBN2612_FE_OCPN857_n_7802), .b(n_7853), .o(n_7997) );
in01s02 g773211 ( .a(n_7759), .o(n_7760) );
no02s01 g773212 ( .a(n_7730), .b(n_7690), .o(n_7759) );
in01s01 g773213 ( .a(n_8038), .o(n_7993) );
no02s01 g773214 ( .a(FE_OCP_RBN2593_n_7743), .b(n_7885), .o(n_8038) );
in01s01 g773215 ( .a(n_7962), .o(n_8031) );
no02s01 g773216 ( .a(FE_OCPN861_n_7743), .b(n_7945), .o(n_7962) );
in01s01 g773218 ( .a(n_7960), .o(n_7961) );
na02s01 g773219 ( .a(FE_OCP_RBN2612_FE_OCPN857_n_7802), .b(n_7982), .o(n_7960) );
in01s01 g773220 ( .a(n_45887), .o(n_7696) );
oa12m08 g773222 ( .a(FE_OCP_DRV_N3498_n_7233), .b(n_7542), .c(FE_OCP_DRV_N3500_n_7204), .o(n_7636) );
ao12s01 g773224 ( .a(n_7580), .b(n_7579), .c(n_7578), .o(n_8676) );
oa12s01 g773225 ( .a(n_7625), .b(n_7624), .c(n_7623), .o(n_8150) );
in01s01 g773226 ( .a(n_7957), .o(n_7941) );
oa22s02 g773227 ( .a(n_44828), .b(n_45889), .c(n_44829), .d(n_7193), .o(n_7957) );
oa12s01 g773228 ( .a(n_7604), .b(n_7603), .c(n_7602), .o(n_7950) );
na02s01 g773229 ( .a(n_7557), .b(n_7569), .o(n_7570) );
no02s01 g773230 ( .a(n_7571), .b(n_7572), .o(n_7573) );
na02s01 g773231 ( .a(n_7549), .b(n_7556), .o(n_7592) );
no02s01 g773232 ( .a(n_7737), .b(n_7669), .o(n_7738) );
na02s01 g773233 ( .a(n_7709), .b(n_7691), .o(n_7744) );
in01s01 g773234 ( .a(n_7657), .o(n_7658) );
na02s01 g773235 ( .a(n_7621), .b(n_7633), .o(n_7657) );
in01s01 g773236 ( .a(n_7596), .o(n_7597) );
no02s01 g773237 ( .a(n_7572), .b(n_7547), .o(n_7596) );
na02s02 g773238 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_27_), .b(n_8635), .o(n_8699) );
in01s01 g773239 ( .a(n_7639), .o(n_7640) );
no02s01 g773240 ( .a(n_45616), .b(n_8531), .o(n_7639) );
in01s01 g773241 ( .a(n_7600), .o(n_7601) );
no02s01 g773242 ( .a(n_7577), .b(n_8742), .o(n_7600) );
in01s01 g773243 ( .a(n_7735), .o(n_7736) );
na02s01 g773244 ( .a(n_7670), .b(n_7709), .o(n_7735) );
in01s01 g773245 ( .a(n_7605), .o(n_7606) );
no02s01 g773246 ( .a(n_7582), .b(n_8840), .o(n_7605) );
na02s01 g773247 ( .a(n_7624), .b(n_7623), .o(n_7625) );
na02s01 g773248 ( .a(n_7603), .b(n_7602), .o(n_7604) );
no02s01 g773249 ( .a(n_7579), .b(n_7578), .o(n_7580) );
in01s01 g773250 ( .a(n_7631), .o(n_7632) );
na02s01 g773251 ( .a(n_8635), .b(n_7593), .o(n_7631) );
in01s04 g773252 ( .a(n_7615), .o(n_7674) );
in01f02 g773253 ( .a(n_7599), .o(n_7615) );
in01s10 g773279 ( .a(n_7712), .o(n_7730) );
in01s06 g773280 ( .a(n_7617), .o(n_7712) );
in01s03 g773283 ( .a(n_7617), .o(n_7650) );
in01s04 g773285 ( .a(n_7599), .o(n_7617) );
in01m04 g773286 ( .a(n_7612), .o(n_7599) );
in01s01 g773301 ( .a(FE_OCP_RBN4146_n_7743), .o(n_9012) );
in01s02 g773328 ( .a(n_8232), .o(n_8362) );
in01s03 g773335 ( .a(FE_OFN4771_n_8309), .o(n_8232) );
in01s06 g773340 ( .a(n_8189), .o(n_8309) );
in01s06 g773343 ( .a(FE_OCP_RBN4146_n_7743), .o(n_8189) );
in01s01 g773345 ( .a(FE_OCP_RBN4138_n_7743), .o(n_8104) );
in01m03 g773373 ( .a(n_7634), .o(n_7708) );
in01f06 g773377 ( .a(n_7598), .o(n_7634) );
in01m04 g773378 ( .a(n_7612), .o(n_7598) );
no02f08 g773379 ( .a(n_7528), .b(n_7070), .o(n_7612) );
in01s01 g773380 ( .a(n_7590), .o(n_7591) );
oa12s01 g773381 ( .a(n_7557), .b(FE_OCP_RBN4066_n_7558), .c(delay_add_ln22_unr5_stage3_stallmux_q_27_), .o(n_7590) );
in01s01 g773382 ( .a(n_7574), .o(n_7575) );
ao12s01 g773383 ( .a(n_7555), .b(FE_OCP_RBN4066_n_7558), .c(delay_add_ln22_unr5_stage3_stallmux_q_29_), .o(n_7574) );
in01s01 g773384 ( .a(n_7609), .o(n_7610) );
na02s01 g773385 ( .a(n_7581), .b(n_7567), .o(n_7609) );
ao12s01 g773386 ( .a(n_7566), .b(n_7565), .c(n_7564), .o(n_8030) );
in01s01 g773387 ( .a(n_7732), .o(n_7733) );
no02f04 TIMEBOOST_cell_1827 ( .a(n_14524), .b(n_15849), .o(TIMEBOOST_net_528) );
in01s01 g773389 ( .a(n_7660), .o(n_7661) );
no02s01 g773390 ( .a(n_7585), .b(n_7614), .o(n_7660) );
in01s01 g773391 ( .a(n_7764), .o(n_7765) );
oa12s01 g773392 ( .a(n_7695), .b(n_7608), .c(delay_sub_ln21_0_unr5_stage3_stallmux_q_31_), .o(n_7764) );
ao12s01 g773393 ( .a(n_7552), .b(n_7551), .c(n_7550), .o(n_8062) );
in01s01 g773394 ( .a(n_7588), .o(n_7589) );
oa12s01 g773395 ( .a(n_7535), .b(n_7558), .c(delay_add_ln22_unr5_stage3_stallmux_q_31_), .o(n_7588) );
ao22s01 g773396 ( .a(n_7539), .b(n_6922), .c(n_7538), .d(n_6923), .o(n_7945) );
na02s02 g773398 ( .a(n_7562), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_25_), .o(n_7594) );
no02s02 g773399 ( .a(n_7562), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_25_), .o(n_8531) );
na02s02 g773400 ( .a(n_7584), .b(n_7595), .o(n_7633) );
in01s01 g773401 ( .a(n_7621), .o(n_7622) );
na02s01 g773402 ( .a(n_7608), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_), .o(n_7621) );
in01s01 g773403 ( .a(n_7569), .o(n_7577) );
na02s01 g773404 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_26_), .o(n_7569) );
no02s01 g773405 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_26_), .o(n_8742) );
na02s01 g773406 ( .a(n_7608), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_30_), .o(n_7709) );
na02s01 g773407 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_27_), .o(n_7557) );
in01s01 g773408 ( .a(n_7567), .o(n_7568) );
na02s01 g773409 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_25_), .b(n_7518), .o(n_7567) );
no02s01 g773410 ( .a(n_7584), .b(n_7651), .o(n_7671) );
no02s01 g773411 ( .a(FE_OCP_RBN4065_n_7558), .b(n_6681), .o(n_7572) );
in01s01 g773412 ( .a(n_7669), .o(n_7670) );
no02s01 g773413 ( .a(n_7608), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_30_), .o(n_7669) );
na02s01 g773414 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_31_), .o(n_7535) );
na02s01 g773415 ( .a(n_7608), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_31_), .o(n_7695) );
in01s01 g773416 ( .a(n_7593), .o(n_8634) );
na02s01 g773417 ( .a(n_7544), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_26_), .o(n_7593) );
in01s01 g773418 ( .a(n_7547), .o(n_7548) );
no02s01 g773419 ( .a(FE_OCP_RBN4066_n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_30_), .o(n_7547) );
in01s01 g773420 ( .a(n_8840), .o(n_7549) );
no02s01 g773421 ( .a(FE_OCP_RBN4066_n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_28_), .o(n_8840) );
in01s01 g773422 ( .a(n_7586), .o(n_7587) );
na02s01 g773423 ( .a(n_7559), .b(n_7532), .o(n_7586) );
no02s01 g773424 ( .a(n_7565), .b(n_7564), .o(n_7566) );
in01s01 g773425 ( .a(n_7554), .o(n_7582) );
na02s01 g773426 ( .a(FE_OCP_RBN4066_n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_28_), .o(n_7554) );
no02s01 g773427 ( .a(n_7584), .b(n_6680), .o(n_7585) );
in01s01 g773428 ( .a(n_7555), .o(n_7556) );
no02s01 g773429 ( .a(FE_OCP_RBN4066_n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_29_), .o(n_7555) );
na02s02 g773430 ( .a(n_7584), .b(n_6631), .o(n_8635) );
na02s02 g773431 ( .a(n_46992), .b(n_6509), .o(n_7581) );
in01s01 g773432 ( .a(n_7540), .o(n_7541) );
na02s02 g773433 ( .a(n_7530), .b(n_7512), .o(n_7540) );
no02s02 TIMEBOOST_cell_1819 ( .a(FE_OFN756_n_44464), .b(n_10330), .o(TIMEBOOST_net_524) );
no02s01 g773435 ( .a(n_7608), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_27_), .o(n_7614) );
no02s01 g773436 ( .a(n_7551), .b(n_7550), .o(n_7552) );
no02s01 g773437 ( .a(FE_OCP_RBN4064_n_7558), .b(n_6707), .o(n_7571) );
na02f04 TIMEBOOST_cell_6765 ( .a(n_16279), .b(n_14805), .o(TIMEBOOST_net_2140) );
ao12s01 g773439 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_26_), .c(delay_add_ln22_unr5_stage3_stallmux_q_27_), .o(n_7537) );
in01s01 g773440 ( .a(n_7678), .o(n_7737) );
oa12s01 g773441 ( .a(n_7584), .b(n_7595), .c(n_7651), .o(n_7678) );
in01s01 g773442 ( .a(FE_OCPN1210_n_8846), .o(n_7691) );
no02s01 g773443 ( .a(n_7584), .b(n_6784), .o(n_8846) );
ao12f06 g773444 ( .a(n_6904), .b(n_7516), .c(n_6817), .o(n_7528) );
no02s06 TIMEBOOST_cell_5534 ( .a(TIMEBOOST_net_1162), .b(n_36559), .o(TIMEBOOST_net_1715) );
in01s01 g773447 ( .a(n_7542), .o(n_7579) );
oa12m08 g773448 ( .a(n_7207), .b(n_7534), .c(n_7167), .o(n_7542) );
na02s01 TIMEBOOST_cell_7097 ( .a(FE_OCP_RBN4468_n_44267), .b(FE_OCP_RBN3251_n_21312), .o(TIMEBOOST_net_2307) );
no02s01 g773451 ( .a(n_7583), .b(n_7563), .o(n_7881) );
in01s01 g773452 ( .a(n_7925), .o(n_7900) );
oa12s01 g773453 ( .a(n_7524), .b(n_7534), .c(n_7523), .o(n_7925) );
na04s10 TIMEBOOST_cell_7123 ( .a(n_17410), .b(n_17346), .c(n_17561), .d(n_17345), .o(n_17590) );
na02f04 TIMEBOOST_cell_5199 ( .a(TIMEBOOST_net_1547), .b(n_14360), .o(n_14460) );
na02s01 g773456 ( .a(n_7527), .b(n_6830), .o(n_7565) );
in01s01 g773457 ( .a(n_7531), .o(n_7532) );
no02s02 g773458 ( .a(n_7522), .b(n_7521), .o(n_7531) );
in01s01 g773459 ( .a(n_7545), .o(n_7546) );
na02s01 g773460 ( .a(n_7503), .b(n_7536), .o(n_7545) );
in01s01 g773461 ( .a(n_7513), .o(n_7514) );
na02s02 g773462 ( .a(n_7465), .b(n_7501), .o(n_7513) );
na03m02 TIMEBOOST_cell_7366 ( .a(FE_OCP_RBN2639_n_13667), .b(FE_OCP_RBN4099_n_12880), .c(TIMEBOOST_net_1473), .o(n_13836) );
in01s01 g773464 ( .a(n_7511), .o(n_7512) );
no02s02 g773465 ( .a(n_7500), .b(delay_add_ln22_unr5_stage3_stallmux_q_24_), .o(n_7511) );
na02s01 g773466 ( .a(n_7534), .b(n_7523), .o(n_7524) );
no02s01 g773467 ( .a(n_7560), .b(n_7157), .o(n_7563) );
no02s01 g773468 ( .a(n_7543), .b(n_7158), .o(n_7583) );
no02s01 g773469 ( .a(n_7516), .b(n_7515), .o(n_7551) );
na02s02 g773470 ( .a(n_7522), .b(n_7521), .o(n_7559) );
na02s02 g773471 ( .a(n_7500), .b(delay_add_ln22_unr5_stage3_stallmux_q_24_), .o(n_7530) );
na02s02 g773473 ( .a(n_7491), .b(n_7278), .o(n_7558) );
in01s01 g773479 ( .a(n_7584), .o(n_7608) );
in01s02 g773480 ( .a(n_7544), .o(n_7584) );
no02s02 g773481 ( .a(n_7526), .b(n_7256), .o(n_7544) );
in01s01 g773482 ( .a(n_7538), .o(n_7539) );
oa12s01 g773483 ( .a(n_6944), .b(n_7525), .c(n_6756), .o(n_7538) );
in01s01 g773484 ( .a(n_46992), .o(n_7518) );
no02s01 g773486 ( .a(n_7526), .b(n_7497), .o(n_7562) );
ao22s01 g773487 ( .a(n_7525), .b(n_6963), .c(n_7493), .d(n_6962), .o(n_7982) );
na02s01 g773488 ( .a(n_7493), .b(n_6813), .o(n_7527) );
in01s01 g773489 ( .a(n_7502), .o(n_7503) );
no02s02 g773490 ( .a(n_7496), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_23_), .o(n_7502) );
in01s01 g773492 ( .a(n_7498), .o(n_7499) );
na02s01 g773493 ( .a(n_45213), .b(n_8406), .o(n_7498) );
in01s01 g773494 ( .a(n_7465), .o(n_7466) );
na02s01 g773495 ( .a(n_7445), .b(delay_add_ln22_unr5_stage3_stallmux_q_23_), .o(n_7465) );
na02s02 g773496 ( .a(n_7446), .b(n_6413), .o(n_7501) );
in01s01 g773497 ( .a(n_7490), .o(n_7491) );
no02s02 g773498 ( .a(n_7462), .b(n_7292), .o(n_7490) );
in01s01 g773499 ( .a(n_7519), .o(n_7520) );
na02s01 g773500 ( .a(n_8302), .b(n_7484), .o(n_7519) );
no02s01 g773501 ( .a(n_7489), .b(n_7294), .o(n_7526) );
no02s01 g773502 ( .a(n_7488), .b(n_7295), .o(n_7497) );
na02s02 g773503 ( .a(n_7496), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_23_), .o(n_7536) );
in01s01 g773505 ( .a(n_7560), .o(n_7543) );
in01s01 g773507 ( .a(n_7516), .o(n_7510) );
in01s01 g773509 ( .a(n_7676), .o(n_8453) );
oa12s02 g773510 ( .a(n_7506), .b(n_7507), .c(n_7505), .o(n_7676) );
in01s01 g773511 ( .a(n_8568), .o(n_7509) );
ao12s02 g773512 ( .a(n_7471), .b(n_7470), .c(n_7469), .o(n_8568) );
oa12s01 g773513 ( .a(n_7475), .b(n_7474), .c(n_7473), .o(n_7885) );
oa12s01 g773514 ( .a(n_7478), .b(n_7477), .c(n_7476), .o(n_7522) );
na02s01 g773515 ( .a(n_7436), .b(n_7426), .o(n_7500) );
in01s01 g773517 ( .a(n_8303), .o(n_7484) );
no02s02 g773518 ( .a(n_7468), .b(n_7467), .o(n_8303) );
na02s01 g773519 ( .a(n_7435), .b(n_7289), .o(n_7436) );
in01s01 g773520 ( .a(n_7494), .o(n_7495) );
na02s01 g773521 ( .a(n_7461), .b(n_7492), .o(n_7494) );
na02s02 g773522 ( .a(n_7468), .b(n_7467), .o(n_8302) );
na02s01 g773523 ( .a(n_7422), .b(n_7290), .o(n_7426) );
in01s01 g773524 ( .a(n_8406), .o(n_7464) );
na02s02 g773525 ( .a(n_7440), .b(delay_add_ln22_unr5_stage3_stallmux_q_22_), .o(n_8406) );
no02s01 g773527 ( .a(n_7440), .b(delay_add_ln22_unr5_stage3_stallmux_q_22_), .o(n_8405) );
no02s02 g773529 ( .a(n_7271), .b(n_7435), .o(n_7462) );
na02s01 g773530 ( .a(n_7477), .b(n_7476), .o(n_7478) );
na02s01 g773531 ( .a(n_7507), .b(n_7505), .o(n_7506) );
no02s01 g773532 ( .a(n_7470), .b(n_7469), .o(n_7471) );
in01s01 g773533 ( .a(n_7488), .o(n_7489) );
na02s01 g773534 ( .a(n_7477), .b(n_7276), .o(n_7488) );
in01s01 g773535 ( .a(n_7452), .o(n_7453) );
na02s01 g773536 ( .a(n_7412), .b(n_7444), .o(n_7452) );
in01s01 g773538 ( .a(n_7493), .o(n_7525) );
in01s01 g773539 ( .a(n_7480), .o(n_7493) );
oa12f08 g773540 ( .a(n_6783), .b(n_7434), .c(n_6936), .o(n_7480) );
na02s01 g773541 ( .a(n_7474), .b(n_7473), .o(n_7475) );
ao12s01 g773542 ( .a(n_7483), .b(n_45864), .c(n_7481), .o(n_7877) );
ao12s01 g773543 ( .a(n_7451), .b(n_7450), .c(n_7449), .o(n_7915) );
ao12s01 g773544 ( .a(n_7443), .b(n_7442), .c(n_7441), .o(n_7496) );
in01s01 g773545 ( .a(n_7445), .o(n_7446) );
oa12s01 g773546 ( .a(n_7406), .b(n_7405), .c(n_7404), .o(n_7445) );
no02s01 g773547 ( .a(n_7442), .b(n_7441), .o(n_7443) );
na02s01 g773548 ( .a(n_7405), .b(n_7404), .o(n_7406) );
no02s01 g773549 ( .a(n_45864), .b(n_7481), .o(n_7483) );
in01s01 g773550 ( .a(n_7486), .o(n_7487) );
na02s01 g773551 ( .a(n_7472), .b(n_7448), .o(n_7486) );
no02s02 g773552 ( .a(n_7442), .b(n_7254), .o(n_7477) );
in01s01 g773553 ( .a(n_7430), .o(n_7431) );
na02s01 g773554 ( .a(n_7423), .b(n_7385), .o(n_7430) );
na02s02 g773555 ( .a(n_7439), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_21_), .o(n_7492) );
in01s01 g773556 ( .a(n_7422), .o(n_7435) );
no02s02 g773557 ( .a(n_7405), .b(n_7257), .o(n_7422) );
na02s02 g773558 ( .a(n_7402), .b(n_7401), .o(n_7444) );
in01s01 g773559 ( .a(n_7411), .o(n_7412) );
no02s02 g773560 ( .a(n_7402), .b(n_7401), .o(n_7411) );
in01s01 g773561 ( .a(n_7460), .o(n_7461) );
no02s02 g773562 ( .a(n_7439), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_21_), .o(n_7460) );
no02s01 g773563 ( .a(n_7450), .b(n_7449), .o(n_7451) );
oa12s01 g773567 ( .a(n_7410), .b(n_7409), .c(n_7408), .o(n_7812) );
in01s01 g773568 ( .a(n_7683), .o(n_8389) );
ao12s01 g773569 ( .a(n_7457), .b(n_7456), .c(n_7455), .o(n_7683) );
ao12s01 g773570 ( .a(n_7429), .b(n_45865), .c(n_7428), .o(n_7908) );
in01s01 g773571 ( .a(n_8444), .o(n_7458) );
oa12s01 g773572 ( .a(n_7418), .b(n_7417), .c(n_7416), .o(n_8444) );
oa12s01 g773573 ( .a(n_45861), .b(n_7427), .c(n_6877), .o(n_7474) );
oa12s01 g773574 ( .a(n_7421), .b(n_7420), .c(n_7419), .o(n_7468) );
no03m02 TIMEBOOST_cell_2512 ( .a(n_42420), .b(n_42469), .c(n_42470), .o(FE_RN_686_0) );
in01s01 g773576 ( .a(n_7384), .o(n_7385) );
no02s02 g773577 ( .a(n_7372), .b(delay_add_ln22_unr5_stage3_stallmux_q_20_), .o(n_7384) );
no02s01 g773578 ( .a(n_7456), .b(n_7455), .o(n_7457) );
na02s01 g773579 ( .a(n_7420), .b(n_7419), .o(n_7421) );
no02s01 g773580 ( .a(n_45865), .b(n_7428), .o(n_7429) );
in01s01 g773581 ( .a(n_7437), .o(n_7438) );
na02s01 g773582 ( .a(n_7396), .b(n_7432), .o(n_7437) );
na02s01 g773583 ( .a(n_7409), .b(n_7408), .o(n_7410) );
na02s01 g773585 ( .a(n_7417), .b(n_7416), .o(n_7418) );
na03s08 TIMEBOOST_cell_8198 ( .a(TIMEBOOST_net_700), .b(n_32843), .c(n_32826), .o(n_32966) );
na02s02 g773587 ( .a(n_7420), .b(n_7224), .o(n_7442) );
na02s01 g773588 ( .a(n_7425), .b(n_7424), .o(n_7472) );
na02s02 g773589 ( .a(n_7372), .b(delay_add_ln22_unr5_stage3_stallmux_q_20_), .o(n_7423) );
in01s01 g773590 ( .a(n_7447), .o(n_7448) );
no02s01 g773591 ( .a(n_7425), .b(n_7424), .o(n_7447) );
na02s01 g773592 ( .a(n_7363), .b(n_7251), .o(n_7373) );
in01s01 g773593 ( .a(n_7399), .o(n_7400) );
na02s01 g773594 ( .a(FE_OCP_RBN2494_n_7349), .b(n_7382), .o(n_7399) );
na02s02 g773595 ( .a(n_7363), .b(n_7197), .o(n_7405) );
no02f08 g773596 ( .a(n_45865), .b(n_6943), .o(n_7434) );
na02s01 g773597 ( .a(n_7427), .b(n_45863), .o(n_7450) );
ao12s01 g773598 ( .a(n_7394), .b(n_7393), .c(n_7392), .o(n_7923) );
ao12s01 g773600 ( .a(n_7375), .b(n_7381), .c(n_7374), .o(n_7439) );
ao12s01 g773601 ( .a(n_7329), .b(n_7347), .c(n_7328), .o(n_7402) );
oa22s01 g773602 ( .a(n_7351), .b(n_6921), .c(n_7352), .d(n_6920), .o(n_7853) );
no02s01 g773604 ( .a(n_7347), .b(n_7328), .o(n_7329) );
no02s01 g773605 ( .a(n_7381), .b(n_7374), .o(n_7375) );
na02s01 g773606 ( .a(n_47176), .b(n_6942), .o(n_7427) );
in01s01 g773607 ( .a(n_7414), .o(n_7415) );
na02s01 g773608 ( .a(n_7403), .b(n_7369), .o(n_7414) );
in01s01 g773609 ( .a(n_7361), .o(n_7362) );
na02s02 g773610 ( .a(n_7360), .b(n_7308), .o(n_7361) );
no02s01 g773611 ( .a(n_7377), .b(n_6863), .o(n_7413) );
na02s02 g773612 ( .a(n_7376), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_19_), .o(n_7432) );
na02s02 g773613 ( .a(n_7345), .b(n_7344), .o(n_7382) );
in01s01 g773614 ( .a(n_7395), .o(n_7396) );
no02s02 g773615 ( .a(n_7376), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_19_), .o(n_7395) );
in01s01 g773616 ( .a(n_7363), .o(n_7348) );
no02s02 g773617 ( .a(n_7347), .b(n_7195), .o(n_7363) );
no02s02 g773618 ( .a(n_7381), .b(n_7173), .o(n_7420) );
no02s02 g773620 ( .a(n_7345), .b(n_7344), .o(n_7349) );
no02s01 g773621 ( .a(n_7393), .b(n_7392), .o(n_7394) );
oa12m08 g773624 ( .a(n_7102), .b(n_7380), .c(n_7068), .o(n_7417) );
in01s02 g773625 ( .a(n_7702), .o(n_7728) );
ao22m01 g773626 ( .a(n_7380), .b(n_7109), .c(n_7346), .d(n_7108), .o(FE_RN_2569_0) );
in01s01 g773627 ( .a(n_7726), .o(n_7725) );
oa12s01 g773628 ( .a(n_7387), .b(n_7389), .c(n_7386), .o(n_7726) );
ao12s01 g773629 ( .a(n_6858), .b(n_47180), .c(n_6887), .o(n_7409) );
no02m06 TIMEBOOST_cell_8758 ( .a(n_29400), .b(n_29407), .o(TIMEBOOST_net_2866) );
oa22s01 g773631 ( .a(n_7306), .b(n_7199), .c(n_7277), .d(n_7198), .o(n_7372) );
na02s01 g773632 ( .a(n_7358), .b(n_7178), .o(n_7359) );
na02s01 g773633 ( .a(n_7288), .b(delay_add_ln22_unr5_stage3_stallmux_q_18_), .o(n_7360) );
na02s02 g773634 ( .a(n_7354), .b(n_7353), .o(n_7403) );
na02s01 g773635 ( .a(n_7389), .b(n_7386), .o(n_7387) );
in01s01 g773637 ( .a(n_7330), .o(n_7331) );
na02s06 g773638 ( .a(n_7300), .b(n_7326), .o(n_7330) );
na02s02 g773639 ( .a(n_7358), .b(n_7124), .o(n_7381) );
na02s01 g773640 ( .a(n_47181), .b(n_6895), .o(n_7393) );
in01s01 g773641 ( .a(n_7378), .o(n_7379) );
na02s01 g773642 ( .a(n_7342), .b(n_7371), .o(n_7378) );
na02s02 g773643 ( .a(n_7169), .b(n_7306), .o(n_7347) );
no02s02 TIMEBOOST_cell_4892 ( .a(n_6723), .b(n_6653), .o(TIMEBOOST_net_1394) );
in01s01 g773645 ( .a(n_7307), .o(n_7308) );
no02s02 g773646 ( .a(n_7288), .b(delay_add_ln22_unr5_stage3_stallmux_q_18_), .o(n_7307) );
in01s01 g773647 ( .a(n_7368), .o(n_7369) );
no02s02 g773648 ( .a(n_7354), .b(n_7353), .o(n_7368) );
in01s01 g773649 ( .a(n_47176), .o(n_7377) );
in01s01 g773651 ( .a(n_7351), .o(n_7352) );
oa12s01 g773652 ( .a(n_6864), .b(n_7332), .c(n_6940), .o(n_7351) );
oa12s01 g773653 ( .a(n_7315), .b(n_7314), .c(n_7313), .o(n_7794) );
in01s01 g773654 ( .a(n_7848), .o(n_7356) );
oa12s01 g773655 ( .a(n_7299), .b(n_7298), .c(n_7297), .o(n_7848) );
ao12s01 g773656 ( .a(n_7324), .b(n_7323), .c(n_7322), .o(n_7376) );
ao12s01 g773657 ( .a(n_7317), .b(n_7332), .c(n_7316), .o(n_7888) );
ao12s01 g773658 ( .a(n_7266), .b(n_7267), .c(n_7265), .o(n_7345) );
ao12s01 g773659 ( .a(n_7304), .b(n_7303), .c(n_7302), .o(n_7771) );
ao22s01 g773660 ( .a(n_7282), .b(n_6892), .c(n_7281), .d(n_6893), .o(n_7723) );
no02s01 g773661 ( .a(n_7267), .b(n_7265), .o(n_7266) );
no02s01 g773662 ( .a(n_7323), .b(n_7322), .o(n_7324) );
in01s01 g773663 ( .a(n_7358), .o(n_7343) );
no02s04 g773664 ( .a(n_7323), .b(n_7143), .o(n_7358) );
na02s01 g773665 ( .a(n_7298), .b(n_7297), .o(n_7299) );
in01s01 g773666 ( .a(n_7300), .o(n_7301) );
na02m01 g773667 ( .a(n_7238), .b(delay_add_ln22_unr5_stage3_stallmux_q_17_), .o(n_7300) );
in01s01 g773668 ( .a(n_7341), .o(n_7342) );
no02s02 g773669 ( .a(n_7320), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_17_), .o(n_7341) );
na02s06 g773670 ( .a(n_7237), .b(n_6167), .o(n_7326) );
no02s01 g773671 ( .a(n_7303), .b(n_7302), .o(n_7304) );
in01s01 g773672 ( .a(n_7306), .o(n_7277) );
no02s02 g773673 ( .a(n_7267), .b(n_7141), .o(n_7306) );
na02s02 g773674 ( .a(n_7320), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_17_), .o(n_7371) );
na02s01 g773675 ( .a(n_7314), .b(n_7313), .o(n_7315) );
in01s01 g773676 ( .a(n_7365), .o(n_7366) );
na02s01 g773677 ( .a(n_7355), .b(n_7337), .o(n_7365) );
no02s02 g773679 ( .a(n_7269), .b(n_7291), .o(n_7318) );
no02s01 g773680 ( .a(n_7332), .b(n_7316), .o(n_7317) );
na02s01 g773681 ( .a(n_7933), .b(n_7795), .o(n_7407) );
no02s01 g773682 ( .a(n_7933), .b(n_7795), .o(n_7388) );
in01m06 g773688 ( .a(n_7346), .o(n_7380) );
in01s01 g773690 ( .a(n_7611), .o(n_8226) );
ao12s01 g773691 ( .a(n_7334), .b(n_7335), .c(n_7333), .o(n_7611) );
oa22s01 g773692 ( .a(n_7321), .b(n_6730), .c(n_8135), .d(n_7286), .o(n_9391) );
oa12s01 g773693 ( .a(n_7357), .b(n_8174), .c(n_7364), .o(n_9331) );
oa22s01 g773696 ( .a(n_7226), .b(n_7161), .c(n_7236), .d(n_7162), .o(n_7288) );
oa22s01 g773697 ( .a(n_7287), .b(n_7155), .c(n_7261), .d(n_7154), .o(n_7354) );
no02s02 g773698 ( .a(n_7244), .b(delay_add_ln22_unr5_stage3_stallmux_q_16_), .o(n_7291) );
na02s01 g773700 ( .a(n_7284), .b(n_7283), .o(n_7285) );
in01s01 g773701 ( .a(n_7309), .o(n_7310) );
na02s01 g773702 ( .a(n_7263), .b(n_7305), .o(n_7309) );
in01s01 g773703 ( .a(n_7337), .o(n_7338) );
na02s01 g773704 ( .a(n_7273), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_16_), .o(n_7337) );
na02s02 g773705 ( .a(n_7272), .b(n_6123), .o(n_7355) );
in01s01 g773707 ( .a(n_7268), .o(n_7269) );
na02s02 g773708 ( .a(n_7244), .b(delay_add_ln22_unr5_stage3_stallmux_q_16_), .o(n_7268) );
na02s04 g773710 ( .a(n_7236), .b(n_7122), .o(n_7267) );
no02s01 g773711 ( .a(n_7335), .b(n_7333), .o(n_7334) );
na02s04 g773712 ( .a(n_7287), .b(n_7098), .o(n_7323) );
in01s01 g773713 ( .a(n_7311), .o(n_7896) );
na02s01 g773714 ( .a(n_7321), .b(n_7286), .o(n_7311) );
na02s01 g773715 ( .a(n_7327), .b(n_7364), .o(n_7933) );
ao12s01 g773716 ( .a(n_6733), .b(n_7270), .c(n_6717), .o(n_7298) );
in01s01 g773717 ( .a(n_7281), .o(n_7282) );
oa12s01 g773718 ( .a(n_6667), .b(n_7264), .c(n_6741), .o(n_7281) );
oa12s01 g773719 ( .a(n_6938), .b(n_7270), .c(n_6878), .o(n_7303) );
na02s01 g773720 ( .a(n_8174), .b(n_7364), .o(n_7357) );
in01s01 g773722 ( .a(n_7801), .o(n_7296) );
oa12s01 g773723 ( .a(n_7243), .b(n_7264), .c(n_7242), .o(n_7801) );
in01s02 g773724 ( .a(n_7237), .o(n_7238) );
ao12s02 g773725 ( .a(n_7191), .b(n_7194), .c(n_7190), .o(n_7237) );
ao12s01 g773726 ( .a(n_7247), .b(n_7246), .c(n_7245), .o(n_7320) );
ao12s01 g773727 ( .a(n_6718), .b(n_7280), .c(n_6767), .o(n_7314) );
ao22s01 g773728 ( .a(n_7270), .b(n_6977), .c(n_7280), .d(n_6976), .o(n_7828) );
no02s01 g773729 ( .a(n_7246), .b(n_7245), .o(n_7247) );
no02s02 g773730 ( .a(n_7194), .b(n_7190), .o(n_7191) );
in01s01 g773731 ( .a(n_7227), .o(n_7228) );
na02s01 g773732 ( .a(n_7225), .b(n_45844), .o(n_7227) );
na02s01 g773733 ( .a(n_7264), .b(n_7242), .o(n_7243) );
in01s01 g773735 ( .a(n_7262), .o(n_7263) );
no02s02 g773736 ( .a(n_7240), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_15_), .o(n_7262) );
na02s01 g773739 ( .a(n_7252), .b(n_7234), .o(n_7628) );
in01s01 g773740 ( .a(n_7287), .o(n_7261) );
no02s04 g773741 ( .a(n_7246), .b(n_7099), .o(n_7287) );
na02s02 g773742 ( .a(n_7240), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_15_), .o(n_7305) );
in01s01 g773743 ( .a(n_7236), .o(n_7226) );
no02s04 g773744 ( .a(n_7194), .b(n_7100), .o(n_7236) );
oa12s01 g773748 ( .a(n_7231), .b(n_7230), .c(n_7229), .o(n_7700) );
in01s01 g773749 ( .a(n_7321), .o(n_8135) );
oa12s01 g773750 ( .a(n_7223), .b(n_7222), .c(n_7221), .o(n_7321) );
in01s01 g773751 ( .a(n_8174), .o(n_7327) );
no02s02 g773752 ( .a(n_7279), .b(n_7260), .o(n_8174) );
in01s01 g773753 ( .a(n_7272), .o(n_7273) );
na02s06 TIMEBOOST_cell_8620 ( .a(n_16328), .b(FE_OCPN1733_n_14524), .o(TIMEBOOST_net_2797) );
no03s02 TIMEBOOST_cell_3658 ( .a(FE_OCP_RBN6715_n_3604), .b(n_3663), .c(n_3699), .o(n_3832) );
na02s01 g773756 ( .a(n_7218), .b(n_7041), .o(n_7219) );
in01s01 g773757 ( .a(n_45889), .o(n_7193) );
na02s02 g773759 ( .a(n_7156), .b(delay_add_ln22_unr5_stage3_stallmux_q_14_), .o(n_7225) );
no02s01 g773760 ( .a(n_7258), .b(n_7045), .o(n_7260) );
no02s01 g773761 ( .a(n_7241), .b(n_7046), .o(n_7279) );
in01s01 g773762 ( .a(n_7234), .o(n_7235) );
na02s01 g773763 ( .a(n_7201), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_14_), .o(n_7234) );
na02s02 g773766 ( .a(n_7202), .b(n_5999), .o(n_7252) );
na02f04 TIMEBOOST_cell_7905 ( .a(TIMEBOOST_net_2583), .b(n_20687), .o(n_20853) );
na02s06 g773768 ( .a(n_7159), .b(n_7030), .o(n_7194) );
na02s06 g773769 ( .a(n_7218), .b(n_6999), .o(n_7246) );
na02s01 g773770 ( .a(FE_OCP_DRV_N3499_n_7204), .b(n_7233), .o(n_7578) );
no02f02 TIMEBOOST_cell_7893 ( .a(TIMEBOOST_net_2577), .b(n_4140), .o(n_47007) );
na02s01 g773772 ( .a(n_7222), .b(n_7221), .o(n_7223) );
na02s01 g773775 ( .a(n_7159), .b(n_7078), .o(n_7160) );
ao12s01 g773776 ( .a(n_6753), .b(n_7206), .c(n_6705), .o(n_7264) );
in01s01 g773777 ( .a(n_7270), .o(n_7280) );
na02f08 g773778 ( .a(n_7181), .b(n_6743), .o(n_7270) );
na02s01 g773779 ( .a(n_7230), .b(n_7229), .o(n_7231) );
ao12s01 g773780 ( .a(n_7189), .b(n_7188), .c(n_7187), .o(n_7240) );
ao12s01 g773781 ( .a(n_7120), .b(n_7137), .c(n_7119), .o(n_7212) );
no02s01 g773782 ( .a(n_7137), .b(n_7119), .o(n_7120) );
no02s01 g773783 ( .a(n_7188), .b(n_7187), .o(n_7189) );
na02s01 g773784 ( .a(n_7207), .b(n_7166), .o(n_7523) );
in01s01 g773785 ( .a(n_7157), .o(n_7158) );
na02s01 g773786 ( .a(n_7147), .b(n_7146), .o(n_7157) );
no02s01 g773787 ( .a(n_7206), .b(n_6688), .o(n_7230) );
no02s01 g773792 ( .a(n_7182), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_13_), .o(n_7204) );
in01s01 g773793 ( .a(n_7159), .o(n_7150) );
no02s06 g773794 ( .a(n_7137), .b(n_7033), .o(n_7159) );
na02s01 g773795 ( .a(n_7182), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_13_), .o(n_7233) );
in01s01 g773796 ( .a(n_7218), .o(n_7203) );
no02s06 g773797 ( .a(n_7188), .b(n_7006), .o(n_7218) );
oa12f08 g773798 ( .a(n_6754), .b(n_7180), .c(n_6706), .o(n_7181) );
in01s01 g773799 ( .a(n_7258), .o(n_7241) );
na02s01 TIMEBOOST_cell_4902 ( .a(n_1741), .b(n_1714), .o(TIMEBOOST_net_1399) );
na02f08 TIMEBOOST_cell_6936 ( .a(TIMEBOOST_net_2226), .b(n_19973), .o(TIMEBOOST_net_818) );
in01s01 g773802 ( .a(n_7715), .o(n_7215) );
ao12s01 g773803 ( .a(n_7171), .b(n_7180), .c(n_7170), .o(n_7715) );
oa12s01 g773804 ( .a(n_7210), .b(n_7209), .c(n_7208), .o(n_8114) );
oa12s01 g773805 ( .a(n_7139), .b(n_7144), .c(n_7138), .o(n_8099) );
in01s01 g773806 ( .a(n_7201), .o(n_7202) );
ao22s01 g773807 ( .a(n_7153), .b(n_7025), .c(n_7131), .d(n_7024), .o(n_7201) );
oa22s01 g773808 ( .a(n_7072), .b(n_7034), .c(n_7101), .d(n_7035), .o(n_7156) );
no02s01 g773809 ( .a(n_7180), .b(n_6687), .o(n_7206) );
na02s01 g773810 ( .a(n_7117), .b(n_7116), .o(n_7505) );
na02s02 g773811 ( .a(n_7091), .b(delay_add_ln22_unr5_stage3_stallmux_q_12_), .o(n_7147) );
na02s01 TIMEBOOST_cell_4259 ( .a(n_37493), .b(n_37965), .o(TIMEBOOST_net_1220) );
in01s01 g773813 ( .a(n_7166), .o(n_7167) );
na02s01 g773814 ( .a(n_7129), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_12_), .o(n_7166) );
na02s01 g773815 ( .a(n_7209), .b(n_7208), .o(n_7210) );
na02s01 g773816 ( .a(n_7144), .b(n_7138), .o(n_7139) );
no02s02 TIMEBOOST_cell_6929 ( .a(n_2288), .b(n_2794), .o(TIMEBOOST_net_2223) );
na02s06 g773818 ( .a(n_7101), .b(n_6986), .o(n_7137) );
na02s02 g773819 ( .a(FE_OCP_RBN2464_n_7129), .b(n_5884), .o(n_7207) );
na02s06 g773820 ( .a(n_7153), .b(n_6925), .o(n_7188) );
na02s01 g773821 ( .a(FE_RN_839_0), .b(n_7165), .o(n_7469) );
na02s01 g773822 ( .a(n_7090), .b(n_5777), .o(n_7146) );
no02s01 g773823 ( .a(n_7180), .b(n_7170), .o(n_7171) );
ao12s01 g773824 ( .a(n_7114), .b(n_7118), .c(n_7113), .o(n_7182) );
ao12s02 g773825 ( .a(n_7066), .b(n_7065), .c(n_7064), .o(n_7136) );
no02s01 g773826 ( .a(n_7118), .b(n_7113), .o(n_7114) );
no02s01 g773827 ( .a(n_7065), .b(n_7064), .o(n_7066) );
na02s01 g773828 ( .a(n_7093), .b(n_7092), .o(n_7455) );
in01s01 g773829 ( .a(n_7101), .o(n_7072) );
no02s06 g773830 ( .a(n_7065), .b(n_6964), .o(n_7101) );
na02s01 g773831 ( .a(FE_RN_837_0), .b(n_7134), .o(n_7416) );
no02s01 g773833 ( .a(n_7103), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_11_), .o(n_7132) );
na02s02 g773834 ( .a(n_7053), .b(n_5671), .o(n_7116) );
na02s01 g773835 ( .a(n_7103), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_11_), .o(n_7165) );
in01s01 g773836 ( .a(n_7153), .o(n_7131) );
no02s06 g773837 ( .a(n_7118), .b(n_6951), .o(n_7153) );
na02s01 g773838 ( .a(n_7054), .b(delay_add_ln22_unr5_stage3_stallmux_q_11_), .o(n_7117) );
na02s08 g773839 ( .a(n_7089), .b(n_6993), .o(n_7144) );
no02s02 TIMEBOOST_cell_8133 ( .a(TIMEBOOST_net_2697), .b(n_32501), .o(n_32533) );
ao12f08 g773841 ( .a(n_7087), .b(n_7084), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_8_), .o(n_7180) );
in01s01 g773842 ( .a(n_7163), .o(n_7164) );
oa12s01 g773843 ( .a(n_7112), .b(n_7111), .c(n_7110), .o(n_7163) );
ao12s01 g773844 ( .a(n_7128), .b(n_7127), .c(n_7126), .o(n_8050) );
ao12s01 g773845 ( .a(n_7080), .b(n_7088), .c(n_7079), .o(n_8016) );
in01s01 g773846 ( .a(n_7090), .o(n_7091) );
ao22s01 g773847 ( .a(n_7028), .b(n_6927), .c(n_7015), .d(n_6926), .o(n_7090) );
ao22s01 g773849 ( .a(n_7073), .b(n_6929), .c(n_7067), .d(n_6928), .o(n_7129) );
na02s01 g773850 ( .a(n_7111), .b(n_7110), .o(n_7112) );
na02s01 g773851 ( .a(n_7022), .b(n_5619), .o(n_7092) );
na02s01 g773852 ( .a(n_7049), .b(n_7048), .o(n_7386) );
in01s01 g773853 ( .a(n_7108), .o(n_7109) );
na02s02 g773854 ( .a(n_7069), .b(n_7102), .o(n_7108) );
no02s01 g773855 ( .a(n_7127), .b(n_7126), .o(n_7128) );
na02s06 g773856 ( .a(n_7088), .b(n_6992), .o(n_7089) );
no02s01 g773857 ( .a(n_7088), .b(n_7079), .o(n_7080) );
na02s06 g773858 ( .a(n_7073), .b(n_6869), .o(n_7118) );
na02s06 g773859 ( .a(n_7028), .b(n_6871), .o(n_7065) );
na02s04 TIMEBOOST_cell_8732 ( .a(n_13726), .b(FE_OCP_RBN2540_n_12880), .o(TIMEBOOST_net_2853) );
na02s01 g773861 ( .a(n_7071), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_10_), .o(n_7134) );
na02s01 g773862 ( .a(n_7023), .b(delay_add_ln22_unr5_stage3_stallmux_q_10_), .o(n_7093) );
no02s01 g773864 ( .a(n_7071), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_10_), .o(n_7095) );
in01s01 g773865 ( .a(n_7053), .o(n_7054) );
ao12s02 g773866 ( .a(n_6989), .b(n_6997), .c(n_6988), .o(n_7053) );
ao12s01 g773867 ( .a(n_7043), .b(n_7052), .c(n_7042), .o(n_7103) );
no02s02 g773868 ( .a(n_6997), .b(n_6988), .o(n_6989) );
no02s01 g773869 ( .a(n_7052), .b(n_7042), .o(n_7043) );
na02s02 g773870 ( .a(n_6953), .b(delay_add_ln22_unr5_stage3_stallmux_q_9_), .o(n_7049) );
na02s02 g773871 ( .a(n_7044), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_9_), .o(n_7102) );
no02f06 g773872 ( .a(n_7083), .b(n_6521), .o(n_7087) );
in01s01 g773873 ( .a(n_7073), .o(n_7067) );
no02s06 g773874 ( .a(n_7052), .b(n_6880), .o(n_7073) );
na02s01 g773875 ( .a(n_7107), .b(n_7106), .o(n_7283) );
in01s01 g773876 ( .a(n_7028), .o(n_7015) );
no02s06 g773877 ( .a(n_6997), .b(n_6873), .o(n_7028) );
in01s01 g773878 ( .a(n_7068), .o(n_7069) );
no02s02 g773879 ( .a(n_7044), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_9_), .o(n_7068) );
na02s01 g773880 ( .a(n_6952), .b(n_5511), .o(n_7048) );
na02s01 g773881 ( .a(n_7086), .b(n_7085), .o(n_7333) );
na02m08 g773882 ( .a(n_7083), .b(n_6695), .o(n_7084) );
ao12s01 g773883 ( .a(n_6683), .b(n_7094), .c(n_6626), .o(n_7111) );
na02f02 TIMEBOOST_cell_5198 ( .a(n_14269), .b(n_14266), .o(TIMEBOOST_net_1547) );
oa12s06 g773885 ( .a(n_6987), .b(n_7055), .c(n_6930), .o(n_7088) );
oa22s01 g773886 ( .a(n_7008), .b(n_7004), .c(n_7009), .d(n_7055), .o(n_7973) );
in01s01 g773887 ( .a(n_7769), .o(n_7105) );
ao12s01 g773888 ( .a(n_7057), .b(n_7094), .c(n_7056), .o(n_7769) );
oa12s01 g773889 ( .a(n_7059), .b(n_7058), .c(n_7060), .o(n_7991) );
in01s01 g773890 ( .a(n_7022), .o(n_7023) );
ao22s01 g773891 ( .a(n_6916), .b(n_6852), .c(n_6941), .d(n_6853), .o(n_7022) );
ao22s01 g773892 ( .a(n_7007), .b(n_6856), .c(n_6996), .d(n_6855), .o(n_7071) );
na02s02 g773894 ( .a(n_7020), .b(n_5430), .o(n_7085) );
na02s06 g773895 ( .a(n_6941), .b(n_6748), .o(n_6997) );
na02s01 g773896 ( .a(n_7058), .b(n_7060), .o(n_7059) );
in01s01 g773897 ( .a(n_7045), .o(n_7046) );
na02s01 g773898 ( .a(n_7037), .b(n_7036), .o(n_7045) );
na02s01 g773900 ( .a(n_7082), .b(n_7081), .o(n_7221) );
na02s08 g773901 ( .a(n_7007), .b(n_6771), .o(n_7052) );
no02m02 TIMEBOOST_cell_8632 ( .a(n_4127), .b(FE_OCP_RBN4291_n_3909), .o(TIMEBOOST_net_2803) );
na02s06 g773903 ( .a(n_7051), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_8_), .o(n_7106) );
na02s06 g773904 ( .a(n_7021), .b(delay_add_ln22_unr5_stage3_stallmux_q_8_), .o(n_7086) );
no02s01 g773905 ( .a(n_7094), .b(n_7056), .o(n_7057) );
in01s01 g773906 ( .a(n_6952), .o(n_6953) );
ao12s01 g773907 ( .a(n_6884), .b(n_6883), .c(n_6882), .o(n_6952) );
oa12s01 g773908 ( .a(n_7014), .b(n_7013), .c(n_7012), .o(n_7714) );
ao12s01 g773909 ( .a(n_6981), .b(n_6980), .c(n_6979), .o(n_7044) );
no02s01 g773910 ( .a(n_6883), .b(n_6882), .o(n_6884) );
no02s01 g773911 ( .a(n_6980), .b(n_6979), .o(n_6981) );
na02s02 g773912 ( .a(n_7002), .b(n_5393), .o(n_7082) );
na02s06 g773913 ( .a(n_7003), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_7_), .o(n_7081) );
na02s01 g773914 ( .a(n_7063), .b(n_7062), .o(n_7138) );
na02s01 g773915 ( .a(n_6934), .b(n_5362), .o(n_7036) );
na02s02 g773916 ( .a(n_6935), .b(delay_add_ln22_unr5_stage3_stallmux_q_7_), .o(n_7037) );
na02s01 g773917 ( .a(n_7017), .b(n_7016), .o(n_7208) );
in01s01 g773918 ( .a(n_6941), .o(n_6916) );
no02s06 g773919 ( .a(n_6883), .b(n_6758), .o(n_6941) );
in01s01 g773920 ( .a(n_7007), .o(n_6996) );
no02m08 g773921 ( .a(n_6772), .b(n_6980), .o(n_7007) );
in01s01 g773922 ( .a(n_7031), .o(n_7094) );
na02s01 g773924 ( .a(n_7013), .b(n_7012), .o(n_7014) );
in01s01 g773925 ( .a(n_7294), .o(n_7295) );
oa12s01 g773926 ( .a(n_7255), .b(n_7217), .c(delay_xor_ln21_unr6_stage3_stallmux_q_25_), .o(n_7294) );
oa12s01 g773928 ( .a(n_7278), .b(n_7217), .c(delay_xor_ln22_unr6_stage3_stallmux_q_25_), .o(n_7292) );
in01s01 g773930 ( .a(n_7055), .o(n_7004) );
ao12s06 g773931 ( .a(n_6843), .b(n_6984), .c(n_6891), .o(n_7055) );
ao12s01 g773932 ( .a(n_6971), .b(n_6970), .c(n_6984), .o(n_7874) );
ao12s01 g773933 ( .a(n_6995), .b(n_6994), .c(n_7000), .o(n_7883) );
in01s01 g773934 ( .a(n_7020), .o(n_7021) );
ao22s02 g773935 ( .a(n_6908), .b(n_6731), .c(n_6909), .d(n_6732), .o(n_7020) );
in01s01 g773936 ( .a(n_7050), .o(n_7051) );
na02s01 g773938 ( .a(n_6993), .b(n_6992), .o(n_7079) );
no02s01 g773939 ( .a(n_6994), .b(n_7000), .o(n_6995) );
na02s01 g773940 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_25_), .b(n_7217), .o(n_7278) );
in01s01 g773941 ( .a(n_7255), .o(n_7256) );
na02s01 g773942 ( .a(n_7217), .b(delay_xor_ln21_unr6_stage3_stallmux_q_25_), .o(n_7255) );
na02s01 TIMEBOOST_cell_1582 ( .a(TIMEBOOST_net_405), .b(n_25409), .o(n_25580) );
no02s01 g773944 ( .a(n_6959), .b(n_6621), .o(n_7013) );
na02s06 g773945 ( .a(n_6915), .b(delay_add_ln22_unr5_stage3_stallmux_q_6_), .o(n_7017) );
na02s01 g773947 ( .a(n_7011), .b(n_7010), .o(n_7126) );
na02s02 g773950 ( .a(n_6991), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_6_), .o(n_7062) );
no02s01 g773951 ( .a(n_6970), .b(n_6984), .o(n_6971) );
na02s01 g773952 ( .a(n_6914), .b(n_5312), .o(n_7016) );
ao12s01 g773953 ( .a(n_7254), .b(n_7217), .c(delay_xor_ln21_unr6_stage3_stallmux_q_23_), .o(n_7441) );
in01s01 g773954 ( .a(n_7289), .o(n_7290) );
ao12s01 g773955 ( .a(n_7271), .b(n_7217), .c(delay_xor_ln22_unr6_stage3_stallmux_q_24_), .o(n_7289) );
na02s01 g773956 ( .a(n_7239), .b(n_7276), .o(n_7476) );
ao12s01 g773958 ( .a(n_7257), .b(n_7217), .c(delay_xor_ln22_unr6_stage3_stallmux_q_23_), .o(n_7404) );
oa12s01 g773959 ( .a(n_6901), .b(n_6900), .c(n_6899), .o(n_7690) );
in01s01 g773960 ( .a(n_7002), .o(n_7003) );
in01s01 g773962 ( .a(n_6934), .o(n_6935) );
ao22s02 g773963 ( .a(n_6822), .b(n_6660), .c(n_6881), .d(n_6661), .o(n_6934) );
no03m08 TIMEBOOST_cell_8207 ( .a(n_17890), .b(FE_RN_2345_0), .c(FE_RN_2344_0), .o(n_17996) );
no02f08 g773967 ( .a(n_6900), .b(n_6620), .o(n_6959) );
in01s02 g773968 ( .a(n_6960), .o(n_6961) );
no02s06 g773969 ( .a(n_6651), .b(n_6937), .o(n_6960) );
in01s01 g773970 ( .a(n_7008), .o(n_7009) );
na02s01 g773971 ( .a(n_6931), .b(n_6987), .o(n_7008) );
na02s01 g773972 ( .a(n_6969), .b(n_6968), .o(n_7058) );
no02s01 g773973 ( .a(n_7217), .b(delay_xor_ln22_unr6_stage3_stallmux_q_24_), .o(n_7271) );
na02s02 g773974 ( .a(n_6918), .b(n_5139), .o(n_7010) );
na02s01 g773975 ( .a(n_7217), .b(delay_xor_ln21_unr6_stage3_stallmux_q_24_), .o(n_7239) );
na02m01 g773976 ( .a(n_6875), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_5_), .o(n_6993) );
no02s01 g773977 ( .a(n_7217), .b(delay_xor_ln22_unr6_stage3_stallmux_q_23_), .o(n_7257) );
in01s01 g773978 ( .a(n_6908), .o(n_6909) );
na02m01 g773979 ( .a(n_6881), .b(n_6831), .o(n_6908) );
no02s01 g773980 ( .a(n_7172), .b(delay_xor_ln21_unr6_stage3_stallmux_q_23_), .o(n_7254) );
na02s01 g773981 ( .a(FE_OCP_RBN3997_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n_6809), .o(n_7276) );
na02s06 g773982 ( .a(n_6919), .b(delay_add_ln22_unr5_stage3_stallmux_q_5_), .o(n_7011) );
na02s01 g773984 ( .a(n_6900), .b(n_6899), .o(n_6901) );
oa12m06 g773985 ( .a(n_6847), .b(n_6973), .c(n_6910), .o(n_7000) );
oa12s06 g773986 ( .a(n_6824), .b(n_6885), .c(n_6945), .o(n_6984) );
oa12s01 g773987 ( .a(n_6975), .b(n_6974), .c(n_6973), .o(n_7819) );
in01s01 g773988 ( .a(n_7026), .o(n_7027) );
ao12s01 g773989 ( .a(n_6947), .b(n_6946), .c(n_6945), .o(n_7026) );
oa12s01 g773990 ( .a(n_6898), .b(n_6897), .c(n_6896), .o(n_7795) );
ao12s01 g773991 ( .a(n_6950), .b(n_6949), .c(n_6948), .o(n_7788) );
in01s01 g773992 ( .a(n_6914), .o(n_6915) );
no02m04 TIMEBOOST_cell_2965 ( .a(TIMEBOOST_net_773), .b(n_18871), .o(n_18901) );
in01s01 g773994 ( .a(n_6990), .o(n_6991) );
na03f08 TIMEBOOST_cell_8343 ( .a(n_38964), .b(FE_OCP_RBN5895_n_38806), .c(n_38921), .o(n_39059) );
in01s01 g773997 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_24_), .o(n_6809) );
na02s02 TIMEBOOST_cell_8702 ( .a(FE_OCP_RBN5530_n_1541), .b(n_1446), .o(TIMEBOOST_net_2838) );
na02f02 TIMEBOOST_cell_5158 ( .a(n_14475), .b(FE_OCP_RBN5046_n_14450), .o(TIMEBOOST_net_1527) );
na02s01 g774003 ( .a(n_6891), .b(n_6842), .o(n_6970) );
na02s03 g774004 ( .a(n_6907), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_4_), .o(n_6987) );
in01s01 g774005 ( .a(n_6930), .o(n_6931) );
no02s06 g774006 ( .a(n_6907), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_4_), .o(n_6930) );
na02s03 g774007 ( .a(n_6860), .b(n_4948), .o(n_6968) );
in01s02 g774008 ( .a(n_6822), .o(n_6881) );
na02s06 g774009 ( .a(n_6802), .b(n_6801), .o(n_6822) );
na02s01 g774010 ( .a(n_6897), .b(n_6896), .o(n_6898) );
na02s04 g774011 ( .a(n_6861), .b(delay_add_ln22_unr5_stage3_stallmux_q_4_), .o(n_6969) );
na02s06 g774012 ( .a(n_6889), .b(n_6597), .o(n_6890) );
na02m03 g774013 ( .a(n_6889), .b(n_6876), .o(n_6937) );
na02s01 g774014 ( .a(n_6903), .b(n_47210), .o(n_6994) );
no02m04 TIMEBOOST_cell_4338 ( .a(TIMEBOOST_net_1259), .b(FE_OCP_RBN5786_n_3421), .o(n_3545) );
no02s01 g774016 ( .a(n_6949), .b(n_6948), .o(n_6950) );
na02s01 g774017 ( .a(n_7224), .b(n_7179), .o(n_7419) );
no02s01 g774018 ( .a(n_6946), .b(n_6945), .o(n_6947) );
na02s01 g774019 ( .a(n_6974), .b(n_6973), .o(n_6975) );
in01s01 g774020 ( .a(n_7250), .o(n_7251) );
ao12s01 g774021 ( .a(n_7196), .b(n_7217), .c(delay_xor_ln22_unr6_stage3_stallmux_q_22_), .o(n_7250) );
oa12s01 g774023 ( .a(n_6958), .b(n_6957), .c(n_6956), .o(n_7707) );
in01s01 g774026 ( .a(n_6918), .o(n_6919) );
no02f08 TIMEBOOST_cell_4384 ( .a(TIMEBOOST_net_1282), .b(n_20150), .o(n_20207) );
in01s01 g774028 ( .a(n_6874), .o(n_6875) );
na02m06 TIMEBOOST_cell_3938 ( .a(TIMEBOOST_net_1059), .b(n_24499), .o(n_24638) );
no02m06 TIMEBOOST_cell_1637 ( .a(n_47256), .b(FE_OCP_RBN4200_n_13796), .o(TIMEBOOST_net_433) );
no02s01 g774034 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_28_), .b(delay_add_ln22_unr5_stage3_stallmux_q_29_), .o(n_6707) );
no02s01 g774035 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_), .o(n_6784) );
no02s01 g774036 ( .a(n_6848), .b(n_6910), .o(n_6974) );
na02s02 g774038 ( .a(n_6780), .b(delay_add_ln22_unr5_stage3_stallmux_q_3_), .o(n_6903) );
in01s01 g774039 ( .a(n_6802), .o(n_6752) );
no02m02 TIMEBOOST_cell_1565 ( .a(n_14479), .b(n_14416), .o(TIMEBOOST_net_397) );
na02s01 g774041 ( .a(n_7172), .b(delay_xor_ln21_unr6_stage3_stallmux_q_22_), .o(n_7179) );
in01s02 g774042 ( .a(n_6842), .o(n_6843) );
na02s03 g774043 ( .a(n_6804), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_3_), .o(n_6842) );
no02s01 g774044 ( .a(n_6885), .b(n_6825), .o(n_6946) );
in01s01 g774046 ( .a(n_7196), .o(n_7197) );
no02s01 g774047 ( .a(n_7172), .b(delay_xor_ln22_unr6_stage3_stallmux_q_22_), .o(n_7196) );
in01s02 g774048 ( .a(n_6889), .o(n_6845) );
no02s20 g774049 ( .a(n_6531), .b(FE_OCP_RBN5527_n_6760), .o(n_6889) );
na02s01 g774050 ( .a(FE_OCP_RBN3997_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n_6746), .o(n_7224) );
na02s01 g774051 ( .a(n_6957), .b(n_6956), .o(n_6958) );
ao12s01 g774052 ( .a(n_7195), .b(n_7172), .c(delay_xor_ln22_unr6_stage3_stallmux_q_21_), .o(n_7328) );
ao12s01 g774053 ( .a(n_7173), .b(n_7172), .c(delay_xor_ln21_unr6_stage3_stallmux_q_21_), .o(n_7374) );
ao12s01 g774059 ( .a(n_6803), .b(n_6835), .c(delay_sub_ln21_0_unr5_stage3_stallmux_q_1_), .o(n_6897) );
ao12s01 g774060 ( .a(n_6834), .b(n_6833), .c(delay_add_ln22_unr5_stage3_stallmux_q_1_), .o(n_6949) );
no02s02 TIMEBOOST_cell_8607 ( .a(TIMEBOOST_net_2790), .b(n_39209), .o(TIMEBOOST_net_1596) );
in01s01 g774063 ( .a(n_6860), .o(n_6861) );
ao12s02 g774064 ( .a(n_6711), .b(n_6729), .c(n_6710), .o(n_6860) );
in01s01 g774066 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_30_), .o(n_6681) );
in01s01 g774068 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_22_), .o(n_6746) );
in01s01 g774072 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_), .o(n_7651) );
na02m08 g774074 ( .a(n_6762), .b(n_6761), .o(n_6763) );
no02s02 g774076 ( .a(n_6724), .b(n_6652), .o(n_6790) );
na02s03 TIMEBOOST_cell_6667 ( .a(FE_OCP_RBN5733_n_19806), .b(n_18230), .o(TIMEBOOST_net_2091) );
in01s01 g774078 ( .a(n_6775), .o(n_6776) );
no02f02 TIMEBOOST_cell_1566 ( .a(TIMEBOOST_net_397), .b(FE_OCP_RBN5045_n_14450), .o(n_14560) );
no02s01 g774082 ( .a(n_7172), .b(delay_xor_ln21_unr6_stage3_stallmux_q_21_), .o(n_7173) );
no02s01 g774083 ( .a(n_6833), .b(delay_add_ln22_unr5_stage3_stallmux_q_1_), .o(n_6834) );
no02s01 g774084 ( .a(n_6835), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_1_), .o(n_6803) );
in01s01 g774085 ( .a(n_6847), .o(n_6848) );
na02s02 g774086 ( .a(n_6832), .b(delay_add_ln22_unr5_stage3_stallmux_q_2_), .o(n_6847) );
no02s02 g774087 ( .a(n_6832), .b(delay_add_ln22_unr5_stage3_stallmux_q_2_), .o(n_6910) );
in01s01 g774088 ( .a(n_6824), .o(n_6825) );
na02s03 g774089 ( .a(n_6798), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_2_), .o(n_6824) );
no02s01 g774090 ( .a(n_7172), .b(delay_xor_ln22_unr6_stage3_stallmux_q_21_), .o(n_7195) );
no02s03 g774091 ( .a(n_6798), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_2_), .o(n_6885) );
na02f08 g774092 ( .a(n_6762), .b(n_6564), .o(n_6957) );
ao12s01 g774097 ( .a(n_6967), .b(n_6966), .c(n_6965), .o(n_7663) );
in01f02 g774101 ( .a(n_6774), .o(n_6725) );
na02m01 g774109 ( .a(FE_OCP_RBN6528_n_6745), .b(n_6547), .o(n_6729) );
in01s02 g774111 ( .a(n_6723), .o(n_6724) );
no02s03 g774112 ( .a(n_6708), .b(n_6734), .o(n_6723) );
no02s01 g774114 ( .a(n_6966), .b(n_6965), .o(n_6967) );
na02s02 g774115 ( .a(n_6867), .b(n_6782), .o(n_6936) );
na02s02 g774116 ( .a(n_6859), .b(n_6829), .o(n_6904) );
in01s01 g774118 ( .a(n_7177), .o(n_7178) );
ao12s01 g774119 ( .a(n_7123), .b(n_6872), .c(delay_xor_ln21_unr6_stage3_stallmux_q_20_), .o(n_7177) );
in01s01 g774120 ( .a(n_7198), .o(n_7199) );
ao12s01 g774121 ( .a(n_7168), .b(n_7172), .c(delay_xor_ln22_unr6_stage3_stallmux_q_20_), .o(n_7198) );
ao12s01 g774122 ( .a(n_7143), .b(n_6872), .c(delay_xor_ln21_unr6_stage3_stallmux_q_19_), .o(n_7322) );
in01s02 g774123 ( .a(n_6719), .o(n_6701) );
oa12s01 g774125 ( .a(n_6675), .b(n_6674), .c(delay_sub_ln21_0_unr5_stage3_stallmux_q_0_), .o(n_7364) );
in01s02 g774126 ( .a(n_6627), .o(n_6589) );
in01s01 g774129 ( .a(n_7286), .o(n_6730) );
oa12s01 g774130 ( .a(n_6655), .b(n_6654), .c(delay_add_ln22_unr5_stage3_stallmux_q_0_), .o(n_7286) );
in01s01 g774132 ( .a(n_6759), .o(n_6833) );
in01s02 g774134 ( .a(n_6739), .o(n_6700) );
in01s02 g774137 ( .a(n_6648), .o(n_6618) );
oa22m04 g774138 ( .a(n_6502), .b(n_6471), .c(n_6488), .d(FE_OCP_RBN3443_n_6471), .o(n_6648) );
in01s01 g774142 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_), .o(n_7595) );
in01s01 g774144 ( .a(n_6866), .o(n_6867) );
na02s01 g774145 ( .a(n_6818), .b(n_6844), .o(n_6866) );
no02s06 g774146 ( .a(n_6590), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_0_), .o(n_6896) );
na02s01 g774147 ( .a(n_6654), .b(delay_add_ln22_unr5_stage3_stallmux_q_0_), .o(n_6655) );
in01s01 g774150 ( .a(n_7168), .o(n_7169) );
no02s01 g774151 ( .a(n_6872), .b(delay_xor_ln22_unr6_stage3_stallmux_q_20_), .o(n_7168) );
in01s01 g774152 ( .a(n_7123), .o(n_7124) );
no02s01 g774153 ( .a(n_6872), .b(delay_xor_ln21_unr6_stage3_stallmux_q_20_), .o(n_7123) );
in01s02 g774154 ( .a(n_6734), .o(n_6679) );
ao12s03 g774157 ( .a(n_6753), .b(n_6676), .c(n_6668), .o(n_6754) );
na02s01 g774158 ( .a(n_6674), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_0_), .o(n_6675) );
no02s01 g774160 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_19_), .o(n_7143) );
in01s02 g774161 ( .a(n_6669), .o(n_6948) );
in01s01 g774163 ( .a(n_7515), .o(n_6859) );
na02s01 g774164 ( .a(n_6769), .b(n_6830), .o(n_7515) );
oa12f10 g774165 ( .a(n_6561), .b(n_6671), .c(n_6593), .o(n_6966) );
no02s04 g774167 ( .a(n_6565), .b(n_6415), .o(n_6576) );
ao12s01 g774168 ( .a(n_7099), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_17_), .o(n_7245) );
ao12s01 g774169 ( .a(n_7141), .b(n_6872), .c(delay_xor_ln22_unr6_stage3_stallmux_q_19_), .o(n_7265) );
na02f02 g774170 ( .a(n_6535), .b(n_6412), .o(n_6558) );
no02f04 g774171 ( .a(FE_OCP_RBN6244_n_6535), .b(n_6396), .o(n_6574) );
oa12s01 g774174 ( .a(n_6673), .b(n_6672), .c(n_6671), .o(n_7673) );
in01s01 g774179 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_27_), .o(n_6680) );
in01s01 g774181 ( .a(n_6639), .o(n_6640) );
na02s01 g774182 ( .a(n_6546), .b(n_6607), .o(n_6639) );
na02s06 g774184 ( .a(n_6656), .b(n_6619), .o(n_6635) );
na02s01 g774185 ( .a(n_6942), .b(n_6939), .o(n_6943) );
na02s01 g774186 ( .a(n_6672), .b(n_6671), .o(n_6673) );
no02s01 g774187 ( .a(n_6872), .b(delay_xor_ln22_unr6_stage3_stallmux_q_19_), .o(n_7141) );
no02s02 g774188 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_17_), .b(n_6806), .o(n_7099) );
in01s02 g774190 ( .a(n_6612), .o(n_6613) );
in01s01 g774192 ( .a(n_6616), .o(n_6617) );
ao12s01 g774194 ( .a(n_6772), .b(FE_OCP_RBN6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln21_unr6_stage3_stallmux_q_9_), .o(n_6979) );
in01s01 g774195 ( .a(n_7154), .o(n_7155) );
ao12s01 g774196 ( .a(n_7097), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_18_), .o(n_7154) );
in01s01 g774197 ( .a(n_7040), .o(n_7041) );
ao12s01 g774198 ( .a(n_6998), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_16_), .o(n_7040) );
ao12m01 g774199 ( .a(n_6873), .b(n_6872), .c(delay_xor_ln22_unr6_stage3_stallmux_q_11_), .o(n_6988) );
ao12s01 g774200 ( .a(n_7033), .b(n_6806), .c(delay_xor_ln22_unr6_stage3_stallmux_q_15_), .o(n_7119) );
in01s01 g774201 ( .a(n_7161), .o(n_7162) );
ao12s01 g774202 ( .a(n_7121), .b(n_6872), .c(delay_xor_ln22_unr6_stage3_stallmux_q_18_), .o(n_7161) );
ao12s01 g774203 ( .a(n_6964), .b(n_6806), .c(delay_xor_ln22_unr6_stage3_stallmux_q_13_), .o(n_7064) );
ao12s02 g774204 ( .a(n_6880), .b(n_6872), .c(delay_xor_ln21_unr6_stage3_stallmux_q_11_), .o(n_7042) );
in01s01 g774205 ( .a(n_6928), .o(n_6929) );
ao12s01 g774206 ( .a(n_6868), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_12_), .o(n_6928) );
ao12s01 g774207 ( .a(n_6951), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_13_), .o(n_7113) );
in01s02 g774208 ( .a(n_6598), .o(n_6599) );
in01s01 g774210 ( .a(n_7024), .o(n_7025) );
ao12s01 g774211 ( .a(n_6924), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_14_), .o(n_7024) );
ao12s02 g774212 ( .a(n_6658), .b(n_6591), .c(n_6630), .o(n_6753) );
in01s01 g774214 ( .a(n_7034), .o(n_7035) );
ao12s01 g774215 ( .a(n_6985), .b(n_6806), .c(delay_xor_ln22_unr6_stage3_stallmux_q_14_), .o(n_7034) );
in01s01 g774216 ( .a(n_6689), .o(n_6690) );
ao12s01 g774217 ( .a(n_6633), .b(FE_OCP_RBN2382_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln21_unr6_stage3_stallmux_q_8_), .o(n_6689) );
in01s01 g774218 ( .a(n_6855), .o(n_6856) );
ao12s01 g774219 ( .a(n_6770), .b(FE_OCP_RBN6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln21_unr6_stage3_stallmux_q_10_), .o(n_6855) );
ao12s01 g774220 ( .a(n_7006), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_15_), .o(n_7187) );
in01s01 g774221 ( .a(n_6926), .o(n_6927) );
ao12s01 g774222 ( .a(n_6870), .b(n_6806), .c(delay_xor_ln22_unr6_stage3_stallmux_q_12_), .o(n_6926) );
in01s01 g774223 ( .a(n_6731), .o(n_6732) );
ao12s01 g774224 ( .a(n_6644), .b(FE_OCP_RBN6508_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln22_unr6_stage3_stallmux_q_8_), .o(n_6731) );
in01s01 g774227 ( .a(n_6852), .o(n_6853) );
ao12s01 g774228 ( .a(n_6747), .b(FE_OCP_RBN6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln22_unr6_stage3_stallmux_q_10_), .o(n_6852) );
in01s01 g774229 ( .a(n_6665), .o(n_6666) );
no02s02 g774230 ( .a(n_6578), .b(n_6552), .o(n_6665) );
in01s01 g774231 ( .a(n_6596), .o(n_6597) );
ao12s02 g774232 ( .a(n_6560), .b(FE_OCP_RBN6508_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln21_unr6_stage3_stallmux_q_6_), .o(n_6596) );
ao12s01 g774233 ( .a(n_6758), .b(FE_OCP_RBN6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln22_unr6_stage3_stallmux_q_9_), .o(n_6882) );
in01s01 g774234 ( .a(n_6609), .o(n_6610) );
ao22s01 g774235 ( .a(n_6580), .b(FE_OCP_RBN6507_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(FE_OCP_RBN6508_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .d(delay_xor_ln22_unr6_stage3_stallmux_q_6_), .o(n_6609) );
ao12s02 g774236 ( .a(n_7100), .b(n_6806), .c(delay_xor_ln22_unr6_stage3_stallmux_q_17_), .o(n_7190) );
in01s01 g774237 ( .a(n_6594), .o(n_6595) );
ao22s01 g774238 ( .a(FE_OCP_RBN6439_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_5_), .c(n_6496), .d(FE_OCP_RBN5504_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6594) );
ao12s01 g774239 ( .a(n_6651), .b(FE_OCP_RBN6508_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln21_unr6_stage3_stallmux_q_7_), .o(n_6932) );
in01s04 g774240 ( .a(n_6637), .o(n_6638) );
in01s01 g774242 ( .a(n_6652), .o(n_6653) );
na02s03 TIMEBOOST_cell_7948 ( .a(FE_OCP_RBN6086_n_10852), .b(FE_OCPN4844_FE_OFN4779_n_44490), .o(TIMEBOOST_net_2605) );
ao22s01 g774245 ( .a(n_6506), .b(FE_OCP_RBN5503_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(FE_OCP_RBN6439_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .d(delay_xor_ln21_unr6_stage3_stallmux_q_5_), .o(n_6601) );
in01s01 g774246 ( .a(n_6660), .o(n_6661) );
ao12s01 g774247 ( .a(n_6570), .b(FE_OCP_RBN6508_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln22_unr6_stage3_stallmux_q_7_), .o(n_6660) );
na03f08 TIMEBOOST_cell_7195 ( .a(n_13406), .b(n_13334), .c(n_13386), .o(n_13496) );
in01s01 g774249 ( .a(n_7077), .o(n_7078) );
ao12s01 g774250 ( .a(n_7029), .b(n_6806), .c(delay_xor_ln22_unr6_stage3_stallmux_q_16_), .o(n_7077) );
oa12s01 g774251 ( .a(n_6585), .b(n_6664), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_28_), .o(n_6769) );
oa12s01 g774252 ( .a(n_6624), .b(n_6828), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_30_), .o(n_6829) );
in01s01 g774253 ( .a(n_6818), .o(n_6819) );
oa12s01 g774254 ( .a(FE_RN_2534_0), .b(n_6862), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_22_), .o(n_6818) );
oa12s01 g774255 ( .a(n_6789), .b(n_6773), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_20_), .o(n_6851) );
in01s01 g774256 ( .a(n_6590), .o(n_6674) );
ao12s01 g774260 ( .a(n_6583), .b(n_6582), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_), .o(n_7630) );
ao22m02 g774262 ( .a(n_44711), .b(FE_OCP_RBN6240_n_6438), .c(n_44710), .d(n_6438), .o(n_6567) );
in01s01 g774264 ( .a(n_6670), .o(n_6646) );
oa12s02 g774266 ( .a(n_6341), .b(n_6487), .c(n_6382), .o(n_6488) );
ao12s04 g774267 ( .a(n_6342), .b(n_44711), .c(n_6383), .o(n_6502) );
ao12s02 g774268 ( .a(n_6370), .b(n_6513), .c(n_6394), .o(n_6555) );
oa12s04 g774269 ( .a(n_6395), .b(FE_OCP_RBN3444_n_6513), .c(n_6279), .o(n_6581) );
ao12f04 g774271 ( .a(n_6425), .b(n_6362), .c(n_6491), .o(n_6565) );
oa12s02 g774272 ( .a(n_6414), .b(n_6487), .c(n_6295), .o(n_6493) );
ao12s04 g774273 ( .a(n_6391), .b(n_44711), .c(n_6291), .o(n_6503) );
ao12s02 g774274 ( .a(n_6389), .b(n_6513), .c(n_6380), .o(n_6554) );
oa12s04 g774275 ( .a(n_6390), .b(FE_OCP_RBN3446_n_6513), .c(n_6371), .o(n_6572) );
na02s01 g774278 ( .a(n_6717), .b(n_6737), .o(n_6718) );
na02s01 g774279 ( .a(n_6895), .b(n_6857), .o(n_6858) );
no02s01 g774281 ( .a(n_6733), .b(n_6696), .o(n_6767) );
na02s02 g774282 ( .a(n_6628), .b(n_6705), .o(n_6706) );
no02s01 g774283 ( .a(n_6684), .b(n_6585), .o(n_6695) );
no02s01 g774285 ( .a(n_6863), .b(n_6850), .o(n_6942) );
no02s01 g774286 ( .a(n_6756), .b(n_6755), .o(n_6813) );
na02s01 g774287 ( .a(n_6830), .b(n_6703), .o(n_6704) );
no02s01 g774290 ( .a(n_6815), .b(n_6816), .o(n_6817) );
no02s01 g774291 ( .a(n_6742), .b(n_6741), .o(n_6743) );
no02s01 g774293 ( .a(n_6684), .b(n_6683), .o(n_7056) );
no02s03 g774294 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_4_), .b(FE_OCP_RBN6435_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6600) );
in01s01 g774295 ( .a(n_6642), .o(n_6571) );
na02s01 g774296 ( .a(FE_OCP_RBN5437_delay_xor_ln22_unr6_stage3_stallmux_q_0_), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6546) );
na02s06 g774297 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(FE_OCP_RBN5436_delay_xor_ln22_unr6_stage3_stallmux_q_0_), .o(n_6642) );
no02s01 g774298 ( .a(n_6688), .b(n_6687), .o(n_7170) );
no02s01 g774299 ( .a(n_6621), .b(n_6620), .o(n_6899) );
no02s06 g774300 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_13_), .o(n_6964) );
no02s02 g774301 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_15_), .o(n_7033) );
in01s01 g774302 ( .a(n_6770), .o(n_6771) );
no02s01 g774303 ( .a(FE_OCP_RBN6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_10_), .o(n_6770) );
in01s01 g774305 ( .a(n_6976), .o(n_6977) );
na02s01 g774306 ( .a(n_6938), .b(n_6879), .o(n_6976) );
in01s01 g774307 ( .a(n_6560), .o(n_6876) );
no02s02 g774308 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_6_), .b(FE_OCP_RBN6440_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6560) );
no02s02 g774310 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_15_), .o(n_7006) );
no02s01 g774311 ( .a(n_6863), .b(n_6862), .o(n_7428) );
in01s01 g774313 ( .a(n_6716), .o(n_6547) );
no02m03 g774314 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_3_), .b(FE_OCP_RBN6435_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6716) );
no02s01 g774315 ( .a(n_6551), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6552) );
no02s06 g774316 ( .a(FE_OCP_RBN6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_9_), .o(n_6772) );
no02s06 g774317 ( .a(FE_OCP_RBN6435_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_3_), .o(n_6708) );
in01s01 g774319 ( .a(n_6870), .o(n_6871) );
no02m01 g774320 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_12_), .b(n_6806), .o(n_6870) );
na02s06 g774321 ( .a(n_6580), .b(FE_OCP_RBN6507_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6801) );
in01s01 g774322 ( .a(n_6577), .o(n_6578) );
na02s06 g774323 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n_6551), .o(n_6577) );
no02s03 g774324 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_4_), .b(FE_OCP_RBN6435_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6715) );
in01s01 g774325 ( .a(n_6644), .o(n_6645) );
no02m01 g774326 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_8_), .b(FE_OCP_RBN6508_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6644) );
in01s01 g774327 ( .a(n_6633), .o(n_6634) );
no02s06 g774328 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_8_), .b(FE_OCP_RBN6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6633) );
no02s06 g774329 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_11_), .o(n_6880) );
no02s04 g774330 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_5_), .b(FE_OCP_RBN6440_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6531) );
in01s01 g774331 ( .a(n_6924), .o(n_6925) );
no02s01 g774332 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_14_), .b(n_6806), .o(n_6924) );
na02s02 g774333 ( .a(n_6667), .b(n_5471), .o(n_6668) );
no02s02 g774334 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_17_), .o(n_7100) );
na03m02 TIMEBOOST_cell_4832 ( .a(n_39719), .b(FE_OCP_RBN3285_n_39674), .c(n_39728), .o(n_39764) );
na02m08 TIMEBOOST_cell_3844 ( .a(TIMEBOOST_net_1012), .b(n_32698), .o(n_32775) );
na02s01 g774337 ( .a(n_6697), .b(n_6737), .o(n_7297) );
in01s01 g774338 ( .a(n_7121), .o(n_7122) );
no02s02 g774339 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_18_), .o(n_7121) );
no02s02 g774340 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_13_), .b(n_6806), .o(n_6951) );
no02s02 g774341 ( .a(FE_OCP_RBN6439_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_5_), .o(n_6523) );
in01s02 g774342 ( .a(n_7029), .o(n_7030) );
no02s03 g774343 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_16_), .o(n_7029) );
na02s10 g774344 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n_6507), .o(n_6619) );
no02s01 g774345 ( .a(n_6865), .b(n_6940), .o(n_7316) );
no02s01 g774346 ( .a(n_6582), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_), .o(n_6583) );
no02m01 g774347 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_9_), .b(FE_OCP_RBN6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6758) );
in01s01 g774348 ( .a(n_6998), .o(n_6999) );
no02s01 g774349 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_16_), .o(n_6998) );
no04s03 TIMEBOOST_cell_4714 ( .a(n_42370), .b(FE_RN_663_0), .c(FE_RN_665_0), .d(FE_RN_664_0), .o(FE_RN_668_0) );
in01s01 g774351 ( .a(n_6651), .o(n_6539) );
no02s02 g774352 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_7_), .b(FE_OCP_RBN6440_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6651) );
in01s02 g774353 ( .a(n_6570), .o(n_6831) );
no02m01 g774354 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_7_), .b(FE_OCP_RBN6508_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6570) );
in01s01 g774355 ( .a(n_6747), .o(n_6748) );
no02s01 g774356 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_10_), .b(FE_OCP_RBN6510_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6747) );
in01s01 g774357 ( .a(n_6868), .o(n_6869) );
no02s02 g774358 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_12_), .b(n_6806), .o(n_6868) );
in01s01 g774359 ( .a(n_6985), .o(n_6986) );
no02s01 g774360 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_14_), .o(n_6985) );
no02m10 g774361 ( .a(n_6528), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_), .o(n_6671) );
no02s03 g774362 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_11_), .b(n_6806), .o(n_6873) );
na02s01 g774363 ( .a(n_6844), .b(n_6939), .o(n_7449) );
no02s01 g774364 ( .a(n_6741), .b(n_6625), .o(n_7242) );
in01s02 g774365 ( .a(n_6656), .o(n_6579) );
na02s10 g774366 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n_6510), .o(n_6656) );
in01s01 g774367 ( .a(n_7097), .o(n_7098) );
no02s01 g774368 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_18_), .o(n_7097) );
na02s01 g774369 ( .a(n_6857), .b(n_6887), .o(n_7392) );
na02s01 g774370 ( .a(n_6703), .b(n_6722), .o(n_7564) );
no02s01 g774371 ( .a(n_6641), .b(n_6541), .o(n_7012) );
no02s01 g774372 ( .a(n_6593), .b(n_6562), .o(n_6672) );
na02s01 g774373 ( .a(n_6783), .b(n_6782), .o(n_7473) );
no02s01 g774374 ( .a(n_6816), .b(n_6828), .o(n_7550) );
no02s01 g774375 ( .a(n_6658), .b(n_6592), .o(n_7229) );
in01s01 g774376 ( .a(n_6962), .o(n_6963) );
na02s01 g774377 ( .a(n_6944), .b(n_6721), .o(n_6962) );
in01s01 g774378 ( .a(n_6920), .o(n_6921) );
ao12s01 g774379 ( .a(n_6749), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_18_), .o(n_6920) );
ao12s01 g774380 ( .a(n_6815), .b(n_6624), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_30_), .o(n_7623) );
ao12s01 g774381 ( .a(n_6764), .b(n_6624), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_28_), .o(n_7602) );
in01s01 g774382 ( .a(n_6922), .o(n_6923) );
ao12s01 g774383 ( .a(n_6755), .b(n_6624), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_26_), .o(n_6922) );
ao12s01 g774384 ( .a(n_6826), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_20_), .o(n_7408) );
ao12s01 g774385 ( .a(n_6850), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_22_), .o(n_7481) );
in01s01 g774386 ( .a(n_6892), .o(n_6893) );
ao12s01 g774387 ( .a(n_6742), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_12_), .o(n_6892) );
ao12s01 g774388 ( .a(n_6836), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_16_), .o(n_7313) );
oa22s01 g774389 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_8_), .c(n_6521), .d(n_5104), .o(n_7110) );
in01s02 g774391 ( .a(n_6529), .o(n_6519) );
oa12s01 g774394 ( .a(n_6854), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_), .o(n_7302) );
oa12s01 g774396 ( .a(n_6849), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_), .o(n_6965) );
oa22s01 g774397 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_4_), .c(n_6521), .d(n_6761), .o(n_6956) );
in01s01 g774398 ( .a(n_6643), .o(n_6587) );
in01s01 g774400 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_6_), .o(n_6580) );
in01s01 g774405 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_5_), .o(n_6496) );
in01s01 g774407 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_4_), .o(n_6504) );
in01s06 g774421 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_0_), .o(n_6510) );
in01s06 g774425 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_2_), .o(n_6551) );
in01s01 g774429 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_5_), .o(n_6506) );
in01s01 g774433 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_25_), .o(n_6509) );
in01s01 g774440 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_4_), .o(n_6512) );
in01m06 g774442 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_2_), .o(n_6542) );
in01s01 g774445 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_26_), .o(n_6631) );
in01s06 g774447 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_1_), .o(n_6507) );
na02s01 g774454 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_), .o(n_6849) );
no02s01 g774456 ( .a(FE_RN_2534_0), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_18_), .o(n_6749) );
no02s01 g774458 ( .a(FE_RN_2534_0), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_17_), .o(n_6940) );
in01s01 g774459 ( .a(n_6864), .o(n_6865) );
na02s01 g774460 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_17_), .o(n_6864) );
in01s01 g774461 ( .a(n_6626), .o(n_6684) );
na02s01 g774462 ( .a(n_6563), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_7_), .o(n_6626) );
na02s01 g774463 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_), .o(n_6938) );
na02s01 g774464 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_23_), .o(n_6844) );
no02s01 g774466 ( .a(FE_RN_2534_0), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_20_), .o(n_6826) );
na02s01 g774467 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_), .o(n_6854) );
no02s01 g774468 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_16_), .o(n_6836) );
no02s01 g774469 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_12_), .o(n_6742) );
no02s02 g774470 ( .a(n_6563), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_5_), .o(n_6620) );
in01s01 g774471 ( .a(n_6630), .o(n_6688) );
na02s01 g774472 ( .a(n_6586), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_9_), .o(n_6630) );
in01s01 g774474 ( .a(n_6857), .o(n_6773) );
na02s02 g774475 ( .a(FE_RN_2534_0), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_19_), .o(n_6857) );
na02s06 g774476 ( .a(n_6563), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_), .o(n_6564) );
no02s01 g774477 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_22_), .o(n_6850) );
no02s01 g774478 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_11_), .o(n_6741) );
in01s01 g774479 ( .a(n_6687), .o(n_6628) );
no02s01 g774480 ( .a(n_6586), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_9_), .o(n_6687) );
no02s01 g774481 ( .a(FE_RN_2534_0), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_21_), .o(n_6863) );
in01s01 g774482 ( .a(n_6569), .o(n_6621) );
na02m01 g774483 ( .a(n_6563), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_5_), .o(n_6569) );
in01s01 g774484 ( .a(n_6667), .o(n_6625) );
na02s01 g774485 ( .a(n_6586), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_11_), .o(n_6667) );
in01s01 g774486 ( .a(n_6878), .o(n_6879) );
no02s01 g774487 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_), .o(n_6878) );
no02s01 g774489 ( .a(n_6563), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_7_), .o(n_6683) );
no02s01 g774490 ( .a(n_6556), .b(n_6061), .o(n_6862) );
na02s01 g774491 ( .a(n_6586), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_15_), .o(n_6737) );
in01s01 g774492 ( .a(n_6696), .o(n_6697) );
no02s01 g774493 ( .a(n_6586), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_15_), .o(n_6696) );
na02s01 g774494 ( .a(n_6556), .b(n_5984), .o(n_6887) );
in01s01 g774495 ( .a(n_6877), .o(n_6939) );
no02s01 g774496 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_23_), .o(n_6877) );
no02s01 g774497 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_29_), .o(n_6816) );
in01s01 g774498 ( .a(n_6561), .o(n_6562) );
na02s10 g774499 ( .a(n_6524), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_2_), .o(n_6561) );
no02s06 g774500 ( .a(n_6585), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_6_), .o(n_6641) );
in01s01 g774501 ( .a(n_6591), .o(n_6592) );
na02s01 g774502 ( .a(n_6585), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_10_), .o(n_6591) );
na02s02 g774503 ( .a(n_6521), .b(n_6142), .o(n_6783) );
no02s10 g774504 ( .a(n_6524), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_2_), .o(n_6593) );
in01s01 g774505 ( .a(n_6756), .o(n_6721) );
no02s01 g774506 ( .a(n_6585), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_25_), .o(n_6756) );
na02s01 g774507 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_25_), .o(n_6944) );
in01s01 g774508 ( .a(n_6703), .o(n_6664) );
na02s01 g774509 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_27_), .o(n_6703) );
no02s01 g774510 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_30_), .o(n_6815) );
no02s01 g774511 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_28_), .o(n_6764) );
no02s01 g774512 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_26_), .o(n_6755) );
in01s01 g774513 ( .a(n_6658), .o(n_6705) );
no02s01 g774514 ( .a(n_6585), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_10_), .o(n_6658) );
in01s01 g774515 ( .a(n_6540), .o(n_6541) );
na02s01 g774516 ( .a(n_6524), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_6_), .o(n_6540) );
in01s01 g774517 ( .a(n_6765), .o(n_6722) );
no02s01 g774518 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_27_), .o(n_6765) );
na02s01 g774519 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_24_), .o(n_6782) );
no02s01 g774520 ( .a(n_6521), .b(n_6473), .o(n_6828) );
oa12s01 g774521 ( .a(FE_RN_2534_0), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_18_), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_17_), .o(n_6895) );
ao12s01 g774522 ( .a(n_6586), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_), .o(n_6733) );
oa12s01 g774523 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_26_), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_25_), .o(n_6830) );
oa12s01 g774525 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_), .o(n_6717) );
no02m06 TIMEBOOST_cell_4474 ( .a(TIMEBOOST_net_1327), .b(FE_OCP_RBN7055_FE_OCPN1068_n_21973), .o(FE_RN_938_0) );
no02m06 TIMEBOOST_cell_8560 ( .a(n_29545), .b(n_29630), .o(TIMEBOOST_net_2767) );
in01s01 g774529 ( .a(n_6528), .o(n_6582) );
in01m06 g774534 ( .a(n_6491), .o(n_6513) );
na02f08 g774538 ( .a(n_6416), .b(n_6387), .o(n_6491) );
in01s01 g774544 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_29_), .o(n_6473) );
in01s01 g774547 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_23_), .o(n_6413) );
no02s01 g774549 ( .a(n_6806), .b(n_6505), .o(n_7070) );
in01f01 g774561 ( .a(n_6521), .o(n_6624) );
in01s06 g774563 ( .a(n_6521), .o(n_6585) );
in01s06 g774564 ( .a(n_6524), .o(n_6521) );
na02s20 g774565 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n_6505), .o(n_6524) );
in01s02 g774571 ( .a(n_6556), .o(n_6789) );
in01s02 g774579 ( .a(n_6556), .o(n_6676) );
in01s02 g774582 ( .a(n_6556), .o(n_6586) );
in01s02 g774584 ( .a(n_6563), .o(n_6556) );
in01s06 g774585 ( .a(n_6517), .o(n_6563) );
no02s10 g774586 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n_6505), .o(n_6517) );
no03s20 TIMEBOOST_cell_3433 ( .a(n_17084), .b(FE_OCP_RBN7108_n_44365), .c(FE_RN_2347_0), .o(n_17072) );
no02f08 TIMEBOOST_cell_1150 ( .a(n_18237), .b(TIMEBOOST_net_189), .o(n_45524) );
na02s01 TIMEBOOST_cell_3339 ( .a(TIMEBOOST_net_960), .b(n_36343), .o(n_36424) );
oa12m01 g774603 ( .a(n_6222), .b(n_6373), .c(n_6244), .o(n_6388) );
na03s02 TIMEBOOST_cell_8708 ( .a(n_6932), .b(n_6937), .c(FE_RN_249_0), .o(TIMEBOOST_net_2841) );
in01s02 g774605 ( .a(n_46993), .o(n_6479) );
na02m04 g774608 ( .a(n_6359), .b(n_6320), .o(n_6404) );
oa12s02 g774618 ( .a(FE_OCP_RBN3404_n_6205), .b(n_6485), .c(n_6213), .o(n_6489) );
no02s02 g774619 ( .a(FE_OCP_RBN3405_n_6205), .b(n_6486), .o(n_6499) );
ao22f04 g774627 ( .a(n_6356), .b(n_6334), .c(n_6357), .d(n_6335), .o(n_6477) );
ao22s02 g774635 ( .a(FE_OCP_RBN3436_n_6485), .b(n_6308), .c(n_6485), .d(n_6309), .o(n_6557) );
in01s40 g774638 ( .a(delay_xor_ln23_unr6_stage3_stallmux_q), .o(n_6505) );
in01s01 g774657 ( .a(FE_OCP_RBN3997_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_7217) );
in01s01 g774662 ( .a(FE_OCP_RBN3997_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_7172) );
in01s01 g774665 ( .a(FE_OCP_RBN3998_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6872) );
in01s06 g774686 ( .a(FE_OCP_RBN3998_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6806) );
no03f04 TIMEBOOST_cell_3517 ( .a(FE_OCP_RBN2508_n_37720), .b(n_38047), .c(n_37723), .o(n_37801) );
no02s02 g774710 ( .a(n_6485), .b(n_6213), .o(n_6486) );
in01f02 g774712 ( .a(n_6358), .o(n_6359) );
no02s01 TIMEBOOST_cell_1493 ( .a(n_8550), .b(n_7965), .o(TIMEBOOST_net_361) );
oa22s01 g774715 ( .a(n_6346), .b(n_5403), .c(n_6345), .d(n_5404), .o(n_6405) );
oa22s01 g774716 ( .a(n_6317), .b(n_5416), .c(n_6316), .d(n_5415), .o(n_6384) );
no02s06 TIMEBOOST_cell_1149 ( .a(FE_RN_23_0), .b(n_17533), .o(TIMEBOOST_net_189) );
in01s02 g774719 ( .a(n_6376), .o(n_6365) );
no02s02 TIMEBOOST_cell_1490 ( .a(TIMEBOOST_net_359), .b(FE_OCP_RBN2798_n_8817), .o(n_8921) );
in01s01 g774721 ( .a(n_6500), .o(n_6490) );
na02f08 TIMEBOOST_cell_4005 ( .a(n_35000), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(TIMEBOOST_net_1093) );
in01s01 g774723 ( .a(n_6382), .o(n_6383) );
in01s02 g774724 ( .a(n_6363), .o(n_6382) );
no03s20 TIMEBOOST_cell_3432 ( .a(n_11919), .b(FE_RN_141_0), .c(FE_OCP_RBN6309_n_45224), .o(n_11772) );
na02m04 g774726 ( .a(n_6348), .b(n_6329), .o(n_6393) );
in01s01 g774728 ( .a(n_6371), .o(n_6380) );
no02f06 g774729 ( .a(n_6228), .b(n_6294), .o(n_6371) );
in01s01 g774730 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_21_), .o(n_7401) );
in01s01 g774735 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_24_), .o(n_7521) );
na02s02 g774739 ( .a(n_6239), .b(n_6169), .o(n_6277) );
in01s01 g774740 ( .a(n_6408), .o(n_6409) );
na02s02 g774741 ( .a(n_6395), .b(n_6394), .o(n_6408) );
in01s01 g774742 ( .a(n_6350), .o(n_6351) );
no02m01 g774743 ( .a(n_6321), .b(FE_OCP_RBN4488_n_6299), .o(n_6350) );
na02s02 g774745 ( .a(n_6414), .b(n_6265), .o(n_6438) );
no02s02 g774746 ( .a(n_6319), .b(n_6328), .o(n_6329) );
no03s10 TIMEBOOST_cell_3431 ( .a(FE_OCP_RBN6313_n_45224), .b(n_11882), .c(FE_RN_138_0), .o(n_11763) );
no02f06 g774748 ( .a(n_6287), .b(n_6213), .o(n_6288) );
no02m06 g774749 ( .a(n_6272), .b(FE_OCP_RBN3286_n_5656), .o(n_6294) );
no02m08 TIMEBOOST_cell_5535 ( .a(TIMEBOOST_net_1715), .b(n_36608), .o(n_36667) );
no02s01 TIMEBOOST_cell_1489 ( .a(n_7737), .b(n_8846), .o(TIMEBOOST_net_359) );
no02s02 g774752 ( .a(FE_OCP_RBN4489_n_6299), .b(n_6319), .o(n_6320) );
na02s06 g774755 ( .a(n_6355), .b(n_6262), .o(n_6485) );
na02m08 TIMEBOOST_cell_2891 ( .a(n_2158), .b(TIMEBOOST_net_736), .o(n_2222) );
in01s01 g774757 ( .a(n_6398), .o(n_6399) );
no02s02 g774758 ( .a(n_6310), .b(n_6287), .o(n_6398) );
oa12s04 g774760 ( .a(n_6220), .b(n_45217), .c(n_6173), .o(n_6332) );
in01s04 g774761 ( .a(n_6356), .o(n_6357) );
in01m04 g774762 ( .a(n_6373), .o(n_6356) );
na02f06 g774763 ( .a(n_6253), .b(n_6230), .o(n_6373) );
in01s01 g774764 ( .a(n_6465), .o(n_6466) );
no02m02 TIMEBOOST_cell_6626 ( .a(TIMEBOOST_net_2070), .b(n_12590), .o(TIMEBOOST_net_1437) );
na02s02 g774767 ( .a(n_6412), .b(n_6326), .o(n_6471) );
ao22f01 g774769 ( .a(n_6328), .b(n_6226), .c(n_45216), .d(n_6225), .o(n_6379) );
in01m02 g774770 ( .a(n_6347), .o(n_6348) );
na02m06 g774771 ( .a(n_6241), .b(n_6299), .o(n_6347) );
in01s02 g774772 ( .a(n_6447), .o(n_6448) );
na02s02 g774773 ( .a(n_6340), .b(n_6353), .o(n_6447) );
in01s01 g774774 ( .a(n_6476), .o(n_6436) );
no02s01 TIMEBOOST_cell_1416 ( .a(n_24671), .b(TIMEBOOST_net_322), .o(n_24816) );
in01s02 g774776 ( .a(n_6442), .o(n_6443) );
no02s02 g774777 ( .a(n_6415), .b(n_6330), .o(n_6442) );
no02f02 TIMEBOOST_cell_5558 ( .a(FE_OCP_RBN1850_n_25898), .b(n_23317), .o(TIMEBOOST_net_1727) );
in01s01 g774780 ( .a(n_6453), .o(n_6454) );
na02s02 g774781 ( .a(n_6352), .b(n_6325), .o(n_6453) );
in01s01 g774782 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_22_), .o(n_7467) );
in01s01 g774784 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_19_), .o(n_7344) );
na02s01 g774786 ( .a(n_45474), .b(n_5693), .o(n_6340) );
no02m04 g774787 ( .a(n_45479), .b(FE_OCPN7087_n_6263), .o(n_6321) );
na02s01 g774788 ( .a(n_45474), .b(FE_OCP_RBN3319_n_5555), .o(n_6327) );
no02m06 g774789 ( .a(n_6230), .b(n_6240), .o(n_6231) );
in01s02 g774790 ( .a(n_6354), .o(n_6355) );
no02m08 g774791 ( .a(n_6324), .b(n_6219), .o(n_6354) );
in01s01 g774792 ( .a(n_6295), .o(n_6291) );
in01s01 g774794 ( .a(n_6265), .o(n_6295) );
na02s02 g774795 ( .a(n_6214), .b(n_5523), .o(n_6265) );
na02m06 g774796 ( .a(n_6261), .b(n_6205), .o(n_6298) );
na02s02 g774797 ( .a(n_45475), .b(n_5732), .o(n_6353) );
na02s06 g774798 ( .a(n_45214), .b(n_6192), .o(n_6253) );
na02s06 g774801 ( .a(n_45479), .b(FE_OCPN7087_n_6263), .o(n_6299) );
no02s02 TIMEBOOST_cell_7042 ( .a(TIMEBOOST_net_2279), .b(n_5130), .o(TIMEBOOST_net_1659) );
in01s02 g774803 ( .a(n_6334), .o(n_6335) );
no02s02 g774804 ( .a(n_6244), .b(n_6240), .o(n_6334) );
na02s01 g774805 ( .a(n_45474), .b(n_5609), .o(n_6326) );
in01s01 g774806 ( .a(n_6394), .o(n_6279) );
in01s01 g774807 ( .a(n_6272), .o(n_6394) );
no02m06 g774808 ( .a(n_6228), .b(FE_OCP_RBN3281_n_5614), .o(n_6272) );
na02s02 g774809 ( .a(n_6290), .b(FE_OCP_RBN3286_n_5656), .o(n_6352) );
na02s01 g774810 ( .a(n_6228), .b(n_5703), .o(n_6325) );
na02s02 TIMEBOOST_cell_5523 ( .a(TIMEBOOST_net_1709), .b(n_11586), .o(n_11739) );
in01s01 g774812 ( .a(n_6368), .o(n_6369) );
na02s01 g774813 ( .a(n_6324), .b(n_6234), .o(n_6368) );
no02s01 TIMEBOOST_cell_1415 ( .a(n_24047), .b(n_24063), .o(TIMEBOOST_net_322) );
na02s02 g774815 ( .a(n_6312), .b(n_6171), .o(n_6360) );
in01s01 g774816 ( .a(n_6395), .o(n_6370) );
na02s02 g774817 ( .a(n_6228), .b(FE_OCP_RBN3281_n_5614), .o(n_6395) );
in01s01 g774818 ( .a(n_6308), .o(n_6309) );
no02s02 g774819 ( .a(FE_OCP_RBN3405_n_6205), .b(n_6213), .o(n_6308) );
no02m04 g774820 ( .a(n_6240), .b(n_6191), .o(n_6241) );
no02s01 g774821 ( .a(n_6228), .b(n_5780), .o(n_6330) );
in01s01 g774822 ( .a(n_6414), .o(n_6391) );
na02s02 g774823 ( .a(n_45475), .b(FE_OCP_RBN6113_n_5444), .o(n_6414) );
no02s02 g774825 ( .a(n_6290), .b(n_5754), .o(n_6415) );
na02s01 g774826 ( .a(n_6228), .b(FE_OCP_RBN3326_n_5813), .o(n_6338) );
in01s01 g774827 ( .a(n_6386), .o(n_6310) );
na02s08 g774828 ( .a(n_6228), .b(FE_OCPN6289_FE_OCP_RBN3263_n_5531), .o(n_6386) );
no02f08 g774829 ( .a(n_6228), .b(FE_OCPN6289_FE_OCP_RBN3263_n_5531), .o(n_6287) );
in01s01 g774830 ( .a(n_6412), .o(n_6396) );
na02s02 g774831 ( .a(n_45475), .b(n_5648), .o(n_6412) );
no03s40 TIMEBOOST_cell_4197 ( .a(FE_RN_105_0), .b(n_40624), .c(n_44610), .o(TIMEBOOST_net_1189) );
in01s01 g774833 ( .a(n_6345), .o(n_6346) );
no02s01 g774834 ( .a(n_6315), .b(n_5439), .o(n_6345) );
in01s01 g774835 ( .a(n_6316), .o(n_6317) );
ao12s01 g774836 ( .a(n_5260), .b(n_6266), .c(n_5329), .o(n_6316) );
in01s01 g774837 ( .a(n_6389), .o(n_6390) );
in01s01 g774838 ( .a(n_6362), .o(n_6389) );
na02s02 g774839 ( .a(n_6228), .b(n_5706), .o(n_6362) );
oa22s01 g774840 ( .a(n_6209), .b(n_5380), .c(n_6210), .d(n_5381), .o(n_6286) );
oa22s01 g774841 ( .a(n_6259), .b(n_5333), .c(n_6260), .d(n_5334), .o(n_6323) );
in01s01 g774842 ( .a(n_6435), .o(n_6407) );
no02f06 TIMEBOOST_cell_1418 ( .a(n_24791), .b(TIMEBOOST_net_323), .o(n_24906) );
in01s02 g774844 ( .a(n_6313), .o(n_6285) );
no02s01 TIMEBOOST_cell_1478 ( .a(n_42007), .b(TIMEBOOST_net_353), .o(n_42079) );
in01m01 g774846 ( .a(n_6238), .o(n_6239) );
oa12s01 g774847 ( .a(n_6012), .b(n_6178), .c(n_6080), .o(n_6238) );
in01s01 g774848 ( .a(n_6341), .o(n_6342) );
in01s01 g774849 ( .a(n_6319), .o(n_6341) );
no02s06 g774850 ( .a(n_45474), .b(n_5637), .o(n_6319) );
in01s02 g774851 ( .a(n_46994), .o(n_6318) );
na02s06 TIMEBOOST_cell_8711 ( .a(TIMEBOOST_net_2842), .b(n_11999), .o(n_12100) );
no02m08 g774857 ( .a(n_6266), .b(n_6250), .o(n_6315) );
no02m08 g774861 ( .a(n_6177), .b(n_5320), .o(n_6244) );
in01s01 g774862 ( .a(n_6222), .o(n_6223) );
in01s01 g774863 ( .a(n_6240), .o(n_6222) );
no02s08 g774864 ( .a(FE_OCP_RBN3276_n_5284), .b(n_6176), .o(n_6240) );
no02s01 TIMEBOOST_cell_1477 ( .a(n_41600), .b(n_41614), .o(TIMEBOOST_net_353) );
no02m04 g774869 ( .a(n_6196), .b(FE_OCPN6287_FE_OCP_RBN6082_n_5454), .o(n_6213) );
na02s02 g774870 ( .a(n_6178), .b(n_6119), .o(n_6224) );
na02m06 g774875 ( .a(n_6196), .b(FE_OCPN6287_FE_OCP_RBN6082_n_5454), .o(n_6205) );
no02f08 g774881 ( .a(n_6145), .b(n_6158), .o(n_6328) );
na02f06 g774882 ( .a(n_6270), .b(n_6186), .o(n_6324) );
na02s01 g774883 ( .a(n_6282), .b(n_6203), .o(n_6343) );
no02s04 TIMEBOOST_cell_1417 ( .a(n_24193), .b(n_24354), .o(TIMEBOOST_net_323) );
na02s02 g774885 ( .a(n_6182), .b(n_6033), .o(n_6208) );
in01s01 g774894 ( .a(n_6419), .o(n_6392) );
no02f10 TIMEBOOST_cell_1502 ( .a(n_34572), .b(TIMEBOOST_net_365), .o(n_34820) );
in01s01 g774896 ( .a(n_6311), .o(n_6312) );
oa12s02 g774897 ( .a(n_6187), .b(n_6237), .c(n_6087), .o(n_6311) );
in01s02 g774898 ( .a(n_6297), .o(n_6254) );
no02f10 TIMEBOOST_cell_1364 ( .a(n_24723), .b(TIMEBOOST_net_296), .o(n_24799) );
oa12m04 g774900 ( .a(n_6197), .b(n_6149), .c(n_6153), .o(n_6230) );
in01s01 g774901 ( .a(n_6261), .o(n_6262) );
ao12f04 g774902 ( .a(n_6198), .b(n_6235), .c(n_6234), .o(n_6261) );
in01s01 g774908 ( .a(n_6228), .o(n_6290) );
na02f10 g774911 ( .a(n_6151), .b(n_6122), .o(n_6228) );
na02f08 g774914 ( .a(n_6101), .b(n_6102), .o(n_6151) );
na02f06 g774915 ( .a(n_6100), .b(FE_OCP_RBN4455_n_6102), .o(n_6122) );
na02m04 g774918 ( .a(n_6144), .b(n_6040), .o(n_6178) );
no02m08 TIMEBOOST_cell_1501 ( .a(n_34413), .b(n_34462), .o(TIMEBOOST_net_365) );
no02m08 TIMEBOOST_cell_1363 ( .a(FE_RN_2361_0), .b(n_24646), .o(TIMEBOOST_net_296) );
na02s01 g774921 ( .a(n_6257), .b(n_6141), .o(n_6276) );
in01s01 g774922 ( .a(n_6281), .o(n_6282) );
in01s01 g774923 ( .a(n_6270), .o(n_6281) );
na02f04 g774924 ( .a(n_6201), .b(n_6189), .o(n_6270) );
na02s01 g774926 ( .a(n_6150), .b(n_6197), .o(n_6215) );
in01s02 g774927 ( .a(n_6191), .o(n_6192) );
na02s04 g774928 ( .a(n_6197), .b(n_6148), .o(n_6191) );
na02s04 g774929 ( .a(n_6139), .b(n_5900), .o(n_6190) );
in01s01 g774930 ( .a(n_6268), .o(n_6269) );
na02s01 g774931 ( .a(n_6235), .b(n_6218), .o(n_6268) );
in01s01 g774932 ( .a(n_6259), .o(n_6260) );
in01s01 g774933 ( .a(n_6266), .o(n_6259) );
no02f08 TIMEBOOST_cell_7914 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(FE_OCP_RBN6810_n_39551), .o(TIMEBOOST_net_2588) );
in01s01 g774935 ( .a(n_6209), .o(n_6210) );
ao12s01 g774936 ( .a(n_5241), .b(n_6160), .c(n_5368), .o(n_6209) );
in01s04 g774937 ( .a(n_6176), .o(n_6177) );
na02m08 g774938 ( .a(n_6110), .b(n_6104), .o(n_6176) );
in01m02 g774939 ( .a(n_6267), .o(n_6245) );
na02s01 TIMEBOOST_cell_1378 ( .a(TIMEBOOST_net_303), .b(n_24077), .o(n_24238) );
oa22s01 g774941 ( .a(n_6185), .b(n_5386), .c(n_6184), .d(n_5385), .o(n_6229) );
no02m06 g774942 ( .a(n_6144), .b(n_6114), .o(n_6145) );
in01m02 g774943 ( .a(n_6301), .o(n_6280) );
na02s01 TIMEBOOST_cell_6663 ( .a(FE_OCP_RBN6601_n_7708), .b(FE_RN_298_0), .o(TIMEBOOST_net_2089) );
in01m01 g774945 ( .a(n_6181), .o(n_6182) );
oa12s02 g774946 ( .a(n_6007), .b(n_6118), .c(n_5982), .o(n_6181) );
no02f08 TIMEBOOST_cell_7053 ( .a(n_45739), .b(n_39692), .o(TIMEBOOST_net_2285) );
in01s01 g774948 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_17_), .o(n_6167) );
in01s01 g774951 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_20_), .o(n_7424) );
na02m06 g774953 ( .a(n_6059), .b(n_6055), .o(n_6110) );
na02m04 g774954 ( .a(FE_OCP_RBN6171_n_6059), .b(n_6054), .o(n_6104) );
na02m06 g774955 ( .a(n_6135), .b(FE_OCP_RBN3236_n_5130), .o(n_6197) );
na02s01 TIMEBOOST_cell_1377 ( .a(n_23808), .b(n_24110), .o(TIMEBOOST_net_303) );
no02m08 TIMEBOOST_cell_7024 ( .a(TIMEBOOST_net_2270), .b(n_26044), .o(n_26194) );
in01s01 g774958 ( .a(n_6225), .o(n_6226) );
na02s02 g774959 ( .a(n_6220), .b(n_6148), .o(n_6225) );
in01s01 g774960 ( .a(n_6149), .o(n_6150) );
no02m04 g774961 ( .a(n_6135), .b(FE_OCP_RBN3236_n_5130), .o(n_6149) );
in01m04 g774962 ( .a(n_6218), .o(n_6219) );
in01m02 g774963 ( .a(n_6198), .o(n_6218) );
no02m04 g774964 ( .a(n_6165), .b(FE_OCP_RBN3239_n_5307), .o(n_6198) );
in01s01 g774965 ( .a(n_6203), .o(n_6204) );
na02s01 g774966 ( .a(n_6186), .b(n_6234), .o(n_6203) );
na02f04 TIMEBOOST_cell_7723 ( .a(TIMEBOOST_net_2492), .b(n_15504), .o(n_15584) );
na02s02 g774968 ( .a(n_6125), .b(n_5980), .o(n_6156) );
in01s01 g774970 ( .a(n_6237), .o(n_6257) );
na02s02 g774971 ( .a(n_6163), .b(n_6127), .o(n_6237) );
na02s02 g774972 ( .a(n_6180), .b(n_6117), .o(n_6207) );
na02m04 g774973 ( .a(n_6165), .b(FE_OCP_RBN3239_n_5307), .o(n_6235) );
no03f04 TIMEBOOST_cell_2749 ( .a(FE_OCP_RBN3174_n_26158), .b(FE_OCP_RBN6088_n_26181), .c(n_26302), .o(n_26327) );
oa12f04 g774975 ( .a(FE_OCP_RBN3357_n_6013), .b(n_6090), .c(n_6089), .o(n_6115) );
no02m08 TIMEBOOST_cell_1350 ( .a(n_24146), .b(TIMEBOOST_net_289), .o(n_24231) );
no02s10 TIMEBOOST_cell_4865 ( .a(n_169), .b(TIMEBOOST_net_1380), .o(n_170) );
in01f04 g774978 ( .a(n_6100), .o(n_6101) );
oa12f06 g774979 ( .a(n_5965), .b(n_5923), .c(n_6041), .o(n_6100) );
in01s02 g774981 ( .a(n_6138), .o(n_6139) );
oa12s04 g774982 ( .a(n_5823), .b(n_6082), .c(n_5681), .o(n_6138) );
in01s01 g774983 ( .a(n_6243), .o(n_6217) );
no02s01 TIMEBOOST_cell_1342 ( .a(n_41757), .b(TIMEBOOST_net_285), .o(n_41836) );
in01s02 g774985 ( .a(n_6233), .o(n_6212) );
no02s01 TIMEBOOST_cell_1332 ( .a(TIMEBOOST_net_280), .b(n_29175), .o(n_29287) );
na02m06 g774987 ( .a(n_6083), .b(n_5983), .o(n_6144) );
ao12f06 g774988 ( .a(n_6094), .b(n_6081), .c(n_6157), .o(n_6158) );
in01s01 g774990 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_18_), .o(n_7353) );
no02s04 TIMEBOOST_cell_1349 ( .a(n_24102), .b(FE_OFN743_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(TIMEBOOST_net_289) );
na02f08 TIMEBOOST_cell_1062 ( .a(FE_RN_1982_0), .b(TIMEBOOST_net_145), .o(FE_RN_1715_0) );
na02f10 g775000 ( .a(n_5965), .b(n_5924), .o(n_6102) );
in01s02 g775001 ( .a(n_6153), .o(n_6220) );
no02m06 g775002 ( .a(FE_OCP_RBN3216_n_5003), .b(n_6132), .o(n_6153) );
na02s02 g775003 ( .a(n_6108), .b(FE_OCP_RBN3209_n_5221), .o(n_6234) );
in01s01 g775005 ( .a(n_6148), .o(n_6173) );
na02s06 g775006 ( .a(n_6132), .b(FE_OCP_RBN3216_n_5003), .o(n_6148) );
na02s03 g775007 ( .a(n_6109), .b(n_5265), .o(n_6186) );
no02s01 TIMEBOOST_cell_1341 ( .a(n_41574), .b(n_41440), .o(TIMEBOOST_net_285) );
na02s02 g775009 ( .a(n_6113), .b(n_5898), .o(n_6143) );
no02s01 TIMEBOOST_cell_1331 ( .a(n_28877), .b(n_28902), .o(TIMEBOOST_net_280) );
na02s02 g775011 ( .a(n_6098), .b(n_5844), .o(n_6133) );
in01s02 g775012 ( .a(n_6162), .o(n_6163) );
no02f04 g775013 ( .a(n_6147), .b(n_6044), .o(n_6162) );
in01s01 g775014 ( .a(n_6179), .o(n_6180) );
na02s02 g775015 ( .a(n_6147), .b(n_6001), .o(n_6179) );
in01s01 g775016 ( .a(n_6184), .o(n_6185) );
in01s01 g775017 ( .a(n_6160), .o(n_6184) );
oa12f06 g775018 ( .a(n_5287), .b(n_6076), .c(n_5186), .o(n_6160) );
oa22s01 g775019 ( .a(n_6097), .b(n_5342), .c(n_6096), .d(n_5343), .o(n_6183) );
in01s01 g775020 ( .a(n_6154), .o(n_6124) );
no02m04 TIMEBOOST_cell_1328 ( .a(TIMEBOOST_net_278), .b(n_19639), .o(n_19784) );
oa12m04 g775022 ( .a(n_6188), .b(n_6128), .c(n_6106), .o(n_6201) );
in01s02 g775023 ( .a(n_6248), .o(n_6206) );
no02f04 TIMEBOOST_cell_6646 ( .a(TIMEBOOST_net_2080), .b(n_13558), .o(n_13689) );
in01s02 g775027 ( .a(n_6118), .o(n_6125) );
in01m02 g775028 ( .a(n_6083), .o(n_6118) );
oa12f04 g775029 ( .a(n_5919), .b(n_6019), .c(n_5887), .o(n_6083) );
in01s01 g775031 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_24_), .o(n_6142) );
na02m08 TIMEBOOST_cell_1061 ( .a(n_32878), .b(FE_RN_2167_0), .o(TIMEBOOST_net_145) );
no02s06 g775035 ( .a(n_5977), .b(n_4675), .o(n_6089) );
na02m08 g775036 ( .a(n_5893), .b(n_4875), .o(n_5965) );
in01m06 g775037 ( .a(n_5923), .o(n_5924) );
no02m08 g775038 ( .a(n_5893), .b(n_4675), .o(n_5923) );
in01s04 g775039 ( .a(FE_OCP_RBN3357_n_6013), .o(n_6028) );
no02m08 g775041 ( .a(n_5976), .b(n_4759), .o(n_6013) );
na02s02 g775042 ( .a(n_6009), .b(n_5726), .o(n_6048) );
no02m02 TIMEBOOST_cell_1327 ( .a(n_19561), .b(FE_OCPN1727_n_18099), .o(TIMEBOOST_net_278) );
na02m04 g775044 ( .a(n_6086), .b(n_6012), .o(n_6114) );
in01s01 g775045 ( .a(n_6169), .o(n_6170) );
na02s01 g775046 ( .a(n_6157), .b(n_6086), .o(n_6169) );
na02f06 g775047 ( .a(n_5930), .b(n_6077), .o(n_6147) );
in01s01 g775049 ( .a(n_6082), .o(n_6098) );
no02s06 g775050 ( .a(n_6020), .b(n_5740), .o(n_6082) );
in01s01 g775051 ( .a(n_6171), .o(n_6172) );
na02s01 g775052 ( .a(n_6107), .b(n_6188), .o(n_6171) );
na02s02 g775053 ( .a(n_6092), .b(n_5967), .o(n_6136) );
no02m04 TIMEBOOST_cell_1389 ( .a(n_18982), .b(n_18547), .o(TIMEBOOST_net_309) );
na02m08 g775055 ( .a(n_5979), .b(n_6038), .o(n_6090) );
in01m02 g775056 ( .a(n_6054), .o(n_6055) );
ao12s04 g775057 ( .a(n_5969), .b(n_6038), .c(n_5963), .o(n_6054) );
in01s04 g775058 ( .a(n_6064), .o(n_6065) );
in01m04 g775059 ( .a(n_6041), .o(n_6064) );
oa12f06 g775060 ( .a(n_5878), .b(n_5970), .c(n_5871), .o(n_6041) );
no02m06 TIMEBOOST_cell_986 ( .a(n_28298), .b(TIMEBOOST_net_107), .o(n_28328) );
no02f04 TIMEBOOST_cell_1344 ( .a(TIMEBOOST_net_286), .b(n_19859), .o(n_19884) );
in01s02 g775063 ( .a(n_6146), .o(n_6137) );
no02s01 TIMEBOOST_cell_1282 ( .a(TIMEBOOST_net_255), .b(n_7510), .o(n_7624) );
in01s01 g775065 ( .a(n_46995), .o(n_6175) );
ao12m04 g775067 ( .a(n_6080), .b(n_6039), .c(n_6012), .o(n_6081) );
in01s02 g775068 ( .a(n_6108), .o(n_6109) );
in01s01 g775070 ( .a(n_6112), .o(n_6113) );
oa12s01 g775071 ( .a(n_47270), .b(n_6036), .c(FE_OCP_RBN4441_n_5891), .o(n_6112) );
in01s01 g775072 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_15_), .o(n_7211) );
in01s01 g775074 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_16_), .o(n_6123) );
na02s02 TIMEBOOST_cell_6885 ( .a(FE_RN_348_0), .b(n_17973), .o(TIMEBOOST_net_2201) );
no02s02 TIMEBOOST_cell_985 ( .a(n_27929), .b(n_28280), .o(TIMEBOOST_net_107) );
na02m06 g775079 ( .a(n_5962), .b(n_5968), .o(n_5979) );
no02m04 g775080 ( .a(n_5948), .b(n_5986), .o(n_6037) );
no02m02 TIMEBOOST_cell_1343 ( .a(n_18140), .b(FE_OCP_RBN2746_n_19747), .o(TIMEBOOST_net_286) );
in01s02 g775082 ( .a(n_6019), .o(n_6020) );
na02s06 g775083 ( .a(n_5987), .b(n_5710), .o(n_6019) );
in01s01 g775084 ( .a(n_6106), .o(n_6107) );
no02s04 g775085 ( .a(n_6074), .b(n_5049), .o(n_6106) );
na02m06 g775086 ( .a(FE_OCP_RBN3380_n_6034), .b(n_4904), .o(n_6157) );
in01s04 g775088 ( .a(n_6086), .o(n_6094) );
na02f06 g775089 ( .a(n_6034), .b(FE_OCP_RBN3144_n_4858), .o(n_6086) );
in01s01 g775090 ( .a(n_6009), .o(n_6010) );
no02s01 g775091 ( .a(n_5987), .b(n_5709), .o(n_6009) );
na02s02 g775093 ( .a(n_6012), .b(n_6006), .o(n_6119) );
na02s04 g775094 ( .a(n_6026), .b(n_5792), .o(n_6053) );
na02s02 g775096 ( .a(n_6036), .b(n_5889), .o(n_6121) );
na03m04 TIMEBOOST_cell_6483 ( .a(FE_OCP_RBN5838_n_44563), .b(n_8990), .c(n_9053), .o(n_9234) );
na02m04 g775098 ( .a(n_6074), .b(n_5049), .o(n_6188) );
in01s01 g775099 ( .a(n_6096), .o(n_6097) );
in01s01 g775100 ( .a(n_6076), .o(n_6096) );
oa12f04 g775101 ( .a(n_5247), .b(n_6062), .c(n_5111), .o(n_6076) );
ao12f02 g775103 ( .a(n_5926), .b(n_5955), .c(n_5815), .o(n_6021) );
in01m03 g775104 ( .a(n_6067), .o(n_6068) );
oa12f04 g775105 ( .a(n_5788), .b(n_5996), .c(n_5769), .o(n_6067) );
oa12f04 g775106 ( .a(n_6066), .b(n_6127), .c(n_6069), .o(n_6128) );
in01s01 g775108 ( .a(n_6077), .o(n_6092) );
in01s02 g775110 ( .a(n_6063), .o(n_6043) );
oa22s02 g775111 ( .a(n_5941), .b(n_5599), .c(n_5927), .d(n_5598), .o(n_6063) );
in01s02 g775112 ( .a(n_5976), .o(n_5977) );
in01m04 g775113 ( .a(n_5946), .o(n_5976) );
no02s01 TIMEBOOST_cell_1058 ( .a(n_33073), .b(TIMEBOOST_net_143), .o(n_33193) );
no02s10 TIMEBOOST_cell_1004 ( .a(n_12333), .b(TIMEBOOST_net_116), .o(n_12361) );
oa22s01 g775116 ( .a(n_6024), .b(n_5258), .c(n_6062), .d(n_5259), .o(n_6085) );
in01s01 g775117 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_21_), .o(n_6061) );
no02m06 g775120 ( .a(n_5964), .b(n_5925), .o(n_6038) );
in01m03 g775121 ( .a(n_5968), .o(n_5969) );
no02m10 TIMEBOOST_cell_1178 ( .a(FE_OCP_RBN2509_n_41215), .b(TIMEBOOST_net_203), .o(n_41294) );
na02m06 g775123 ( .a(n_5870), .b(n_5766), .o(n_5871) );
no02f06 g775124 ( .a(n_5839), .b(n_5769), .o(n_5878) );
in01s02 g775125 ( .a(n_5947), .o(n_5948) );
no02s04 g775126 ( .a(n_5926), .b(n_5925), .o(n_5947) );
na02s04 TIMEBOOST_cell_4518 ( .a(TIMEBOOST_net_1349), .b(n_10952), .o(n_11061) );
no02s01 TIMEBOOST_cell_1057 ( .a(n_32608), .b(n_33146), .o(TIMEBOOST_net_143) );
no02f04 TIMEBOOST_cell_8820 ( .a(n_15423), .b(n_15469), .o(TIMEBOOST_net_2897) );
no02s06 TIMEBOOST_cell_4509 ( .a(FE_OCPN1705_n_14730), .b(n_16333), .o(TIMEBOOST_net_1345) );
in01s02 g775131 ( .a(n_5997), .o(n_5998) );
no02s04 g775132 ( .a(n_5943), .b(n_5964), .o(n_5997) );
na02s02 g775133 ( .a(n_5870), .b(n_5868), .o(n_5904) );
no02s02 g775134 ( .a(n_5839), .b(FE_OCP_RBN4451_n_5870), .o(n_5921) );
na02s02 g775135 ( .a(n_5788), .b(n_5801), .o(n_5910) );
no02s02 g775136 ( .a(n_5787), .b(n_5769), .o(n_5907) );
in01m01 g775137 ( .a(n_6080), .o(n_6006) );
no02s03 g775138 ( .a(n_5989), .b(FE_OCP_RBN3121_n_4751), .o(n_6080) );
no02s06 g775139 ( .a(n_5927), .b(n_5577), .o(n_5987) );
in01s01 g775140 ( .a(n_6140), .o(n_6141) );
na02s01 g775141 ( .a(n_6187), .b(n_6066), .o(n_6140) );
no02s04 g775144 ( .a(n_6015), .b(FE_OCP_RBN4444_n_5849), .o(n_6036) );
na02s06 g775148 ( .a(n_5989), .b(FE_OCP_RBN3121_n_4751), .o(n_6012) );
in01s01 g775149 ( .a(n_6051), .o(n_6052) );
no02m04 TIMEBOOST_cell_3178 ( .a(n_25676), .b(n_25379), .o(TIMEBOOST_net_880) );
ao22f04 g775152 ( .a(n_5939), .b(n_5918), .c(n_5938), .d(n_5917), .o(n_6034) );
in01m02 g775153 ( .a(n_6105), .o(n_6071) );
no02s01 TIMEBOOST_cell_1280 ( .a(TIMEBOOST_net_254), .b(FE_RN_1667_0), .o(n_23859) );
oa22f04 g775155 ( .a(FE_OCP_RBN6149_n_5974), .b(n_5782), .c(n_5974), .d(n_5779), .o(n_6074) );
in01s02 g775156 ( .a(n_6039), .o(n_6040) );
ao12f04 g775157 ( .a(n_46427), .b(n_6008), .c(n_6007), .o(n_6039) );
in01s01 g775158 ( .a(n_6047), .o(n_6005) );
no02m04 TIMEBOOST_cell_1314 ( .a(TIMEBOOST_net_271), .b(n_13726), .o(n_13728) );
oa12s01 g775160 ( .a(n_5991), .b(n_5994), .c(n_5990), .o(n_6042) );
in01s02 g775161 ( .a(n_6025), .o(n_6026) );
oa12s02 g775162 ( .a(n_5727), .b(n_5959), .c(n_5657), .o(n_6025) );
no02m03 TIMEBOOST_cell_3177 ( .a(TIMEBOOST_net_879), .b(n_4161), .o(n_4376) );
na02s01 g775166 ( .a(n_5994), .b(n_5990), .o(n_5991) );
no02s06 TIMEBOOST_cell_1177 ( .a(n_41229), .b(n_40932), .o(TIMEBOOST_net_203) );
no02s04 g775168 ( .a(n_5818), .b(n_4759), .o(n_5926) );
no02m04 g775169 ( .a(n_5881), .b(FE_OCPN3584_n_4556), .o(n_5943) );
in01s01 g775173 ( .a(n_5769), .o(n_5801) );
no02s06 g775174 ( .a(n_5750), .b(n_4875), .o(n_5769) );
na02f06 g775176 ( .a(n_5802), .b(n_4875), .o(n_5870) );
no02m08 g775177 ( .a(n_5800), .b(FE_OCP_RBN2962_n_4046), .o(n_5925) );
na02s02 g775178 ( .a(n_5818), .b(FE_OCPN3584_n_4556), .o(n_5815) );
no02s06 g775179 ( .a(n_5882), .b(FE_OCP_RBN2962_n_4046), .o(n_5964) );
in01s01 g775181 ( .a(n_5839), .o(n_5868) );
no02m06 g775182 ( .a(n_5802), .b(n_4875), .o(n_5839) );
in01s03 g775183 ( .a(n_5787), .o(n_5788) );
in01m02 g775186 ( .a(n_5766), .o(n_5787) );
na02m04 g775187 ( .a(n_5750), .b(n_4675), .o(n_5766) );
in01s01 g775189 ( .a(n_6066), .o(n_6087) );
na02s06 g775190 ( .a(n_46996), .b(FE_OCP_RBN3155_n_4925), .o(n_6066) );
na02s02 g775191 ( .a(n_5958), .b(n_5689), .o(n_6023) );
in01s03 g775192 ( .a(n_6069), .o(n_6187) );
no02f06 g775193 ( .a(n_46996), .b(FE_OCP_RBN3155_n_4925), .o(n_6069) );
no02s01 TIMEBOOST_cell_1279 ( .a(FE_RN_1666_0), .b(n_23542), .o(TIMEBOOST_net_254) );
in01s01 g775196 ( .a(n_5927), .o(n_5941) );
oa12m06 g775197 ( .a(n_5589), .b(n_5811), .c(n_5566), .o(n_5927) );
in01s01 g775198 ( .a(n_6032), .o(n_6033) );
na02s02 g775199 ( .a(n_6008), .b(n_5961), .o(n_6032) );
no02s02 TIMEBOOST_cell_1313 ( .a(n_13661), .b(FE_OCP_RBN2540_n_12880), .o(TIMEBOOST_net_271) );
na02s01 g775201 ( .a(n_5896), .b(n_5620), .o(n_5953) );
no02s04 g775202 ( .a(n_46427), .b(n_5982), .o(n_5983) );
in01f04 g775204 ( .a(n_5962), .o(n_5963) );
in01m02 g775205 ( .a(n_5963), .o(n_5986) );
in01f04 g775207 ( .a(n_5955), .o(n_5962) );
na02m06 TIMEBOOST_cell_6659 ( .a(n_19339), .b(n_19406), .o(TIMEBOOST_net_2087) );
in01s01 g775209 ( .a(n_6062), .o(n_6024) );
no02s01 TIMEBOOST_cell_4872 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .o(TIMEBOOST_net_1384) );
oa12s01 g775211 ( .a(n_5951), .b(n_5950), .c(n_5949), .o(n_5992) );
in01s01 g775212 ( .a(FE_OCP_RBN3326_n_5813), .o(n_5852) );
oa22m04 g775215 ( .a(n_5674), .b(n_5556), .c(n_5675), .d(n_5557), .o(n_5813) );
in01f02 g775217 ( .a(n_5693), .o(n_5732) );
no02s06 g775220 ( .a(n_5959), .b(n_5784), .o(n_6015) );
in01s02 g775221 ( .a(n_46997), .o(n_6004) );
in01s02 g775224 ( .a(n_5996), .o(n_6017) );
in01s04 g775225 ( .a(n_5970), .o(n_5996) );
no02f06 g775226 ( .a(n_5905), .b(n_5707), .o(n_5970) );
na02f04 g775228 ( .a(n_6011), .b(n_6003), .o(n_6127) );
in01s01 g775230 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_14_), .o(n_5999) );
in01s01 g775232 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_19_), .o(n_5984) );
na02s01 g775234 ( .a(n_5944), .b(n_4973), .o(n_5994) );
na02s02 g775235 ( .a(n_5691), .b(n_5667), .o(n_5782) );
no02s04 g775236 ( .a(n_5692), .b(n_5714), .o(n_5779) );
na02s01 g775237 ( .a(n_5950), .b(n_5949), .o(n_5951) );
in01s02 g775238 ( .a(n_5917), .o(n_5918) );
na02m02 g775239 ( .a(n_5857), .b(n_5837), .o(n_5917) );
na02f04 g775240 ( .a(n_5952), .b(n_5940), .o(n_6008) );
na02m01 g775241 ( .a(n_5902), .b(n_5761), .o(n_5928) );
in01s02 g775243 ( .a(n_5957), .o(n_5958) );
in01s02 g775244 ( .a(n_5959), .o(n_5957) );
na02s06 g775245 ( .a(n_5883), .b(n_5736), .o(n_5959) );
na02m04 g775246 ( .a(n_6002), .b(n_6001), .o(n_6003) );
in01s01 g775247 ( .a(n_6116), .o(n_6117) );
na02s01 g775248 ( .a(n_6011), .b(n_6002), .o(n_6116) );
in01s01 g775249 ( .a(n_46427), .o(n_5961) );
in01m04 g775252 ( .a(n_5938), .o(n_5939) );
no02m06 g775253 ( .a(n_5867), .b(FE_OCP_RBN6854_n_5735), .o(n_5938) );
no02m04 TIMEBOOST_cell_3966 ( .a(TIMEBOOST_net_1073), .b(n_8275), .o(FE_RN_975_0) );
no02f04 TIMEBOOST_cell_6638 ( .a(TIMEBOOST_net_2076), .b(FE_RN_961_0), .o(n_23315) );
na02m04 g775256 ( .a(n_5857), .b(n_5778), .o(n_5858) );
na02m04 g775257 ( .a(n_5667), .b(n_5655), .o(n_5707) );
in01s01 g775259 ( .a(n_5895), .o(n_5896) );
no02s04 TIMEBOOST_cell_6020 ( .a(n_33411), .b(TIMEBOOST_net_1861), .o(n_33504) );
no02s02 TIMEBOOST_cell_3284 ( .a(n_26716), .b(n_26454), .o(TIMEBOOST_net_933) );
in01s02 g775262 ( .a(n_5972), .o(n_5937) );
na02m06 TIMEBOOST_cell_1308 ( .a(TIMEBOOST_net_268), .b(FE_RN_2419_0), .o(n_13726) );
in01s04 g775264 ( .a(n_5881), .o(n_5882) );
na02m06 TIMEBOOST_cell_7611 ( .a(TIMEBOOST_net_2436), .b(n_9140), .o(n_9342) );
in01s04 g775267 ( .a(n_5818), .o(n_5800) );
na02s01 TIMEBOOST_cell_5498 ( .a(n_22288), .b(FE_OCP_RBN1869_n_21358), .o(TIMEBOOST_net_1697) );
na02s01 TIMEBOOST_cell_3268 ( .a(n_31287), .b(n_31351), .o(TIMEBOOST_net_925) );
in01s01 g775271 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_13_), .o(n_7135) );
na02s01 TIMEBOOST_cell_1123 ( .a(n_33276), .b(n_33274), .o(TIMEBOOST_net_176) );
no02m04 g775277 ( .a(n_5816), .b(n_5808), .o(n_5867) );
no02m04 g775278 ( .a(n_5808), .b(n_5743), .o(n_5778) );
no02s01 TIMEBOOST_cell_6588 ( .a(TIMEBOOST_net_2051), .b(n_28080), .o(n_28177) );
na02m02 g775280 ( .a(n_5751), .b(n_5735), .o(n_5773) );
in01m01 g775281 ( .a(n_5836), .o(n_5837) );
no02m04 g775282 ( .a(n_5810), .b(n_4759), .o(n_5836) );
no02m06 TIMEBOOST_cell_5497 ( .a(TIMEBOOST_net_1696), .b(n_10585), .o(n_10707) );
no02s06 TIMEBOOST_cell_6593 ( .a(n_17133), .b(n_17084), .o(TIMEBOOST_net_2054) );
na02m06 TIMEBOOST_cell_3267 ( .a(TIMEBOOST_net_924), .b(n_30468), .o(n_30582) );
na02f04 TIMEBOOST_cell_5625 ( .a(TIMEBOOST_net_1760), .b(n_26620), .o(n_26797) );
na02f02 g775287 ( .a(n_5656), .b(n_4875), .o(n_5669) );
no02f04 TIMEBOOST_cell_7657 ( .a(TIMEBOOST_net_2459), .b(n_13552), .o(n_13597) );
in01s01 g775290 ( .a(n_5667), .o(n_5714) );
na02s04 g775291 ( .a(n_5644), .b(FE_OCPN3584_n_4556), .o(n_5667) );
no02m08 TIMEBOOST_cell_6302 ( .a(TIMEBOOST_net_2002), .b(n_35746), .o(TIMEBOOST_net_561) );
na02m04 g775293 ( .a(n_5810), .b(n_4759), .o(n_5857) );
na02f06 g775294 ( .a(n_5894), .b(n_5005), .o(n_5944) );
in01s02 g775295 ( .a(n_5832), .o(n_5833) );
no02s04 g775296 ( .a(FE_OCP_RBN6855_n_5735), .b(n_5808), .o(n_5832) );
no02s01 g775297 ( .a(n_5894), .b(n_4864), .o(n_5950) );
in01s01 g775298 ( .a(n_5691), .o(n_5692) );
in01s02 g775299 ( .a(n_5672), .o(n_5691) );
no02f04 g775300 ( .a(n_5644), .b(FE_OCPN3584_n_4556), .o(n_5672) );
na02s02 g775301 ( .a(n_5806), .b(n_5607), .o(n_5866) );
no02s03 g775302 ( .a(n_5798), .b(n_5516), .o(n_5811) );
oa12f02 g775303 ( .a(n_5886), .b(n_5825), .c(n_5763), .o(n_5919) );
in01s01 g775304 ( .a(n_5980), .o(n_5981) );
na02s02 g775305 ( .a(n_6007), .b(n_5916), .o(n_5980) );
in01m02 g775306 ( .a(n_5561), .o(n_5562) );
oa12f04 g775307 ( .a(n_5423), .b(n_5446), .c(FE_OCP_RBN4374_n_5048), .o(n_5561) );
no02s01 g775308 ( .a(n_5636), .b(FE_OCP_RBN6114_n_5444), .o(n_5637) );
na02s02 g775309 ( .a(n_46998), .b(FE_OCP_RBN3122_n_4784), .o(n_6002) );
na02s01 g775310 ( .a(FE_OCP_RBN3286_n_5656), .b(n_5614), .o(n_5706) );
na03s08 TIMEBOOST_cell_4576 ( .a(n_1426), .b(delay_xor_ln22_unr3_stage2_stallmux_q_1_), .c(FE_OCP_RBN6409_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1491) );
na02s02 TIMEBOOST_cell_1307 ( .a(FE_OCP_RBN1016_n_13601), .b(FE_RN_462_0), .o(TIMEBOOST_net_268) );
in01s01 g775314 ( .a(n_6011), .o(n_6044) );
na02m03 g775315 ( .a(n_5933), .b(n_4784), .o(n_6011) );
in01s02 g775316 ( .a(n_5674), .o(n_5675) );
oa12f04 g775317 ( .a(n_5530), .b(n_5554), .c(n_5365), .o(n_5674) );
na02s04 g775319 ( .a(n_5901), .b(n_5558), .o(n_5974) );
na02f06 g775320 ( .a(n_5830), .b(n_5835), .o(n_5952) );
oa12s01 g775321 ( .a(n_5864), .b(n_5863), .c(n_5862), .o(n_5922) );
in01s02 g775322 ( .a(n_5971), .o(n_5935) );
no02f08 TIMEBOOST_cell_1318 ( .a(n_41818), .b(TIMEBOOST_net_273), .o(n_41757) );
oa12s01 g775324 ( .a(n_5861), .b(n_5860), .c(n_5859), .o(n_5915) );
oa12s04 g775325 ( .a(n_5701), .b(n_5876), .c(n_5877), .o(n_5883) );
ao12s02 g775327 ( .a(n_5877), .b(n_5876), .c(n_5582), .o(n_5902) );
na02m02 g775328 ( .a(n_5888), .b(FE_OCP_RBN3322_n_5586), .o(n_5901) );
na02f06 g775331 ( .a(FE_OCP_RBN6869_n_5751), .b(FE_OCP_RBN6866_n_5743), .o(n_5816) );
no02m02 g775332 ( .a(n_5586), .b(n_5654), .o(n_5655) );
na02s01 g775333 ( .a(n_5863), .b(n_5862), .o(n_5864) );
na02m02 g775335 ( .a(n_5558), .b(FE_OCP_RBN3322_n_5586), .o(n_5677) );
no02s04 g775336 ( .a(n_5700), .b(n_4875), .o(n_5808) );
na02m04 g775338 ( .a(n_5700), .b(n_4875), .o(n_5735) );
no02f06 g775339 ( .a(n_5814), .b(n_5000), .o(n_5894) );
in01s01 g775340 ( .a(n_5966), .o(n_5967) );
na02s02 g775341 ( .a(n_6001), .b(n_5930), .o(n_5966) );
na02s04 g775342 ( .a(n_5909), .b(FE_OCPN1094_n_4459), .o(n_6007) );
in01s02 g775343 ( .a(n_5982), .o(n_5916) );
no02s04 g775344 ( .a(n_5909), .b(FE_OCPN1094_n_4459), .o(n_5982) );
na02m04 g775345 ( .a(n_5785), .b(n_5768), .o(n_5835) );
na02s01 g775346 ( .a(n_5860), .b(n_5859), .o(n_5861) );
no02f06 TIMEBOOST_cell_1317 ( .a(n_41460), .b(n_41683), .o(TIMEBOOST_net_273) );
na02f03 g775348 ( .a(n_5786), .b(n_5767), .o(n_5830) );
na02s01 g775349 ( .a(n_5807), .b(n_5660), .o(n_5880) );
oa12s01 g775351 ( .a(n_5776), .b(n_5775), .c(n_5774), .o(n_5853) );
in01s01 g775354 ( .a(FE_OCP_RBN3319_n_5555), .o(n_5636) );
in01s01 g775359 ( .a(n_5609), .o(n_5648) );
in01s02 g775360 ( .a(n_5609), .o(n_5610) );
na02f06 g775361 ( .a(n_5528), .b(n_5480), .o(n_5609) );
in01s01 g775362 ( .a(n_5840), .o(n_5789) );
oa22m01 g775363 ( .a(n_5721), .b(n_5463), .c(n_5673), .d(n_5464), .o(n_5840) );
no02s06 TIMEBOOST_cell_3222 ( .a(n_25272), .b(n_25359), .o(TIMEBOOST_net_902) );
oa12s01 g775365 ( .a(n_5875), .b(n_5874), .c(n_5873), .o(n_5929) );
in01s01 g775366 ( .a(n_5805), .o(n_5806) );
in01s01 g775367 ( .a(n_5798), .o(n_5805) );
oa12m04 g775368 ( .a(n_5431), .b(n_5721), .c(n_5372), .o(n_5798) );
in01s01 g775370 ( .a(FE_OCP_RBN3286_n_5656), .o(n_5703) );
in01s01 g775375 ( .a(n_5754), .o(n_5780) );
in01s01 g775376 ( .a(n_5717), .o(n_5754) );
in01s02 g775377 ( .a(n_5717), .o(n_5718) );
na02s01 TIMEBOOST_cell_1042 ( .a(TIMEBOOST_net_135), .b(n_37380), .o(n_37376) );
in01s02 g775379 ( .a(n_5913), .o(n_5906) );
oa22s02 g775380 ( .a(n_5757), .b(n_5563), .c(n_5756), .d(n_5564), .o(n_5913) );
in01s02 g775381 ( .a(n_46998), .o(n_5933) );
na02s02 TIMEBOOST_cell_6602 ( .a(TIMEBOOST_net_2058), .b(n_45145), .o(n_40701) );
in01s01 g775384 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_12_), .o(n_5884) );
in01s01 g775388 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_12_), .o(n_5777) );
na02m04 g775390 ( .a(n_5437), .b(n_5056), .o(n_5528) );
na02s03 g775391 ( .a(n_5436), .b(n_5057), .o(n_5480) );
no02f02 g775392 ( .a(n_5417), .b(n_5422), .o(n_5446) );
no02m04 g775393 ( .a(n_5526), .b(n_5529), .o(n_5554) );
na02s01 g775394 ( .a(n_5874), .b(n_5873), .o(n_5875) );
in01s02 g775396 ( .a(n_5888), .o(n_5911) );
no02f04 g775397 ( .a(n_5796), .b(n_5654), .o(n_5888) );
na02s01 g775398 ( .a(n_5775), .b(n_5774), .o(n_5776) );
no02f02 g775399 ( .a(n_5793), .b(n_5587), .o(n_5838) );
na02m06 g775401 ( .a(n_5712), .b(n_5572), .o(n_5743) );
no02f02 g775404 ( .a(n_5543), .b(FE_OCP_RBN2969_n_4046), .o(n_5586) );
in01s02 g775405 ( .a(n_5767), .o(n_5768) );
na02s04 g775406 ( .a(n_5680), .b(n_5712), .o(n_5767) );
no03s02 TIMEBOOST_cell_7664 ( .a(n_2537), .b(n_3023), .c(n_2473), .o(TIMEBOOST_net_2463) );
no02s04 g775409 ( .a(n_5684), .b(n_5679), .o(n_5751) );
no02s01 TIMEBOOST_cell_4524 ( .a(TIMEBOOST_net_1352), .b(n_17137), .o(n_17386) );
na02f03 g775411 ( .a(n_5444), .b(n_5494), .o(n_5495) );
in01s02 g775413 ( .a(n_5558), .o(n_5601) );
na02m03 g775414 ( .a(n_5543), .b(FE_OCP_RBN2969_n_4046), .o(n_5558) );
no02s01 TIMEBOOST_cell_6305 ( .a(n_43003), .b(n_43002), .o(TIMEBOOST_net_2004) );
na02s01 TIMEBOOST_cell_1041 ( .a(n_37375), .b(n_36962), .o(TIMEBOOST_net_135) );
na02s04 g775417 ( .a(n_5821), .b(n_47008), .o(n_5930) );
no02m04 g775418 ( .a(n_5541), .b(n_5499), .o(n_5605) );
na02f02 g775419 ( .a(n_5824), .b(n_5823), .o(n_5825) );
in01s01 g775420 ( .a(n_5876), .o(n_5807) );
na02f06 g775421 ( .a(n_5690), .b(n_5547), .o(n_5876) );
in01s01 g775422 ( .a(n_5899), .o(n_5900) );
na02s01 g775423 ( .a(n_5824), .b(n_5886), .o(n_5899) );
na02s02 g775424 ( .a(n_5886), .b(n_5702), .o(n_5887) );
na02s03 g775425 ( .a(n_5820), .b(n_4700), .o(n_6001) );
oa12s01 g775426 ( .a(n_4820), .b(n_5741), .c(n_4901), .o(n_5860) );
in01s01 g775427 ( .a(n_5814), .o(n_5863) );
ao12f06 g775428 ( .a(n_4871), .b(n_5711), .c(n_4885), .o(n_5814) );
na02f04 g775429 ( .a(n_5730), .b(n_5771), .o(n_5909) );
no02s01 TIMEBOOST_cell_3212 ( .a(n_5091), .b(n_4972), .o(TIMEBOOST_net_897) );
in01m02 g775432 ( .a(n_5436), .o(n_5437) );
in01m02 g775433 ( .a(n_5417), .o(n_5436) );
na02m02 g775434 ( .a(n_5348), .b(n_5127), .o(n_5417) );
na02s02 g775435 ( .a(n_5349), .b(n_5422), .o(n_5423) );
na02s02 g775436 ( .a(n_5434), .b(n_5529), .o(n_5530) );
no02s01 g775437 ( .a(n_5742), .b(n_4819), .o(n_5874) );
in01s02 g775438 ( .a(n_5796), .o(n_5797) );
no02m08 g775439 ( .a(n_5770), .b(n_47197), .o(n_5796) );
na02s04 g775440 ( .a(n_5568), .b(n_5581), .o(n_5654) );
no02m08 TIMEBOOST_cell_4526 ( .a(TIMEBOOST_net_1353), .b(n_25967), .o(n_26112) );
in01m02 g775442 ( .a(n_5785), .o(n_5786) );
no02s04 g775443 ( .a(n_5685), .b(n_5596), .o(n_5785) );
na02m04 g775444 ( .a(n_5651), .b(FE_OCPN1663_n_4556), .o(n_5712) );
in01s02 g775445 ( .a(n_5679), .o(n_5680) );
no02s04 g775446 ( .a(n_5651), .b(FE_OCPN1663_n_4556), .o(n_5679) );
na02s03 g775448 ( .a(n_5524), .b(n_5568), .o(n_5587) );
no02s02 TIMEBOOST_cell_4425 ( .a(n_47015), .b(FE_OCP_RBN6771_n_3700), .o(TIMEBOOST_net_1303) );
na02s02 g775450 ( .a(n_5642), .b(n_5719), .o(n_5730) );
in01m02 g775451 ( .a(n_5540), .o(n_5541) );
in01s02 g775452 ( .a(n_5526), .o(n_5540) );
na02m04 g775453 ( .a(n_5433), .b(n_5336), .o(n_5526) );
na02s04 g775456 ( .a(n_5723), .b(n_4376), .o(n_5886) );
na02m02 g775457 ( .a(n_46999), .b(FE_OCP_RBN3050_n_4376), .o(n_5824) );
na02s04 g775458 ( .a(n_5641), .b(n_5720), .o(n_5771) );
in01s02 g775459 ( .a(n_5428), .o(n_5429) );
ao12m04 g775460 ( .a(n_4998), .b(n_45323), .c(n_5061), .o(n_5428) );
in01s01 g775461 ( .a(n_5897), .o(n_5898) );
na02s01 g775462 ( .a(n_5879), .b(n_5842), .o(n_5897) );
oa12s01 g775463 ( .a(n_4746), .b(n_5716), .c(n_4921), .o(n_5775) );
oa12s02 g775464 ( .a(n_5382), .b(n_5486), .c(n_5440), .o(n_5487) );
no02m02 g775465 ( .a(n_5441), .b(n_5340), .o(n_5503) );
oa12s01 g775466 ( .a(n_5666), .b(n_5716), .c(n_5665), .o(n_5753) );
in01s02 g775467 ( .a(n_5820), .o(n_5821) );
in01s01 g775470 ( .a(FE_OCP_RBN6115_n_5444), .o(n_5523) );
in01s02 g775473 ( .a(n_5756), .o(n_5757) );
oa12s02 g775474 ( .a(n_5475), .b(n_5755), .c(n_5534), .o(n_5756) );
in01s01 g775475 ( .a(n_5724), .o(n_5708) );
oa12s01 g775476 ( .a(n_5617), .b(n_5624), .c(n_5616), .o(n_5724) );
na02m06 g775481 ( .a(n_5505), .b(n_5496), .o(n_5614) );
in01s02 g775482 ( .a(n_5841), .o(n_5795) );
oa12s02 g775483 ( .a(n_5698), .b(n_5755), .c(n_5697), .o(n_5841) );
oa12f04 g775485 ( .a(n_5535), .b(n_5622), .c(n_5412), .o(n_5690) );
in01s01 g775486 ( .a(n_5721), .o(n_5673) );
oa12f04 g775487 ( .a(n_5274), .b(n_5624), .c(n_5353), .o(n_5721) );
in01s01 g775488 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_11_), .o(n_5671) );
na02m02 g775492 ( .a(n_5770), .b(n_5581), .o(n_5793) );
in01s02 g775493 ( .a(n_5684), .o(n_5685) );
na02f04 g775494 ( .a(n_5608), .b(n_5650), .o(n_5684) );
in01s02 g775495 ( .a(n_5719), .o(n_5720) );
na02m02 g775496 ( .a(n_5650), .b(n_5572), .o(n_5719) );
na02f04 g775497 ( .a(n_5457), .b(FE_OCPN1663_n_4556), .o(n_5568) );
na02s01 g775498 ( .a(n_5716), .b(n_5665), .o(n_5666) );
na02s04 g775500 ( .a(n_5456), .b(n_4316), .o(n_5524) );
na02s02 g775501 ( .a(n_5486), .b(n_5442), .o(n_5496) );
in01s02 g775502 ( .a(n_5812), .o(n_5879) );
no02s03 g775503 ( .a(n_5759), .b(FE_OCP_RBN3087_n_4458), .o(n_5812) );
in01s01 g775504 ( .a(n_5844), .o(n_5845) );
na02s02 g775505 ( .a(n_5823), .b(n_5702), .o(n_5844) );
no02m02 g775506 ( .a(n_5486), .b(n_5440), .o(n_5441) );
in01s02 g775507 ( .a(n_5433), .o(n_5434) );
na02m04 g775508 ( .a(n_5375), .b(n_5301), .o(n_5433) );
na02s01 g775509 ( .a(n_5755), .b(n_5697), .o(n_5698) );
no02s02 g775510 ( .a(n_5739), .b(n_5681), .o(n_5763) );
na02m01 g775511 ( .a(n_5624), .b(n_5616), .o(n_5617) );
na02s04 g775512 ( .a(FE_OCP_RBN6081_n_5486), .b(n_5443), .o(n_5505) );
na02s02 g775513 ( .a(n_5759), .b(FE_OCP_RBN3087_n_4458), .o(n_5842) );
in01s01 g775515 ( .a(n_5348), .o(n_5349) );
in01s01 g775517 ( .a(n_5741), .o(n_5742) );
in01s01 g775518 ( .a(n_5711), .o(n_5741) );
no02f08 g775519 ( .a(n_5716), .b(n_4874), .o(n_5711) );
na02m06 TIMEBOOST_cell_4246 ( .a(n_18190), .b(TIMEBOOST_net_1213), .o(n_18242) );
oa12s01 g775524 ( .a(n_5595), .b(n_5594), .c(n_5593), .o(n_5664) );
in01s02 g775525 ( .a(n_46999), .o(n_5723) );
na02s01 g775528 ( .a(n_5594), .b(n_5593), .o(n_5595) );
na02m02 g775530 ( .a(n_5506), .b(n_5559), .o(n_5592) );
na02f04 g775531 ( .a(n_5663), .b(n_5451), .o(n_5770) );
in01s02 g775533 ( .a(n_5572), .o(n_5596) );
na02s06 g775534 ( .a(n_5485), .b(n_5494), .o(n_5572) );
na02s02 g775535 ( .a(n_5454), .b(n_4759), .o(n_5488) );
na02f04 TIMEBOOST_cell_6252 ( .a(TIMEBOOST_net_1977), .b(n_4814), .o(n_4946) );
na02s04 g775538 ( .a(n_5581), .b(n_5451), .o(n_5465) );
na02s04 g775539 ( .a(n_5484), .b(n_4316), .o(n_5650) );
in01s02 g775541 ( .a(n_5375), .o(n_5486) );
ao12f04 g775542 ( .a(n_5248), .b(n_5232), .c(n_5185), .o(n_5375) );
no02s01 g775544 ( .a(FE_OCP_RBN4441_n_5891), .b(n_5765), .o(n_5889) );
na02f08 g775545 ( .a(n_5553), .b(n_4862), .o(n_5716) );
na02s04 g775546 ( .a(n_5632), .b(FE_OCP_RBN3024_n_47011), .o(n_5823) );
in01s02 g775549 ( .a(n_5681), .o(n_5702) );
no02s06 g775550 ( .a(n_5632), .b(FE_OCP_RBN3024_n_47011), .o(n_5681) );
ao22m02 g775551 ( .a(n_5612), .b(n_5378), .c(n_5611), .d(n_5377), .o(n_5759) );
in01s02 g775552 ( .a(n_5456), .o(n_5457) );
no02s01 TIMEBOOST_cell_3158 ( .a(n_30171), .b(n_30172), .o(TIMEBOOST_net_870) );
in01s01 g775554 ( .a(n_5645), .o(n_5613) );
oa12s01 g775555 ( .a(n_5521), .b(n_5551), .c(n_5520), .o(n_5645) );
oa12f02 g775558 ( .a(n_5134), .b(n_5138), .c(n_5041), .o(n_5272) );
in01m01 g775559 ( .a(n_5622), .o(n_5755) );
oa12f04 g775560 ( .a(n_5394), .b(n_5590), .c(n_5288), .o(n_5622) );
in01s01 g775561 ( .a(n_5739), .o(n_5740) );
oa12f02 g775562 ( .a(n_5710), .b(n_5638), .c(n_5709), .o(n_5739) );
in01s02 g775563 ( .a(n_5641), .o(n_5642) );
in01s01 g775564 ( .a(n_5608), .o(n_5641) );
oa12f06 g775566 ( .a(n_5216), .b(n_5551), .c(n_5153), .o(n_5624) );
in01s01 g775567 ( .a(n_5676), .o(n_5748) );
ao12s01 g775568 ( .a(n_5580), .b(n_5590), .c(n_5579), .o(n_5676) );
in01s01 g775569 ( .a(n_5397), .o(n_6263) );
oa22f04 g775571 ( .a(n_5236), .b(n_5169), .c(n_5206), .d(n_5170), .o(n_5397) );
in01s01 g775575 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_10_), .o(n_5619) );
na02m04 g775579 ( .a(FE_OCP_RBN4399_n_5308), .b(n_4759), .o(n_5581) );
na02f04 TIMEBOOST_cell_6296 ( .a(TIMEBOOST_net_1999), .b(n_10908), .o(n_11005) );
no02m02 g775582 ( .a(n_5473), .b(n_5512), .o(n_5559) );
no02m08 TIMEBOOST_cell_3157 ( .a(TIMEBOOST_net_869), .b(n_45185), .o(n_34908) );
na02s04 g775584 ( .a(n_5308), .b(FE_OCP_RBN2969_n_4046), .o(n_5451) );
in01s02 g775587 ( .a(n_5791), .o(n_5792) );
na02s02 g775588 ( .a(n_5783), .b(n_5728), .o(n_5791) );
na02s02 g775589 ( .a(n_5783), .b(n_5658), .o(n_5784) );
na02s01 g775590 ( .a(n_5551), .b(n_5520), .o(n_5521) );
no02m01 g775591 ( .a(n_5590), .b(n_5579), .o(n_5580) );
in01s01 g775592 ( .a(n_5725), .o(n_5726) );
na02s01 g775593 ( .a(n_5639), .b(n_5710), .o(n_5725) );
in01s01 g775594 ( .a(n_47270), .o(n_5765) );
ao12s01 g775597 ( .a(n_5548), .b(n_5552), .c(n_4702), .o(n_5594) );
oa12f06 g775598 ( .a(n_4788), .b(n_5552), .c(n_5548), .o(n_5553) );
in01s01 g775599 ( .a(n_5695), .o(n_5696) );
in01s01 g775600 ( .a(n_5663), .o(n_5695) );
ao12s04 g775601 ( .a(n_5266), .b(n_5571), .c(n_5358), .o(n_5663) );
oa22f02 g775604 ( .a(FE_OCP_RBN6830_n_45484), .b(n_5315), .c(n_45484), .d(n_5316), .o(n_5454) );
in01s02 g775605 ( .a(n_5484), .o(n_5485) );
no03f02 TIMEBOOST_cell_7570 ( .a(n_29154), .b(n_29055), .c(FE_OCP_RBN3709_n_29055), .o(TIMEBOOST_net_2416) );
oa12m02 g775607 ( .a(n_5152), .b(FE_OCP_RBN6830_n_45484), .c(n_5149), .o(n_5361) );
ao12s02 g775608 ( .a(FE_OCP_RBN6820_n_5152), .b(n_45484), .c(n_5177), .o(n_5389) );
na02f04 g775609 ( .a(n_5497), .b(n_5504), .o(n_5632) );
oa12s01 g775610 ( .a(n_5518), .b(n_5552), .c(n_5517), .o(n_5578) );
na02s01 g775613 ( .a(n_5552), .b(n_5517), .o(n_5518) );
no02s02 g775615 ( .a(n_5477), .b(n_5476), .o(n_5506) );
no02m06 TIMEBOOST_cell_5483 ( .a(TIMEBOOST_net_1689), .b(n_16072), .o(n_16216) );
no02s02 TIMEBOOST_cell_5107 ( .a(TIMEBOOST_net_1501), .b(n_8817), .o(TIMEBOOST_net_1063) );
in01m01 g775618 ( .a(n_5472), .o(n_5473) );
na02s02 g775619 ( .a(n_5458), .b(n_4606), .o(n_5472) );
no02s02 g775620 ( .a(n_5458), .b(n_4606), .o(n_5512) );
in01s02 g775621 ( .a(n_5377), .o(n_5378) );
na02s02 g775622 ( .a(n_5267), .b(n_5358), .o(n_5377) );
na02s01 g775624 ( .a(n_5736), .b(n_5662), .o(n_5761) );
na02m03 g775625 ( .a(n_5460), .b(n_5425), .o(n_5504) );
no02s02 g775626 ( .a(n_5661), .b(n_5626), .o(n_5701) );
na02m03 g775627 ( .a(n_5628), .b(n_47012), .o(n_5783) );
na02s02 g775628 ( .a(n_5627), .b(FE_OCP_RBN5956_n_47012), .o(n_5728) );
na02s03 g775629 ( .a(n_47001), .b(FE_OCPN4830_n_5603), .o(n_5710) );
na02s02 g775630 ( .a(n_5459), .b(n_5424), .o(n_5497) );
in01s01 g775631 ( .a(n_5638), .o(n_5639) );
no02s02 g775632 ( .a(n_47001), .b(FE_OCPN4830_n_5603), .o(n_5638) );
na02s04 g775633 ( .a(n_5192), .b(n_5152), .o(n_5232) );
oa12f06 g775634 ( .a(n_5116), .b(n_5455), .c(n_5203), .o(n_5551) );
in01s01 g775635 ( .a(FE_OCP_RBN3276_n_5284), .o(n_5320) );
ao12m02 g775639 ( .a(n_4956), .b(n_5031), .c(n_4966), .o(n_5138) );
no02s01 TIMEBOOST_cell_1114 ( .a(TIMEBOOST_net_171), .b(n_23535), .o(n_23619) );
in01s01 g775641 ( .a(n_5618), .o(n_5567) );
oa12s01 g775642 ( .a(n_5482), .b(n_5510), .c(n_5481), .o(n_5618) );
in01s01 g775643 ( .a(n_5538), .o(n_5569) );
ao12s01 g775644 ( .a(n_5406), .b(n_5455), .c(n_5405), .o(n_5538) );
na02s02 TIMEBOOST_cell_4260 ( .a(TIMEBOOST_net_1220), .b(n_44867), .o(n_38000) );
oa12f06 g775647 ( .a(n_5226), .b(n_5510), .c(n_5325), .o(n_5590) );
oa12s04 g775648 ( .a(n_4966), .b(FE_OCP_RBN6821_n_45319), .c(n_4956), .o(n_5206) );
ao12s02 g775649 ( .a(n_5035), .b(n_45319), .c(FE_OCP_RBN4378_n_4956), .o(n_5236) );
in01s01 g775650 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_9_), .o(n_5511) );
no02m02 g775652 ( .a(n_5409), .b(n_5313), .o(n_5477) );
na02s04 g775653 ( .a(n_5345), .b(n_5344), .o(n_5476) );
in01s02 g775654 ( .a(n_5424), .o(n_5425) );
na02s02 g775655 ( .a(n_5314), .b(n_5345), .o(n_5424) );
no02m08 TIMEBOOST_cell_3149 ( .a(TIMEBOOST_net_865), .b(n_15770), .o(n_15948) );
na02s04 g775657 ( .a(n_5215), .b(n_4556), .o(n_5358) );
no02s04 TIMEBOOST_cell_4434 ( .a(TIMEBOOST_net_1307), .b(n_4520), .o(n_4726) );
in01s02 g775659 ( .a(n_5266), .o(n_5267) );
no02s04 g775660 ( .a(n_5215), .b(n_4759), .o(n_5266) );
na02f02 TIMEBOOST_cell_6999 ( .a(TIMEBOOST_net_1297), .b(n_10369), .o(TIMEBOOST_net_2258) );
na02s03 g775662 ( .a(n_5565), .b(n_5584), .o(n_5566) );
na02m02 g775663 ( .a(n_47000), .b(n_5629), .o(n_5736) );
in01s01 g775664 ( .a(n_5661), .o(n_5662) );
no02f02 g775665 ( .a(n_47000), .b(n_5629), .o(n_5661) );
in01s02 g775666 ( .a(n_5442), .o(n_5443) );
no02m02 g775667 ( .a(n_5440), .b(n_5340), .o(n_5442) );
no02s01 TIMEBOOST_cell_1113 ( .a(n_22850), .b(n_22980), .o(TIMEBOOST_net_171) );
in01s01 g775669 ( .a(n_5598), .o(n_5599) );
no02s01 g775670 ( .a(n_5709), .b(n_5577), .o(n_5598) );
in01s01 g775671 ( .a(n_5688), .o(n_5689) );
na02s02 g775672 ( .a(n_5658), .b(n_5727), .o(n_5688) );
no02s01 g775673 ( .a(n_5455), .b(n_5405), .o(n_5406) );
na02s01 g775674 ( .a(n_5510), .b(n_5481), .o(n_5482) );
in01s01 g775675 ( .a(n_5620), .o(n_5621) );
na02s01 g775676 ( .a(n_5565), .b(n_5589), .o(n_5620) );
oa12f08 g775677 ( .a(n_4739), .b(n_5432), .c(n_4598), .o(n_5552) );
in01s01 g775678 ( .a(n_5611), .o(n_5612) );
in01s01 g775679 ( .a(n_5571), .o(n_5611) );
ao12m04 g775680 ( .a(n_5160), .b(n_5539), .c(n_5204), .o(n_5571) );
na02s02 TIMEBOOST_cell_3174 ( .a(n_34538), .b(n_34481), .o(TIMEBOOST_net_878) );
oa12m04 g775688 ( .a(n_5108), .b(n_5084), .c(n_5032), .o(n_5192) );
in01s01 g775689 ( .a(n_5527), .o(n_5489) );
oa22s01 g775690 ( .a(n_5410), .b(n_5224), .c(n_5332), .d(n_5225), .o(n_5527) );
in01s02 g775691 ( .a(n_5627), .o(n_5628) );
ao22m02 g775695 ( .a(n_5129), .b(n_5172), .c(n_5128), .d(n_5171), .o(n_5307) );
oa12s01 g775696 ( .a(n_5414), .b(n_5432), .c(n_5413), .o(n_5498) );
na02s02 g775698 ( .a(n_5357), .b(n_5402), .o(n_5478) );
in01s01 g775699 ( .a(n_5499), .o(n_5500) );
oa22s02 g775700 ( .a(n_5365), .b(FE_OCP_RBN4296_n_4080), .c(n_5335), .d(n_5529), .o(n_5499) );
in01s02 g775701 ( .a(n_5556), .o(n_5557) );
na02s02 g775702 ( .a(n_5450), .b(n_5411), .o(n_5556) );
in01s01 g775703 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_12_), .o(n_5471) );
na02s01 g775705 ( .a(n_5365), .b(FE_OCP_RBN4266_FE_RN_998_0), .o(n_5450) );
na02s01 g775706 ( .a(n_5335), .b(FE_OCP_RBN5860_FE_RN_998_0), .o(n_5411) );
na02s01 g775707 ( .a(n_5432), .b(n_5413), .o(n_5414) );
in01s01 g775708 ( .a(n_5545), .o(n_5546) );
no02s02 g775709 ( .a(n_5539), .b(n_5072), .o(n_5545) );
no02s01 TIMEBOOST_cell_1135 ( .a(n_41120), .b(n_40816), .o(TIMEBOOST_net_182) );
na02s04 g775712 ( .a(n_5159), .b(n_5071), .o(n_5160) );
in01s01 g775713 ( .a(n_5459), .o(n_5460) );
na02s02 g775714 ( .a(n_5409), .b(n_5344), .o(n_5459) );
na02m04 g775715 ( .a(n_5255), .b(n_4556), .o(n_5345) );
na02m08 TIMEBOOST_cell_4422 ( .a(TIMEBOOST_net_1301), .b(n_16044), .o(n_16220) );
in01s01 g775717 ( .a(n_5313), .o(n_5314) );
no02f02 g775718 ( .a(n_5255), .b(n_4556), .o(n_5313) );
no02s01 TIMEBOOST_cell_4501 ( .a(FE_OCP_RBN4472_n_31819), .b(n_30711), .o(TIMEBOOST_net_1341) );
in01s01 g775720 ( .a(n_5212), .o(n_5213) );
na02s02 g775721 ( .a(n_5159), .b(n_5204), .o(n_5212) );
na02s02 g775722 ( .a(n_5335), .b(n_4009), .o(n_5357) );
na02s02 g775723 ( .a(n_5365), .b(n_4069), .o(n_5402) );
na02s02 g775724 ( .a(n_5490), .b(n_3867), .o(n_5565) );
no02s04 g775725 ( .a(n_5462), .b(FE_OCP_RBN2990_n_4041), .o(n_5577) );
na02f08 g775726 ( .a(n_5410), .b(n_5150), .o(n_5510) );
in01s01 g775727 ( .a(n_5658), .o(n_5657) );
na02s02 g775728 ( .a(n_5550), .b(FE_OCP_RBN2939_n_47013), .o(n_5658) );
in01s01 g775729 ( .a(n_5659), .o(n_5660) );
no02s01 g775730 ( .a(n_5877), .b(n_5626), .o(n_5659) );
in01s01 g775732 ( .a(n_5340), .o(n_5382) );
no02s02 g775733 ( .a(n_5300), .b(FE_OCP_RBN4281_n_3848), .o(n_5340) );
na02s03 g775734 ( .a(n_5491), .b(FE_OCP_RBN2952_n_3867), .o(n_5589) );
no02m01 g775735 ( .a(n_5461), .b(n_4041), .o(n_5709) );
na02s02 g775736 ( .a(n_5549), .b(n_47013), .o(n_5727) );
no02s04 g775737 ( .a(n_5335), .b(n_3922), .o(n_5440) );
oa22m02 g775740 ( .a(n_4964), .b(n_4938), .c(n_4965), .d(n_4939), .o(n_5130) );
na02s02 g775741 ( .a(n_5335), .b(n_4163), .o(n_5336) );
no02s06 TIMEBOOST_cell_7408 ( .a(n_37093), .b(n_37100), .o(TIMEBOOST_net_2335) );
oa12f06 g775743 ( .a(n_5052), .b(n_5367), .c(n_4980), .o(n_5455) );
in01s01 g775745 ( .a(n_5418), .o(n_5483) );
ao12s01 g775746 ( .a(n_5291), .b(n_5367), .c(n_5290), .o(n_5418) );
na02s02 g775747 ( .a(n_5300), .b(n_4078), .o(n_5301) );
oa12f02 g775753 ( .a(n_4917), .b(n_4907), .c(n_4825), .o(n_5031) );
in01s01 g775757 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_8_), .o(n_5430) );
na02s02 g775759 ( .a(n_5452), .b(n_4908), .o(n_5468) );
na02s02 g775761 ( .a(n_5304), .b(n_5251), .o(n_5409) );
no02s04 g775763 ( .a(n_5421), .b(n_5051), .o(n_5532) );
na02s02 g775765 ( .a(n_5305), .b(n_5125), .o(n_5426) );
no02s03 g775766 ( .a(n_5420), .b(n_5050), .o(n_5539) );
no02s02 g775767 ( .a(n_5198), .b(n_5087), .o(n_5344) );
na02s04 g775769 ( .a(n_5251), .b(n_5199), .o(n_5310) );
na02s02 g775770 ( .a(n_5003), .b(FE_OCP_RBN2966_n_4046), .o(n_5045) );
na02s01 TIMEBOOST_cell_5444 ( .a(FE_OCPN1663_n_4556), .b(n_4675), .o(TIMEBOOST_net_1670) );
na02s02 g775772 ( .a(n_5028), .b(FE_OCP_RBN2966_n_4046), .o(n_5159) );
na02s04 g775773 ( .a(FE_OCP_RBN4380_n_5028), .b(n_4316), .o(n_5204) );
na02f06 g775774 ( .a(n_5332), .b(n_5145), .o(n_5410) );
in01s01 g775775 ( .a(n_5606), .o(n_5607) );
na02s02 g775776 ( .a(n_5584), .b(n_5583), .o(n_5606) );
in01s01 g775777 ( .a(n_5563), .o(n_5564) );
na02s01 g775778 ( .a(n_5547), .b(n_5502), .o(n_5563) );
in01s01 g775779 ( .a(n_5626), .o(n_5582) );
no02s02 g775780 ( .a(n_5508), .b(FE_OCP_RBN4289_n_47014), .o(n_5626) );
no02s06 g775781 ( .a(n_5509), .b(FE_OCP_RBN4290_n_47014), .o(n_5877) );
no02s01 g775782 ( .a(n_5367), .b(n_5290), .o(n_5291) );
no02s02 g775783 ( .a(n_5501), .b(n_5534), .o(n_5535) );
oa12f08 g775784 ( .a(n_4612), .b(n_5339), .c(n_4685), .o(n_5432) );
in01s01 g775785 ( .a(n_5490), .o(n_5491) );
in01s01 g775787 ( .a(n_5128), .o(n_5129) );
in01s01 g775788 ( .a(n_5084), .o(n_5128) );
ao12s04 g775789 ( .a(n_4975), .b(n_4916), .c(n_5026), .o(n_5084) );
oa12s01 g775790 ( .a(n_5295), .b(n_5339), .c(n_5294), .o(n_5399) );
in01s01 g775791 ( .a(FE_OCP_RBN3209_n_5221), .o(n_5265) );
no02s06 TIMEBOOST_cell_6300 ( .a(TIMEBOOST_net_2001), .b(n_35736), .o(n_35783) );
in01s04 g775802 ( .a(n_5335), .o(n_5365) );
in01m04 g775803 ( .a(n_5300), .o(n_5335) );
in01s02 g775805 ( .a(n_5549), .o(n_5550) );
no02f04 TIMEBOOST_cell_4251 ( .a(n_13273), .b(n_13310), .o(TIMEBOOST_net_1216) );
in01m02 g775807 ( .a(n_5461), .o(n_5462) );
no02m04 TIMEBOOST_cell_1130 ( .a(TIMEBOOST_net_179), .b(n_33297), .o(n_33361) );
in01s01 g775809 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_7_), .o(n_5393) );
in01s01 g775811 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_7_), .o(n_5362) );
in01s02 g775813 ( .a(n_5420), .o(n_5421) );
na02s06 g775814 ( .a(n_5359), .b(n_5013), .o(n_5420) );
in01s01 g775815 ( .a(n_5304), .o(n_5305) );
no02s02 g775816 ( .a(n_5233), .b(n_5200), .o(n_5304) );
na02s01 TIMEBOOST_cell_8579 ( .a(TIMEBOOST_net_2776), .b(n_42520), .o(n_42521) );
no02s02 TIMEBOOST_cell_7458 ( .a(FE_OCP_RBN2389_n_23227), .b(n_23226), .o(TIMEBOOST_net_2360) );
no02s02 TIMEBOOST_cell_1129 ( .a(FE_OCP_RBN6561_n_33208), .b(n_33240), .o(TIMEBOOST_net_179) );
in01s01 g775820 ( .a(n_5071), .o(n_5072) );
no02s04 g775821 ( .a(n_5030), .b(n_5051), .o(n_5071) );
na02f04 TIMEBOOST_cell_5509 ( .a(TIMEBOOST_net_1702), .b(n_16371), .o(n_16469) );
na02s02 g775823 ( .a(n_5163), .b(FE_OCP_RBN2962_n_4046), .o(n_5251) );
na02f04 TIMEBOOST_cell_7502 ( .a(n_23216), .b(FE_RN_72_0), .o(TIMEBOOST_net_2382) );
no02f06 TIMEBOOST_cell_6278 ( .a(TIMEBOOST_net_1990), .b(n_26519), .o(n_26580) );
in01s01 g775826 ( .a(n_5136), .o(n_5137) );
no02s02 g775827 ( .a(n_5050), .b(n_5030), .o(n_5136) );
na02s01 g775828 ( .a(n_5339), .b(n_5294), .o(n_5295) );
in01s01 g775829 ( .a(n_5198), .o(n_5199) );
no02s02 g775830 ( .a(n_5163), .b(FE_OCP_RBN2962_n_4046), .o(n_5198) );
in01s01 g775831 ( .a(n_5516), .o(n_5583) );
no02s02 g775832 ( .a(n_5493), .b(n_47015), .o(n_5516) );
na02s02 g775833 ( .a(n_47002), .b(n_5447), .o(n_5547) );
na02s02 g775834 ( .a(n_5493), .b(n_47015), .o(n_5584) );
in01s01 g775835 ( .a(n_5463), .o(n_5464) );
na02s01 g775836 ( .a(n_5373), .b(n_5431), .o(n_5463) );
in01s01 g775837 ( .a(n_5501), .o(n_5502) );
no02s02 g775838 ( .a(n_47002), .b(n_5447), .o(n_5501) );
ao12m02 g775840 ( .a(n_4676), .b(n_5364), .c(n_4716), .o(n_5452) );
oa12s01 g775841 ( .a(n_5263), .b(n_5262), .c(n_5261), .o(n_5371) );
oa22s02 g775843 ( .a(FE_OCP_RBN6025_n_4858), .b(FE_OCP_RBN2967_n_4046), .c(n_4858), .d(FE_OCP_RBN2964_n_4046), .o(n_5028) );
in01s01 g775844 ( .a(n_4964), .o(n_4965) );
in01s01 g775845 ( .a(n_4907), .o(n_4964) );
ao12s02 g775846 ( .a(n_4578), .b(n_4776), .c(n_4659), .o(n_4907) );
ao12f04 g775847 ( .a(n_4962), .b(n_5283), .c(n_5017), .o(n_5332) );
oa12f06 g775848 ( .a(n_4823), .b(n_5240), .c(n_4919), .o(n_5367) );
in01s01 g775849 ( .a(n_5350), .o(n_5408) );
ao12s01 g775850 ( .a(n_5229), .b(n_5283), .c(n_5228), .o(n_5350) );
in01s02 g775851 ( .a(n_5508), .o(n_5509) );
oa22m02 g775852 ( .a(n_5400), .b(n_4789), .c(n_5364), .d(n_4790), .o(n_5508) );
in01s01 g775856 ( .a(n_5286), .o(n_5379) );
ao12s01 g775857 ( .a(n_5195), .b(n_5240), .c(n_5194), .o(n_5286) );
na02s01 g775859 ( .a(n_5262), .b(n_5261), .o(n_5263) );
oa12f08 g775860 ( .a(n_4577), .b(n_5193), .c(n_4460), .o(n_5339) );
in01s01 g775861 ( .a(n_5230), .o(n_5231) );
no02s02 g775862 ( .a(n_5200), .b(n_5087), .o(n_5230) );
no02s02 g775863 ( .a(n_4922), .b(n_4316), .o(n_5030) );
in01s02 g775864 ( .a(n_5142), .o(n_5143) );
no02s04 g775865 ( .a(FE_OCP_RBN4387_n_5013), .b(n_5051), .o(n_5142) );
no02s03 g775866 ( .a(n_4923), .b(FE_OCP_RBN2964_n_4046), .o(n_5050) );
in01s01 g775867 ( .a(n_5249), .o(n_5250) );
no02s02 g775868 ( .a(n_5248), .b(n_5184), .o(n_5249) );
no02s01 g775869 ( .a(n_5283), .b(n_5228), .o(n_5229) );
no02s01 g775870 ( .a(n_5240), .b(n_5194), .o(n_5195) );
no02s04 g775871 ( .a(n_5184), .b(n_5149), .o(n_5185) );
na02s01 g775872 ( .a(n_5475), .b(n_5374), .o(n_5697) );
in01s01 g775873 ( .a(n_5372), .o(n_5373) );
no02s03 g775874 ( .a(n_47003), .b(n_47016), .o(n_5372) );
na02s02 g775875 ( .a(n_47003), .b(n_47016), .o(n_5431) );
oa12s02 g775877 ( .a(n_4802), .b(n_5217), .c(n_4842), .o(n_5346) );
in01s01 g775879 ( .a(n_5359), .o(n_5395) );
oa12m04 g775880 ( .a(n_4844), .b(n_5234), .c(n_4808), .o(n_5359) );
in01s02 g775881 ( .a(n_5276), .o(n_5277) );
in01s02 g775882 ( .a(n_5233), .o(n_5276) );
ao12f02 g775883 ( .a(n_5002), .b(n_5140), .c(n_4979), .o(n_5233) );
in01s01 g775885 ( .a(n_5323), .o(n_5285) );
oa12s01 g775886 ( .a(n_5158), .b(n_5157), .c(n_5156), .o(n_5323) );
in01s02 g775888 ( .a(n_5049), .o(n_5076) );
in01s02 g775890 ( .a(n_4968), .o(n_4969) );
in01m01 g775891 ( .a(n_4916), .o(n_4968) );
in01s01 g775893 ( .a(n_5363), .o(n_5324) );
oa12s01 g775894 ( .a(n_5209), .b(n_5208), .c(n_5207), .o(n_5363) );
no02m10 TIMEBOOST_cell_8471 ( .a(TIMEBOOST_net_2722), .b(n_22972), .o(n_22998) );
no02f08 TIMEBOOST_cell_8880 ( .a(n_45050), .b(FE_OCP_RBN1159_n_20763), .o(TIMEBOOST_net_2927) );
no02m10 TIMEBOOST_cell_838 ( .a(TIMEBOOST_net_33), .b(n_1547), .o(n_1602) );
in01s01 g775899 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_6_), .o(n_5312) );
no02s01 g775904 ( .a(n_5193), .b(n_4503), .o(n_5262) );
ao12m02 g775905 ( .a(n_4848), .b(n_4853), .c(n_4841), .o(n_5011) );
no03m08 TIMEBOOST_cell_8354 ( .a(n_14215), .b(FE_OCP_RBN5993_n_15387), .c(n_15503), .o(n_15623) );
na02s02 g775907 ( .a(n_5217), .b(n_4868), .o(n_5351) );
in01s01 g775909 ( .a(n_5364), .o(n_5400) );
no02m06 g775910 ( .a(n_5235), .b(n_4603), .o(n_5364) );
in01s01 g775912 ( .a(n_5087), .o(n_5125) );
no02m04 g775913 ( .a(FE_OCP_RBN3180_n_4959), .b(FE_OCP_RBN2962_n_4046), .o(n_5087) );
na02s06 TIMEBOOST_cell_3161 ( .a(TIMEBOOST_net_871), .b(n_45185), .o(n_34906) );
no02s02 g775915 ( .a(n_4959), .b(FE_OCP_RBN2966_n_4046), .o(n_5200) );
no02s03 g775916 ( .a(n_4936), .b(n_4316), .o(n_5051) );
na02m03 g775918 ( .a(n_4936), .b(n_4316), .o(n_5013) );
no02s03 TIMEBOOST_cell_6980 ( .a(TIMEBOOST_net_2248), .b(n_24254), .o(TIMEBOOST_net_1556) );
na02f06 g775920 ( .a(n_5023), .b(FE_OCPN4547_n_4727), .o(n_5240) );
in01s01 g775921 ( .a(n_5315), .o(n_5316) );
na02s02 g775922 ( .a(n_5177), .b(n_5152), .o(n_5315) );
na02s02 g775923 ( .a(n_5218), .b(n_4647), .o(n_5279) );
na02s01 g775925 ( .a(n_5157), .b(n_5156), .o(n_5158) );
no02s01 g775926 ( .a(n_5275), .b(n_5353), .o(n_5616) );
in01s01 g775927 ( .a(n_5412), .o(n_5475) );
no02s03 g775928 ( .a(n_5322), .b(n_3817), .o(n_5412) );
na02s01 g775929 ( .a(n_5289), .b(n_5394), .o(n_5579) );
no02s02 g775930 ( .a(n_5085), .b(FE_OCP_RBN6745_n_3746), .o(n_5184) );
no02s06 g775931 ( .a(FE_OCP_RBN3145_n_5085), .b(FE_OCP_RBN6744_n_3746), .o(n_5248) );
in01s01 g775932 ( .a(n_5534), .o(n_5374) );
no02s02 g775933 ( .a(n_5321), .b(n_3819), .o(n_5534) );
ao12f04 g775934 ( .a(n_4949), .b(n_5020), .c(n_4935), .o(n_5283) );
na02s01 g775935 ( .a(n_5208), .b(n_5207), .o(n_5209) );
in01s01 g775936 ( .a(n_4849), .o(n_4850) );
in01s01 g775937 ( .a(n_4776), .o(n_4849) );
oa12m02 g775938 ( .a(n_4474), .b(n_4605), .c(n_4411), .o(n_4776) );
oa12s01 g775939 ( .a(n_5132), .b(n_5144), .c(n_5131), .o(n_5211) );
in01s02 g775941 ( .a(n_4922), .o(n_4923) );
ao22m02 g775942 ( .a(FE_OCP_RBN3120_n_4751), .b(n_4316), .c(n_4751), .d(FE_OCP_RBN2964_n_4046), .o(n_4922) );
in01s01 g775943 ( .a(FE_OCP_RBN3144_n_4858), .o(n_4904) );
oa22s02 g775946 ( .a(FE_OCP_RBN6009_n_4683), .b(n_4533), .c(n_4683), .d(n_4532), .o(n_4858) );
no02f08 g775947 ( .a(n_5144), .b(n_4504), .o(n_5193) );
na02s01 g775948 ( .a(n_5144), .b(n_5131), .o(n_5132) );
na02s02 g775949 ( .a(n_4807), .b(n_4717), .o(n_4808) );
in01s01 g775951 ( .a(n_5217), .o(n_5280) );
na02s04 g775952 ( .a(n_5141), .b(n_4658), .o(n_5217) );
no02m02 g775953 ( .a(n_4978), .b(n_4843), .o(n_4979) );
na02s02 g775955 ( .a(n_4807), .b(FE_OCP_RBN6040_n_4800), .o(n_4908) );
in01s01 g775956 ( .a(n_5065), .o(n_5066) );
no02s01 g775957 ( .a(n_4978), .b(n_4958), .o(n_5065) );
no02s02 g775959 ( .a(n_5181), .b(n_4549), .o(n_5218) );
in01s04 g775960 ( .a(n_5234), .o(n_5235) );
na02f04 g775961 ( .a(n_5181), .b(n_4507), .o(n_5234) );
in01s02 g775964 ( .a(n_5149), .o(n_5177) );
no02s04 g775965 ( .a(n_5101), .b(FE_OCPN3576_n_3625), .o(n_5149) );
no02s02 g775966 ( .a(n_5243), .b(n_5242), .o(n_5353) );
na02s03 g775971 ( .a(n_5101), .b(FE_OCPN3576_n_3625), .o(n_5152) );
in01s02 g775972 ( .a(n_5171), .o(n_5172) );
na02s02 g775973 ( .a(n_5108), .b(FE_OCP_RBN4371_n_5032), .o(n_5171) );
no02s01 g775974 ( .a(n_5325), .b(n_5227), .o(n_5481) );
na02s01 g775975 ( .a(n_5216), .b(n_5154), .o(n_5520) );
no02s04 g775976 ( .a(n_4729), .b(n_4601), .o(n_4730) );
na02s02 g775977 ( .a(n_5253), .b(n_47019), .o(n_5394) );
in01s02 g775978 ( .a(n_5169), .o(n_5170) );
na02s04 g775979 ( .a(n_5134), .b(FE_OCP_RBN4381_n_5041), .o(n_5169) );
no02m02 g775980 ( .a(n_5123), .b(n_4723), .o(n_5161) );
in01s01 g775982 ( .a(n_5274), .o(n_5275) );
na02s02 g775983 ( .a(n_5243), .b(n_5242), .o(n_5274) );
in01s01 g775984 ( .a(n_5288), .o(n_5289) );
no02m02 g775985 ( .a(n_5253), .b(n_47019), .o(n_5288) );
na02s02 g775986 ( .a(n_5048), .b(n_5036), .o(n_5127) );
no02s02 g775987 ( .a(n_4800), .b(n_4669), .o(n_4844) );
na02m02 g775988 ( .a(n_4957), .b(n_4763), .o(n_5002) );
oa12f04 g775992 ( .a(n_4767), .b(n_4942), .c(n_4689), .o(n_5023) );
ao12s01 g775993 ( .a(n_4918), .b(n_5107), .c(n_4821), .o(n_5208) );
in01s01 g775994 ( .a(n_4815), .o(n_4816) );
oa12s02 g775995 ( .a(n_4688), .b(n_4624), .c(n_4601), .o(n_4815) );
no02s02 g775996 ( .a(n_4729), .b(n_4591), .o(n_4736) );
no02m01 TIMEBOOST_cell_8476 ( .a(n_12055), .b(n_11975), .o(TIMEBOOST_net_2725) );
oa12s01 g776001 ( .a(n_5081), .b(n_5080), .c(n_5079), .o(n_5151) );
in01s01 g776002 ( .a(n_5196), .o(n_5273) );
ao12s01 g776003 ( .a(n_5060), .b(n_5059), .c(n_5058), .o(n_5196) );
in01s02 g776004 ( .a(n_5321), .o(n_5322) );
no03s02 TIMEBOOST_cell_5506 ( .a(n_5142), .b(n_5359), .c(n_5143), .o(TIMEBOOST_net_1701) );
no02f06 TIMEBOOST_cell_5313 ( .a(TIMEBOOST_net_1604), .b(n_20320), .o(n_20420) );
oa12s01 g776007 ( .a(n_4644), .b(n_4986), .c(n_4765), .o(n_5157) );
in01s01 g776008 ( .a(n_5244), .o(n_5210) );
oa12s01 g776009 ( .a(n_5054), .b(n_5107), .c(n_5053), .o(n_5244) );
in01s01 g776010 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_8_), .o(n_5104) );
in01s01 g776014 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_5_), .o(n_5139) );
na02s02 g776017 ( .a(n_5061), .b(n_5009), .o(n_5036) );
in01s02 g776018 ( .a(n_5098), .o(n_5099) );
na02s04 g776019 ( .a(n_5061), .b(n_5018), .o(n_5098) );
na02s01 g776020 ( .a(n_5080), .b(n_5079), .o(n_5081) );
na02s02 g776021 ( .a(n_4872), .b(n_4878), .o(n_4898) );
na02s01 TIMEBOOST_cell_4374 ( .a(TIMEBOOST_net_1277), .b(n_15403), .o(n_15449) );
no02s01 TIMEBOOST_cell_3877 ( .a(n_7), .b(TIMEBOOST_net_603), .o(TIMEBOOST_net_1029) );
in01s01 g776024 ( .a(n_5140), .o(n_5141) );
no02s03 g776025 ( .a(n_5055), .b(n_4616), .o(n_5140) );
na02s02 g776026 ( .a(n_4726), .b(n_4316), .o(n_4807) );
no02s02 g776027 ( .a(n_4915), .b(FE_OCP_RBN6783_n_4046), .o(n_4978) );
na02f06 TIMEBOOST_cell_3119 ( .a(TIMEBOOST_net_850), .b(n_14772), .o(n_14886) );
no02s04 g776030 ( .a(n_4726), .b(n_4316), .o(n_4800) );
in01s01 g776031 ( .a(n_4957), .o(n_4958) );
na02s02 g776032 ( .a(n_4915), .b(FE_OCP_RBN6783_n_4046), .o(n_4957) );
na02s03 g776034 ( .a(n_5055), .b(n_4625), .o(n_5123) );
no02s02 TIMEBOOST_cell_4410 ( .a(TIMEBOOST_net_1295), .b(n_15396), .o(n_15569) );
no02f04 g776036 ( .a(n_5077), .b(n_4428), .o(n_5181) );
na02s01 TIMEBOOST_cell_6364 ( .a(TIMEBOOST_net_2033), .b(n_17221), .o(n_17378) );
in01s02 g776039 ( .a(n_5082), .o(n_5083) );
na02s02 g776040 ( .a(n_5026), .b(n_4976), .o(n_5082) );
na02m02 g776041 ( .a(n_4837), .b(n_4517), .o(n_4853) );
no02m04 g776043 ( .a(n_47005), .b(FE_OCP_RBN2847_n_47018), .o(n_5032) );
in01s01 g776044 ( .a(n_5226), .o(n_5227) );
na02s03 g776045 ( .a(n_47004), .b(n_5178), .o(n_5226) );
na02s02 g776046 ( .a(n_4989), .b(FE_OCP_RBN2900_n_3807), .o(n_5134) );
na02s01 g776047 ( .a(n_5107), .b(n_5053), .o(n_5054) );
no02s03 g776048 ( .a(n_47004), .b(n_5178), .o(n_5325) );
na02m02 g776049 ( .a(n_5115), .b(n_4496), .o(n_5176) );
na02s03 g776050 ( .a(n_47005), .b(FE_OCP_RBN2846_n_47018), .o(n_5108) );
na02s02 g776051 ( .a(n_5110), .b(n_5109), .o(n_5216) );
no02s01 g776052 ( .a(n_5224), .b(n_5146), .o(n_5225) );
no02s06 g776053 ( .a(n_4581), .b(n_4544), .o(n_4729) );
in01s01 g776054 ( .a(n_5153), .o(n_5154) );
no02s03 g776055 ( .a(n_5110), .b(n_5109), .o(n_5153) );
no02m02 g776057 ( .a(n_4989), .b(FE_OCP_RBN2900_n_3807), .o(n_5041) );
no02s01 g776058 ( .a(n_5117), .b(n_5203), .o(n_5405) );
no02s01 g776059 ( .a(n_5059), .b(n_5058), .o(n_5060) );
na02f04 g776060 ( .a(n_4990), .b(n_4787), .o(n_5020) );
no02m02 g776062 ( .a(n_4559), .b(FE_OCP_RBN3043_n_4296), .o(n_4683) );
oa22s02 g776065 ( .a(n_4531), .b(n_4452), .c(n_4530), .d(n_4451), .o(n_4751) );
in01s01 g776066 ( .a(n_5095), .o(n_5096) );
na02s02 g776067 ( .a(n_4994), .b(n_4940), .o(n_5095) );
no02s06 TIMEBOOST_cell_6346 ( .a(TIMEBOOST_net_2024), .b(n_31869), .o(TIMEBOOST_net_968) );
no02s02 TIMEBOOST_cell_5360 ( .a(n_3905), .b(n_3835), .o(TIMEBOOST_net_1628) );
na03f06 TIMEBOOST_cell_2497 ( .a(TIMEBOOST_net_389), .b(n_8528), .c(n_8578), .o(n_8641) );
in01s02 g776071 ( .a(n_5093), .o(n_5094) );
no02s03 TIMEBOOST_cell_3254 ( .a(n_44853), .b(n_10413), .o(TIMEBOOST_net_918) );
ao12s02 g776073 ( .a(n_4557), .b(n_4558), .c(n_4296), .o(n_4605) );
in01s01 g776074 ( .a(n_5056), .o(n_5057) );
oa22s02 g776075 ( .a(n_5048), .b(n_5422), .c(FE_OCP_RBN4372_n_5048), .d(FE_OCP_RBN2987_n_4238), .o(n_5056) );
in01s02 g776078 ( .a(n_4998), .o(n_5018) );
no02s04 g776079 ( .a(n_5048), .b(FE_OCP_RBN2942_n_4101), .o(n_4998) );
na02s04 g776080 ( .a(n_5048), .b(FE_OCP_RBN2942_n_4101), .o(n_5061) );
no02s01 g776081 ( .a(n_4928), .b(n_4292), .o(n_5080) );
in01s01 g776082 ( .a(n_4878), .o(n_4879) );
oa12m02 g776083 ( .a(n_4666), .b(n_4656), .c(n_4804), .o(n_4878) );
no02m02 g776084 ( .a(n_4840), .b(n_4804), .o(n_4841) );
in01s02 g776085 ( .a(FE_OCP_RBN3089_n_4872), .o(n_4900) );
no02s02 g776088 ( .a(n_4840), .b(n_4848), .o(n_4872) );
no02s02 g776089 ( .a(n_4842), .b(n_4657), .o(n_4763) );
na02s02 g776090 ( .a(n_4716), .b(n_4602), .o(n_4669) );
na02f04 g776091 ( .a(n_4946), .b(n_4546), .o(n_5055) );
in01s02 g776092 ( .a(n_4789), .o(n_4790) );
na02s02 g776093 ( .a(n_4717), .b(n_4716), .o(n_4789) );
in01s01 g776094 ( .a(n_4867), .o(n_4868) );
no02s02 g776095 ( .a(n_4843), .b(n_4842), .o(n_4867) );
na02s01 g776096 ( .a(n_4981), .b(n_5052), .o(n_5290) );
no02s02 g776097 ( .a(n_5048), .b(FE_OCP_RBN2950_n_4158), .o(n_5021) );
na02s01 g776098 ( .a(n_4946), .b(n_4595), .o(n_5064) );
no02f06 TIMEBOOST_cell_7817 ( .a(TIMEBOOST_net_2539), .b(FE_OCP_RBN2673_n_38534), .o(n_38596) );
in01s01 g776100 ( .a(n_5116), .o(n_5117) );
na02s02 g776101 ( .a(n_5063), .b(n_5062), .o(n_5116) );
in01s01 g776102 ( .a(n_4975), .o(n_4976) );
no02m04 g776103 ( .a(n_4906), .b(FE_OCP_RBN2853_n_4905), .o(n_4975) );
na02s02 g776104 ( .a(n_4906), .b(FE_OCP_RBN2853_n_4905), .o(n_5026) );
in01s02 g776105 ( .a(n_5105), .o(n_5106) );
na02s02 g776106 ( .a(FE_OCP_RBN4379_n_4956), .b(n_4966), .o(n_5105) );
in01s01 g776107 ( .a(n_5145), .o(n_5146) );
na02s02 g776108 ( .a(n_5015), .b(n_3697), .o(n_5145) );
no02s02 g776109 ( .a(n_5063), .b(n_5062), .o(n_5203) );
no02s02 TIMEBOOST_cell_6345 ( .a(n_31864), .b(n_31835), .o(TIMEBOOST_net_2024) );
na02s01 g776111 ( .a(n_5048), .b(n_4467), .o(n_4940) );
no02s06 TIMEBOOST_cell_1089 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_19_), .b(n_32860), .o(TIMEBOOST_net_159) );
na02s01 g776113 ( .a(FE_OCP_RBN4372_n_5048), .b(n_4466), .o(n_4994) );
no02m01 g776114 ( .a(n_4558), .b(n_4557), .o(n_4559) );
no02s02 TIMEBOOST_cell_8149 ( .a(TIMEBOOST_net_2705), .b(n_12796), .o(TIMEBOOST_net_764) );
no02f06 TIMEBOOST_cell_5359 ( .a(TIMEBOOST_net_1627), .b(n_15039), .o(n_15343) );
in01s01 g776117 ( .a(n_5150), .o(n_5224) );
na02s04 g776118 ( .a(n_5016), .b(n_3663), .o(n_5150) );
na02m02 g776119 ( .a(n_4742), .b(n_4855), .o(n_4920) );
in01s01 g776120 ( .a(n_4837), .o(n_4838) );
no02m04 g776121 ( .a(n_4848), .b(n_4620), .o(n_4837) );
oa12s01 g776122 ( .a(n_4892), .b(n_4891), .c(n_4890), .o(n_4997) );
in01s01 g776124 ( .a(FE_OCP_RBN4366_n_4692), .o(n_5940) );
oa12s01 g776128 ( .a(n_4912), .b(n_4911), .c(n_4910), .o(n_4987) );
na02s04 g776129 ( .a(n_4660), .b(n_45463), .o(n_4915) );
no03s08 TIMEBOOST_cell_8420 ( .a(n_39905), .b(n_39812), .c(n_39982), .o(TIMEBOOST_net_983) );
in01s01 g776133 ( .a(n_4624), .o(n_4690) );
in01s01 g776134 ( .a(n_4581), .o(n_4624) );
oa12s02 g776135 ( .a(n_4484), .b(n_4454), .c(n_4394), .o(n_4581) );
no02s04 g776139 ( .a(n_4611), .b(n_4639), .o(n_4784) );
in01s01 g776140 ( .a(n_4990), .o(n_5107) );
ao12f04 g776141 ( .a(n_4799), .b(n_4951), .c(n_4673), .o(n_4990) );
in01s02 g776143 ( .a(n_5114), .o(n_5115) );
in01s01 g776144 ( .a(n_5077), .o(n_5114) );
in01s01 g776146 ( .a(n_4986), .o(n_5059) );
in01s01 g776147 ( .a(n_4942), .o(n_4986) );
oa12f04 g776148 ( .a(n_4649), .b(n_4806), .c(n_4735), .o(n_4942) );
oa22f02 g776149 ( .a(n_4782), .b(FE_OCP_RBN4266_FE_RN_998_0), .c(n_4783), .d(FE_OCP_RBN5860_FE_RN_998_0), .o(n_4989) );
no02s02 TIMEBOOST_cell_1122 ( .a(TIMEBOOST_net_175), .b(n_33359), .o(n_33360) );
oa12s01 g776151 ( .a(n_4930), .b(n_4929), .c(n_4951), .o(n_4992) );
in01s01 g776152 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_4_), .o(n_4948) );
in01s01 g776156 ( .a(n_4927), .o(n_4928) );
na02f06 g776157 ( .a(n_4851), .b(n_4217), .o(n_4927) );
na02s01 g776158 ( .a(n_4911), .b(n_4910), .o(n_4912) );
no02m02 TIMEBOOST_cell_3087 ( .a(TIMEBOOST_net_834), .b(n_3418), .o(TIMEBOOST_net_392) );
no02s02 g776161 ( .a(n_4653), .b(FE_OFN4765_n_3029), .o(n_4840) );
no02s06 g776162 ( .a(n_4652), .b(n_3082), .o(n_4848) );
no02s02 g776163 ( .a(n_4933), .b(n_4348), .o(n_5012) );
no02s02 TIMEBOOST_cell_1121 ( .a(n_33311), .b(n_33313), .o(TIMEBOOST_net_175) );
no02s02 g776165 ( .a(n_4861), .b(n_4476), .o(n_4941) );
na02s02 g776167 ( .a(n_47008), .b(n_4316), .o(n_4660) );
na02s02 g776169 ( .a(n_4554), .b(FE_OCP_RBN6778_n_4046), .o(n_4716) );
in01s01 g776170 ( .a(n_4843), .o(n_4802) );
no02s02 g776171 ( .a(FE_OCP_RBN6816_n_4654), .b(FE_OCP_RBN6783_n_4046), .o(n_4843) );
na02f04 TIMEBOOST_cell_6085 ( .a(n_24968), .b(FE_OCP_RBN5718_n_24718), .o(TIMEBOOST_net_1894) );
in01s01 g776173 ( .a(n_4717), .o(n_4676) );
na02s03 g776174 ( .a(n_4555), .b(n_4316), .o(n_4717) );
na03s20 TIMEBOOST_cell_4574 ( .a(n_16899), .b(delay_xor_ln21_unr12_stage5_stallmux_q_2_), .c(FE_OCP_RBN7112_n_44365), .o(n_16984) );
no02s02 TIMEBOOST_cell_6303 ( .a(n_10890), .b(n_10834), .o(TIMEBOOST_net_2003) );
no02s03 g776177 ( .a(n_4654), .b(FE_OCP_RBN6767_n_3704), .o(n_4842) );
in01s01 g776178 ( .a(n_5024), .o(n_5025) );
no02s02 g776179 ( .a(n_4895), .b(n_4424), .o(n_5024) );
no02s02 g776180 ( .a(n_4505), .b(FE_OCP_RBN6809_n_4563), .o(n_4639) );
na02s02 g776181 ( .a(n_4462), .b(n_4236), .o(n_4524) );
in01s01 g776182 ( .a(n_4966), .o(n_5035) );
na02m06 g776186 ( .a(n_4887), .b(n_4886), .o(n_4966) );
na02s01 g776187 ( .a(n_4891), .b(n_4890), .o(n_4892) );
na02s01 g776188 ( .a(n_4929), .b(n_4951), .o(n_4930) );
in01s01 g776189 ( .a(n_4980), .o(n_4981) );
no02s03 g776190 ( .a(n_4954), .b(n_4953), .o(n_4980) );
no02f06 g776194 ( .a(n_4887), .b(n_4886), .o(n_4956) );
na02s03 g776195 ( .a(n_4954), .b(n_4953), .o(n_5052) );
no02m08 TIMEBOOST_cell_5057 ( .a(TIMEBOOST_net_1476), .b(TIMEBOOST_net_309), .o(n_19101) );
na02s01 g776197 ( .a(n_4963), .b(n_5017), .o(n_5228) );
in01s02 g776198 ( .a(n_4938), .o(n_4939) );
na02s02 g776199 ( .a(n_4917), .b(n_4826), .o(n_4938) );
no02s02 g776200 ( .a(n_4506), .b(n_4563), .o(n_4611) );
in01s01 g776201 ( .a(n_4855), .o(n_4856) );
oa12s02 g776202 ( .a(n_4535), .b(n_4630), .c(n_4568), .o(n_4855) );
in01s01 g776204 ( .a(n_4946), .o(n_4995) );
na02f02 TIMEBOOST_cell_7722 ( .a(n_15384), .b(n_14452), .o(TIMEBOOST_net_2492) );
in01s01 g776206 ( .a(n_4530), .o(n_4531) );
in01s01 g776207 ( .a(n_4558), .o(n_4530) );
na02m04 g776208 ( .a(n_4338), .b(n_4264), .o(n_4558) );
na02f08 g776210 ( .a(n_4740), .b(n_4795), .o(n_5048) );
in01s01 g776212 ( .a(n_5015), .o(n_5016) );
no02s01 TIMEBOOST_cell_1076 ( .a(TIMEBOOST_net_152), .b(FE_OCP_RBN7021_n_33330), .o(n_33381) );
na02s02 TIMEBOOST_cell_6342 ( .a(TIMEBOOST_net_2022), .b(n_6327), .o(n_6456) );
na02s03 g776215 ( .a(n_4667), .b(FE_OCP_RBN5860_FE_RN_998_0), .o(n_4740) );
na02m06 g776216 ( .a(n_4668), .b(FE_OCP_RBN4266_FE_RN_998_0), .o(n_4795) );
no02s02 g776217 ( .a(n_4583), .b(n_4592), .o(n_4656) );
na02s03 g776218 ( .a(n_4666), .b(n_4535), .o(n_4620) );
na02s03 g776220 ( .a(n_4630), .b(FE_OCP_RBN4339_n_4403), .o(n_4743) );
in01s01 g776221 ( .a(n_4741), .o(n_4742) );
na02s03 g776222 ( .a(n_4666), .b(n_4665), .o(n_4741) );
na02s02 g776224 ( .a(n_4830), .b(n_4516), .o(n_4876) );
na02s01 TIMEBOOST_cell_6341 ( .a(n_45475), .b(n_5636), .o(TIMEBOOST_net_2022) );
in01s01 g776226 ( .a(n_4860), .o(n_4861) );
no02s02 g776227 ( .a(n_4814), .b(n_4487), .o(n_4860) );
no02m08 TIMEBOOST_cell_8519 ( .a(TIMEBOOST_net_2746), .b(n_13759), .o(n_13860) );
na02s02 g776230 ( .a(n_4812), .b(n_4345), .o(n_4933) );
in01s01 g776231 ( .a(n_4657), .o(n_4658) );
na02s02 g776232 ( .a(n_4626), .b(n_4625), .o(n_4657) );
in01s02 g776233 ( .a(n_4602), .o(n_4603) );
no02m02 g776234 ( .a(n_4550), .b(n_4549), .o(n_4602) );
na02m02 g776236 ( .a(n_4626), .b(n_4617), .o(n_4723) );
no02s02 g776238 ( .a(n_4508), .b(n_4550), .o(n_4647) );
in01s01 g776239 ( .a(n_4894), .o(n_4895) );
na02m04 g776240 ( .a(n_4811), .b(n_4287), .o(n_4894) );
in01s01 g776241 ( .a(n_4962), .o(n_4963) );
no02s02 g776242 ( .a(n_47006), .b(n_47341), .o(n_4962) );
in01s01 g776243 ( .a(n_4462), .o(n_4463) );
na02s02 g776244 ( .a(n_4320), .b(n_4175), .o(n_4462) );
na02s02 g776245 ( .a(n_4319), .b(n_4263), .o(n_4338) );
in01s01 g776246 ( .a(n_4851), .o(n_4911) );
na02f06 TIMEBOOST_cell_4237 ( .a(n_37534), .b(n_37709), .o(TIMEBOOST_net_1209) );
in01s01 g776248 ( .a(n_4825), .o(n_4826) );
no02s02 g776249 ( .a(n_4792), .b(FE_OFN4816_n_47017), .o(n_4825) );
no02s04 TIMEBOOST_cell_7521 ( .a(TIMEBOOST_net_2391), .b(n_13165), .o(n_13313) );
na02s02 g776251 ( .a(n_47006), .b(n_47341), .o(n_5017) );
na02m02 g776252 ( .a(n_4792), .b(FE_OFN4816_n_47017), .o(n_4917) );
no02s01 g776253 ( .a(n_4824), .b(n_4919), .o(n_5194) );
no02s04 g776254 ( .a(n_4931), .b(n_4774), .o(n_4935) );
na02s01 g776255 ( .a(n_4950), .b(n_4932), .o(n_5207) );
no02s01 TIMEBOOST_cell_1075 ( .a(n_33380), .b(n_33160), .o(TIMEBOOST_net_152) );
na02s04 g776257 ( .a(n_4536), .b(n_4665), .o(n_4804) );
in01s02 g776258 ( .a(n_4782), .o(n_4783) );
no02m02 TIMEBOOST_cell_6149 ( .a(TIMEBOOST_net_1094), .b(n_35092), .o(TIMEBOOST_net_1926) );
oa12s01 g776260 ( .a(n_4696), .b(n_4697), .c(n_4695), .o(n_4775) );
oa12s01 g776261 ( .a(n_4757), .b(n_4786), .c(n_4756), .o(n_4828) );
in01s01 g776262 ( .a(n_4806), .o(n_4891) );
oa12f04 g776263 ( .a(n_4480), .b(n_4786), .c(n_4582), .o(n_4806) );
in01s01 g776264 ( .a(n_4505), .o(n_4506) );
in01s01 g776265 ( .a(n_4454), .o(n_4505) );
oa12s04 g776266 ( .a(n_4365), .b(n_4323), .c(n_4248), .o(n_4454) );
na02f04 TIMEBOOST_cell_8735 ( .a(TIMEBOOST_net_2854), .b(n_18757), .o(n_18893) );
na02s01 TIMEBOOST_cell_1116 ( .a(n_33273), .b(TIMEBOOST_net_172), .o(n_33275) );
ao12f04 g776269 ( .a(n_4482), .b(n_4827), .c(n_4594), .o(n_4951) );
in01s02 g776270 ( .a(n_4554), .o(n_4555) );
in01s01 g776273 ( .a(n_4459), .o(n_4520) );
oa22s02 g776274 ( .a(n_4271), .b(n_4226), .c(n_4272), .d(FE_OCP_RBN5991_n_4226), .o(n_4459) );
oa12s01 g776275 ( .a(n_4781), .b(n_4827), .c(n_4780), .o(n_4857) );
in01s01 g776276 ( .a(n_4652), .o(n_4653) );
no02m04 TIMEBOOST_cell_8545 ( .a(TIMEBOOST_net_2759), .b(n_38530), .o(TIMEBOOST_net_2430) );
ao22m02 g776279 ( .a(FE_OCP_RBN3088_n_4458), .b(FE_OCP_RBN2921_n_3878), .c(n_4458), .d(FE_OCP_RBN6767_n_3704), .o(n_4654) );
in01s01 g776281 ( .a(n_47008), .o(n_4700) );
no02s01 TIMEBOOST_cell_4193 ( .a(n_36750), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_1187) );
na02s01 g776290 ( .a(n_4697), .b(n_4695), .o(n_4696) );
no02m03 g776291 ( .a(n_4635), .b(n_5529), .o(n_4713) );
na02m06 TIMEBOOST_cell_8017 ( .a(TIMEBOOST_net_2639), .b(n_45474), .o(n_6363) );
no02s04 g776293 ( .a(n_4468), .b(n_4568), .o(n_4536) );
na02m08 g776296 ( .a(n_4592), .b(n_4397), .o(n_4630) );
no03f10 TIMEBOOST_cell_6421 ( .a(TIMEBOOST_net_1847), .b(FE_RN_286_0), .c(FE_RN_285_0), .o(n_28125) );
in01m01 g776299 ( .a(n_4535), .o(n_4583) );
no02s04 g776300 ( .a(n_4475), .b(n_4403), .o(n_4535) );
na02s06 g776301 ( .a(n_4472), .b(FE_OFN4765_n_3029), .o(n_4666) );
na02s02 g776302 ( .a(n_4396), .b(n_4093), .o(n_4439) );
no02s01 TIMEBOOST_cell_6391 ( .a(FE_OCPN5113_n_22249), .b(n_21393), .o(TIMEBOOST_net_2047) );
no02s04 g776305 ( .a(n_4568), .b(n_4475), .o(n_4609) );
na02s06 g776306 ( .a(n_4473), .b(n_3297), .o(n_4665) );
in01s01 g776307 ( .a(n_4830), .o(n_4831) );
no02s02 g776308 ( .a(n_4704), .b(n_4274), .o(n_4830) );
na02s01 TIMEBOOST_cell_1115 ( .a(n_33274), .b(n_32944), .o(TIMEBOOST_net_172) );
no02s01 TIMEBOOST_cell_6955 ( .a(FE_OCP_RBN2661_n_9304), .b(FE_OCP_RBN6635_n_9304), .o(TIMEBOOST_net_2236) );
no02s03 g776311 ( .a(n_4703), .b(FE_OCPN3572_n_4374), .o(n_4814) );
in01s02 g776312 ( .a(n_4616), .o(n_4617) );
no02s04 g776313 ( .a(n_4552), .b(FE_OCP_RBN2920_n_3878), .o(n_4616) );
na02s02 g776314 ( .a(n_4552), .b(FE_OCP_RBN2920_n_3878), .o(n_4626) );
in01s01 g776315 ( .a(n_4507), .o(n_4508) );
na02s02 g776316 ( .a(n_4429), .b(n_4316), .o(n_4507) );
no02s02 g776317 ( .a(n_4429), .b(FE_OCP_RBN6774_n_4046), .o(n_4550) );
in01s01 g776318 ( .a(n_4811), .o(n_4812) );
no02f04 g776319 ( .a(n_4771), .b(n_4310), .o(n_4811) );
in01s01 g776320 ( .a(n_4846), .o(n_4847) );
na02s02 g776321 ( .a(n_4771), .b(n_4171), .o(n_4846) );
no02m04 g776322 ( .a(n_4766), .b(n_4765), .o(n_4767) );
no02s02 g776323 ( .a(n_4762), .b(n_4761), .o(n_4919) );
na02s01 g776324 ( .a(n_4786), .b(n_4756), .o(n_4757) );
no02s01 g776325 ( .a(n_4766), .b(FE_OCPN4546_n_4727), .o(n_5156) );
in01s01 g776326 ( .a(n_4823), .o(n_4824) );
na02s02 g776327 ( .a(n_4762), .b(n_4761), .o(n_4823) );
na03f02 TIMEBOOST_cell_7252 ( .a(n_9970), .b(n_9927), .c(n_9963), .o(TIMEBOOST_net_2149) );
in01s01 g776329 ( .a(n_4931), .o(n_4932) );
no02m02 g776330 ( .a(n_4809), .b(n_3717), .o(n_4931) );
na02s01 g776331 ( .a(n_4827), .b(n_4780), .o(n_4781) );
no02s01 g776333 ( .a(n_4918), .b(n_4774), .o(n_5053) );
in01s01 g776334 ( .a(n_4319), .o(n_4320) );
no02m04 g776335 ( .a(n_4197), .b(n_4065), .o(n_4319) );
in01s01 g776336 ( .a(n_4949), .o(n_4950) );
no02s03 g776337 ( .a(n_4810), .b(n_3715), .o(n_4949) );
in01m02 g776338 ( .a(n_4667), .o(n_4668) );
na02f04 g776339 ( .a(n_4560), .b(n_4548), .o(n_4667) );
in01m02 g776342 ( .a(n_4880), .o(n_4881) );
na02s04 g776343 ( .a(n_4750), .b(n_4672), .o(n_4880) );
na02m02 TIMEBOOST_cell_8023 ( .a(TIMEBOOST_net_2642), .b(n_16424), .o(TIMEBOOST_net_1759) );
na02s02 g776346 ( .a(n_4494), .b(n_4398), .o(n_4565) );
no02m08 g776348 ( .a(n_4517), .b(n_4422), .o(n_4592) );
no02s06 g776349 ( .a(n_4347), .b(n_3106), .o(n_4568) );
no02s02 g776351 ( .a(n_4543), .b(n_4465), .o(n_4560) );
no02m04 g776352 ( .a(n_4346), .b(n_4093), .o(n_4475) );
in01s01 g776353 ( .a(n_4703), .o(n_4704) );
na02f04 g776354 ( .a(n_4634), .b(n_4186), .o(n_4703) );
in01s01 g776355 ( .a(n_4680), .o(n_4681) );
no02s02 g776356 ( .a(n_4634), .b(n_4222), .o(n_4680) );
in01s02 g776357 ( .a(n_4496), .o(n_4497) );
no02s02 g776358 ( .a(n_4549), .b(n_4428), .o(n_4496) );
in01s01 g776359 ( .a(n_4595), .o(n_4596) );
na02s02 g776360 ( .a(n_4546), .b(n_4625), .o(n_4595) );
na02m04 g776361 ( .a(n_4661), .b(n_4172), .o(n_4771) );
in01s01 g776362 ( .a(n_4714), .o(n_4715) );
na02s02 g776363 ( .a(n_4579), .b(n_4659), .o(n_4714) );
na02s02 g776365 ( .a(n_47007), .b(n_4662), .o(n_4727) );
in01s01 g776367 ( .a(n_4774), .o(n_4821) );
no02s03 g776368 ( .a(n_4720), .b(n_4719), .o(n_4774) );
no02s01 g776369 ( .a(n_4735), .b(n_4650), .o(n_4890) );
na02s02 g776370 ( .a(n_4661), .b(n_4267), .o(n_4664) );
no02f02 g776371 ( .a(n_47007), .b(n_4662), .o(n_4766) );
no02s01 g776372 ( .a(n_4689), .b(n_4765), .o(n_5058) );
na02s02 g776373 ( .a(n_4646), .b(FE_OCP_RBN5811_n_3645), .o(n_4750) );
in01s01 g776374 ( .a(n_4787), .o(n_4918) );
na02s02 g776375 ( .a(n_4720), .b(n_4719), .o(n_4787) );
no02s01 g776376 ( .a(n_4799), .b(n_4674), .o(n_4929) );
na02s02 g776378 ( .a(n_4671), .b(FE_OCP_RBN2850_n_3645), .o(n_4672) );
oa12f06 g776379 ( .a(n_4106), .b(n_4608), .c(n_4170), .o(n_4697) );
in01m02 g776380 ( .a(n_4635), .o(n_4636) );
in01f02 g776381 ( .a(n_4604), .o(n_4635) );
na02s10 TIMEBOOST_cell_4212 ( .a(n_32928), .b(TIMEBOOST_net_1196), .o(n_33015) );
in01s01 TIMEBOOST_cell_8890 ( .a(n_1189), .o(TIMEBOOST_net_2934) );
in01s01 g776384 ( .a(n_4271), .o(n_4272) );
in01s01 g776385 ( .a(n_4197), .o(n_4271) );
ao12m04 g776386 ( .a(n_3841), .b(n_4054), .c(n_3928), .o(n_4197) );
oa12m04 g776387 ( .a(n_4501), .b(n_4619), .c(n_4382), .o(n_4786) );
no02s01 TIMEBOOST_cell_5466 ( .a(FE_OCP_RBN4462_n_44267), .b(n_21413), .o(TIMEBOOST_net_1681) );
in01m01 g776390 ( .a(n_4323), .o(n_4363) );
ao12m04 g776391 ( .a(n_4019), .b(n_4154), .c(n_4149), .o(n_4323) );
oa12s01 g776392 ( .a(n_4615), .b(n_4614), .c(n_4619), .o(n_4679) );
in01s01 g776399 ( .a(n_4466), .o(n_4467) );
in01s01 g776400 ( .a(n_4396), .o(n_4466) );
in01s01 g776401 ( .a(n_4396), .o(n_4388) );
ao12f04 g776403 ( .a(n_4589), .b(n_4710), .c(n_4492), .o(n_4827) );
in01s01 g776404 ( .a(n_4809), .o(n_4810) );
na03s02 TIMEBOOST_cell_6571 ( .a(n_11107), .b(n_11106), .c(n_11159), .o(n_11178) );
oa12s01 g776406 ( .a(n_4562), .b(n_4608), .c(n_4561), .o(n_4631) );
na02s04 TIMEBOOST_cell_918 ( .a(TIMEBOOST_net_73), .b(n_46413), .o(n_32714) );
oa12s01 g776410 ( .a(n_4709), .b(n_4708), .c(n_4710), .o(n_4793) );
in01s02 g776411 ( .a(n_4472), .o(n_4473) );
na02s02 TIMEBOOST_cell_2930 ( .a(n_18787), .b(n_18706), .o(TIMEBOOST_net_756) );
na02s01 g776416 ( .a(n_4608), .b(n_4561), .o(n_4562) );
no02s02 TIMEBOOST_cell_3045 ( .a(TIMEBOOST_net_813), .b(n_3681), .o(n_3812) );
na02s04 g776418 ( .a(n_4358), .b(n_4457), .o(n_4543) );
no02s06 g776420 ( .a(n_4343), .b(n_4093), .o(n_4403) );
in01s01 g776421 ( .a(n_4494), .o(n_4495) );
na02s02 g776422 ( .a(n_4366), .b(n_4457), .o(n_4494) );
in01s01 g776424 ( .a(n_4397), .o(n_4468) );
na02s06 g776425 ( .a(n_4343), .b(n_4093), .o(n_4397) );
no02s01 TIMEBOOST_cell_8478 ( .a(n_37136), .b(n_37190), .o(TIMEBOOST_net_2726) );
no02m06 TIMEBOOST_cell_2929 ( .a(TIMEBOOST_net_755), .b(n_29240), .o(n_29477) );
na02s03 g776428 ( .a(n_4585), .b(n_4198), .o(n_4641) );
no02s01 TIMEBOOST_cell_4483 ( .a(n_4875), .b(n_4759), .o(TIMEBOOST_net_1332) );
no02f04 g776430 ( .a(n_4538), .b(n_4176), .o(n_4634) );
na02s02 g776431 ( .a(n_4538), .b(n_4254), .o(n_4539) );
in01s01 TIMEBOOST_cell_8913 ( .a(TIMEBOOST_net_2956), .o(TIMEBOOST_net_2957) );
no02s03 g776433 ( .a(n_4266), .b(FE_OCP_RBN6775_n_4046), .o(n_4428) );
no02s02 g776434 ( .a(n_4265), .b(FE_OCP_RBN6774_n_4046), .o(n_4549) );
na02s02 g776435 ( .a(FE_OCP_RBN4345_n_4378), .b(FE_OCP_RBN6767_n_3704), .o(n_4546) );
na02s02 g776436 ( .a(n_4378), .b(FE_OCP_RBN2920_n_3878), .o(n_4625) );
na02s02 TIMEBOOST_cell_3993 ( .a(n_2502), .b(n_2898), .o(TIMEBOOST_net_1087) );
no02m02 g776438 ( .a(n_4103), .b(n_4007), .o(n_4161) );
na03s08 TIMEBOOST_cell_917 ( .a(FE_OCPN1902_n_32712), .b(n_32709), .c(FE_OCP_RBN3984_n_32791), .o(TIMEBOOST_net_73) );
no02s02 g776440 ( .a(n_4485), .b(n_3563), .o(n_4765) );
na02s01 g776441 ( .a(n_4529), .b(n_4528), .o(n_4659) );
in01s01 g776442 ( .a(n_4689), .o(n_4644) );
no02s02 g776443 ( .a(n_4486), .b(FE_OCPN6921_n_3580), .o(n_4689) );
in01s01 g776444 ( .a(n_4578), .o(n_4579) );
no02s02 g776445 ( .a(n_4529), .b(n_4528), .o(n_4578) );
no02s02 g776446 ( .a(n_4588), .b(n_4587), .o(n_4735) );
no02s02 g776447 ( .a(n_4643), .b(n_4642), .o(n_4799) );
na02s01 g776448 ( .a(n_4614), .b(n_4619), .o(n_4615) );
no02s02 g776449 ( .a(n_4178), .b(n_4202), .o(n_4324) );
na02s01 g776450 ( .a(n_4708), .b(n_4710), .o(n_4709) );
in01s01 g776451 ( .a(n_4649), .o(n_4650) );
na02s02 g776452 ( .a(n_4588), .b(n_4587), .o(n_4649) );
na02s02 g776453 ( .a(n_4542), .b(FE_OCP_RBN2850_n_3645), .o(n_4591) );
in01s02 g776454 ( .a(n_4753), .o(n_4754) );
na02m02 g776455 ( .a(n_4688), .b(n_4542), .o(n_4753) );
in01s01 g776456 ( .a(n_4673), .o(n_4674) );
na02s02 g776457 ( .a(n_4643), .b(n_4642), .o(n_4673) );
na02s02 g776458 ( .a(n_4464), .b(n_4327), .o(n_4465) );
in01s02 g776459 ( .a(n_4346), .o(n_4347) );
oa22m04 g776460 ( .a(n_4158), .b(FE_OFN4765_n_3029), .c(FE_OCP_RBN5929_n_4158), .d(n_4093), .o(n_4346) );
na02m04 g776462 ( .a(n_4502), .b(n_4230), .o(n_4661) );
na02m06 g776463 ( .a(n_4325), .b(n_4242), .o(n_4517) );
na02m04 TIMEBOOST_cell_934 ( .a(TIMEBOOST_net_81), .b(n_32721), .o(n_32792) );
in01s01 g776465 ( .a(n_4671), .o(n_4646) );
na02s03 g776466 ( .a(n_4443), .b(n_4511), .o(n_4671) );
in01s01 g776468 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_1_), .o(n_6698) );
in01s01 g776472 ( .a(n_4398), .o(n_4399) );
na02s02 g776473 ( .a(n_4385), .b(n_4358), .o(n_4398) );
na02s02 g776474 ( .a(n_4392), .b(n_4317), .o(n_4511) );
na02s02 g776475 ( .a(n_4391), .b(n_4318), .o(n_4443) );
in01s01 g776476 ( .a(n_4422), .o(n_4423) );
no02m04 g776477 ( .a(n_4234), .b(n_3837), .o(n_4422) );
na02s02 g776478 ( .a(n_4313), .b(n_3297), .o(n_4464) );
in01s01 g776480 ( .a(n_4366), .o(n_4405) );
na02s02 g776481 ( .a(n_4252), .b(n_3106), .o(n_4366) );
na02m04 g776482 ( .a(n_4314), .b(FE_OFN4765_n_3029), .o(n_4547) );
na02s02 g776483 ( .a(n_4253), .b(n_3082), .o(n_4457) );
na02m04 g776484 ( .a(n_4233), .b(FE_OCP_RBN6762_n_3790), .o(n_4325) );
na02m04 g776486 ( .a(FE_OCP_RBN3044_n_4449), .b(n_4174), .o(n_4585) );
no02s01 TIMEBOOST_cell_8491 ( .a(TIMEBOOST_net_2732), .b(n_37474), .o(n_37542) );
no02s01 TIMEBOOST_cell_8463 ( .a(TIMEBOOST_net_2718), .b(n_32441), .o(n_32535) );
na02m04 g776490 ( .a(n_4425), .b(n_4393), .o(n_4490) );
no02s02 g776491 ( .a(n_4487), .b(n_4350), .o(n_4488) );
na02m04 TIMEBOOST_cell_933 ( .a(FE_RN_224_0), .b(FE_OCP_RBN2423_n_32554), .o(TIMEBOOST_net_81) );
in01s01 g776493 ( .a(n_4476), .o(n_4477) );
na02s01 g776494 ( .a(n_4447), .b(n_4351), .o(n_4476) );
na02s04 g776495 ( .a(n_4449), .b(n_4128), .o(n_4502) );
in01s01 g776496 ( .a(n_4538), .o(n_4525) );
na02s02 TIMEBOOST_cell_6322 ( .a(TIMEBOOST_net_2012), .b(n_16977), .o(n_17130) );
in01s01 g776498 ( .a(n_4441), .o(n_4442) );
na02s02 g776499 ( .a(n_4322), .b(n_4393), .o(n_4441) );
in01s01 g776500 ( .a(n_4544), .o(n_4688) );
no02m04 g776501 ( .a(n_4479), .b(FE_OCP_RBN2808_n_3338), .o(n_4544) );
no02s01 g776502 ( .a(n_4481), .b(n_4582), .o(n_4756) );
oa12s02 g776503 ( .a(n_2927), .b(n_4131), .c(n_4073), .o(n_4132) );
na03s02 TIMEBOOST_cell_7349 ( .a(n_2873), .b(n_2679), .c(n_2890), .o(n_3024) );
in01s01 g776505 ( .a(n_4532), .o(n_4533) );
na02s02 g776506 ( .a(n_4474), .b(FE_OCP_RBN6806_n_4411), .o(n_4532) );
na02s01 g776507 ( .a(n_4483), .b(n_4594), .o(n_4780) );
in01s01 g776510 ( .a(n_4542), .o(n_4601) );
na02s03 g776511 ( .a(n_4479), .b(FE_OCP_RBN2808_n_3338), .o(n_4542) );
oa12f06 g776512 ( .a(n_4090), .b(n_4432), .c(n_3990), .o(n_4608) );
na02m06 TIMEBOOST_cell_6693 ( .a(n_34459), .b(n_34491), .o(TIMEBOOST_net_2104) );
in01s01 g776514 ( .a(n_4103), .o(n_4104) );
in01s01 g776515 ( .a(n_4054), .o(n_4103) );
oa12f04 g776516 ( .a(n_3782), .b(n_3896), .c(n_3692), .o(n_4054) );
no02s01 TIMEBOOST_cell_3042 ( .a(n_24053), .b(n_24039), .o(TIMEBOOST_net_812) );
oa12m04 g776518 ( .a(n_4334), .b(n_4572), .c(n_4446), .o(n_4619) );
in01s01 g776519 ( .a(FE_OCP_RBN2987_n_4238), .o(n_5422) );
ao12m04 g776524 ( .a(n_4331), .b(n_4553), .c(n_4404), .o(n_4710) );
in01s01 g776525 ( .a(n_4177), .o(n_4178) );
in01s01 g776526 ( .a(n_4154), .o(n_4177) );
oa12s04 g776527 ( .a(n_3873), .b(n_3992), .c(n_3983), .o(n_4154) );
oa12s01 g776528 ( .a(n_4519), .b(n_4518), .c(n_4553), .o(n_4590) );
na02s01 TIMEBOOST_cell_4494 ( .a(TIMEBOOST_net_1337), .b(n_5953), .o(n_6047) );
oa22s06 g776530 ( .a(n_4101), .b(FE_OFN4765_n_3029), .c(FE_OCP_RBN5917_n_4101), .d(n_3862), .o(n_4343) );
no02s01 TIMEBOOST_cell_8546 ( .a(FE_OCP_RBN6612_n_2289), .b(n_2674), .o(TIMEBOOST_net_2760) );
in01s01 g776535 ( .a(n_4485), .o(n_4486) );
ao22s02 g776536 ( .a(n_4302), .b(n_4146), .c(n_4303), .d(n_4145), .o(n_4485) );
oa12s01 g776537 ( .a(n_4574), .b(n_4573), .c(n_4572), .o(n_4623) );
oa22m02 g776542 ( .a(n_47012), .b(FE_OCP_RBN6774_n_4046), .c(FE_OCP_RBN5957_n_47012), .d(FE_OCP_RBN6776_n_4046), .o(n_4378) );
in01s02 g776543 ( .a(n_4265), .o(n_4266) );
oa12s01 g776545 ( .a(n_4420), .b(n_4432), .c(n_4419), .o(n_4526) );
in01s01 g776546 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_4_), .o(n_6761) );
na02s01 g776548 ( .a(n_4432), .b(n_4419), .o(n_4420) );
in01s01 TIMEBOOST_cell_5905 ( .a(FE_OFN1_n_43918), .o(TIMEBOOST_net_1794) );
na02s02 TIMEBOOST_cell_4186 ( .a(n_27620), .b(TIMEBOOST_net_1183), .o(FE_RN_347_0) );
na02f08 TIMEBOOST_cell_5373 ( .a(TIMEBOOST_net_1634), .b(n_26025), .o(n_26176) );
in01s01 g776552 ( .a(n_4317), .o(n_4318) );
na02s02 g776553 ( .a(n_4112), .b(n_4167), .o(n_4317) );
no03s02 TIMEBOOST_cell_8175 ( .a(FE_RN_765_0), .b(FE_RN_764_0), .c(n_11707), .o(FE_RN_767_0) );
na02s02 g776555 ( .a(n_4307), .b(n_3297), .o(n_4327) );
no02m04 TIMEBOOST_cell_3275 ( .a(n_16541), .b(TIMEBOOST_net_928), .o(n_16632) );
no02m04 TIMEBOOST_cell_6325 ( .a(FE_OCP_RBN4408_n_26394), .b(n_26555), .o(TIMEBOOST_net_2014) );
na02s04 g776558 ( .a(n_4387), .b(n_4273), .o(n_4487) );
in01m02 g776559 ( .a(n_4424), .o(n_4425) );
na02m04 g776560 ( .a(n_4286), .b(n_4345), .o(n_4424) );
in01s01 g776561 ( .a(n_4515), .o(n_4516) );
na02s01 g776562 ( .a(FE_OCPN3571_n_4374), .b(n_4387), .o(n_4515) );
na02s02 g776564 ( .a(n_4287), .b(n_4286), .o(n_4348) );
na02s02 g776566 ( .a(n_4355), .b(n_4210), .o(n_4407) );
na02s01 g776567 ( .a(n_4283), .b(FE_OCP_RBN5870_n_3704), .o(n_4447) );
na02s04 g776568 ( .a(n_4225), .b(FE_OCP_RBN6778_n_4046), .o(n_4393) );
in01s01 g776569 ( .a(n_4350), .o(n_4351) );
no02m02 g776570 ( .a(n_4283), .b(FE_OCP_RBN5870_n_3704), .o(n_4350) );
in01s01 g776571 ( .a(n_4321), .o(n_4322) );
no02s02 g776572 ( .a(n_4225), .b(n_4046), .o(n_4321) );
no02m04 g776574 ( .a(n_4389), .b(n_3959), .o(n_4449) );
in01s01 g776575 ( .a(n_4480), .o(n_4481) );
na02s02 g776576 ( .a(n_4434), .b(n_4433), .o(n_4480) );
na02s02 g776577 ( .a(n_4360), .b(FE_OCP_RBN5787_n_3421), .o(n_4474) );
no02s02 g776579 ( .a(n_4360), .b(FE_OCP_RBN5787_n_3421), .o(n_4411) );
no02m04 TIMEBOOST_cell_7687 ( .a(TIMEBOOST_net_2474), .b(n_8587), .o(n_8732) );
no03f08 TIMEBOOST_cell_4680 ( .a(n_19277), .b(TIMEBOOST_net_824), .c(n_19213), .o(n_19358) );
na02s01 g776582 ( .a(n_4573), .b(n_4572), .o(n_4574) );
in01s01 g776583 ( .a(n_4451), .o(n_4452) );
no02s02 g776584 ( .a(n_4557), .b(FE_OCP_RBN3042_n_4296), .o(n_4451) );
no02s02 g776585 ( .a(n_4051), .b(n_4032), .o(n_4125) );
no02s01 g776587 ( .a(n_4589), .b(n_4493), .o(n_4708) );
no02s02 g776589 ( .a(n_4434), .b(n_4433), .o(n_4582) );
na02s01 g776590 ( .a(n_4383), .b(n_4501), .o(n_4614) );
na02s01 g776591 ( .a(n_4518), .b(n_4553), .o(n_4519) );
in01s01 g776592 ( .a(n_4482), .o(n_4483) );
no02s02 g776593 ( .a(n_4438), .b(n_4437), .o(n_4482) );
na02s02 TIMEBOOST_cell_5408 ( .a(n_3867), .b(FE_OCP_RBN5869_n_3704), .o(TIMEBOOST_net_1652) );
na02s03 g776595 ( .a(n_4438), .b(n_4437), .o(n_4594) );
na02s02 g776597 ( .a(n_4484), .b(n_4395), .o(n_4563) );
na02s06 g776598 ( .a(n_4218), .b(n_4092), .o(n_4385) );
in01s01 g776599 ( .a(n_4391), .o(n_4392) );
na03m08 TIMEBOOST_cell_8297 ( .a(n_14751), .b(FE_OCP_RBN5853_n_14750), .c(n_14678), .o(n_14829) );
in01s02 g776601 ( .a(n_4233), .o(n_4234) );
no02m06 g776602 ( .a(n_4111), .b(n_4091), .o(n_4233) );
no02s04 g776603 ( .a(n_4129), .b(n_4166), .o(n_4242) );
na02s02 TIMEBOOST_cell_6321 ( .a(FE_OCP_RBN3179_n_16088), .b(n_16943), .o(TIMEBOOST_net_2012) );
in01s01 g776605 ( .a(n_4430), .o(n_4431) );
na02s02 g776606 ( .a(n_4389), .b(n_4122), .o(n_4430) );
oa12s01 g776607 ( .a(n_4500), .b(n_4499), .c(n_4498), .o(n_4600) );
na02f04 TIMEBOOST_cell_8734 ( .a(n_18717), .b(n_18277), .o(TIMEBOOST_net_2854) );
oa12s01 g776609 ( .a(n_4402), .b(n_4401), .c(n_4400), .o(n_4491) );
in01s01 g776610 ( .a(FE_OCP_RBN2950_n_4158), .o(n_5009) );
in01s01 g776614 ( .a(n_4252), .o(n_4253) );
no02s04 TIMEBOOST_cell_2852 ( .a(n_37311), .b(n_37154), .o(TIMEBOOST_net_717) );
in01m02 g776616 ( .a(n_4313), .o(n_4314) );
na03s02 TIMEBOOST_cell_8426 ( .a(FE_OCP_RBN6874_n_31520), .b(FE_OCP_RBN3231_n_31107), .c(n_31721), .o(n_31827) );
na02m04 TIMEBOOST_cell_3081 ( .a(TIMEBOOST_net_831), .b(n_8213), .o(n_8243) );
na02s03 g776620 ( .a(n_4012), .b(n_3082), .o(n_4358) );
in01s01 g776621 ( .a(n_4111), .o(n_4112) );
no02m04 g776622 ( .a(n_3963), .b(n_3082), .o(n_4111) );
no02s01 TIMEBOOST_cell_4200 ( .a(TIMEBOOST_net_1190), .b(n_37172), .o(n_37821) );
na02f04 TIMEBOOST_cell_2851 ( .a(n_37369), .b(TIMEBOOST_net_716), .o(n_37401) );
na02s02 g776625 ( .a(n_4011), .b(FE_OFN4765_n_3029), .o(n_4092) );
in01s01 g776626 ( .a(n_4166), .o(n_4167) );
no02s04 g776627 ( .a(n_3964), .b(n_3106), .o(n_4166) );
no02f08 TIMEBOOST_cell_8567 ( .a(TIMEBOOST_net_2770), .b(TIMEBOOST_net_1258), .o(n_14774) );
in01s01 g776629 ( .a(n_4302), .o(n_4303) );
no02s02 g776630 ( .a(n_4235), .b(n_4209), .o(n_4302) );
na02s04 g776631 ( .a(n_4235), .b(n_4208), .o(n_4355) );
na02m03 g776632 ( .a(n_4285), .b(n_4071), .o(n_4389) );
na02s02 g776633 ( .a(n_4082), .b(FE_OCPN4828_FE_OCP_RBN4275_n_3700), .o(n_4287) );
na02s02 g776634 ( .a(n_4300), .b(FE_OCP_RBN6765_n_3704), .o(n_4387) );
in01s01 g776635 ( .a(n_4352), .o(n_4353) );
no02s02 g776636 ( .a(n_4285), .b(n_4121), .o(n_4352) );
na02s02 g776637 ( .a(n_4081), .b(n_4046), .o(n_4286) );
no02s02 g776639 ( .a(n_4300), .b(FE_OCP_RBN6765_n_3704), .o(n_4374) );
na02s01 g776640 ( .a(n_4009), .b(n_3922), .o(n_4078) );
na02s01 g776641 ( .a(n_4401), .b(n_4400), .o(n_4402) );
na02s01 g776642 ( .a(n_4499), .b(n_4498), .o(n_4500) );
na02s02 g776644 ( .a(n_4229), .b(n_4228), .o(n_4296) );
in01s01 g776645 ( .a(n_4492), .o(n_4493) );
na02s04 g776646 ( .a(n_4436), .b(n_4435), .o(n_4492) );
na02s02 g776647 ( .a(n_47009), .b(FE_OCP_RBN2771_n_4336), .o(n_4484) );
no02s03 g776648 ( .a(n_4436), .b(n_4435), .o(n_4589) );
no02s02 g776649 ( .a(n_4229), .b(n_4228), .o(n_4557) );
na02s01 g776650 ( .a(n_4069), .b(FE_OCP_RBN4281_n_3848), .o(n_4163) );
in01s01 g776651 ( .a(n_4382), .o(n_4383) );
no02s02 g776652 ( .a(n_4340), .b(n_4339), .o(n_4382) );
na02s02 g776653 ( .a(n_4340), .b(n_4339), .o(n_4501) );
in01s01 g776654 ( .a(n_4394), .o(n_4395) );
no02s04 g776655 ( .a(n_47009), .b(FE_OCP_RBN2771_n_4336), .o(n_4394) );
no02s04 TIMEBOOST_cell_4257 ( .a(n_29485), .b(n_25859), .o(TIMEBOOST_net_1219) );
oa12f06 g776659 ( .a(n_3997), .b(n_4108), .c(n_4297), .o(n_4432) );
in01s02 g776660 ( .a(n_4131), .o(n_4057) );
na02s06 g776661 ( .a(n_3860), .b(n_2982), .o(n_4131) );
in01s01 g776663 ( .a(n_4218), .o(n_4243) );
na02m04 g776664 ( .a(n_4029), .b(n_4039), .o(n_4218) );
in01s01 g776665 ( .a(n_4305), .o(n_4306) );
ao12s02 g776666 ( .a(n_3970), .b(n_4213), .c(n_4035), .o(n_4305) );
no02m08 TIMEBOOST_cell_6288 ( .a(TIMEBOOST_net_1995), .b(n_10216), .o(n_10375) );
no02f06 TIMEBOOST_cell_8512 ( .a(n_29266), .b(n_29161), .o(TIMEBOOST_net_2743) );
in01s01 g776672 ( .a(n_4050), .o(n_4051) );
in01s01 g776673 ( .a(n_3992), .o(n_4050) );
oa12m04 g776674 ( .a(n_3651), .b(n_3822), .c(n_3749), .o(n_3992) );
in01s01 g776677 ( .a(n_3896), .o(n_3905) );
oa12f04 g776678 ( .a(n_3701), .b(n_3786), .c(n_3648), .o(n_3896) );
oa12s01 g776679 ( .a(n_4270), .b(n_4297), .c(n_4269), .o(n_4380) );
no02s06 TIMEBOOST_cell_3032 ( .a(n_34224), .b(n_34037), .o(TIMEBOOST_net_807) );
in01s02 g776682 ( .a(n_5603), .o(n_3971) );
no02s06 TIMEBOOST_cell_788 ( .a(TIMEBOOST_net_8), .b(n_37097), .o(n_37164) );
na02m03 g776684 ( .a(n_4042), .b(n_3953), .o(n_4225) );
oa22s02 g776685 ( .a(FE_OCP_RBN5857_FE_RN_998_0), .b(n_3106), .c(FE_OCP_RBN5860_FE_RN_998_0), .d(n_3082), .o(n_4307) );
na02s06 g776688 ( .a(n_3858), .b(n_2975), .o(n_3860) );
na02s02 g776689 ( .a(n_3915), .b(n_2962), .o(n_3935) );
no02s01 g776690 ( .a(n_3858), .b(n_3857), .o(n_3859) );
na02m02 TIMEBOOST_cell_4256 ( .a(TIMEBOOST_net_1218), .b(n_29039), .o(n_29097) );
na02s01 g776692 ( .a(n_4297), .b(n_4269), .o(n_4270) );
na02s02 g776693 ( .a(n_4134), .b(n_4083), .o(n_4129) );
na02s04 g776694 ( .a(n_4133), .b(n_3954), .o(n_4091) );
in01s02 g776695 ( .a(n_4220), .o(n_4221) );
na02m02 g776696 ( .a(n_4134), .b(n_4133), .o(n_4220) );
no02s04 g776697 ( .a(n_4256), .b(n_4072), .o(n_4345) );
in01s01 g776698 ( .a(n_4273), .o(n_4274) );
no02s04 g776699 ( .a(n_4115), .b(n_4222), .o(n_4273) );
na02s02 g776700 ( .a(FE_OCP_RBN2991_n_4041), .b(FE_OCP_RBN6765_n_3704), .o(n_3953) );
no02m02 g776701 ( .a(n_4152), .b(n_4025), .o(n_4285) );
in01s01 g776702 ( .a(n_4368), .o(n_4369) );
no02s02 g776703 ( .a(n_4310), .b(n_4256), .o(n_4368) );
na02m02 TIMEBOOST_cell_5441 ( .a(TIMEBOOST_net_1668), .b(n_9893), .o(n_10136) );
na02s02 g776706 ( .a(n_4186), .b(n_4116), .o(n_4245) );
no02s02 TIMEBOOST_cell_5300 ( .a(n_4177), .b(n_4203), .o(TIMEBOOST_net_1598) );
na02s01 g776708 ( .a(n_4041), .b(FE_OCPN4828_FE_OCP_RBN4275_n_3700), .o(n_4042) );
no02s01 g776709 ( .a(n_4335), .b(n_4446), .o(n_4573) );
na02s02 g776710 ( .a(n_4015), .b(FE_OCP_RBN6743_n_3746), .o(n_4068) );
no02s02 g776711 ( .a(n_3731), .b(n_3728), .o(n_3838) );
na02s06 TIMEBOOST_cell_3031 ( .a(TIMEBOOST_net_806), .b(n_2528), .o(n_2638) );
in01s02 g776715 ( .a(FE_OCP_RBN4294_n_4080), .o(n_5529) );
na02s02 g776718 ( .a(FE_OCP_RBN5858_FE_RN_998_0), .b(n_3872), .o(n_4080) );
na02s02 g776720 ( .a(n_4249), .b(n_4365), .o(n_4416) );
na02s02 g776721 ( .a(n_4075), .b(n_4088), .o(n_4247) );
no02s01 TIMEBOOST_cell_8515 ( .a(TIMEBOOST_net_2744), .b(n_38087), .o(n_38110) );
no02s01 g776724 ( .a(n_4304), .b(n_4277), .o(n_4401) );
no02s01 g776725 ( .a(n_4330), .b(n_4276), .o(n_4499) );
no02m01 g776726 ( .a(n_3894), .b(n_3792), .o(n_3942) );
no02s06 TIMEBOOST_cell_787 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_21_), .o(TIMEBOOST_net_8) );
na02s01 g776730 ( .a(n_4332), .b(n_4404), .o(n_4518) );
na02s04 g776732 ( .a(n_3956), .b(n_4083), .o(n_4165) );
in01s02 g776734 ( .a(n_3963), .o(n_3964) );
no02m08 TIMEBOOST_cell_7026 ( .a(TIMEBOOST_net_2271), .b(n_16080), .o(n_16172) );
na03m06 TIMEBOOST_cell_8360 ( .a(n_44165), .b(n_38730), .c(n_38793), .o(n_38811) );
na02s02 g776738 ( .a(n_4156), .b(n_4263), .o(n_4264) );
in01s01 g776739 ( .a(n_4081), .o(n_4082) );
na02s01 TIMEBOOST_cell_4373 ( .a(n_15103), .b(n_14439), .o(TIMEBOOST_net_1277) );
na02s06 TIMEBOOST_cell_6310 ( .a(TIMEBOOST_net_2006), .b(FE_OCP_RBN4480_n_11439), .o(n_11698) );
oa12s02 g776742 ( .a(n_3917), .b(n_4028), .c(n_3862), .o(n_4029) );
ao12s02 g776744 ( .a(n_3856), .b(n_4028), .c(n_3862), .o(n_4039) );
na02s02 TIMEBOOST_cell_3030 ( .a(n_2084), .b(n_2085), .o(TIMEBOOST_net_806) );
in01s01 g776746 ( .a(n_4011), .o(n_4012) );
in01s01 g776750 ( .a(n_4009), .o(n_4069) );
in01s01 g776751 ( .a(n_3981), .o(n_4009) );
in01s01 g776752 ( .a(n_3981), .o(n_3982) );
na02s02 g776757 ( .a(n_3830), .b(n_2791), .o(n_3872) );
in01s02 g776768 ( .a(n_3858), .o(n_3915) );
no02s06 g776769 ( .a(n_3737), .b(n_2988), .o(n_3858) );
na02s02 g776771 ( .a(n_4026), .b(n_4000), .o(n_4095) );
na02s02 g776772 ( .a(n_3955), .b(n_3954), .o(n_3956) );
no02s02 TIMEBOOST_cell_5361 ( .a(TIMEBOOST_net_1628), .b(FE_RN_1926_0), .o(n_47011) );
no02m10 TIMEBOOST_cell_3029 ( .a(n_34124), .b(TIMEBOOST_net_805), .o(n_34164) );
na02s04 g776775 ( .a(n_3934), .b(n_3862), .o(n_4134) );
na02s03 g776776 ( .a(n_3933), .b(n_3106), .o(n_4133) );
no02s01 g776777 ( .a(n_4061), .b(n_3967), .o(n_4110) );
no02s02 g776778 ( .a(n_4126), .b(n_3909), .o(n_4179) );
no02s06 TIMEBOOST_cell_7025 ( .a(n_14452), .b(n_16007), .o(TIMEBOOST_net_2271) );
na02s04 TIMEBOOST_cell_6309 ( .a(n_11459), .b(n_11007), .o(TIMEBOOST_net_2006) );
no02s01 TIMEBOOST_cell_4358 ( .a(TIMEBOOST_net_1269), .b(n_20713), .o(n_20714) );
in01s01 g776783 ( .a(n_4115), .o(n_4116) );
no02s02 g776784 ( .a(n_4030), .b(FE_OCP_RBN5870_n_3704), .o(n_4115) );
na02m04 TIMEBOOST_cell_5330 ( .a(n_15853), .b(n_15374), .o(TIMEBOOST_net_1613) );
no02s02 g776786 ( .a(n_4114), .b(n_4046), .o(n_4310) );
na02s02 g776787 ( .a(n_5629), .b(FE_OCPN4828_FE_OCP_RBN4275_n_3700), .o(n_4024) );
no02s03 g776788 ( .a(n_4113), .b(FE_OCPN4828_FE_OCP_RBN4275_n_3700), .o(n_4256) );
na02s01 g776789 ( .a(n_4030), .b(FE_OCP_RBN5870_n_3704), .o(n_4186) );
in01s01 g776790 ( .a(n_4331), .o(n_4332) );
no02s02 g776791 ( .a(n_47010), .b(n_4231), .o(n_4331) );
na02s03 g776792 ( .a(n_4212), .b(FE_OCP_RBN5731_n_4211), .o(n_4365) );
in01s01 g776793 ( .a(n_4329), .o(n_4330) );
na02s02 g776794 ( .a(n_4169), .b(n_2584), .o(n_4329) );
in01m01 g776795 ( .a(n_4248), .o(n_4249) );
no02s06 g776796 ( .a(n_4212), .b(FE_OCP_RBN5731_n_4211), .o(n_4248) );
no02s02 g776797 ( .a(n_4281), .b(n_4280), .o(n_4446) );
na02s02 g776798 ( .a(n_47010), .b(n_4231), .o(n_4404) );
na02s02 g776799 ( .a(n_4155), .b(n_4175), .o(n_4156) );
in01s01 g776800 ( .a(n_4236), .o(n_4237) );
na02s02 g776801 ( .a(n_4263), .b(n_4155), .o(n_4236) );
no02s02 g776802 ( .a(n_4099), .b(n_2531), .o(n_4277) );
in01s01 g776803 ( .a(n_4334), .o(n_4335) );
na02s02 g776804 ( .a(n_4281), .b(n_4280), .o(n_4334) );
no02s02 g776805 ( .a(n_4100), .b(n_2532), .o(n_4304) );
in01s01 g776806 ( .a(n_4275), .o(n_4276) );
na02s04 g776807 ( .a(n_4168), .b(n_2583), .o(n_4275) );
no02s01 TIMEBOOST_cell_6831 ( .a(n_30757), .b(n_30729), .o(TIMEBOOST_net_2173) );
ao12f06 g776809 ( .a(n_3815), .b(n_4139), .c(n_3940), .o(n_4297) );
in01s01 g776810 ( .a(n_4015), .o(n_4016) );
in01s02 g776813 ( .a(n_4075), .o(n_4213) );
ao12s04 g776814 ( .a(n_3880), .b(n_3987), .c(n_3943), .o(n_4075) );
in01s01 g776815 ( .a(n_4190), .o(n_4191) );
in01s01 g776816 ( .a(n_4152), .o(n_4190) );
no02s02 TIMEBOOST_cell_3250 ( .a(n_21346), .b(n_45024), .o(TIMEBOOST_net_916) );
oa12s01 g776818 ( .a(n_4085), .b(n_4139), .c(n_4084), .o(n_4192) );
no02s04 TIMEBOOST_cell_6742 ( .a(TIMEBOOST_net_2128), .b(n_38981), .o(TIMEBOOST_net_1584) );
in01s01 g776824 ( .a(n_3822), .o(n_3894) );
oa12s04 g776825 ( .a(n_3586), .b(n_3724), .c(n_3539), .o(n_3822) );
in01s01 g776826 ( .a(n_3786), .o(n_3731) );
oa12m06 g776827 ( .a(n_3568), .b(n_3630), .c(n_3535), .o(n_3786) );
in01s01 g776829 ( .a(n_3737), .o(n_3738) );
oa12s06 g776830 ( .a(n_2874), .b(n_3600), .c(n_2818), .o(n_3737) );
na02s01 g776831 ( .a(n_4139), .b(n_4084), .o(n_4085) );
na02s02 TIMEBOOST_cell_8018 ( .a(n_11236), .b(n_11237), .o(TIMEBOOST_net_2640) );
no02s04 g776833 ( .a(n_3851), .b(n_3754), .o(n_3954) );
in01s01 g776834 ( .a(n_3913), .o(n_3914) );
na02s02 g776835 ( .a(n_3864), .b(n_3863), .o(n_3913) );
no02s02 g776836 ( .a(n_3918), .b(n_3919), .o(n_4083) );
na02s02 g776837 ( .a(n_3855), .b(n_3863), .o(n_3871) );
no02s04 g776839 ( .a(n_3919), .b(n_3851), .o(n_4000) );
na02s01 g776840 ( .a(n_3855), .b(n_3765), .o(n_3856) );
no02s02 g776841 ( .a(n_4058), .b(n_4173), .o(n_4230) );
in01s01 g776842 ( .a(n_4061), .o(n_4062) );
no02s02 g776843 ( .a(n_3987), .b(n_3931), .o(n_4061) );
na02m02 TIMEBOOST_cell_8760 ( .a(n_8238), .b(FE_OCP_RBN6629_n_8269), .o(TIMEBOOST_net_2867) );
in01s01 g776845 ( .a(n_4126), .o(n_4127) );
no02f06 TIMEBOOST_cell_6328 ( .a(TIMEBOOST_net_2015), .b(n_16497), .o(n_16588) );
in01s01 g776847 ( .a(n_4254), .o(n_4255) );
no02s01 g776848 ( .a(n_4176), .b(n_4222), .o(n_4254) );
na02s02 g776850 ( .a(n_4172), .b(n_4171), .o(n_4267) );
oa12s02 g776852 ( .a(n_2948), .b(n_3633), .c(n_2887), .o(n_3830) );
in01s01 g776853 ( .a(n_4202), .o(n_4203) );
na02s02 g776854 ( .a(n_4149), .b(n_4020), .o(n_4202) );
na02s02 g776855 ( .a(n_3744), .b(n_3613), .o(n_3775) );
na02s02 g776856 ( .a(n_3968), .b(FE_OCP_RBN5768_n_3498), .o(n_4155) );
no02s01 g776857 ( .a(n_3656), .b(n_3623), .o(n_3722) );
oa12s02 g776858 ( .a(n_4208), .b(n_4209), .c(n_4037), .o(n_4204) );
na02s02 g776860 ( .a(n_4175), .b(FE_OCP_RBN3025_n_4065), .o(n_4226) );
na02s04 g776862 ( .a(n_3969), .b(FE_OCP_RBN6688_n_3498), .o(n_4263) );
no02s02 TIMEBOOST_cell_6741 ( .a(FE_OCP_RBN5736_n_38569), .b(n_44925), .o(TIMEBOOST_net_2128) );
no02s04 TIMEBOOST_cell_5301 ( .a(TIMEBOOST_net_1598), .b(n_4324), .o(n_4458) );
no02s02 TIMEBOOST_cell_6634 ( .a(TIMEBOOST_net_2074), .b(FE_RN_202_0), .o(n_28534) );
ao12s04 g776867 ( .a(n_3918), .b(n_3955), .c(n_3753), .o(n_4026) );
no02s02 g776868 ( .a(n_3887), .b(n_3847), .o(n_3917) );
ao12s01 g776869 ( .a(n_3975), .b(n_4209), .c(n_4208), .o(n_4210) );
no02s01 TIMEBOOST_cell_5450 ( .a(n_5090), .b(n_5091), .o(TIMEBOOST_net_1673) );
oa12s01 g776871 ( .a(n_4119), .b(n_4118), .c(FE_OFN82_n_4117), .o(n_4180) );
in01s01 g776874 ( .a(FE_OCP_RBN4281_n_3848), .o(n_3922) );
oa22s02 g776878 ( .a(n_3681), .b(n_2918), .c(n_3655), .d(n_2919), .o(n_3848) );
in01s01 g776879 ( .a(n_4099), .o(n_4100) );
in01s02 g776881 ( .a(n_3933), .o(n_3934) );
no02m02 TIMEBOOST_cell_5502 ( .a(n_10993), .b(n_10927), .o(TIMEBOOST_net_1699) );
no02s06 TIMEBOOST_cell_3056 ( .a(FE_OCP_RBN5745_n_24618), .b(n_22207), .o(TIMEBOOST_net_819) );
oa12s01 g776884 ( .a(n_3977), .b(n_3945), .c(n_3944), .o(n_4157) );
in01s02 g776885 ( .a(n_4168), .o(n_4169) );
no02s06 TIMEBOOST_cell_3206 ( .a(n_39586), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(TIMEBOOST_net_894) );
in01s01 g776887 ( .a(n_4113), .o(n_4114) );
no02s02 TIMEBOOST_cell_4341 ( .a(n_7894), .b(n_7941), .o(TIMEBOOST_net_1261) );
na02s04 g776891 ( .a(n_3607), .b(n_3642), .o(n_3867) );
in01s01 g776892 ( .a(n_5629), .o(n_3994) );
na02s01 TIMEBOOST_cell_874 ( .a(TIMEBOOST_net_51), .b(n_37020), .o(n_37136) );
oa22s02 g776899 ( .a(FE_OCP_RBN6742_n_3746), .b(FE_OFN4763_n_3029), .c(n_3746), .d(n_3862), .o(n_4028) );
na03s08 TIMEBOOST_cell_8303 ( .a(n_4439), .b(n_4388), .c(FE_OFN4765_n_3029), .o(n_4652) );
no02f04 TIMEBOOST_cell_8117 ( .a(TIMEBOOST_net_2689), .b(n_20759), .o(n_20872) );
na02f08 TIMEBOOST_cell_4350 ( .a(TIMEBOOST_net_1265), .b(n_42135), .o(n_42147) );
na02f08 TIMEBOOST_cell_3055 ( .a(TIMEBOOST_net_818), .b(FE_RN_19_0), .o(n_20127) );
na02s02 g776905 ( .a(n_3811), .b(FE_OCP_RBN5914_n_3750), .o(n_3847) );
na02s02 g776906 ( .a(n_3811), .b(FE_OCP_RBN2901_n_3643), .o(n_3864) );
na02m06 TIMEBOOST_cell_2921 ( .a(TIMEBOOST_net_751), .b(n_13409), .o(n_13513) );
in01s01 TIMEBOOST_cell_5906 ( .a(TIMEBOOST_net_1794), .o(TIMEBOOST_net_1795) );
no02s06 g776909 ( .a(n_3762), .b(FE_OFN4764_n_3029), .o(n_3919) );
no02s02 g776910 ( .a(n_3761), .b(n_3082), .o(n_3851) );
no02s01 g776911 ( .a(n_3776), .b(n_3862), .o(n_3887) );
na02s02 g776912 ( .a(n_3776), .b(n_3862), .o(n_3855) );
na02s04 g776913 ( .a(n_3778), .b(n_3854), .o(n_3950) );
na02m06 TIMEBOOST_cell_8580 ( .a(n_34996), .b(FE_OCPN1681_n_30614), .o(TIMEBOOST_net_2777) );
na02s02 g776915 ( .a(n_3948), .b(n_3920), .o(n_3949) );
no02s02 TIMEBOOST_cell_5449 ( .a(TIMEBOOST_net_1672), .b(n_5531), .o(TIMEBOOST_net_1324) );
na02s02 g776917 ( .a(n_3884), .b(n_3773), .o(n_3850) );
no02f04 TIMEBOOST_cell_3229 ( .a(TIMEBOOST_net_905), .b(n_20383), .o(n_20510) );
no02s04 g776919 ( .a(n_3852), .b(n_3849), .o(n_3987) );
na02s02 g776920 ( .a(n_3849), .b(n_3979), .o(n_4010) );
no02s02 g776922 ( .a(n_3995), .b(n_4046), .o(n_4176) );
na02m02 TIMEBOOST_cell_8497 ( .a(TIMEBOOST_net_2735), .b(FE_RN_1585_0), .o(FE_RN_1586_0) );
na02s06 TIMEBOOST_cell_4340 ( .a(TIMEBOOST_net_1260), .b(n_8008), .o(n_8136) );
na02s02 g776925 ( .a(n_4014), .b(FE_OCPN4828_FE_OCP_RBN4275_n_3700), .o(n_4172) );
no02s06 g776926 ( .a(n_3996), .b(FE_OCP_RBN5870_n_3704), .o(n_4222) );
no02s02 TIMEBOOST_cell_7545 ( .a(TIMEBOOST_net_2403), .b(n_24164), .o(TIMEBOOST_net_1873) );
in01s01 g776928 ( .a(n_4072), .o(n_4171) );
no02s02 g776929 ( .a(n_4014), .b(FE_OCPN4828_FE_OCP_RBN4275_n_3700), .o(n_4072) );
no02s02 g776930 ( .a(n_3764), .b(n_3710), .o(n_3863) );
no02s02 g776931 ( .a(n_3759), .b(n_3528), .o(n_3821) );
na02s02 g776932 ( .a(n_4023), .b(FE_OCP_RBN5754_n_4022), .o(n_4175) );
in01s01 g776934 ( .a(n_3724), .o(n_3744) );
oa12f04 g776935 ( .a(n_3511), .b(n_3572), .c(n_3459), .o(n_3724) );
no02s04 g776937 ( .a(n_4023), .b(FE_OCP_RBN5754_n_4022), .o(n_4065) );
in01s01 g776938 ( .a(n_4019), .o(n_4020) );
no02m02 g776939 ( .a(n_3973), .b(FE_OCP_RBN5724_n_47022), .o(n_4019) );
na02s01 g776940 ( .a(n_4118), .b(FE_OFN82_n_4117), .o(n_4119) );
na02s02 g776941 ( .a(n_3973), .b(FE_OCP_RBN5724_n_47022), .o(n_4149) );
na02s01 g776942 ( .a(n_3583), .b(n_3509), .o(n_3607) );
na02s02 g776943 ( .a(n_4008), .b(FE_OFN82_n_4117), .o(n_4400) );
in01s01 g776945 ( .a(n_3977), .o(n_4498) );
na02s02 g776946 ( .a(n_3945), .b(n_3944), .o(n_3977) );
na02s02 g776947 ( .a(n_3584), .b(n_3510), .o(n_3642) );
in01s01 g776949 ( .a(n_3630), .o(n_3656) );
na02m08 g776950 ( .a(n_3558), .b(n_3488), .o(n_3630) );
na02s01 TIMEBOOST_cell_873 ( .a(n_37022), .b(n_36916), .o(TIMEBOOST_net_51) );
oa12f06 g776952 ( .a(n_3768), .b(n_3883), .c(n_3985), .o(n_4139) );
in01s01 g776953 ( .a(n_4173), .o(n_4174) );
na02s03 TIMEBOOST_cell_2021 ( .a(n_13954), .b(n_13375), .o(TIMEBOOST_net_625) );
oa12s01 g776955 ( .a(n_3986), .b(n_3985), .c(n_3984), .o(n_4089) );
in01s01 g776956 ( .a(n_3968), .o(n_3969) );
in01s01 g776958 ( .a(n_3681), .o(n_3655) );
in01s01 g776960 ( .a(n_3633), .o(n_3681) );
no02s06 g776962 ( .a(n_3561), .b(n_2797), .o(n_3633) );
na02s01 g776963 ( .a(n_3985), .b(n_3984), .o(n_3986) );
in01s04 g776964 ( .a(n_3955), .o(n_3877) );
na02f06 g776965 ( .a(n_3837), .b(n_3790), .o(n_3955) );
no02s01 g776966 ( .a(n_5356), .b(n_6250), .o(n_5439) );
na02s02 g776967 ( .a(n_3879), .b(n_3840), .o(n_3880) );
na02s02 g776968 ( .a(n_3885), .b(n_3886), .o(n_3891) );
in01s01 g776970 ( .a(n_3849), .o(n_3897) );
na02s04 g776971 ( .a(n_3743), .b(n_3813), .o(n_3849) );
no02s02 g776974 ( .a(n_3760), .b(n_3846), .o(n_3773) );
no02s02 g776975 ( .a(n_3774), .b(n_3846), .o(n_3948) );
na02s02 g776976 ( .a(n_3957), .b(n_4034), .o(n_4209) );
na02s02 g776977 ( .a(n_3941), .b(n_4036), .o(n_4037) );
na02s02 g776978 ( .a(n_5355), .b(n_5356), .o(n_6304) );
no02s01 g776979 ( .a(n_4049), .b(n_4121), .o(n_4122) );
in01s01 g776980 ( .a(n_4087), .o(n_4088) );
na02s01 g776981 ( .a(n_4035), .b(n_4034), .o(n_4087) );
in01s01 g776982 ( .a(n_3966), .o(n_3967) );
na02s02 g776983 ( .a(n_3943), .b(n_3879), .o(n_3966) );
in01s01 g776984 ( .a(n_4044), .o(n_4045) );
na02s01 g776985 ( .a(n_3958), .b(n_3957), .o(n_4044) );
in01s01 g776986 ( .a(n_3979), .o(n_3980) );
no02s02 g776987 ( .a(n_3852), .b(n_3931), .o(n_3979) );
in01s01 g776988 ( .a(n_4147), .o(n_4148) );
na02s01 g776989 ( .a(n_4071), .b(n_4070), .o(n_4147) );
in01s01 g776990 ( .a(n_5403), .o(n_5404) );
na02s01 g776991 ( .a(n_5384), .b(n_5355), .o(n_5403) );
na02s02 g776993 ( .a(n_3885), .b(n_3884), .o(n_3920) );
na02s01 g776995 ( .a(n_3810), .b(n_3886), .o(n_3909) );
in01s01 g776996 ( .a(n_4145), .o(n_4146) );
na02s01 g776997 ( .a(n_4208), .b(n_3941), .o(n_4145) );
na02s02 g776999 ( .a(n_4128), .b(n_4059), .o(n_4198) );
in01s01 g777000 ( .a(n_4143), .o(n_4144) );
na02s01 g777001 ( .a(n_3960), .b(n_4098), .o(n_4143) );
in01s02 g777002 ( .a(n_4096), .o(n_4097) );
no02s03 g777003 ( .a(n_4025), .b(n_4121), .o(n_4096) );
na02s01 g777005 ( .a(n_4063), .b(n_4036), .o(n_4140) );
in01s01 g777006 ( .a(n_4032), .o(n_4033) );
no02s02 g777007 ( .a(n_3983), .b(n_3874), .o(n_4032) );
in01s01 g777008 ( .a(n_4006), .o(n_4007) );
na02s02 g777009 ( .a(FE_OCP_RBN2953_n_3841), .b(n_3928), .o(n_4006) );
ao12s06 g777010 ( .a(n_3592), .b(n_3593), .c(n_3594), .o(n_3600) );
ao12s02 g777011 ( .a(n_2728), .b(n_3635), .c(n_2790), .o(n_3636) );
oa12s01 g777012 ( .a(n_3594), .b(n_3593), .c(n_3592), .o(n_3595) );
in01s01 g777013 ( .a(n_3764), .o(n_3765) );
oa12s02 g777014 ( .a(n_3668), .b(n_3689), .c(FE_OFN4763_n_3029), .o(n_3764) );
ao12s02 g777015 ( .a(n_3659), .b(n_3689), .c(FE_OFN4763_n_3029), .o(n_3811) );
in01s02 g777016 ( .a(n_3853), .o(n_3854) );
na02s02 g777019 ( .a(n_3813), .b(n_3735), .o(n_3875) );
in01s02 g777020 ( .a(n_3995), .o(n_3996) );
oa22m02 g777021 ( .a(n_5447), .b(FE_OCP_RBN5872_n_3700), .c(n_3620), .d(FE_OCP_RBN6772_n_3700), .o(n_3995) );
na02m02 g777022 ( .a(n_3770), .b(n_3802), .o(n_3973) );
oa12m06 g777023 ( .a(n_3431), .b(n_3557), .c(n_3556), .o(n_3558) );
in01s01 g777026 ( .a(n_3583), .o(n_3584) );
ao12s01 g777027 ( .a(n_3556), .b(n_3557), .c(n_3388), .o(n_3583) );
ao22s01 g777028 ( .a(n_3686), .b(FE_OCP_RBN4256_n_3705), .c(n_3687), .d(n_3704), .o(n_3945) );
in01s01 g777029 ( .a(n_4008), .o(n_4118) );
na02f08 TIMEBOOST_cell_6725 ( .a(n_19637), .b(TIMEBOOST_net_292), .o(TIMEBOOST_net_2120) );
na02s02 g777036 ( .a(n_3608), .b(n_3632), .o(n_3746) );
in01s01 g777037 ( .a(n_3758), .o(n_3759) );
no02f04 TIMEBOOST_cell_5289 ( .a(TIMEBOOST_net_1592), .b(n_20881), .o(n_21029) );
ao22s02 g777039 ( .a(FE_OCP_RBN5869_n_3704), .b(n_3609), .c(FE_OCP_RBN5872_n_3700), .d(n_47016), .o(n_4014) );
in01s01 g777040 ( .a(FE_OCP_RBN5862_n_3718), .o(n_4886) );
oa12s01 g777043 ( .a(n_3904), .b(n_3903), .c(delay_sub_ln23_0_unr1_stage2_stallmux_q_0_), .o(n_4031) );
in01s01 g777044 ( .a(n_47015), .o(n_3678) );
na03f06 TIMEBOOST_cell_8258 ( .a(TIMEBOOST_net_2221), .b(n_19806), .c(FE_OCP_RBN5732_n_19806), .o(n_19942) );
na02s06 TIMEBOOST_cell_1974 ( .a(TIMEBOOST_net_601), .b(n_47246), .o(n_18478) );
in01s02 g777048 ( .a(n_3761), .o(n_3762) );
ao12s02 g777051 ( .a(n_2798), .b(n_3484), .c(n_2663), .o(n_3561) );
na02s02 g777052 ( .a(n_3582), .b(n_2848), .o(n_3632) );
na02s01 g777053 ( .a(n_3903), .b(delay_sub_ln23_0_unr1_stage2_stallmux_q_0_), .o(n_3904) );
na02s02 g777054 ( .a(n_3560), .b(n_2847), .o(n_3608) );
na03f06 TIMEBOOST_cell_8273 ( .a(n_19076), .b(n_19153), .c(n_19213), .o(n_19277) );
no02m04 TIMEBOOST_cell_8573 ( .a(TIMEBOOST_net_2773), .b(TIMEBOOST_net_2498), .o(n_4479) );
no02s03 g777057 ( .a(n_3720), .b(FE_OFN4764_n_3029), .o(n_3918) );
in01s01 g777058 ( .a(n_3753), .o(n_3754) );
na02s04 g777059 ( .a(n_3720), .b(FE_OFN4764_n_3029), .o(n_3753) );
no02s01 g777060 ( .a(n_4819), .b(n_4818), .o(n_4820) );
no02s01 g777061 ( .a(n_4973), .b(n_4972), .o(n_4974) );
na02s02 g777062 ( .a(n_5328), .b(n_5387), .o(n_6250) );
no02s01 g777063 ( .a(n_5191), .b(n_5188), .o(n_5356) );
in01s01 g777064 ( .a(n_4034), .o(n_3970) );
na02s02 g777065 ( .a(n_3604), .b(n_3833), .o(n_4034) );
na02s03 g777066 ( .a(n_3882), .b(FE_OCP_RBN2915_n_3878), .o(n_4063) );
na02s02 g777068 ( .a(FE_OCP_RBN6719_n_3604), .b(FE_OCP_RBN5867_n_3661), .o(n_3735) );
in01s01 g777069 ( .a(n_5333), .o(n_5334) );
na02s01 g777070 ( .a(n_5329), .b(n_5328), .o(n_5333) );
in01s01 g777072 ( .a(n_3941), .o(n_3975) );
na02s02 g777073 ( .a(n_3824), .b(FE_OCP_RBN4255_n_3705), .o(n_3941) );
na02s02 g777074 ( .a(n_3638), .b(n_3755), .o(n_3884) );
na02s02 g777075 ( .a(n_3806), .b(FE_OCP_RBN5875_n_3700), .o(n_3957) );
na02s04 g777076 ( .a(n_3825), .b(FE_OCP_RBN5863_n_3705), .o(n_4208) );
na02s02 g777077 ( .a(n_3661), .b(n_3705), .o(n_3813) );
in01s01 g777078 ( .a(n_4070), .o(n_4049) );
na02s02 g777079 ( .a(n_3900), .b(FE_OCP_RBN5868_n_3704), .o(n_4070) );
in01s01 g777081 ( .a(n_3743), .o(n_3799) );
na02s04 g777082 ( .a(n_3677), .b(n_3705), .o(n_3743) );
in01s02 g777083 ( .a(n_3795), .o(n_3885) );
no02s02 g777085 ( .a(n_3755), .b(FE_OCP_RBN6716_n_3604), .o(n_3795) );
na02s02 g777086 ( .a(n_3881), .b(FE_OCP_RBN4255_n_3705), .o(n_4036) );
no02s02 g777087 ( .a(n_3803), .b(n_3698), .o(n_3852) );
na02s02 g777088 ( .a(n_3733), .b(FE_OCP_RBN4256_n_3705), .o(n_3886) );
na02s01 g777089 ( .a(n_3805), .b(n_3704), .o(n_3958) );
no02s01 g777090 ( .a(n_3890), .b(n_3698), .o(n_4025) );
in01m02 g777091 ( .a(n_3926), .o(n_4121) );
na02s01 g777092 ( .a(n_3890), .b(n_3604), .o(n_3926) );
na02s02 g777093 ( .a(n_3751), .b(FE_OCP_RBN6719_n_3604), .o(n_3879) );
na02s01 g777094 ( .a(n_3929), .b(FE_OCP_RBN5868_n_3704), .o(n_4098) );
na02s01 g777095 ( .a(n_3899), .b(FE_OCP_RBN4274_n_3700), .o(n_4071) );
na02s02 g777096 ( .a(n_3832), .b(FE_OCP_RBN5863_n_3705), .o(n_4035) );
na02s01 g777097 ( .a(n_3605), .b(n_4759), .o(n_5355) );
in01s01 g777098 ( .a(n_3809), .o(n_3810) );
no02s02 g777099 ( .a(n_3733), .b(n_3604), .o(n_3809) );
in01s02 g777100 ( .a(n_3778), .o(n_3774) );
in01s02 g777102 ( .a(n_3760), .o(n_3778) );
no02s02 g777103 ( .a(n_3650), .b(n_3604), .o(n_3760) );
na02s03 g777104 ( .a(FE_OCP_RBN4274_n_3700), .b(n_3752), .o(n_3943) );
in01s01 g777105 ( .a(n_5384), .o(n_5341) );
na02s02 g777106 ( .a(n_3606), .b(n_4675), .o(n_5384) );
no02s02 g777107 ( .a(n_3698), .b(n_3666), .o(n_3846) );
no02s01 g777108 ( .a(n_3677), .b(FE_OCP_RBN5868_n_3704), .o(n_3777) );
no02f08 TIMEBOOST_cell_5986 ( .a(TIMEBOOST_net_1844), .b(n_28150), .o(n_28228) );
in01s01 g777110 ( .a(n_3959), .o(n_3960) );
no02s02 g777111 ( .a(n_3929), .b(FE_OCP_RBN5868_n_3704), .o(n_3959) );
na02s01 g777112 ( .a(n_3989), .b(FE_OCP_RBN2915_n_3878), .o(n_4128) );
in01s01 g777113 ( .a(n_4058), .o(n_4059) );
no02s01 g777114 ( .a(n_3989), .b(FE_OCP_RBN2915_n_3878), .o(n_4058) );
in01s01 g777115 ( .a(n_3840), .o(n_3931) );
na02s02 g777116 ( .a(n_3803), .b(n_3604), .o(n_3840) );
no02s04 TIMEBOOST_cell_4332 ( .a(TIMEBOOST_net_1256), .b(n_46417), .o(n_38577) );
no02m03 g777119 ( .a(n_3784), .b(FE_OCPN902_n_47020), .o(n_3841) );
na02s02 g777120 ( .a(n_3670), .b(n_3696), .o(n_3802) );
no02s03 g777122 ( .a(n_3828), .b(FE_OCPN4933_n_47023), .o(n_3983) );
in01m01 g777124 ( .a(n_3873), .o(n_3874) );
na02f03 g777125 ( .a(n_3828), .b(FE_OCPN4933_n_47023), .o(n_3873) );
na02s02 g777126 ( .a(n_3575), .b(n_3460), .o(n_3683) );
na02s02 g777127 ( .a(n_3784), .b(FE_OCPN902_n_47020), .o(n_3928) );
no02m04 g777128 ( .a(n_3547), .b(n_3396), .o(n_3572) );
na02s01 g777129 ( .a(n_3557), .b(n_3444), .o(n_3569) );
na02m02 g777130 ( .a(n_3671), .b(n_3695), .o(n_3770) );
no02f04 g777131 ( .a(n_3767), .b(n_3756), .o(n_3985) );
na02m04 g777133 ( .a(n_3654), .b(n_3679), .o(n_3790) );
na02s01 g777134 ( .a(n_4779), .b(n_4796), .o(n_4871) );
in01s02 g777136 ( .a(n_3780), .o(n_3781) );
no02s03 g777137 ( .a(n_3669), .b(n_3660), .o(n_3780) );
no02f02 g777138 ( .a(n_3725), .b(n_151), .o(n_3767) );
no02s02 g777139 ( .a(n_3659), .b(n_3643), .o(n_3660) );
no02s06 g777141 ( .a(FE_OCP_RBN2901_n_3643), .b(n_3710), .o(n_3750) );
na02s06 g777142 ( .a(n_3629), .b(n_3679), .o(n_3837) );
na02s04 g777143 ( .a(n_3653), .b(n_3570), .o(n_3654) );
na02s02 g777144 ( .a(n_3668), .b(n_3631), .o(n_3669) );
in01s02 g777145 ( .a(n_3695), .o(n_3696) );
na02s02 g777146 ( .a(n_3679), .b(n_3653), .o(n_3695) );
no02s01 g777147 ( .a(n_4721), .b(n_4818), .o(n_4796) );
na02s01 g777148 ( .a(n_5001), .b(n_5069), .o(n_5113) );
na02s01 g777149 ( .a(n_4852), .b(n_4873), .o(n_4874) );
no02s01 g777150 ( .a(n_4773), .b(n_4731), .o(n_4788) );
no02s01 g777151 ( .a(n_4834), .b(n_4901), .o(n_4885) );
in01s01 g777152 ( .a(n_4819), .o(n_4779) );
na02s01 g777153 ( .a(n_4746), .b(n_4745), .o(n_4819) );
na02s01 g777154 ( .a(n_5330), .b(n_5368), .o(n_5331) );
no02s01 g777155 ( .a(n_4863), .b(n_4864), .o(n_4973) );
na02s01 g777156 ( .a(n_5297), .b(n_5298), .o(n_5299) );
no02s01 g777157 ( .a(n_4685), .b(n_4613), .o(n_5294) );
in01s01 g777158 ( .a(n_5258), .o(n_5259) );
na02s01 g777159 ( .a(n_5112), .b(n_5247), .o(n_5258) );
in01s01 g777160 ( .a(n_5328), .o(n_5260) );
na02s01 g777161 ( .a(n_5166), .b(n_4675), .o(n_5328) );
in01s01 g777162 ( .a(n_5385), .o(n_5386) );
na02s01 g777163 ( .a(n_5368), .b(n_5298), .o(n_5385) );
na02s01 g777164 ( .a(n_4862), .b(n_4732), .o(n_5593) );
no02s01 g777165 ( .a(n_4216), .b(n_4292), .o(n_4910) );
na02s01 g777166 ( .a(n_4999), .b(n_4817), .o(n_5862) );
no02s01 g777167 ( .a(n_4901), .b(n_4818), .o(n_5873) );
no02s01 g777168 ( .a(n_4362), .b(n_4576), .o(n_5261) );
na02s01 g777169 ( .a(n_4201), .b(n_4193), .o(n_4695) );
no02s01 g777170 ( .a(n_4504), .b(n_4503), .o(n_5131) );
na02s01 g777171 ( .a(n_5001), .b(n_4884), .o(n_5990) );
no02s01 g777172 ( .a(n_4371), .b(n_4262), .o(n_5079) );
na02s02 g777173 ( .a(n_4426), .b(n_4361), .o(n_4460) );
in01s01 g777174 ( .a(n_5191), .o(n_5329) );
no02s01 g777175 ( .a(n_5166), .b(n_4675), .o(n_5191) );
na02s01 g777176 ( .a(n_4599), .b(n_4739), .o(n_5413) );
na02s01 g777177 ( .a(n_3940), .b(n_3816), .o(n_4084) );
no02s01 g777178 ( .a(n_4622), .b(n_4921), .o(n_5665) );
in01s01 g777179 ( .a(n_5380), .o(n_5381) );
na02s01 g777180 ( .a(n_5330), .b(n_5297), .o(n_5380) );
na02s01 g777181 ( .a(n_4833), .b(n_4722), .o(n_5859) );
in01s01 g777182 ( .a(n_5174), .o(n_5175) );
no02s01 g777183 ( .a(n_5147), .b(n_5090), .o(n_5174) );
no02s01 g777184 ( .a(n_3769), .b(n_3883), .o(n_3984) );
no02s01 g777185 ( .a(n_3998), .b(n_4108), .o(n_4269) );
na02s01 g777186 ( .a(n_3757), .b(n_3726), .o(n_3903) );
no02s01 g777187 ( .a(n_4170), .b(n_4107), .o(n_4561) );
no02s01 g777188 ( .a(n_5006), .b(n_4863), .o(n_5949) );
in01s01 g777189 ( .a(n_5342), .o(n_5343) );
na02s01 g777190 ( .a(n_5187), .b(n_5287), .o(n_5342) );
na02s01 g777191 ( .a(n_4873), .b(n_4745), .o(n_5774) );
na02s01 g777192 ( .a(n_3991), .b(n_4090), .o(n_4419) );
no02s01 g777193 ( .a(n_5548), .b(n_4773), .o(n_5517) );
in01s01 g777194 ( .a(n_5415), .o(n_5416) );
na02s01 g777195 ( .a(n_5189), .b(n_5387), .o(n_5415) );
na02s02 g777197 ( .a(n_3782), .b(n_3693), .o(n_3835) );
in01s01 g777198 ( .a(n_3635), .o(n_3579) );
in01s02 g777199 ( .a(n_3593), .o(n_3635) );
ao12s06 g777200 ( .a(n_2734), .b(n_3492), .c(n_2656), .o(n_3593) );
oa12s01 g777201 ( .a(n_3483), .b(n_3533), .c(n_3532), .o(n_3560) );
na02f04 TIMEBOOST_cell_7000 ( .a(TIMEBOOST_net_2258), .b(FE_OCP_RBN3146_n_10369), .o(n_10537) );
in01s01 g777204 ( .a(n_3677), .o(n_3706) );
in01s01 g777206 ( .a(n_47016), .o(n_3609) );
in01s01 g777211 ( .a(n_3547), .o(n_3575) );
oa12f04 g777212 ( .a(n_3356), .b(n_3507), .c(n_3309), .o(n_3547) );
no02s01 TIMEBOOST_cell_5931 ( .a(n_1367), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(TIMEBOOST_net_1817) );
in01s01 g777214 ( .a(n_3605), .o(n_3606) );
oa12s01 g777215 ( .a(n_3527), .b(n_3526), .c(n_3525), .o(n_3605) );
na02s01 TIMEBOOST_cell_4361 ( .a(n_42459), .b(n_42367), .o(TIMEBOOST_net_1271) );
in01s02 g777218 ( .a(n_47017), .o(n_3591) );
in01s02 g777220 ( .a(n_3824), .o(n_3825) );
in01s01 g777222 ( .a(n_3832), .o(n_3833) );
no02m04 TIMEBOOST_cell_8862 ( .a(n_11403), .b(FE_OCP_RBN3135_n_10274), .o(TIMEBOOST_net_2918) );
oa22s01 g777224 ( .a(n_3564), .b(n_3195), .c(n_3596), .d(n_4761), .o(n_3733) );
in01s01 g777226 ( .a(n_3751), .o(n_3752) );
in01s01 g777228 ( .a(n_3899), .o(n_3900) );
no02s01 TIMEBOOST_cell_5241 ( .a(TIMEBOOST_net_1568), .b(n_35968), .o(n_35969) );
no02s06 g777232 ( .a(n_3417), .b(n_3424), .o(n_3557) );
in01s01 g777235 ( .a(n_3686), .o(n_3687) );
in01s01 g777236 ( .a(n_3650), .o(n_3686) );
na02s02 g777237 ( .a(n_3566), .b(n_3590), .o(n_3650) );
no02f04 TIMEBOOST_cell_8873 ( .a(TIMEBOOST_net_2923), .b(n_26222), .o(n_26358) );
na02s02 TIMEBOOST_cell_6396 ( .a(TIMEBOOST_net_2049), .b(n_27144), .o(n_27273) );
in01s01 g777240 ( .a(n_3805), .o(n_3806) );
ao22s02 g777241 ( .a(FE_OCP_RBN6718_n_3604), .b(n_5178), .c(FE_OCP_RBN6715_n_3604), .d(n_3380), .o(n_3805) );
in01s02 g777242 ( .a(n_5447), .o(n_3620) );
no02s02 TIMEBOOST_cell_5975 ( .a(n_23308), .b(n_23307), .o(TIMEBOOST_net_1839) );
in01s01 g777244 ( .a(n_3881), .o(n_3882) );
oa22s02 g777245 ( .a(n_3704), .b(n_3819), .c(FE_OCP_RBN4255_n_3705), .d(n_3817), .o(n_3881) );
in01s01 g777248 ( .a(n_3616), .o(n_3625) );
in01s02 g777249 ( .a(n_3616), .o(n_3610) );
na02s06 g777250 ( .a(n_3504), .b(n_3518), .o(n_3616) );
na02s02 g777252 ( .a(n_3565), .b(n_3581), .o(n_3666) );
no02m04 TIMEBOOST_cell_8587 ( .a(TIMEBOOST_net_2780), .b(n_9462), .o(n_9621) );
ao22s02 g777255 ( .a(n_47018), .b(FE_OFN4763_n_3029), .c(FE_OCP_RBN5804_n_47018), .d(n_2913), .o(n_3689) );
na02m08 TIMEBOOST_cell_2901 ( .a(n_18758), .b(TIMEBOOST_net_741), .o(n_18951) );
na02s06 g777257 ( .a(n_3533), .b(n_2771), .o(n_3518) );
na02s02 g777258 ( .a(n_3450), .b(n_3483), .o(n_3484) );
na02s02 g777259 ( .a(n_3492), .b(n_2764), .o(n_3493) );
na02s01 g777260 ( .a(n_3485), .b(n_2770), .o(n_3504) );
na02s01 g777262 ( .a(n_3525), .b(n_3526), .o(n_3527) );
no02f03 g777263 ( .a(n_3577), .b(FE_OCP_RBN5811_n_3645), .o(n_3646) );
na02s03 TIMEBOOST_cell_6939 ( .a(n_34350), .b(n_34351), .o(TIMEBOOST_net_2228) );
no02s06 TIMEBOOST_cell_8494 ( .a(n_32897), .b(TIMEBOOST_net_159), .o(TIMEBOOST_net_2734) );
no02f03 g777266 ( .a(n_3543), .b(n_3601), .o(n_3640) );
na02s02 g777267 ( .a(n_3578), .b(n_2913), .o(n_3668) );
na02s04 g777268 ( .a(n_3546), .b(n_2913), .o(n_3653) );
na02s06 g777269 ( .a(n_3545), .b(FE_OFN4764_n_3029), .o(n_3679) );
in01s02 g777270 ( .a(n_3670), .o(n_3671) );
no02s04 g777271 ( .a(n_3629), .b(n_3571), .o(n_3670) );
no02s02 g777272 ( .a(n_3578), .b(n_2913), .o(n_3659) );
na02s01 g777273 ( .a(n_4759), .b(n_3265), .o(n_4873) );
na02s01 g777274 ( .a(FE_OCP_RBN6714_n_3604), .b(n_4953), .o(n_3685) );
in01s01 g777275 ( .a(n_5111), .o(n_5112) );
no02s01 g777276 ( .a(n_5067), .b(n_4875), .o(n_5111) );
no02s01 g777277 ( .a(n_3698), .b(n_3697), .o(n_3699) );
no02s02 g777278 ( .a(n_4316), .b(n_4537), .o(n_4685) );
na02s03 g777279 ( .a(FE_OCP_RBN5870_n_3704), .b(FE_OFN802_n_3911), .o(n_4090) );
in01s01 g777280 ( .a(n_4731), .o(n_4732) );
no02s01 g777281 ( .a(FE_OCP_RBN6778_n_4046), .b(FE_OFN807_n_4686), .o(n_4731) );
in01s01 g777282 ( .a(n_4361), .o(n_4362) );
na02s01 g777283 ( .a(FE_OCP_RBN6765_n_3704), .b(n_4298), .o(n_4361) );
no02s02 g777284 ( .a(FE_OCPN4828_FE_OCP_RBN4275_n_3700), .b(FE_OFN4815_n_4018), .o(n_4170) );
in01s01 g777285 ( .a(n_5091), .o(n_4884) );
no02s01 g777286 ( .a(n_4760), .b(FE_OCPN3584_n_4556), .o(n_5091) );
in01s01 g777287 ( .a(n_3815), .o(n_3816) );
no02m06 g777288 ( .a(FE_OCP_RBN6768_n_3700), .b(FE_OFN800_n_3771), .o(n_3815) );
no02s01 TIMEBOOST_cell_5932 ( .a(TIMEBOOST_net_1817), .b(n_1435), .o(n_1485) );
no02s02 g777290 ( .a(n_4606), .b(n_4632), .o(n_5548) );
no02s01 g777291 ( .a(n_3564), .b(n_4662), .o(n_3612) );
no02s01 g777292 ( .a(n_3604), .b(n_5062), .o(n_3714) );
in01s01 g777293 ( .a(n_5188), .o(n_5189) );
no02s01 g777294 ( .a(n_5165), .b(n_4675), .o(n_5188) );
na02s02 TIMEBOOST_cell_7613 ( .a(TIMEBOOST_net_2437), .b(n_2347), .o(n_2467) );
in01s01 g777296 ( .a(n_4864), .o(n_4817) );
no02s01 g777297 ( .a(n_4777), .b(FE_OCP_RBN2964_n_4046), .o(n_4864) );
in01s01 g777298 ( .a(n_5186), .o(n_5187) );
no02s02 g777299 ( .a(n_5168), .b(n_4675), .o(n_5186) );
na02s01 g777300 ( .a(n_4606), .b(FE_OFN808_n_3264), .o(n_4745) );
in01s01 g777301 ( .a(n_4576), .o(n_4577) );
no02s01 g777302 ( .a(FE_OCP_RBN6778_n_4046), .b(n_4298), .o(n_4576) );
na02s02 g777303 ( .a(n_3564), .b(n_3563), .o(n_3565) );
in01s01 g777304 ( .a(n_4200), .o(n_4201) );
no02s02 g777305 ( .a(FE_OCPN4828_FE_OCP_RBN4275_n_3700), .b(n_4136), .o(n_4200) );
na02s02 g777306 ( .a(n_3562), .b(FE_OCPN6921_n_3580), .o(n_3581) );
in01s01 g777307 ( .a(n_4612), .o(n_4613) );
na02s02 g777308 ( .a(n_4537), .b(FE_OCP_RBN6782_n_4046), .o(n_4612) );
na02s01 g777309 ( .a(n_3470), .b(n_4675), .o(n_5297) );
in01s01 g777310 ( .a(n_4106), .o(n_4107) );
na02s02 g777311 ( .a(FE_OCP_RBN5870_n_3704), .b(FE_OFN4815_n_4018), .o(n_4106) );
no02s02 g777312 ( .a(FE_OCP_RBN5872_n_3700), .b(FE_OFN801_n_3902), .o(n_4108) );
in01s01 g777313 ( .a(n_4215), .o(n_4292) );
na02s01 g777314 ( .a(FE_OCP_RBN5870_n_3704), .b(FE_OFN803_n_4142), .o(n_4215) );
in01s01 g777315 ( .a(n_3756), .o(n_3757) );
no02s03 g777316 ( .a(n_3604), .b(n_2360), .o(n_3756) );
na02s02 g777317 ( .a(n_4316), .b(FE_OFN804_n_4575), .o(n_4739) );
in01s01 g777318 ( .a(n_5001), .o(n_4972) );
na02s01 g777319 ( .a(n_5494), .b(n_4760), .o(n_5001) );
no02f02 TIMEBOOST_cell_4326 ( .a(n_38340), .b(TIMEBOOST_net_1253), .o(n_38418) );
no02s02 g777321 ( .a(FE_OCP_RBN6765_n_3704), .b(n_4207), .o(n_4371) );
na02s01 g777322 ( .a(n_5197), .b(n_4759), .o(n_5368) );
in01s01 g777323 ( .a(n_4598), .o(n_4599) );
no02s02 g777324 ( .a(FE_OCP_RBN6782_n_4046), .b(FE_OFN804_n_4575), .o(n_4598) );
na02s01 TIMEBOOST_cell_4113 ( .a(n_35980), .b(FE_OCP_RBN4910_n_44222), .o(TIMEBOOST_net_1147) );
no02s02 g777326 ( .a(FE_OCP_RBN6774_n_4046), .b(n_4333), .o(n_4504) );
in01s01 g777327 ( .a(n_3768), .o(n_3769) );
na02s02 g777328 ( .a(n_3604), .b(n_3721), .o(n_3768) );
no02s01 g777329 ( .a(n_4675), .b(n_3501), .o(n_4901) );
in01s01 g777330 ( .a(n_4426), .o(n_4503) );
na02s01 g777331 ( .a(n_4316), .b(n_4333), .o(n_4426) );
na02s01 g777332 ( .a(n_3564), .b(n_4587), .o(n_3566) );
na02s04 TIMEBOOST_cell_5433 ( .a(TIMEBOOST_net_1664), .b(n_26216), .o(n_26292) );
in01s01 g777334 ( .a(n_5241), .o(n_5298) );
no02s01 g777335 ( .a(n_5197), .b(n_4759), .o(n_5241) );
no02m04 g777336 ( .a(FE_OCP_RBN4255_n_3705), .b(n_3721), .o(n_3883) );
in01s01 g777337 ( .a(n_4216), .o(n_4217) );
no02s01 g777338 ( .a(FE_OCP_RBN5870_n_3704), .b(FE_OFN803_n_4142), .o(n_4216) );
no02s01 g777339 ( .a(n_4556), .b(n_3500), .o(n_4818) );
in01s01 g777340 ( .a(n_4852), .o(n_4921) );
na02s01 g777341 ( .a(n_4759), .b(n_4597), .o(n_4852) );
in01s01 g777342 ( .a(n_5005), .o(n_5006) );
na02s01 g777343 ( .a(FE_OCPN3584_n_4556), .b(n_4797), .o(n_5005) );
na02s02 g777344 ( .a(n_3562), .b(n_3012), .o(n_3590) );
na02s01 g777345 ( .a(n_5165), .b(n_4675), .o(n_5387) );
in01s01 g777346 ( .a(n_4702), .o(n_4773) );
na02s01 g777347 ( .a(n_4316), .b(n_4632), .o(n_4702) );
in01s01 g777348 ( .a(n_5069), .o(n_5147) );
na02s01 g777349 ( .a(n_4970), .b(n_4759), .o(n_5069) );
in01s01 g777350 ( .a(n_3990), .o(n_3991) );
no02s06 g777351 ( .a(FE_OCPN4828_FE_OCP_RBN4275_n_3700), .b(FE_OFN802_n_3911), .o(n_3990) );
na02s02 g777352 ( .a(n_5168), .b(n_4675), .o(n_5287) );
no02s01 g777353 ( .a(n_4970), .b(n_4759), .o(n_5090) );
na02m06 g777354 ( .a(FE_OCP_RBN5869_n_3704), .b(FE_OFN800_n_3771), .o(n_3940) );
in01s01 g777355 ( .a(n_4622), .o(n_4746) );
no02s01 g777356 ( .a(n_4556), .b(n_4597), .o(n_4622) );
in01s01 g777357 ( .a(n_4999), .o(n_5000) );
na02s01 g777358 ( .a(n_4759), .b(n_4777), .o(n_4999) );
na02s02 g777359 ( .a(FE_OCP_RBN6778_n_4046), .b(FE_OFN807_n_4686), .o(n_4862) );
na02s01 g777360 ( .a(n_3471), .b(n_4759), .o(n_5330) );
in01s01 g777361 ( .a(n_4721), .o(n_4722) );
no02s01 g777362 ( .a(FE_OCPN1663_n_4556), .b(n_4693), .o(n_4721) );
no02s03 TIMEBOOST_cell_4314 ( .a(TIMEBOOST_net_1247), .b(n_2344), .o(n_2430) );
in01s01 g777364 ( .a(n_4833), .o(n_4834) );
na02s01 g777365 ( .a(n_5494), .b(n_4693), .o(n_4833) );
in01s01 g777366 ( .a(n_4193), .o(n_4194) );
na02s01 g777367 ( .a(FE_OCP_RBN6774_n_4046), .b(n_4136), .o(n_4193) );
in01s01 g777368 ( .a(n_3725), .o(n_3726) );
no02f02 g777369 ( .a(n_3638), .b(n_2359), .o(n_3725) );
in01s01 g777370 ( .a(n_3997), .o(n_3998) );
na02s03 g777371 ( .a(FE_OCP_RBN6761_n_3705), .b(FE_OFN801_n_3902), .o(n_3997) );
no02s01 g777372 ( .a(n_4797), .b(n_5494), .o(n_4863) );
in01s01 g777373 ( .a(n_4261), .o(n_4262) );
na02s02 g777374 ( .a(FE_OCP_RBN6778_n_4046), .b(n_4207), .o(n_4261) );
na02s01 g777375 ( .a(n_5067), .b(n_4675), .o(n_5247) );
na02m02 g777376 ( .a(n_3674), .b(n_3673), .o(n_3782) );
in01s02 g777377 ( .a(n_3692), .o(n_3693) );
no02m04 g777378 ( .a(n_3674), .b(n_3673), .o(n_3692) );
no02m01 g777380 ( .a(n_3652), .b(n_3749), .o(n_3792) );
no02s02 g777381 ( .a(n_3475), .b(n_3248), .o(n_3496) );
ao12s04 g777382 ( .a(n_3218), .b(n_3416), .c(n_3179), .o(n_3417) );
no02s01 g777384 ( .a(n_3507), .b(n_3363), .o(n_3508) );
na03s08 TIMEBOOST_cell_2295 ( .a(n_28062), .b(n_28270), .c(n_28271), .o(n_28307) );
na02s04 g777387 ( .a(n_3551), .b(n_3549), .o(n_3643) );
in01s02 g777388 ( .a(n_3631), .o(n_3710) );
ao12s04 g777389 ( .a(n_3548), .b(n_3522), .c(n_3615), .o(n_3631) );
ao12s01 g777390 ( .a(n_3467), .b(n_3466), .c(n_3465), .o(n_5166) );
ao12s04 g777391 ( .a(n_3217), .b(n_3416), .c(n_3199), .o(n_3424) );
no02s01 g777392 ( .a(n_3466), .b(n_3465), .o(n_3467) );
in01m02 g777393 ( .a(n_3576), .o(n_3577) );
no02s04 g777394 ( .a(n_3549), .b(n_3548), .o(n_3576) );
no02s06 g777395 ( .a(n_3519), .b(n_3573), .o(n_3629) );
in01s02 g777396 ( .a(n_3601), .o(n_3602) );
no02m06 g777397 ( .a(n_3559), .b(n_3573), .o(n_3601) );
na02s02 g777398 ( .a(n_3521), .b(FE_OCP_RBN2629_n_2737), .o(n_3551) );
in01s02 g777399 ( .a(n_3570), .o(n_3571) );
no02s04 g777400 ( .a(n_3559), .b(n_3478), .o(n_3570) );
no02m02 g777401 ( .a(n_3627), .b(n_3626), .o(n_3749) );
in01m01 g777402 ( .a(n_3651), .o(n_3652) );
na02m03 g777403 ( .a(n_3627), .b(n_3626), .o(n_3651) );
in01s01 g777404 ( .a(n_3727), .o(n_3728) );
na02s02 g777405 ( .a(n_3649), .b(n_3701), .o(n_3727) );
in01s02 g777406 ( .a(n_3485), .o(n_3533) );
in01s02 g777408 ( .a(n_3450), .o(n_3485) );
ao12s02 g777409 ( .a(n_2601), .b(n_3386), .c(n_2666), .o(n_3450) );
ao12m06 g777411 ( .a(n_2631), .b(n_3400), .c(n_2658), .o(n_3492) );
ao12s01 g777412 ( .a(n_2937), .b(n_3456), .c(n_2877), .o(n_3526) );
in01s02 g777413 ( .a(n_3564), .o(n_3639) );
in01m06 g777422 ( .a(n_3596), .o(n_3705) );
in01m04 g777423 ( .a(n_3564), .o(n_3596) );
in01s06 g777459 ( .a(n_3564), .o(n_3604) );
in01s06 g777460 ( .a(FE_OCP_RBN6717_n_3604), .o(n_3704) );
in01s06 g777487 ( .a(FE_OCP_RBN6777_n_4046), .o(n_4316) );
in01s03 g777506 ( .a(n_4556), .o(n_4875) );
in01s01 g777514 ( .a(n_4675), .o(n_5494) );
in01s10 g777539 ( .a(n_4759), .o(n_4675) );
in01s10 g777544 ( .a(n_4606), .o(n_4759) );
in01s10 g777545 ( .a(n_4556), .o(n_4606) );
in01s10 g777550 ( .a(FE_OCP_RBN2962_n_4046), .o(n_4556) );
in01s10 g777567 ( .a(FE_OCP_RBN5872_n_3700), .o(n_4046) );
in01m08 g777582 ( .a(n_3698), .o(n_3700) );
in01s08 g777583 ( .a(n_3638), .o(n_3698) );
in01f08 g777586 ( .a(n_3562), .o(n_3638) );
in01f08 g777587 ( .a(n_3564), .o(n_3562) );
in01s01 g777590 ( .a(n_3507), .o(n_3477) );
oa12f04 g777591 ( .a(n_3165), .b(n_3414), .c(n_3123), .o(n_3507) );
no02s02 g777593 ( .a(n_3394), .b(n_3151), .o(n_3475) );
in01s02 g777594 ( .a(n_3817), .o(n_3819) );
na02s03 g777595 ( .a(n_3415), .b(n_3452), .o(n_3817) );
in01s01 g777601 ( .a(n_5242), .o(n_3472) );
na02s02 g777602 ( .a(n_3395), .b(n_3387), .o(n_5242) );
in01s02 g777603 ( .a(n_3545), .o(n_3546) );
na02m04 TIMEBOOST_cell_2920 ( .a(n_12847), .b(n_12848), .o(TIMEBOOST_net_751) );
in01m02 g777605 ( .a(n_4528), .o(n_3641) );
na02s02 TIMEBOOST_cell_5286 ( .a(n_3457), .b(FE_OCP_RBN5820_n_3396), .o(TIMEBOOST_net_1591) );
na02m02 TIMEBOOST_cell_4363 ( .a(n_15394), .b(n_15267), .o(TIMEBOOST_net_1272) );
ao12s01 g777608 ( .a(n_3449), .b(n_3456), .c(n_3448), .o(n_5165) );
oa22s02 g777609 ( .a(FE_OCP_RBN2851_n_4905), .b(n_2913), .c(n_4905), .d(FE_OFN4763_n_3029), .o(n_3578) );
no02s01 g777611 ( .a(FE_OCP_RBN4213_n_3386), .b(n_2695), .o(n_3412) );
no03f06 TIMEBOOST_cell_7170 ( .a(n_24360), .b(n_24288), .c(TIMEBOOST_net_316), .o(n_24484) );
no02s02 TIMEBOOST_cell_2917 ( .a(TIMEBOOST_net_749), .b(n_18931), .o(FE_RN_858_0) );
no02s01 g777615 ( .a(n_3456), .b(n_3448), .o(n_3449) );
na02s01 g777616 ( .a(n_3505), .b(FE_OCP_RBN5771_n_3338), .o(n_3530) );
na02s01 TIMEBOOST_cell_4362 ( .a(TIMEBOOST_net_1271), .b(n_42503), .o(n_42504) );
in01m02 g777618 ( .a(n_3542), .o(n_3543) );
na02m04 g777619 ( .a(n_3519), .b(n_3479), .o(n_3542) );
na02s01 TIMEBOOST_cell_2919 ( .a(TIMEBOOST_net_750), .b(n_38022), .o(n_38094) );
no02s06 g777621 ( .a(n_3482), .b(n_2913), .o(n_3573) );
na02f06 TIMEBOOST_cell_6086 ( .a(TIMEBOOST_net_1894), .b(n_24985), .o(n_25095) );
no02s04 g777623 ( .a(n_3481), .b(FE_OCP_RBN2629_n_2737), .o(n_3559) );
na02s02 g777624 ( .a(n_3389), .b(n_3190), .o(n_3452) );
na02s02 g777626 ( .a(n_3586), .b(FE_OCP_RBN2880_n_3539), .o(n_3613) );
na02s01 g777627 ( .a(n_3372), .b(n_3211), .o(n_3387) );
na02s01 g777628 ( .a(n_3393), .b(n_3210), .o(n_3395) );
na02m01 g777629 ( .a(n_3414), .b(n_3191), .o(n_3415) );
na02s06 g777630 ( .a(n_3334), .b(n_3200), .o(n_3416) );
in01m01 g777631 ( .a(n_3648), .o(n_3649) );
no02s04 g777632 ( .a(n_3598), .b(n_3597), .o(n_3648) );
na02s03 g777633 ( .a(n_3598), .b(n_3597), .o(n_3701) );
no02s01 g777634 ( .a(n_3393), .b(n_3154), .o(n_3394) );
oa12s01 g777635 ( .a(n_2954), .b(n_3423), .c(FE_RN_889_0), .o(n_3466) );
no02s04 g777636 ( .a(n_3429), .b(n_3474), .o(n_3549) );
na02s04 g777637 ( .a(n_3433), .b(n_3473), .o(n_3548) );
in01s01 g777638 ( .a(n_3470), .o(n_3471) );
ao12s01 g777639 ( .a(n_3398), .b(n_3423), .c(n_3397), .o(n_3470) );
na02f02 g777640 ( .a(n_3538), .b(n_3499), .o(n_3627) );
oa12s01 g777641 ( .a(n_3491), .b(n_3490), .c(n_3489), .o(n_5067) );
in01s02 g777642 ( .a(n_3521), .o(n_3522) );
ao22s02 g777643 ( .a(n_3645), .b(n_2913), .c(FE_OCP_RBN5809_n_3645), .d(FE_OFN4764_n_3029), .o(n_3521) );
in01s01 g777644 ( .a(n_3418), .o(n_3419) );
in01s01 g777645 ( .a(n_3400), .o(n_3418) );
oa12m06 g777646 ( .a(n_2569), .b(n_3320), .c(n_2499), .o(n_3400) );
na02s01 g777647 ( .a(n_3490), .b(n_3489), .o(n_3491) );
na02f02 g777648 ( .a(FE_OCP_RBN2863_n_3468), .b(FE_OCP_RBN5767_n_3498), .o(n_3538) );
na02s02 g777649 ( .a(n_3468), .b(FE_OCP_RBN6688_n_3498), .o(n_3499) );
no02s01 g777650 ( .a(n_3397), .b(n_3423), .o(n_3398) );
in01s01 g777651 ( .a(n_3505), .o(n_3506) );
na02s02 g777652 ( .a(n_3474), .b(n_3473), .o(n_3505) );
na02s02 g777653 ( .a(n_3428), .b(n_2913), .o(n_3433) );
no02s02 g777654 ( .a(n_3428), .b(n_2913), .o(n_3429) );
in01s01 g777655 ( .a(n_3623), .o(n_3624) );
na02s02 g777656 ( .a(n_3568), .b(n_3536), .o(n_3623) );
in01s01 g777657 ( .a(n_3528), .o(n_3529) );
na02s01 g777658 ( .a(n_3511), .b(n_3458), .o(n_3528) );
no02m02 g777660 ( .a(n_3495), .b(FE_OCP_RBN4167_n_3494), .o(n_3539) );
na02s04 g777661 ( .a(n_3458), .b(n_3457), .o(n_3459) );
na02s02 g777662 ( .a(n_3495), .b(FE_OCP_RBN4167_n_3494), .o(n_3586) );
ao12m04 g777665 ( .a(n_2541), .b(n_3313), .c(n_2582), .o(n_3386) );
na02f04 g777667 ( .a(n_3447), .b(n_3408), .o(n_3519) );
in01s02 g777668 ( .a(n_3478), .o(n_3479) );
oa12s04 g777669 ( .a(n_3368), .b(n_3407), .c(FE_OCP_RBN2629_n_2737), .o(n_3478) );
in01s01 g777670 ( .a(n_3414), .o(n_3389) );
no02s04 g777671 ( .a(n_3357), .b(n_3346), .o(n_3414) );
na02s01 TIMEBOOST_cell_4353 ( .a(FE_OCP_RBN6791_n_20242), .b(n_20124), .o(TIMEBOOST_net_1267) );
in01s02 g777676 ( .a(n_3481), .o(n_3482) );
no02s06 TIMEBOOST_cell_2060 ( .a(TIMEBOOST_net_644), .b(n_24272), .o(n_24372) );
in01s01 g777680 ( .a(n_5109), .o(n_3381) );
na02s01 TIMEBOOST_cell_3835 ( .a(FE_RN_782_0), .b(n_45685), .o(TIMEBOOST_net_1008) );
in01s02 g777682 ( .a(n_47019), .o(n_3439) );
in01s01 g777684 ( .a(n_3372), .o(n_3393) );
in01s01 g777685 ( .a(n_3334), .o(n_3372) );
oa12f06 g777686 ( .a(n_3102), .b(n_3303), .c(n_3140), .o(n_3334) );
oa12s01 g777687 ( .a(n_3355), .b(n_3354), .c(n_3353), .o(n_5197) );
no02s03 g777688 ( .a(n_3332), .b(n_2640), .o(n_3377) );
na02m06 TIMEBOOST_cell_2063 ( .a(n_34328), .b(FE_RN_2251_0), .o(TIMEBOOST_net_646) );
no02f02 TIMEBOOST_cell_8521 ( .a(TIMEBOOST_net_2747), .b(n_24155), .o(n_24259) );
no02s02 TIMEBOOST_cell_5355 ( .a(TIMEBOOST_net_1625), .b(FE_OCP_RBN4372_n_5048), .o(n_5093) );
no02m04 g777693 ( .a(n_3447), .b(n_3369), .o(n_3468) );
na02s01 g777694 ( .a(n_2880), .b(n_3365), .o(n_3423) );
na02s02 g777695 ( .a(n_3407), .b(FE_OCP_RBN2629_n_2737), .o(n_3408) );
na02s02 g777696 ( .a(n_3503), .b(n_3502), .o(n_3568) );
in01s01 g777697 ( .a(n_3535), .o(n_3536) );
no02s04 g777698 ( .a(n_3503), .b(n_3502), .o(n_3535) );
na02s03 g777699 ( .a(n_3403), .b(n_3006), .o(n_3458) );
no02s01 g777700 ( .a(n_3303), .b(n_3172), .o(n_3304) );
na02s04 g777701 ( .a(n_3404), .b(n_2978), .o(n_3511) );
no02f06 TIMEBOOST_cell_2118 ( .a(TIMEBOOST_net_673), .b(n_9934), .o(n_10030) );
na02s01 g777703 ( .a(n_3353), .b(n_3354), .o(n_3355) );
no02s02 g777704 ( .a(n_3340), .b(n_3152), .o(n_3360) );
ao12m02 g777706 ( .a(n_3126), .b(n_3345), .c(n_3059), .o(n_3346) );
ao12s01 g777707 ( .a(n_2803), .b(n_3367), .c(n_2745), .o(n_3490) );
na02m04 g777709 ( .a(n_3413), .b(n_3384), .o(n_3474) );
ao12s02 g777710 ( .a(n_3383), .b(n_3335), .c(n_2913), .o(n_3473) );
ao12s01 g777711 ( .a(n_3352), .b(n_3367), .c(n_3351), .o(n_4970) );
ao12m02 g777712 ( .a(n_3125), .b(n_3345), .c(n_3329), .o(n_3357) );
ao12s01 g777714 ( .a(n_3315), .b(n_3326), .c(n_3314), .o(n_5168) );
ao12s01 g777715 ( .a(n_3436), .b(n_3435), .c(n_3434), .o(n_4760) );
na02s04 g777717 ( .a(n_3337), .b(n_3358), .o(n_3645) );
no02s02 TIMEBOOST_cell_4161 ( .a(n_31809), .b(n_31854), .o(TIMEBOOST_net_1171) );
in01s02 g777719 ( .a(n_3331), .o(n_3332) );
in01m01 g777720 ( .a(n_3313), .o(n_3331) );
ao12m04 g777721 ( .a(n_2546), .b(n_3246), .c(n_2522), .o(n_3313) );
na02s02 g777722 ( .a(n_3324), .b(n_2567), .o(n_3358) );
na02s01 g777723 ( .a(n_3296), .b(n_2566), .o(n_3337) );
no02m04 g777725 ( .a(n_3413), .b(n_3383), .o(n_3437) );
no02s01 g777726 ( .a(n_3367), .b(n_3351), .o(n_3352) );
no02s01 g777727 ( .a(n_3434), .b(n_3435), .o(n_3436) );
no02s01 g777728 ( .a(n_3326), .b(n_3314), .o(n_3315) );
na02s01 g777729 ( .a(n_3338), .b(FE_OCP_RBN2629_n_2737), .o(n_3339) );
na02s02 g777730 ( .a(n_3336), .b(FE_OCP_RBN2629_n_2737), .o(n_3384) );
no02f04 TIMEBOOST_cell_4160 ( .a(TIMEBOOST_net_1170), .b(n_26666), .o(n_26748) );
in01s01 g777732 ( .a(n_3509), .o(n_3510) );
na02s01 g777733 ( .a(n_3426), .b(n_3488), .o(n_3509) );
no02s06 g777734 ( .a(n_3425), .b(n_3406), .o(n_3431) );
na02s02 g777736 ( .a(FE_OCP_RBN5820_n_3396), .b(n_3457), .o(n_3460) );
ao12m06 g777737 ( .a(FE_OCPN4533_n_3319), .b(n_3318), .c(FE_OCPN3562_n_3317), .o(n_3320) );
oa12s02 g777739 ( .a(FE_OCPN3562_n_3317), .b(n_3318), .c(n_3319), .o(n_3343) );
no02f04 g777740 ( .a(n_3405), .b(n_3349), .o(n_3447) );
oa12s01 g777741 ( .a(n_2909), .b(n_3291), .c(n_2838), .o(n_3354) );
in01s01 g777743 ( .a(n_3403), .o(n_3404) );
no02s04 TIMEBOOST_cell_8872 ( .a(FE_OCP_RBN4388_n_26173), .b(n_23398), .o(TIMEBOOST_net_2923) );
ao12s01 g777745 ( .a(n_3282), .b(n_3281), .c(n_3280), .o(n_4693) );
in01s01 g777746 ( .a(n_3303), .o(n_3279) );
in01s02 g777748 ( .a(n_5178), .o(n_3380) );
na02s03 g777749 ( .a(n_3294), .b(n_3322), .o(n_5178) );
ao12s01 g777750 ( .a(n_3455), .b(n_3454), .c(n_3453), .o(n_4777) );
in01m02 g777751 ( .a(n_4228), .o(n_3385) );
no02m06 g777752 ( .a(n_3316), .b(n_3298), .o(n_4228) );
no02f06 TIMEBOOST_cell_6224 ( .a(TIMEBOOST_net_1963), .b(n_16077), .o(n_16218) );
ao12s01 g777754 ( .a(n_3307), .b(n_3306), .c(n_3305), .o(n_4797) );
ao12s02 g777756 ( .a(n_3043), .b(n_3293), .c(n_3329), .o(n_3340) );
in01s01 g777757 ( .a(n_3500), .o(n_3501) );
ao12s01 g777758 ( .a(n_3411), .b(n_3410), .c(n_3409), .o(n_3500) );
in01s01 g777759 ( .a(n_5062), .o(n_3323) );
na02s01 g777760 ( .a(n_3254), .b(n_3233), .o(n_5062) );
no02s04 g777761 ( .a(n_3312), .b(n_3333), .o(n_3407) );
no02s02 g777762 ( .a(n_3318), .b(n_2485), .o(n_3298) );
no02m04 g777763 ( .a(n_3270), .b(n_2486), .o(n_3316) );
no02s01 g777764 ( .a(n_3410), .b(n_3409), .o(n_3411) );
no02s01 g777765 ( .a(n_3454), .b(n_3453), .o(n_3455) );
no02m04 TIMEBOOST_cell_6223 ( .a(n_16000), .b(n_15984), .o(TIMEBOOST_net_1963) );
na02s02 g777767 ( .a(n_3375), .b(FE_OCP_RBN5729_n_4211), .o(n_3376) );
no02s01 g777768 ( .a(n_3281), .b(n_3280), .o(n_3282) );
na02f08 g777769 ( .a(n_3291), .b(n_2840), .o(n_3326) );
na02m01 TIMEBOOST_cell_4282 ( .a(TIMEBOOST_net_1231), .b(n_13924), .o(n_14023) );
no02s01 TIMEBOOST_cell_6899 ( .a(n_18737), .b(n_18765), .o(TIMEBOOST_net_2208) );
in01s02 g777772 ( .a(n_3368), .o(n_3369) );
na02m04 g777773 ( .a(n_3347), .b(n_2913), .o(n_3368) );
no02m04 g777774 ( .a(n_3347), .b(n_2913), .o(n_3349) );
no02s02 g777775 ( .a(n_3498), .b(FE_OCP_RBN2629_n_2737), .o(n_3312) );
no02s04 g777776 ( .a(FE_OCP_RBN6686_n_3498), .b(n_2913), .o(n_3333) );
no02s01 g777777 ( .a(n_3306), .b(n_3305), .o(n_3307) );
no02m02 g777779 ( .a(n_3379), .b(FE_OCP_RBN5644_n_2674), .o(n_3396) );
na02s01 g777780 ( .a(n_3232), .b(n_3130), .o(n_3233) );
na02m02 g777781 ( .a(n_3379), .b(FE_OCP_RBN5644_n_2674), .o(n_3457) );
in01s01 g777782 ( .a(n_3425), .o(n_3426) );
no02s03 g777783 ( .a(n_3391), .b(FE_OCP_RBN4164_n_3390), .o(n_3425) );
na02s04 g777784 ( .a(n_3255), .b(n_3101), .o(n_3345) );
na02m02 g777785 ( .a(n_3391), .b(FE_OCP_RBN4164_n_3390), .o(n_3488) );
na02s02 g777786 ( .a(n_3293), .b(n_3105), .o(n_3294) );
no02s01 g777788 ( .a(n_3406), .b(n_3556), .o(n_3444) );
na02s01 g777789 ( .a(n_3255), .b(n_3104), .o(n_3322) );
na02s01 g777790 ( .a(n_3202), .b(n_3131), .o(n_3254) );
oa12s02 g777791 ( .a(n_3245), .b(FE_OCP_RBN2769_n_3238), .c(n_3286), .o(n_3296) );
no02f10 TIMEBOOST_cell_3095 ( .a(n_29744), .b(TIMEBOOST_net_838), .o(n_29800) );
no02m04 g777793 ( .a(n_3375), .b(n_3308), .o(n_3413) );
ao12s01 g777794 ( .a(n_2821), .b(n_3225), .c(n_2730), .o(n_3367) );
in01m01 g777795 ( .a(n_3405), .o(n_3373) );
no02f04 g777796 ( .a(n_3328), .b(n_3321), .o(n_3405) );
ao12s01 g777797 ( .a(n_2687), .b(n_3227), .c(n_2701), .o(n_3435) );
na02s01 TIMEBOOST_cell_4178 ( .a(TIMEBOOST_net_1179), .b(n_36327), .o(n_36412) );
in01s02 g777800 ( .a(n_3335), .o(n_3336) );
na02s02 g777801 ( .a(n_3285), .b(n_3257), .o(n_3335) );
na02s10 TIMEBOOST_cell_3256 ( .a(n_43287), .b(n_43530), .o(TIMEBOOST_net_919) );
no02s01 TIMEBOOST_cell_6061 ( .a(n_29157), .b(n_29364), .o(TIMEBOOST_net_1882) );
no03s02 TIMEBOOST_cell_6793 ( .a(n_4044), .b(n_4305), .c(n_4045), .o(TIMEBOOST_net_2154) );
na02m06 g777805 ( .a(n_3222), .b(n_3245), .o(n_3246) );
na02s01 g777806 ( .a(n_3224), .b(n_2735), .o(n_3306) );
no02s02 g777807 ( .a(FE_OCP_RBN2796_n_3250), .b(n_2913), .o(n_3308) );
na02s02 g777808 ( .a(FE_OCP_RBN5740_n_4336), .b(n_2913), .o(n_3285) );
na02s02 g777809 ( .a(n_4336), .b(FE_OCP_RBN2629_n_2737), .o(n_3257) );
no02s02 g777810 ( .a(n_3250), .b(FE_OCP_RBN2630_n_2737), .o(n_3383) );
no02s03 g777811 ( .a(n_3362), .b(FE_OCPN1620_n_3361), .o(n_3556) );
in01s02 g777812 ( .a(n_3388), .o(n_3406) );
na02s04 g777813 ( .a(n_3362), .b(FE_OCPN1620_n_3361), .o(n_3388) );
in01s01 g777814 ( .a(n_3318), .o(n_3270) );
oa12s01 g777816 ( .a(n_2710), .b(n_3212), .c(n_2651), .o(n_3410) );
in01s01 g777817 ( .a(n_3375), .o(n_3370) );
na02m08 TIMEBOOST_cell_6810 ( .a(TIMEBOOST_net_2162), .b(n_5669), .o(n_5818) );
no03s04 TIMEBOOST_cell_8260 ( .a(FE_OCP_RBN2706_n_47023), .b(FE_OCP_RBN5658_n_2438), .c(n_3037), .o(n_3142) );
ao12s01 g777820 ( .a(n_3229), .b(n_3228), .c(n_2712), .o(n_3281) );
in01s01 g777821 ( .a(n_3299), .o(n_3300) );
oa12m02 g777822 ( .a(n_3243), .b(n_3239), .c(n_3241), .o(n_3299) );
oa12m02 g777824 ( .a(n_3242), .b(FE_OCP_RBN2627_n_2737), .c(n_3260), .o(n_3321) );
no02m08 TIMEBOOST_cell_2110 ( .a(n_16223), .b(TIMEBOOST_net_669), .o(n_16398) );
na02s01 TIMEBOOST_cell_4281 ( .a(n_13442), .b(n_13471), .o(TIMEBOOST_net_1231) );
in01s01 g777827 ( .a(n_3697), .o(n_3663) );
oa22s01 g777828 ( .a(n_3192), .b(n_3004), .c(n_3236), .d(n_3005), .o(n_3697) );
in01s01 g777830 ( .a(n_3255), .o(n_3293) );
ao12m04 g777831 ( .a(n_2922), .b(n_3236), .c(n_2977), .o(n_3255) );
no02s02 TIMEBOOST_cell_6679 ( .a(TIMEBOOST_net_1509), .b(n_3981), .o(TIMEBOOST_net_2097) );
no02m02 TIMEBOOST_cell_4325 ( .a(n_38164), .b(n_38220), .o(TIMEBOOST_net_1253) );
in01s01 g777835 ( .a(FE_OFN808_n_3264), .o(n_3265) );
oa22s01 g777836 ( .a(n_3186), .b(n_2733), .c(n_3228), .d(n_2732), .o(n_3264) );
in01s01 g777837 ( .a(n_3232), .o(n_3202) );
ao12m04 g777838 ( .a(n_2964), .b(n_3176), .c(n_2999), .o(n_3232) );
in01s01 g777839 ( .a(n_4953), .o(n_3258) );
no02m06 TIMEBOOST_cell_7812 ( .a(TIMEBOOST_net_2146), .b(n_24656), .o(TIMEBOOST_net_2537) );
oa22s04 g777841 ( .a(n_4022), .b(n_2913), .c(FE_OCP_RBN5752_n_4022), .d(FE_OCP_RBN2627_n_2737), .o(n_3347) );
no02f04 TIMEBOOST_cell_6377 ( .a(n_21078), .b(n_21039), .o(TIMEBOOST_net_2040) );
no02m01 g777843 ( .a(n_3204), .b(n_2425), .o(n_3205) );
no02s04 TIMEBOOST_cell_2109 ( .a(n_16146), .b(FE_OCPN1733_n_14524), .o(TIMEBOOST_net_669) );
no02m08 TIMEBOOST_cell_5273 ( .a(TIMEBOOST_net_1584), .b(n_39157), .o(n_39253) );
na02s08 TIMEBOOST_cell_4280 ( .a(TIMEBOOST_net_1230), .b(n_13924), .o(n_14021) );
no02s02 g777848 ( .a(n_3272), .b(FE_OCP_RBN5723_n_47022), .o(n_3302) );
na02s04 TIMEBOOST_cell_8828 ( .a(n_4355), .b(n_4063), .o(TIMEBOOST_net_2901) );
no02m04 TIMEBOOST_cell_5178 ( .a(n_29672), .b(n_45758), .o(TIMEBOOST_net_1537) );
no02s01 g777851 ( .a(n_3176), .b(n_3027), .o(n_3177) );
in01s01 g777852 ( .a(n_3363), .o(n_3364) );
na02s02 g777853 ( .a(n_3356), .b(n_3310), .o(n_3363) );
in01s02 g777855 ( .a(n_3222), .o(n_3238) );
oa12m06 g777856 ( .a(n_2413), .b(n_3120), .c(n_2367), .o(n_3222) );
no02s02 TIMEBOOST_cell_1912 ( .a(TIMEBOOST_net_570), .b(n_22313), .o(n_22420) );
in01s01 g777859 ( .a(n_3224), .o(n_3225) );
in01s01 g777860 ( .a(n_3227), .o(n_3224) );
no02s06 TIMEBOOST_cell_5971 ( .a(n_40816), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_13_), .o(TIMEBOOST_net_1837) );
oa12s02 g777864 ( .a(n_3196), .b(n_3215), .c(FE_OCP_RBN2627_n_2737), .o(n_3271) );
no02s01 TIMEBOOST_cell_5318 ( .a(n_35842), .b(FE_OCP_RBN3299_n_35539), .o(TIMEBOOST_net_1607) );
ao12s01 g777866 ( .a(n_3158), .b(n_3157), .c(n_3156), .o(n_4597) );
ao22s02 g777868 ( .a(n_4211), .b(n_2913), .c(FE_OCP_RBN5729_n_4211), .d(FE_OCP_RBN2630_n_2737), .o(n_3250) );
no02s02 g777869 ( .a(n_3133), .b(n_2450), .o(n_3141) );
no02s06 TIMEBOOST_cell_2055 ( .a(n_30191), .b(n_29473), .o(TIMEBOOST_net_642) );
no02s01 g777871 ( .a(n_3157), .b(n_3156), .o(n_3158) );
na02s02 g777872 ( .a(n_3220), .b(n_47023), .o(n_3263) );
na02s02 g777873 ( .a(n_3185), .b(n_3243), .o(n_3244) );
na02s02 TIMEBOOST_cell_5317 ( .a(TIMEBOOST_net_1606), .b(n_43110), .o(n_43190) );
na02m04 TIMEBOOST_cell_4278 ( .a(TIMEBOOST_net_1229), .b(n_33765), .o(n_33888) );
no02s02 g777876 ( .a(n_3241), .b(n_3161), .o(n_3242) );
in01s01 g777877 ( .a(n_3228), .o(n_3186) );
in01s01 g777878 ( .a(n_3212), .o(n_3228) );
na02m08 g777879 ( .a(n_3112), .b(n_2736), .o(n_3212) );
in01s02 g777881 ( .a(n_3239), .o(n_3261) );
na02f04 g777882 ( .a(n_3174), .b(n_45190), .o(n_3239) );
na02m02 g777883 ( .a(n_3275), .b(n_3274), .o(n_3356) );
in01s01 g777884 ( .a(n_3309), .o(n_3310) );
no02m03 g777885 ( .a(n_3275), .b(n_3274), .o(n_3309) );
in01s01 g777886 ( .a(n_3204), .o(n_3198) );
oa12m06 g777887 ( .a(n_2271), .b(n_3147), .c(n_2313), .o(n_3204) );
in01s01 g777888 ( .a(n_47341), .o(n_3240) );
in01s01 g777890 ( .a(n_4761), .o(n_3195) );
na02s01 g777891 ( .a(n_3117), .b(n_3115), .o(n_4761) );
in01s01 g777892 ( .a(n_3272), .o(n_3273) );
na02s01 TIMEBOOST_cell_8589 ( .a(TIMEBOOST_net_2781), .b(n_29869), .o(n_29954) );
in01s01 g777894 ( .a(n_3236), .o(n_3192) );
ao12f04 g777895 ( .a(n_2902), .b(n_3149), .c(n_2956), .o(n_3236) );
na02s06 g777897 ( .a(n_3164), .b(n_3148), .o(n_4022) );
in01s01 g777898 ( .a(n_3176), .o(n_3135) );
ao12m04 g777899 ( .a(n_2907), .b(n_3114), .c(n_2963), .o(n_3176) );
in01s01 g777900 ( .a(n_3259), .o(n_3260) );
na02s02 g777902 ( .a(n_3119), .b(n_2329), .o(n_3164) );
na02s02 g777903 ( .a(n_3147), .b(n_2328), .o(n_3148) );
na02s04 g777905 ( .a(FE_OCP_RBN2768_n_3167), .b(n_3216), .o(n_3220) );
na02s02 g777906 ( .a(n_3189), .b(FE_OCP_RBN5657_n_2438), .o(n_3243) );
no02m02 g777907 ( .a(n_3189), .b(FE_OCP_RBN5656_n_2438), .o(n_3241) );
na02s01 TIMEBOOST_cell_4067 ( .a(n_44498), .b(FE_OCP_RBN5954_FE_OFN4772_n_44463), .o(TIMEBOOST_net_1124) );
no02s02 g777909 ( .a(n_3183), .b(n_3122), .o(n_3196) );
na02s04 g777910 ( .a(n_3055), .b(n_3159), .o(n_3174) );
no02s02 g777911 ( .a(FE_OCP_RBN5708_n_3055), .b(n_3160), .o(n_3185) );
na02s01 g777913 ( .a(n_3083), .b(n_2968), .o(n_3117) );
na02s01 g777914 ( .a(n_3114), .b(n_2967), .o(n_3115) );
no02s01 g777915 ( .a(n_3149), .b(n_2983), .o(n_3150) );
in01s04 g777916 ( .a(n_3133), .o(n_3120) );
oa12s06 g777918 ( .a(n_2358), .b(n_3096), .c(n_2314), .o(n_3133) );
ao12s01 g777919 ( .a(n_3108), .b(n_3111), .c(n_2589), .o(n_3157) );
ao12s01 g777920 ( .a(n_3088), .b(n_3111), .c(n_3087), .o(n_4686) );
na02s02 g777922 ( .a(n_3097), .b(n_3107), .o(n_4211) );
na02f02 g777923 ( .a(n_3175), .b(n_3194), .o(n_3275) );
oa12m06 g777924 ( .a(n_2655), .b(n_3111), .c(n_3108), .o(n_3112) );
in01s02 g777925 ( .a(n_3214), .o(n_3215) );
na02s02 TIMEBOOST_cell_2880 ( .a(FE_RN_839_0), .b(n_7165), .o(TIMEBOOST_net_731) );
na02s01 g777927 ( .a(n_3096), .b(n_45194), .o(n_3097) );
na02s01 g777928 ( .a(n_3075), .b(n_2408), .o(n_3107) );
no02s02 g777929 ( .a(n_3122), .b(n_2785), .o(n_3216) );
in01s01 g777930 ( .a(n_3183), .o(n_3184) );
no02s02 g777931 ( .a(n_3142), .b(FE_OCP_RBN2627_n_2737), .o(n_3183) );
na02m08 TIMEBOOST_cell_2879 ( .a(n_7417), .b(TIMEBOOST_net_730), .o(n_7470) );
in01s01 g777933 ( .a(n_3169), .o(n_3170) );
na02s02 g777934 ( .a(n_3142), .b(FE_OCP_RBN2627_n_2737), .o(n_3169) );
na02s02 g777935 ( .a(n_47022), .b(FE_OCP_RBN2627_n_2737), .o(n_3132) );
no02s01 g777936 ( .a(n_3111), .b(n_3087), .o(n_3088) );
no02m02 g777938 ( .a(n_2987), .b(n_3138), .o(n_3167) );
na02s02 g777939 ( .a(n_47021), .b(n_3080), .o(n_3175) );
na02s02 g777940 ( .a(n_3137), .b(n_3597), .o(n_3194) );
in01s01 g777941 ( .a(n_3147), .o(n_3119) );
oa12m06 g777942 ( .a(n_2265), .b(n_3092), .c(n_2244), .o(n_3147) );
in01s02 g777943 ( .a(n_3159), .o(n_3160) );
ao12m04 g777944 ( .a(n_3049), .b(n_3116), .c(FE_OCP_RBN5649_n_2438), .o(n_3159) );
oa12m02 g777946 ( .a(n_3047), .b(n_3116), .c(FE_OCP_RBN5649_n_2438), .o(n_3161) );
oa12s01 g777947 ( .a(n_3046), .b(n_3045), .c(n_3044), .o(n_4537) );
oa12s01 g777948 ( .a(n_3073), .b(n_3072), .c(n_3071), .o(n_4632) );
in01s02 g777949 ( .a(n_47020), .o(n_3231) );
oa22s01 g777952 ( .a(n_3163), .b(FE_OCP_RBN4147_n_3217), .c(n_3218), .d(n_3217), .o(n_3248) );
in01s01 g777953 ( .a(n_3717), .o(n_3715) );
ao12s01 g777954 ( .a(n_3091), .b(n_3090), .c(n_3089), .o(n_3717) );
in01s01 g777955 ( .a(n_4662), .o(n_3118) );
ao12s01 g777956 ( .a(n_3070), .b(n_3069), .c(n_3068), .o(n_4662) );
in01s01 g777959 ( .a(n_3114), .o(n_3083) );
oa12m04 g777960 ( .a(n_2906), .b(n_3030), .c(n_2830), .o(n_3114) );
no02s02 g777963 ( .a(n_3092), .b(n_2286), .o(n_3093) );
na02s01 g777964 ( .a(n_3045), .b(n_3044), .o(n_3046) );
oa12m06 g777965 ( .a(n_2593), .b(n_3022), .c(n_2603), .o(n_3111) );
no02s01 g777966 ( .a(n_3069), .b(n_3068), .o(n_3070) );
in01s01 g777968 ( .a(n_3210), .o(n_3211) );
na02s01 g777969 ( .a(n_3200), .b(n_3199), .o(n_3210) );
no02s01 g777970 ( .a(n_3090), .b(n_3089), .o(n_3091) );
no02s01 g777971 ( .a(n_3154), .b(FE_OCP_RBN4147_n_3217), .o(n_3179) );
in01s01 g777972 ( .a(n_3190), .o(n_3191) );
na02s02 g777973 ( .a(n_3124), .b(n_3165), .o(n_3190) );
na02s01 g777974 ( .a(n_3072), .b(n_3071), .o(n_3073) );
in01s01 g777975 ( .a(n_3096), .o(n_3075) );
oa12s06 g777976 ( .a(n_2324), .b(n_3031), .c(n_2301), .o(n_3096) );
oa12s04 g777977 ( .a(n_2832), .b(n_3057), .c(FE_OCP_RBN5652_n_2438), .o(n_3138) );
oa12s02 g777978 ( .a(n_2866), .b(n_3056), .c(FE_OCP_RBN5658_n_2438), .o(n_3122) );
in01s02 g777979 ( .a(n_47021), .o(n_3137) );
no02s01 TIMEBOOST_cell_2802 ( .a(n_1443), .b(n_1508), .o(TIMEBOOST_net_692) );
no02s01 g777986 ( .a(n_3031), .b(n_2333), .o(n_3032) );
no02s02 g777987 ( .a(n_3048), .b(n_2850), .o(n_3100) );
no02s02 g777988 ( .a(n_47023), .b(FE_OCP_RBN5660_n_2438), .o(n_3037) );
no02s01 g777990 ( .a(n_3022), .b(n_2635), .o(n_3072) );
no02m08 TIMEBOOST_cell_5103 ( .a(n_8746), .b(TIMEBOOST_net_1499), .o(n_8817) );
in01s02 g777993 ( .a(n_3154), .o(n_3199) );
no02s02 g777994 ( .a(n_3128), .b(n_3127), .o(n_3154) );
in01s01 g777995 ( .a(n_3200), .o(n_3151) );
na02s03 g777996 ( .a(n_3128), .b(n_3127), .o(n_3200) );
in01s01 g777997 ( .a(n_3123), .o(n_3124) );
no02s03 g777998 ( .a(n_3067), .b(n_2558), .o(n_3123) );
in01s02 g777999 ( .a(n_3086), .o(n_3165) );
no02s01 g778000 ( .a(n_3066), .b(FE_OCP_RBN2574_n_2558), .o(n_3086) );
in01s01 g778001 ( .a(n_3172), .o(n_3173) );
no02s01 g778002 ( .a(n_3103), .b(n_3140), .o(n_3172) );
oa12s01 g778005 ( .a(n_2389), .b(n_3008), .c(n_2449), .o(n_3045) );
in01s01 g778006 ( .a(n_3580), .o(n_3563) );
oa12s01 g778007 ( .a(n_2970), .b(n_2969), .c(n_3013), .o(n_3580) );
in01s01 g778008 ( .a(n_3218), .o(n_3163) );
no02s02 g778009 ( .a(n_3065), .b(n_3098), .o(n_3218) );
ao12s01 g778010 ( .a(n_2992), .b(n_2991), .c(n_2990), .o(n_4575) );
in01s01 g778011 ( .a(n_3030), .o(n_3069) );
ao12m04 g778012 ( .a(n_2749), .b(n_3013), .c(n_2816), .o(n_3030) );
oa12s01 g778013 ( .a(n_2986), .b(n_3008), .c(n_2985), .o(n_4298) );
in01s01 g778014 ( .a(n_4719), .o(n_3113) );
no02s02 g778015 ( .a(n_3021), .b(n_3051), .o(n_4719) );
oa22s01 g778017 ( .a(n_3076), .b(n_3058), .c(n_3126), .d(n_3125), .o(n_3152) );
in01s02 g778018 ( .a(n_3673), .o(n_3155) );
na02s06 g778019 ( .a(n_3019), .b(n_3009), .o(n_3673) );
oa12s01 g778020 ( .a(n_2856), .b(n_3020), .c(n_3034), .o(n_3090) );
na02s02 g778022 ( .a(n_2996), .b(n_2248), .o(n_3019) );
na02s02 g778023 ( .a(n_3000), .b(n_2247), .o(n_3009) );
na02s01 g778025 ( .a(n_3008), .b(n_2985), .o(n_2986) );
no02m08 g778026 ( .a(n_2991), .b(n_2634), .o(n_3022) );
no02m03 g778028 ( .a(n_3018), .b(FE_OCP_RBN5652_n_2438), .o(n_3049) );
in01s01 g778029 ( .a(n_3047), .o(n_3048) );
na02s02 g778030 ( .a(n_3018), .b(FE_OCP_RBN5653_n_2438), .o(n_3047) );
in01s01 g778031 ( .a(n_3102), .o(n_3103) );
na02m02 g778032 ( .a(n_3085), .b(n_3084), .o(n_3102) );
no02s01 g778033 ( .a(n_3035), .b(n_3626), .o(n_3065) );
no02s02 g778034 ( .a(n_3085), .b(n_3084), .o(n_3140) );
no02s01 g778035 ( .a(n_3038), .b(n_3058), .o(n_3059) );
no02s02 g778036 ( .a(FE_OCP_RBN2767_n_3035), .b(FE_OCP_RBN4175_n_3626), .o(n_3098) );
na02s01 g778037 ( .a(n_2969), .b(n_3013), .o(n_2970) );
no02s01 g778038 ( .a(n_2861), .b(n_3020), .o(n_3021) );
no02s01 g778039 ( .a(n_2991), .b(n_2990), .o(n_2992) );
in01s01 g778040 ( .a(n_3130), .o(n_3131) );
na02s01 g778041 ( .a(FE_RN_16_0), .b(n_3109), .o(n_3130) );
no02s01 g778042 ( .a(n_2862), .b(n_2980), .o(n_3051) );
no02m06 g778043 ( .a(n_2980), .b(n_2777), .o(n_3063) );
in01s01 g778044 ( .a(n_3104), .o(n_3105) );
na02s01 g778045 ( .a(n_3101), .b(n_3329), .o(n_3104) );
na02s06 g778047 ( .a(n_2944), .b(n_2263), .o(n_3031) );
no02f08 TIMEBOOST_cell_4022 ( .a(TIMEBOOST_net_1101), .b(TIMEBOOST_net_657), .o(n_35102) );
oa12s01 g778049 ( .a(n_2961), .b(n_2960), .c(n_2959), .o(n_4333) );
in01s02 g778050 ( .a(n_3066), .o(n_3067) );
oa22s02 g778051 ( .a(n_3055), .b(n_3502), .c(FE_OCP_RBN5709_n_3055), .d(FE_OCP_RBN6641_n_3502), .o(n_3066) );
in01s02 g778054 ( .a(n_3056), .o(n_3057) );
no02s02 g778055 ( .a(n_2953), .b(n_2995), .o(n_3056) );
na02s06 g778056 ( .a(n_2914), .b(n_2264), .o(n_2944) );
na02s01 g778058 ( .a(n_2914), .b(n_2280), .o(n_2915) );
na02s01 g778059 ( .a(n_2960), .b(n_2959), .o(n_2961) );
na02f06 TIMEBOOST_cell_5311 ( .a(TIMEBOOST_net_1603), .b(n_39678), .o(n_39691) );
no02m04 TIMEBOOST_cell_2947 ( .a(TIMEBOOST_net_764), .b(n_12949), .o(n_13290) );
no02s02 g778062 ( .a(FE_OCP_RBN4176_n_3626), .b(FE_OCP_RBN5653_n_2438), .o(n_2995) );
no02s02 g778063 ( .a(n_3626), .b(FE_OCP_RBN5663_n_2438), .o(n_2953) );
in01s01 g778064 ( .a(n_3038), .o(n_3329) );
no02s02 g778065 ( .a(n_3024), .b(n_3023), .o(n_3038) );
no02s02 g778067 ( .a(n_3040), .b(n_3039), .o(n_3061) );
in01s01 g778068 ( .a(n_3101), .o(n_3043) );
na02s02 g778069 ( .a(n_3024), .b(n_3023), .o(n_3101) );
na02s02 g778070 ( .a(n_3040), .b(n_3039), .o(n_3109) );
in01s01 g778071 ( .a(n_3000), .o(n_2996) );
oa12m06 g778072 ( .a(n_2202), .b(FE_OCP_RBN5692_n_2884), .c(n_2181), .o(n_3000) );
ao12s01 g778073 ( .a(n_2375), .b(n_2924), .c(n_2331), .o(n_3008) );
in01s01 TIMEBOOST_cell_5920 ( .a(TIMEBOOST_net_1808), .o(TIMEBOOST_net_1809) );
ao12m06 g778076 ( .a(n_2561), .b(n_2924), .c(n_2501), .o(n_2991) );
oa12m04 g778077 ( .a(n_2724), .b(FE_OCP_RBN2703_FE_RN_984_0), .c(FE_OCP_RBN4174_FE_OCPN1913_n_2669), .o(n_3013) );
in01s01 g778078 ( .a(n_4642), .o(n_3025) );
na02s01 g778079 ( .a(n_2939), .b(n_2949), .o(n_4642) );
in01s01 g778080 ( .a(n_4587), .o(n_3012) );
na03f08 TIMEBOOST_cell_8419 ( .a(FE_OCP_RBN2084_n_19970), .b(n_19804), .c(n_20001), .o(n_20094) );
na02s04 TIMEBOOST_cell_4066 ( .a(TIMEBOOST_net_1123), .b(n_9333), .o(n_9377) );
in01s01 g778084 ( .a(n_2980), .o(n_3020) );
oa12m06 g778085 ( .a(n_2775), .b(n_2938), .c(n_2739), .o(n_2980) );
in01s02 g778086 ( .a(n_3597), .o(n_3080) );
no02s06 g778087 ( .a(n_2897), .b(n_2943), .o(n_3597) );
in01s02 g778088 ( .a(n_3076), .o(n_3126) );
na02s06 TIMEBOOST_cell_6232 ( .a(TIMEBOOST_net_1967), .b(n_30933), .o(TIMEBOOST_net_1651) );
no02s02 g778091 ( .a(n_2884), .b(n_2216), .o(n_2897) );
no02s02 g778092 ( .a(FE_OCP_RBN5691_n_2884), .b(n_2217), .o(n_2943) );
no02s01 g778093 ( .a(n_2924), .b(n_2533), .o(n_2960) );
na02s02 g778094 ( .a(n_2866), .b(n_2865), .o(n_2867) );
na02s06 g778096 ( .a(n_2940), .b(n_2851), .o(n_3055) );
na02s03 g778098 ( .a(n_2987), .b(n_2865), .o(n_3016) );
na02f08 TIMEBOOST_cell_6736 ( .a(TIMEBOOST_net_2125), .b(n_14667), .o(n_14798) );
no02m08 TIMEBOOST_cell_8534 ( .a(n_24458), .b(n_24548), .o(TIMEBOOST_net_2754) );
na02s02 g778101 ( .a(n_2950), .b(n_2978), .o(n_2979) );
na02m08 TIMEBOOST_cell_2943 ( .a(n_2428), .b(TIMEBOOST_net_762), .o(n_2524) );
no03f06 TIMEBOOST_cell_8315 ( .a(n_14798), .b(FE_OCP_RBN4206_n_13796), .c(n_14856), .o(n_14857) );
in01s01 g778104 ( .a(n_3026), .o(n_3027) );
na02s01 g778105 ( .a(n_2965), .b(n_2999), .o(n_3026) );
na02s01 g778106 ( .a(n_2827), .b(n_2896), .o(n_2949) );
na02s01 g778107 ( .a(n_2826), .b(n_2938), .o(n_2939) );
in01s01 g778108 ( .a(n_3004), .o(n_3005) );
na02s01 g778109 ( .a(n_2923), .b(n_2977), .o(n_3004) );
no02s01 g778110 ( .a(n_2761), .b(FE_OCP_RBN2703_FE_RN_984_0), .o(n_2892) );
no02s06 g778113 ( .a(n_2209), .b(n_2820), .o(n_2914) );
no02m08 TIMEBOOST_cell_2908 ( .a(n_33530), .b(n_33081), .o(TIMEBOOST_net_745) );
oa12s01 g778115 ( .a(n_2846), .b(n_2845), .c(n_2844), .o(n_4207) );
na03m10 TIMEBOOST_cell_4758 ( .a(n_20463), .b(n_20764), .c(TIMEBOOST_net_901), .o(n_20910) );
no02f08 TIMEBOOST_cell_8550 ( .a(FE_OCP_RBN5646_n_33785), .b(n_33717), .o(TIMEBOOST_net_2762) );
no02s02 g778119 ( .a(n_2789), .b(n_2226), .o(n_2855) );
no02s06 g778120 ( .a(n_2208), .b(n_2805), .o(n_2820) );
no02s04 TIMEBOOST_cell_5045 ( .a(TIMEBOOST_net_1470), .b(FE_OCP_RBN2674_n_8163), .o(n_8296) );
no02m08 g778122 ( .a(n_2845), .b(n_2534), .o(n_2924) );
na02s01 g778123 ( .a(n_2845), .b(n_2844), .o(n_2846) );
no02s04 TIMEBOOST_cell_8565 ( .a(TIMEBOOST_net_2769), .b(FE_OCP_RBN5861_n_3718), .o(n_3933) );
na02f04 TIMEBOOST_cell_7503 ( .a(n_23346), .b(TIMEBOOST_net_2382), .o(FE_RN_74_0) );
no02m02 TIMEBOOST_cell_2907 ( .a(TIMEBOOST_net_744), .b(n_18379), .o(n_18438) );
na02s02 g778127 ( .a(n_2872), .b(FE_OCPN1620_n_3361), .o(n_2890) );
in01s02 g778128 ( .a(n_2950), .o(n_2951) );
no02m02 g778129 ( .a(n_2932), .b(n_2774), .o(n_2950) );
na02s02 g778131 ( .a(FE_OCP_RBN4166_n_3494), .b(FE_OCP_RBN5658_n_2438), .o(n_2832) );
in01s01 g778132 ( .a(n_2957), .o(n_2958) );
na02s02 g778133 ( .a(n_2886), .b(n_2823), .o(n_2957) );
na02s02 g778134 ( .a(FE_OCP_RBN4167_n_3494), .b(FE_OCP_RBN5653_n_2438), .o(n_2866) );
na02s01 g778135 ( .a(n_2899), .b(n_2898), .o(n_2977) );
in01s01 g778136 ( .a(n_2922), .o(n_2923) );
no02s02 g778137 ( .a(n_2899), .b(n_2898), .o(n_2922) );
in01s01 g778138 ( .a(n_2967), .o(n_2968) );
na02s01 g778139 ( .a(n_2908), .b(n_2963), .o(n_2967) );
na02s02 g778140 ( .a(n_2930), .b(FE_OFN321_n_2929), .o(n_2999) );
in01s01 g778141 ( .a(n_2964), .o(n_2965) );
no02s02 g778142 ( .a(n_2930), .b(FE_OFN321_n_2929), .o(n_2964) );
na02s01 g778144 ( .a(n_2956), .b(n_2903), .o(n_2983) );
oa12m06 g778146 ( .a(n_2180), .b(FE_OCP_RBN2645_n_2747), .c(n_2141), .o(n_2884) );
in01m02 g778147 ( .a(n_2850), .o(n_2851) );
oa12s02 g778148 ( .a(n_2823), .b(FE_OCP_RBN4164_n_3390), .c(FE_OCP_RBN5649_n_2438), .o(n_2850) );
na02s02 g778149 ( .a(n_2932), .b(n_2743), .o(n_2987) );
na02s03 g778151 ( .a(n_2885), .b(n_2813), .o(n_2940) );
ao12s01 g778152 ( .a(n_2716), .b(n_2715), .c(n_2714), .o(n_4136) );
in01s01 g778153 ( .a(FE_OCP_RBN2703_FE_RN_984_0), .o(n_2875) );
na02m06 g778156 ( .a(n_2802), .b(n_2793), .o(n_3502) );
oa12s01 g778157 ( .a(n_2755), .b(n_2754), .c(n_2753), .o(n_4433) );
in01s01 g778158 ( .a(n_2938), .o(n_2896) );
na02m06 g778159 ( .a(n_2824), .b(n_2637), .o(n_2938) );
ao12s01 g778160 ( .a(n_2854), .b(n_2853), .c(n_2852), .o(n_4437) );
na02s03 g778161 ( .a(FE_OCP_RBN2646_n_2747), .b(n_2193), .o(n_2802) );
na02s01 g778162 ( .a(n_2747), .b(n_2192), .o(n_2793) );
no02s01 g778163 ( .a(n_2715), .b(n_2714), .o(n_2716) );
in01s01 g778164 ( .a(n_2888), .o(n_2889) );
na02s06 g778165 ( .a(n_2860), .b(n_2673), .o(n_2888) );
in01s01 g778166 ( .a(n_2872), .o(n_2873) );
na02s02 g778167 ( .a(n_2843), .b(n_2579), .o(n_2872) );
na02s02 g778168 ( .a(FE_OCP_RBN4163_n_3390), .b(FE_OCP_RBN5649_n_2438), .o(n_2813) );
in01s01 g778169 ( .a(n_2907), .o(n_2908) );
no02s02 g778170 ( .a(n_2859), .b(n_2858), .o(n_2907) );
na02s02 g778171 ( .a(n_2859), .b(n_2858), .o(n_2963) );
na02s01 g778172 ( .a(n_2754), .b(n_2753), .o(n_2755) );
in01s01 g778173 ( .a(n_2902), .o(n_2903) );
no02s03 g778174 ( .a(n_2864), .b(n_2863), .o(n_2902) );
na02s03 g778175 ( .a(n_2864), .b(n_2863), .o(n_2956) );
no02s01 g778176 ( .a(n_2853), .b(n_2852), .o(n_2854) );
na02m04 g778178 ( .a(n_2778), .b(n_2624), .o(n_2824) );
na02s01 g778179 ( .a(n_2906), .b(n_2831), .o(n_3068) );
in01s01 g778180 ( .a(n_2805), .o(n_2789) );
no02m08 g778182 ( .a(n_2742), .b(n_2479), .o(n_2845) );
in01s01 g778183 ( .a(n_2865), .o(n_2785) );
ao12s02 g778184 ( .a(n_2774), .b(n_3006), .c(FE_OCP_RBN5653_n_2438), .o(n_2865) );
in01s02 g778185 ( .a(n_2885), .o(n_2886) );
no02s03 g778186 ( .a(n_2843), .b(n_2680), .o(n_2885) );
no02m02 g778187 ( .a(n_2860), .b(n_2675), .o(n_2932) );
oa12s01 g778188 ( .a(n_3209), .b(n_3208), .c(n_3207), .o(n_4018) );
ao12s01 g778189 ( .a(n_2808), .b(n_2871), .c(n_2870), .o(n_3089) );
in01s01 g778191 ( .a(FE_OCP_RBN4166_n_3494), .o(n_2784) );
oa12s01 g778192 ( .a(n_2700), .b(n_2699), .c(n_2698), .o(n_3494) );
oa12s01 g778193 ( .a(n_2693), .b(n_2692), .c(n_2691), .o(n_4142) );
na02s01 g778195 ( .a(n_2699), .b(n_2698), .o(n_2700) );
na02s01 g778196 ( .a(n_3208), .b(n_3207), .o(n_3209) );
na02s01 g778197 ( .a(n_2692), .b(n_2691), .o(n_2693) );
na02s01 g778198 ( .a(n_3006), .b(FE_OCP_RBN5649_n_2438), .o(n_2743) );
no02m06 g778199 ( .a(n_45505), .b(n_2383), .o(n_2742) );
no02s01 g778201 ( .a(n_2871), .b(n_2870), .o(n_2808) );
na02s02 g778202 ( .a(n_2795), .b(n_2794), .o(n_2906) );
in01s01 g778203 ( .a(n_2830), .o(n_2831) );
no02s02 g778204 ( .a(n_2795), .b(n_2794), .o(n_2830) );
na02s01 g778205 ( .a(n_2750), .b(n_2816), .o(n_2969) );
in01s01 g778206 ( .a(n_2861), .o(n_2862) );
na02s01 g778207 ( .a(n_2856), .b(n_2799), .o(n_2861) );
oa12m06 g778209 ( .a(n_2123), .b(n_2711), .c(n_2097), .o(n_2747) );
oa12s01 g778210 ( .a(n_2431), .b(n_2619), .c(n_2274), .o(n_2715) );
ao12s02 g778211 ( .a(n_44059), .b(FE_OCPN1620_n_3361), .c(FE_OCP_RBN6611_n_2289), .o(n_2823) );
na02s06 g778213 ( .a(n_2792), .b(n_2649), .o(n_2843) );
na02m08 g778214 ( .a(n_2829), .b(n_2665), .o(n_2860) );
no02s01 TIMEBOOST_cell_8776 ( .a(n_2784), .b(FE_OCP_RBN4166_n_3494), .o(TIMEBOOST_net_2875) );
in01s01 g778216 ( .a(n_2778), .o(n_2852) );
na02s04 TIMEBOOST_cell_2806 ( .a(n_1656), .b(n_1657), .o(TIMEBOOST_net_694) );
ao12s01 g778218 ( .a(n_2668), .b(n_2667), .c(n_2709), .o(n_4339) );
oa12s01 g778220 ( .a(n_2690), .b(n_2689), .c(n_2688), .o(n_4435) );
oa12m02 g778222 ( .a(n_2505), .b(n_2709), .c(n_2573), .o(n_2753) );
ao22m01 g778224 ( .a(n_2711), .b(n_2155), .c(n_2638), .d(n_2154), .o(n_3390) );
na02s01 g778225 ( .a(n_2619), .b(n_2326), .o(n_3208) );
no02s02 g778226 ( .a(n_2679), .b(FE_OCP_RBN6611_n_2289), .o(n_2680) );
no02s01 g778227 ( .a(n_2674), .b(FE_OCP_RBN6611_n_2289), .o(n_2675) );
na02s02 g778228 ( .a(n_2718), .b(n_2717), .o(n_2816) );
na02s01 g778229 ( .a(n_2689), .b(n_2688), .o(n_2690) );
in01s01 g778230 ( .a(n_2826), .o(n_2827) );
na02s01 g778231 ( .a(n_2775), .b(n_2740), .o(n_2826) );
in01s01 g778232 ( .a(n_2749), .o(n_2750) );
no02s02 g778233 ( .a(n_2718), .b(n_2717), .o(n_2749) );
no02s01 g778234 ( .a(n_2667), .b(n_2709), .o(n_2668) );
no02s02 g778235 ( .a(n_2763), .b(FE_OCP_RBN2573_n_2558), .o(n_2748) );
na02s01 TIMEBOOST_cell_8660 ( .a(n_31730), .b(n_30933), .o(TIMEBOOST_net_2817) );
in01s01 g778237 ( .a(n_2799), .o(n_3034) );
na02s02 g778238 ( .a(n_47025), .b(n_2766), .o(n_2799) );
in01s01 g778239 ( .a(n_2777), .o(n_2856) );
no02s02 g778240 ( .a(n_47025), .b(n_2766), .o(n_2777) );
oa12m06 g778242 ( .a(n_2111), .b(n_2615), .c(n_2153), .o(n_2699) );
no02f06 TIMEBOOST_cell_5237 ( .a(TIMEBOOST_net_1566), .b(n_15352), .o(n_15552) );
in01s01 g778244 ( .a(n_2760), .o(n_2761) );
na02s01 g778245 ( .a(n_2724), .b(FE_OCPN1913_n_2669), .o(n_2760) );
na02s02 g778246 ( .a(n_2725), .b(n_3127), .o(n_2726) );
oa12s01 g778247 ( .a(n_2947), .b(n_2946), .c(delay_sub_ln21_0_unr2_stage2_stallmux_q_29_), .o(n_2948) );
na02s01 g778248 ( .a(n_45506), .b(n_2480), .o(n_2692) );
in01s01 g778250 ( .a(n_2792), .o(n_2756) );
no02s06 g778251 ( .a(n_2725), .b(n_2563), .o(n_2792) );
no02s06 g778253 ( .a(n_2763), .b(n_2565), .o(n_2829) );
no02s02 g778254 ( .a(n_2650), .b(n_2704), .o(n_2871) );
in01s01 g778255 ( .a(n_3006), .o(n_2978) );
oa12s02 g778256 ( .a(n_2588), .b(n_2615), .c(n_2587), .o(n_3006) );
ao12s01 g778257 ( .a(n_2576), .b(n_2575), .c(n_2574), .o(n_3911) );
no02s02 TIMEBOOST_cell_5298 ( .a(n_4050), .b(n_4033), .o(TIMEBOOST_net_1597) );
na02s01 g778259 ( .a(n_2894), .b(n_2836), .o(n_2887) );
na02s01 g778260 ( .a(n_2615), .b(n_2587), .o(n_2588) );
in01s01 g778261 ( .a(n_2918), .o(n_2919) );
na02s02 g778262 ( .a(n_2894), .b(n_2895), .o(n_2918) );
in01s01 g778263 ( .a(n_2997), .o(n_2998) );
no02s01 g778264 ( .a(n_4073), .b(n_2976), .o(n_2997) );
no02s01 g778265 ( .a(n_3857), .b(n_2920), .o(n_2982) );
in01s01 g778266 ( .a(n_3014), .o(n_3015) );
na02s01 g778267 ( .a(n_2921), .b(n_2975), .o(n_3014) );
na02s01 g778268 ( .a(n_2575), .b(n_2325), .o(n_2619) );
no02s01 g778269 ( .a(n_2575), .b(n_2574), .o(n_2576) );
na02s01 g778270 ( .a(n_2633), .b(n_3125), .o(n_2646) );
no02s06 TIMEBOOST_cell_5297 ( .a(TIMEBOOST_net_1596), .b(n_39162), .o(n_39335) );
no02s01 g778272 ( .a(n_2647), .b(n_3084), .o(n_2650) );
no02s01 g778273 ( .a(n_2642), .b(n_2294), .o(n_2704) );
in01s01 g778274 ( .a(n_2739), .o(n_2740) );
no02s03 g778275 ( .a(n_47026), .b(FE_OCPN1052_n_2702), .o(n_2739) );
na02s02 g778276 ( .a(n_2623), .b(n_2622), .o(n_2724) );
no02s01 g778277 ( .a(n_2625), .b(n_2636), .o(n_2853) );
na02s01 g778280 ( .a(n_2535), .b(FE_RN_982_0), .o(n_2754) );
no02s01 g778281 ( .a(n_3857), .b(n_2988), .o(n_2989) );
na02s02 g778282 ( .a(n_47026), .b(FE_OCPN1052_n_2702), .o(n_2775) );
in01s01 g778283 ( .a(n_2911), .o(n_2912) );
ao12s01 g778284 ( .a(n_2835), .b(n_2947), .c(delay_sub_ln21_0_unr2_stage2_stallmux_q_29_), .o(n_2911) );
in01s06 g778285 ( .a(n_2638), .o(n_2711) );
na02f04 TIMEBOOST_cell_5245 ( .a(TIMEBOOST_net_1570), .b(n_14682), .o(n_14736) );
in01s01 g778289 ( .a(n_2725), .o(n_2697) );
na02m04 g778290 ( .a(n_2647), .b(n_2548), .o(n_2725) );
na02m08 g778291 ( .a(FE_OCP_RBN6632_n_2633), .b(n_2543), .o(n_2763) );
ao12s02 g778293 ( .a(n_2525), .b(n_2524), .c(n_2523), .o(n_2674) );
oa12s01 g778294 ( .a(n_2555), .b(n_2554), .c(FE_OCP_RBN2571_n_2430), .o(n_4280) );
no02m04 g778295 ( .a(n_2517), .b(n_2443), .o(n_2709) );
na02m04 g778296 ( .a(n_2559), .b(n_2464), .o(n_2688) );
in01s01 g778297 ( .a(n_2973), .o(n_2974) );
oa12s01 g778298 ( .a(n_2901), .b(n_2910), .c(delay_add_ln22_unr2_stage2_stallmux_q_31_), .o(n_2973) );
in01s01 g778299 ( .a(n_3361), .o(n_2679) );
oa12m01 g778300 ( .a(n_2519), .b(n_2528), .c(n_2518), .o(n_3361) );
ao12s01 g778301 ( .a(n_2600), .b(n_2599), .c(FE_OCP_RBN5626_n_2457), .o(n_4231) );
na02m06 TIMEBOOST_cell_8885 ( .a(TIMEBOOST_net_2929), .b(TIMEBOOST_net_2696), .o(n_22494) );
in01s01 g778304 ( .a(n_44059), .o(n_2579) );
ao22s02 g778306 ( .a(n_2558), .b(FE_OCP_RBN6611_n_2289), .c(n_2664), .d(FE_OCP_RBN6611_n_2289), .o(n_2673) );
in01s01 g778307 ( .a(n_2849), .o(n_2894) );
no02s01 g778308 ( .a(n_2796), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_28_), .o(n_2849) );
in01s01 g778309 ( .a(n_2895), .o(n_2946) );
na02s01 g778310 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_28_), .b(n_2796), .o(n_2895) );
in01s01 g778311 ( .a(n_2835), .o(n_2836) );
no02s01 g778312 ( .a(n_2947), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_29_), .o(n_2835) );
in01s01 g778313 ( .a(n_2847), .o(n_2848) );
no02s01 g778314 ( .a(n_2798), .b(n_2797), .o(n_2847) );
in01s01 g778315 ( .a(n_2904), .o(n_2905) );
na02s01 g778316 ( .a(n_2874), .b(n_2819), .o(n_2904) );
in01s01 g778317 ( .a(n_2927), .o(n_2976) );
na02s01 g778318 ( .a(n_2910), .b(delay_add_ln22_unr2_stage2_stallmux_q_30_), .o(n_2927) );
na02s01 g778319 ( .a(n_2910), .b(delay_add_ln22_unr2_stage2_stallmux_q_31_), .o(n_2901) );
no02s01 g778320 ( .a(n_2524), .b(n_2523), .o(n_2525) );
na02s01 g778321 ( .a(n_2910), .b(delay_add_ln22_unr2_stage2_stallmux_q_29_), .o(n_2975) );
in01s01 g778322 ( .a(n_3857), .o(n_2962) );
no02s01 g778323 ( .a(n_2869), .b(delay_add_ln22_unr2_stage2_stallmux_q_28_), .o(n_3857) );
no02s01 g778324 ( .a(n_2910), .b(delay_add_ln22_unr2_stage2_stallmux_q_30_), .o(n_4073) );
na02s01 g778325 ( .a(n_2528), .b(n_2518), .o(n_2519) );
na02m08 g778326 ( .a(n_2524), .b(n_2066), .o(n_2615) );
no02s01 g778327 ( .a(n_47024), .b(n_1095), .o(n_2988) );
in01s01 g778328 ( .a(n_2920), .o(n_2921) );
no02s01 g778329 ( .a(n_2910), .b(delay_add_ln22_unr2_stage2_stallmux_q_29_), .o(n_2920) );
na02m08 TIMEBOOST_cell_2825 ( .a(n_7209), .b(TIMEBOOST_net_703), .o(n_7258) );
no02s01 g778331 ( .a(n_2841), .b(n_2834), .o(n_2909) );
na02s03 g778332 ( .a(FE_OCP_RBN6617_n_2289), .b(FE_OCP_RBN4147_n_3217), .o(n_2649) );
na02s02 g778333 ( .a(n_2664), .b(FE_OCP_RBN6613_n_2289), .o(n_2665) );
no02m04 TIMEBOOST_cell_6248 ( .a(TIMEBOOST_net_1975), .b(n_5609), .o(TIMEBOOST_net_1662) );
no02s01 g778335 ( .a(n_2604), .b(n_3039), .o(n_2605) );
na02s01 g778336 ( .a(n_2554), .b(FE_OCP_RBN2571_n_2430), .o(n_2555) );
in01s01 g778337 ( .a(n_2624), .o(n_2625) );
na02m02 g778338 ( .a(n_2607), .b(n_2606), .o(n_2624) );
no02s01 g778339 ( .a(n_2506), .b(n_2573), .o(n_2667) );
no02s02 g778341 ( .a(n_2495), .b(n_2494), .o(n_2526) );
no02f08 TIMEBOOST_cell_8551 ( .a(TIMEBOOST_net_2762), .b(FE_OCP_RBN4913_n_33833), .o(n_33962) );
in01s02 g778343 ( .a(n_2636), .o(n_2637) );
no02s02 g778344 ( .a(n_2607), .b(n_2606), .o(n_2636) );
no02s01 g778346 ( .a(n_2599), .b(FE_OCP_RBN5626_n_2457), .o(n_2600) );
na02s01 g778347 ( .a(n_2627), .b(n_2626), .o(n_2689) );
na02s02 g778349 ( .a(n_2495), .b(n_2494), .o(n_2535) );
ao12m06 g778350 ( .a(n_2366), .b(n_2308), .c(n_2508), .o(n_2575) );
na02m08 g778352 ( .a(FE_OCP_RBN6625_n_2537), .b(n_2474), .o(n_2633) );
in01s01 g778353 ( .a(n_2647), .o(n_2642) );
no02s04 g778354 ( .a(n_2604), .b(n_2498), .o(n_2647) );
na02s02 TIMEBOOST_cell_2904 ( .a(n_29017), .b(FE_OCP_RBN2514_n_28699), .o(TIMEBOOST_net_743) );
in01s01 g778357 ( .a(n_2531), .o(n_2532) );
oa12s01 g778358 ( .a(n_2447), .b(n_2446), .c(n_2445), .o(n_2531) );
na03s08 TIMEBOOST_cell_5707 ( .a(n_32699), .b(n_32698), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_6_), .o(n_32708) );
oa12s01 g778360 ( .a(n_2478), .b(n_2508), .c(n_2477), .o(n_3902) );
no02s01 TIMEBOOST_cell_3828 ( .a(TIMEBOOST_net_1004), .b(n_28131), .o(n_28201) );
in01s01 g778362 ( .a(n_2583), .o(n_2584) );
ao12s01 g778363 ( .a(n_2489), .b(n_2488), .c(n_2487), .o(n_2583) );
na02s01 g778364 ( .a(n_2787), .b(n_2115), .o(n_2910) );
in01s01 g778365 ( .a(n_2809), .o(n_2810) );
na02s01 g778366 ( .a(n_2790), .b(n_3594), .o(n_2809) );
no02s02 g778367 ( .a(n_2686), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_27_), .o(n_2798) );
in01s01 g778368 ( .a(n_2818), .o(n_2819) );
no02s02 g778369 ( .a(n_2782), .b(delay_add_ln22_unr2_stage2_stallmux_q_27_), .o(n_2818) );
na02s02 g778370 ( .a(n_2782), .b(delay_add_ln22_unr2_stage2_stallmux_q_27_), .o(n_2874) );
no02s01 g778371 ( .a(n_2685), .b(n_1031), .o(n_2797) );
in01s01 g778372 ( .a(n_2947), .o(n_2791) );
no02s01 g778373 ( .a(n_2751), .b(n_2114), .o(n_2947) );
in01s01 g778374 ( .a(n_2770), .o(n_2771) );
no02s01 g778375 ( .a(n_2731), .b(n_3532), .o(n_2770) );
na02s01 g778376 ( .a(n_2508), .b(n_2477), .o(n_2478) );
na02s02 g778378 ( .a(n_2453), .b(n_2206), .o(n_2469) );
no02s03 g778379 ( .a(n_2510), .b(n_2404), .o(n_2561) );
na02s01 g778380 ( .a(n_2538), .b(FE_OFN321_n_2929), .o(n_2539) );
no02m06 TIMEBOOST_cell_2903 ( .a(n_33508), .b(TIMEBOOST_net_742), .o(n_33595) );
in01s01 g778383 ( .a(n_47024), .o(n_2869) );
no02s02 g778385 ( .a(n_2430), .b(n_2442), .o(n_2443) );
in01s01 g778386 ( .a(n_2840), .o(n_2841) );
no02s02 g778388 ( .a(n_2467), .b(n_2466), .o(n_2573) );
na02s02 g778389 ( .a(n_2511), .b(FE_OCPN1632_n_1835), .o(n_2626) );
ao12s01 g778390 ( .a(n_2751), .b(n_2684), .c(n_2683), .o(n_2796) );
no02s01 TIMEBOOST_cell_3827 ( .a(n_28200), .b(n_28128), .o(TIMEBOOST_net_1004) );
na02s02 TIMEBOOST_cell_6001 ( .a(n_18043), .b(n_17918), .o(TIMEBOOST_net_1852) );
na02s01 g778393 ( .a(n_2446), .b(n_2445), .o(n_2447) );
na02s03 g778394 ( .a(n_2512), .b(n_1836), .o(n_2627) );
in01s01 g778395 ( .a(n_2505), .o(n_2506) );
na02s02 g778396 ( .a(n_2467), .b(n_2466), .o(n_2505) );
no02s01 g778397 ( .a(n_2488), .b(n_2487), .o(n_2489) );
na02s02 g778398 ( .a(n_2457), .b(n_2463), .o(n_2464) );
oa12f08 g778400 ( .a(n_2049), .b(n_45488), .c(n_2017), .o(n_2528) );
na02m04 g778402 ( .a(n_2538), .b(n_2412), .o(n_2604) );
na02m08 g778404 ( .a(n_2502), .b(n_2436), .o(n_2537) );
ao22s04 g778406 ( .a(FE_OCP_RBN4118_n_45487), .b(n_2069), .c(n_45487), .d(n_2068), .o(n_3217) );
oa22s01 g778407 ( .a(n_2410), .b(n_2461), .c(n_2475), .d(n_2442), .o(n_2554) );
ao22s01 g778409 ( .a(n_2458), .b(n_2492), .c(n_2520), .d(n_2463), .o(n_2599) );
in01s01 g778410 ( .a(n_2664), .o(n_3274) );
oa12s02 g778411 ( .a(n_2429), .b(n_2428), .c(n_2427), .o(n_2664) );
na02s01 TIMEBOOST_cell_4133 ( .a(n_36306), .b(n_36305), .o(TIMEBOOST_net_1157) );
no02s01 g778413 ( .a(n_2684), .b(n_2683), .o(n_2751) );
in01s01 g778414 ( .a(n_2786), .o(n_2787) );
no02s01 g778415 ( .a(n_2722), .b(n_2137), .o(n_2786) );
in01s01 g778417 ( .a(n_2790), .o(n_3592) );
na02s01 g778418 ( .a(n_2672), .b(delay_add_ln22_unr2_stage2_stallmux_q_26_), .o(n_2790) );
in01s01 g778419 ( .a(n_2728), .o(n_3594) );
no02s01 g778420 ( .a(n_2672), .b(delay_add_ln22_unr2_stage2_stallmux_q_26_), .o(n_2728) );
na02s01 g778422 ( .a(n_2602), .b(n_2666), .o(n_2695) );
in01s01 g778423 ( .a(n_2731), .o(n_3483) );
no02s01 g778424 ( .a(n_2616), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_26_), .o(n_2731) );
na02s01 g778425 ( .a(n_2428), .b(n_2427), .o(n_2429) );
in01s01 g778426 ( .a(n_2663), .o(n_3532) );
na02s01 g778427 ( .a(n_2616), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_26_), .o(n_2663) );
no02s02 g778429 ( .a(n_2734), .b(n_2657), .o(n_2764) );
na02s01 g778431 ( .a(n_2735), .b(n_2643), .o(n_2687) );
no02s04 g778433 ( .a(FE_OCP_RBN2573_n_2558), .b(FE_OCP_RBN6610_n_2289), .o(n_2565) );
no02s02 g778434 ( .a(n_3127), .b(FE_OCP_RBN6610_n_2289), .o(n_2563) );
no02s01 g778435 ( .a(n_2479), .b(n_2378), .o(n_2480) );
no02m06 TIMEBOOST_cell_4132 ( .a(TIMEBOOST_net_1156), .b(FE_OCP_RBN6118_n_5555), .o(n_5750) );
na02f20 TIMEBOOST_cell_7433 ( .a(TIMEBOOST_net_2347), .b(FE_RN_644_0), .o(n_23044) );
no02f08 TIMEBOOST_cell_2899 ( .a(n_13413), .b(TIMEBOOST_net_740), .o(n_13459) );
no02s01 TIMEBOOST_cell_2856 ( .a(n_37293), .b(n_37247), .o(TIMEBOOST_net_719) );
ao12s01 g778443 ( .a(n_2935), .b(n_2876), .c(n_3297), .o(n_3465) );
oa12s01 g778444 ( .a(n_2882), .b(n_2878), .c(FE_OFN4764_n_3029), .o(n_3525) );
no02m06 g778446 ( .a(n_2460), .b(n_2341), .o(n_2538) );
in01m04 g778447 ( .a(n_2453), .o(n_2502) );
no02f02 TIMEBOOST_cell_4107 ( .a(n_15652), .b(n_14419), .o(TIMEBOOST_net_1144) );
na02s04 TIMEBOOST_cell_8805 ( .a(TIMEBOOST_net_2889), .b(n_15730), .o(n_15795) );
no02s01 TIMEBOOST_cell_4971 ( .a(TIMEBOOST_net_1433), .b(n_33459), .o(TIMEBOOST_net_228) );
ao12s01 g778453 ( .a(n_2398), .b(n_2397), .c(n_2396), .o(n_3771) );
in01s01 g778454 ( .a(n_2685), .o(n_2686) );
oa22s01 g778455 ( .a(n_2629), .b(n_2145), .c(n_2556), .d(n_2146), .o(n_2685) );
in01s02 g778456 ( .a(n_2511), .o(n_2512) );
na02m06 TIMEBOOST_cell_2807 ( .a(TIMEBOOST_net_694), .b(n_1699), .o(n_1795) );
ao12s01 g778458 ( .a(n_2407), .b(n_2406), .c(n_2405), .o(n_2488) );
no03f06 TIMEBOOST_cell_8325 ( .a(n_19511), .b(FE_OCP_RBN3717_n_19535), .c(n_19564), .o(n_19688) );
oa12s01 g778460 ( .a(n_2345), .b(n_2344), .c(n_2343), .o(n_2446) );
oa22s01 g778461 ( .a(n_2694), .b(n_2124), .c(n_2614), .d(n_2125), .o(n_2782) );
no02s02 g778463 ( .a(n_2109), .b(n_2694), .o(n_2722) );
na02s01 g778464 ( .a(n_2344), .b(n_2343), .o(n_2345) );
no02s02 g778465 ( .a(n_2126), .b(n_2629), .o(n_2684) );
in01s01 g778466 ( .a(n_2601), .o(n_2602) );
no02s01 g778467 ( .a(n_2570), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_25_), .o(n_2601) );
no02s02 g778468 ( .a(n_2628), .b(delay_add_ln22_unr2_stage2_stallmux_q_25_), .o(n_2734) );
in01s01 g778469 ( .a(n_2640), .o(n_2641) );
na02s01 g778470 ( .a(n_2542), .b(n_2582), .o(n_2640) );
na02s01 g778471 ( .a(n_2570), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_25_), .o(n_2666) );
in01s01 g778472 ( .a(n_2656), .o(n_2657) );
na02s02 g778473 ( .a(n_2628), .b(delay_add_ln22_unr2_stage2_stallmux_q_25_), .o(n_2656) );
in01s01 g778474 ( .a(n_2681), .o(n_2682) );
na02s01 g778475 ( .a(n_2658), .b(n_2630), .o(n_2681) );
na02s01 TIMEBOOST_cell_4130 ( .a(TIMEBOOST_net_1155), .b(n_35856), .o(n_35976) );
no02s01 g778478 ( .a(n_2397), .b(n_2396), .o(n_2398) );
na02s02 g778479 ( .a(n_2340), .b(FE_OCP_RBN5566_n_2346), .o(n_2347) );
na02s01 g778482 ( .a(n_2878), .b(FE_OCP_RBN2627_n_2737), .o(n_2882) );
no02s02 g778483 ( .a(n_2431), .b(n_2348), .o(n_2479) );
no02s01 g778484 ( .a(n_2876), .b(FE_OCP_RBN5660_n_2438), .o(n_2935) );
na02s06 g778486 ( .a(n_3058), .b(FE_OCP_RBN6606_n_2289), .o(n_2543) );
no03s20 TIMEBOOST_cell_8183 ( .a(FE_OCPN1342_n_11927), .b(n_11919), .c(FE_OCPN1651_n_11918), .o(n_12026) );
na02m02 TIMEBOOST_cell_8798 ( .a(n_24751), .b(FE_OCPN1354_n_22484), .o(TIMEBOOST_net_2886) );
no02s01 TIMEBOOST_cell_2857 ( .a(TIMEBOOST_net_719), .b(n_37543), .o(TIMEBOOST_net_236) );
ao12s02 g778490 ( .a(n_3229), .b(n_2549), .c(FE_OCP_RBN6606_n_2289), .o(n_2735) );
ao12m08 g778492 ( .a(n_2061), .b(n_2369), .c(n_2032), .o(n_2428) );
no02s01 g778493 ( .a(n_2406), .b(n_2405), .o(n_2407) );
na02s06 TIMEBOOST_cell_2855 ( .a(TIMEBOOST_net_718), .b(n_37563), .o(n_37607) );
no02m08 g778498 ( .a(n_2340), .b(n_2282), .o(n_2419) );
in01m04 g778499 ( .a(n_2433), .o(n_2460) );
no02s04 g778500 ( .a(n_2392), .b(n_2290), .o(n_2433) );
oa12s01 g778502 ( .a(n_2817), .b(n_2834), .c(n_2768), .o(n_2880) );
in01s01 g778503 ( .a(n_2520), .o(n_2458) );
no02s04 g778504 ( .a(n_2373), .b(n_2336), .o(n_2520) );
oa12s02 g778506 ( .a(n_2352), .b(n_2369), .c(n_2351), .o(n_2558) );
in01s01 g778507 ( .a(n_3127), .o(n_2393) );
ao12s02 g778508 ( .a(n_2319), .b(n_2318), .c(n_2317), .o(n_3127) );
oa22s01 g778509 ( .a(n_2296), .b(n_2360), .c(n_2295), .d(n_2359), .o(n_3721) );
na03s08 TIMEBOOST_cell_5842 ( .a(n_43046), .b(n_43192), .c(n_43053), .o(TIMEBOOST_net_1649) );
in01s01 g778511 ( .a(n_2475), .o(n_2410) );
no02s04 g778512 ( .a(n_2323), .b(n_2310), .o(n_2475) );
ao22s01 g778513 ( .a(n_2516), .b(n_2116), .c(n_2465), .d(n_2117), .o(n_2616) );
oa22s01 g778514 ( .a(n_2608), .b(n_2090), .c(n_2530), .d(n_2091), .o(n_2672) );
no02s01 g778515 ( .a(n_2521), .b(n_3286), .o(n_2522) );
na02s01 g778516 ( .a(n_2484), .b(n_2483), .o(n_2582) );
in01s01 g778517 ( .a(n_2594), .o(n_2595) );
na02s02 g778518 ( .a(n_2569), .b(n_2500), .o(n_2594) );
in01s01 g778519 ( .a(n_2541), .o(n_2542) );
no02s01 g778520 ( .a(n_2484), .b(n_2483), .o(n_2541) );
in01s02 g778521 ( .a(n_2614), .o(n_2694) );
no02s02 g778522 ( .a(n_2608), .b(n_2083), .o(n_2614) );
in01s01 g778523 ( .a(n_2566), .o(n_2567) );
no02s01 g778524 ( .a(n_2546), .b(n_2521), .o(n_2566) );
na02s01 g778525 ( .a(n_2369), .b(n_2351), .o(n_2352) );
in01s01 g778526 ( .a(n_2630), .o(n_2631) );
na02s01 g778527 ( .a(n_2551), .b(delay_add_ln22_unr2_stage2_stallmux_q_24_), .o(n_2630) );
no02s01 g778528 ( .a(n_2318), .b(n_2317), .o(n_2319) );
in01s01 g778529 ( .a(n_2556), .o(n_2629) );
no02s01 g778530 ( .a(n_2108), .b(n_2516), .o(n_2556) );
na02s02 g778531 ( .a(n_2550), .b(n_1197), .o(n_2658) );
in01s01 g778532 ( .a(n_2729), .o(n_2730) );
na02s01 g778533 ( .a(n_2618), .b(n_2701), .o(n_2729) );
na02s01 g778534 ( .a(n_2954), .b(n_2814), .o(n_3397) );
no02s01 g778536 ( .a(n_2937), .b(n_2842), .o(n_3448) );
na02s01 g778537 ( .a(n_2769), .b(n_2817), .o(n_3353) );
na02m02 g778538 ( .a(FE_OCP_RBN6606_n_2289), .b(n_3084), .o(n_2548) );
no02s02 g778539 ( .a(n_2278), .b(n_2031), .o(n_2323) );
no02s02 g778540 ( .a(n_2299), .b(n_2766), .o(n_2310) );
no02s02 g778541 ( .a(n_2321), .b(n_2717), .o(n_2373) );
no02s02 g778542 ( .a(n_2335), .b(n_2237), .o(n_2336) );
in01s01 g778543 ( .a(n_2332), .o(n_2397) );
na02m06 TIMEBOOST_cell_6683 ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .b(FE_OCP_RBN4192_n_38537), .o(TIMEBOOST_net_2099) );
no02s03 g778545 ( .a(n_2307), .b(n_2348), .o(n_2349) );
oa12s01 g778546 ( .a(n_2720), .b(n_3297), .c(n_2744), .o(n_3489) );
ao12s01 g778547 ( .a(n_2617), .b(FE_OFN798_n_2620), .c(FE_OFN4764_n_3029), .o(n_3434) );
in01s01 g778549 ( .a(n_2374), .o(n_2375) );
oa12s01 g778550 ( .a(n_2331), .b(n_2533), .c(n_2330), .o(n_2374) );
ao12s01 g778551 ( .a(FE_OCP_RBN6610_n_2289), .b(n_2710), .c(n_2577), .o(n_3229) );
in01s01 g778552 ( .a(n_2340), .o(n_2320) );
na02m06 g778553 ( .a(n_2233), .b(n_2299), .o(n_2340) );
in01s01 g778554 ( .a(n_2392), .o(n_2361) );
na02s06 g778555 ( .a(n_2238), .b(n_2335), .o(n_2392) );
no02s02 g778556 ( .a(n_2456), .b(n_2350), .o(n_2501) );
oa12s02 g778557 ( .a(FE_OCP_RBN4072_n_2289), .b(n_2269), .c(n_1871), .o(n_2431) );
oa12s01 g778558 ( .a(n_2497), .b(n_2514), .c(n_2496), .o(n_2628) );
ao12s01 g778560 ( .a(n_2440), .b(n_2441), .c(n_2439), .o(n_2570) );
in01s01 g778561 ( .a(n_3058), .o(n_3125) );
oa12s02 g778562 ( .a(n_2304), .b(n_2303), .c(n_2302), .o(n_3058) );
in01s01 g778563 ( .a(n_2342), .o(n_2406) );
in01s01 g778565 ( .a(FE_OFN797_n_2285), .o(n_2876) );
ao22s01 g778566 ( .a(n_2213), .b(n_1489), .c(n_2212), .d(n_1490), .o(n_2285) );
ao22s01 g778567 ( .a(n_2251), .b(n_1488), .c(n_2252), .d(n_1487), .o(n_2878) );
na02s01 g778568 ( .a(n_2514), .b(n_2496), .o(n_2497) );
no02s01 g778569 ( .a(n_2441), .b(n_2439), .o(n_2440) );
in01s01 g778570 ( .a(n_2503), .o(n_2504) );
na02s01 g778571 ( .a(n_3245), .b(n_2422), .o(n_2503) );
in01s01 g778572 ( .a(n_2465), .o(n_2516) );
no02s01 g778573 ( .a(n_2082), .b(n_2441), .o(n_2465) );
in01s01 g778574 ( .a(n_2499), .o(n_2500) );
no02s02 g778575 ( .a(n_2476), .b(delay_add_ln22_unr2_stage2_stallmux_q_23_), .o(n_2499) );
na02s01 g778576 ( .a(n_2303), .b(n_2302), .o(n_2304) );
no02s01 g778577 ( .a(n_2420), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_23_), .o(n_2546) );
in01s01 g778578 ( .a(n_2485), .o(n_2486) );
na02s01 g778579 ( .a(n_2416), .b(n_3317), .o(n_2485) );
na02s02 g778580 ( .a(n_2476), .b(delay_add_ln22_unr2_stage2_stallmux_q_23_), .o(n_2569) );
na02m08 g778581 ( .a(n_2303), .b(n_1965), .o(n_2369) );
no02s01 g778582 ( .a(n_2421), .b(n_1174), .o(n_2521) );
in01s02 g778583 ( .a(n_2530), .o(n_2608) );
no02s02 g778584 ( .a(n_2514), .b(n_2073), .o(n_2530) );
in01s01 g778585 ( .a(n_2712), .o(n_2706) );
no02s01 g778586 ( .a(n_2591), .b(n_2651), .o(n_2712) );
na02s02 g778587 ( .a(n_2325), .b(n_2306), .o(n_2307) );
in01s01 g778589 ( .a(n_2732), .o(n_2733) );
na02s01 g778590 ( .a(n_2639), .b(n_2710), .o(n_2732) );
no02s01 g778591 ( .a(n_2534), .b(n_2533), .o(n_2844) );
na02s01 g778592 ( .a(n_2384), .b(n_2423), .o(n_2691) );
na02s01 g778593 ( .a(n_2326), .b(n_2325), .o(n_2574) );
no02s01 g778594 ( .a(n_2449), .b(n_2448), .o(n_2985) );
no02s01 g778595 ( .a(n_2366), .b(n_44344), .o(n_2477) );
na02s01 g778596 ( .a(n_2825), .b(n_2758), .o(n_3314) );
no02s02 TIMEBOOST_cell_8674 ( .a(n_36515), .b(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_2824) );
no02s01 g778598 ( .a(n_2652), .b(n_3108), .o(n_3087) );
no02s01 g778599 ( .a(n_2705), .b(n_2803), .o(n_3351) );
na02s02 g778600 ( .a(n_2402), .b(n_2423), .o(n_2424) );
na02s01 g778602 ( .a(FE_OCP_RBN6611_n_2289), .b(n_2744), .o(n_2720) );
no02s01 g778603 ( .a(n_2652), .b(n_2612), .o(n_2655) );
na02s01 g778604 ( .a(n_2701), .b(n_2643), .o(n_3305) );
no02s01 g778605 ( .a(n_2654), .b(n_2661), .o(n_3280) );
na02s02 TIMEBOOST_cell_6707 ( .a(n_13530), .b(n_13535), .o(TIMEBOOST_net_2111) );
na02s01 g778607 ( .a(n_2259), .b(n_2261), .o(n_2396) );
in01s01 g778608 ( .a(n_2877), .o(n_2842) );
na02s01 g778609 ( .a(n_2913), .b(n_2807), .o(n_2877) );
na02s02 g778610 ( .a(n_2388), .b(n_2452), .o(n_2456) );
na02s01 g778612 ( .a(FE_OCP_RBN5655_n_2438), .b(FE_OFN796_n_2719), .o(n_2817) );
na02s01 g778613 ( .a(n_2491), .b(n_2140), .o(n_2549) );
na02s01 g778615 ( .a(FE_OCP_RBN5660_n_2438), .b(n_2752), .o(n_2814) );
no02s01 g778616 ( .a(n_2350), .b(n_2330), .o(n_2959) );
no02s01 g778617 ( .a(n_2635), .b(n_2634), .o(n_2990) );
no02s01 g778618 ( .a(n_2592), .b(n_2545), .o(n_3071) );
in01s01 g778619 ( .a(n_2295), .o(n_2296) );
no02s01 g778620 ( .a(n_2273), .b(n_2266), .o(n_2295) );
na02s02 g778621 ( .a(FE_OCP_RBN6606_n_2289), .b(n_2473), .o(n_2474) );
na02s01 g778622 ( .a(n_2544), .b(n_2571), .o(n_2603) );
in01s01 g778623 ( .a(n_2768), .o(n_2769) );
no02s01 g778624 ( .a(FE_OCP_RBN5655_n_2438), .b(FE_OFN796_n_2719), .o(n_2768) );
na02s01 g778625 ( .a(n_2391), .b(n_2452), .o(n_3044) );
in01s01 g778626 ( .a(n_2617), .o(n_2618) );
no02s01 g778627 ( .a(FE_OFN798_n_2620), .b(FE_OCP_RBN6615_n_2289), .o(n_2617) );
na02s01 g778628 ( .a(n_2745), .b(n_2744), .o(n_2746) );
in01s01 g778629 ( .a(n_2900), .o(n_2954) );
no02s01 g778630 ( .a(FE_OCP_RBN5660_n_2438), .b(n_2752), .o(n_2900) );
na02s01 g778631 ( .a(n_2402), .b(n_2322), .o(n_2714) );
na02s01 g778632 ( .a(n_2613), .b(n_2736), .o(n_3156) );
no02s01 g778633 ( .a(n_2807), .b(n_2913), .o(n_2937) );
ao12s01 g778636 ( .a(n_2660), .b(FE_OFN4764_n_3029), .c(n_2611), .o(n_3453) );
oa12s01 g778637 ( .a(n_2590), .b(n_3297), .c(n_2577), .o(n_3409) );
oa12s01 g778638 ( .a(n_2306), .b(n_3082), .c(n_2255), .o(n_3207) );
in01s01 g778639 ( .a(n_2299), .o(n_2278) );
no02m06 g778640 ( .a(n_2249), .b(n_2211), .o(n_2299) );
in01s01 g778641 ( .a(n_2335), .o(n_2321) );
no02m06 g778642 ( .a(n_2293), .b(n_2219), .o(n_2335) );
in01s01 g778643 ( .a(n_3084), .o(n_2294) );
oa12m01 g778644 ( .a(n_2241), .b(n_2240), .c(n_2239), .o(n_3084) );
in01s01 g778645 ( .a(n_2550), .o(n_2551) );
ao22s01 g778646 ( .a(n_2455), .b(n_2047), .c(n_2434), .d(n_2046), .o(n_2550) );
oa22s01 g778647 ( .a(n_2370), .b(n_2070), .c(n_2382), .d(n_2071), .o(n_2484) );
in01s01 g778648 ( .a(n_2422), .o(n_3286) );
na02s01 g778649 ( .a(n_2387), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_22_), .o(n_2422) );
na02s01 g778650 ( .a(n_2382), .b(n_2027), .o(n_2441) );
na02s04 g778651 ( .a(n_2455), .b(n_2012), .o(n_2514) );
na02s01 g778652 ( .a(n_2380), .b(n_2379), .o(n_3317) );
in01s01 g778653 ( .a(n_2450), .o(n_2451) );
na02s01 g778654 ( .a(n_2368), .b(n_2413), .o(n_2450) );
in01s01 g778655 ( .a(n_2437), .o(n_3245) );
no02s01 g778656 ( .a(n_2387), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_22_), .o(n_2437) );
in01s01 g778657 ( .a(n_3319), .o(n_2416) );
no02s01 g778658 ( .a(n_2380), .b(n_2379), .o(n_3319) );
in01s01 g778659 ( .a(n_2425), .o(n_2426) );
na02s01 g778660 ( .a(n_2385), .b(n_2386), .o(n_2425) );
na02s01 g778661 ( .a(n_2240), .b(n_2239), .o(n_2241) );
in01s01 g778662 ( .a(n_2544), .o(n_2545) );
na02s01 g778663 ( .a(FE_OCP_RBN6610_n_2289), .b(n_2515), .o(n_2544) );
na02s02 g778664 ( .a(FE_OCP_RBN5596_n_45903), .b(n_2237), .o(n_2238) );
na02s01 g778665 ( .a(FE_OCP_RBN5597_n_45903), .b(n_2250), .o(n_2325) );
no02m02 g778666 ( .a(n_45903), .b(n_1565), .o(n_2273) );
in01s01 g778667 ( .a(n_2592), .o(n_2593) );
no02s01 g778668 ( .a(FE_OCP_RBN6610_n_2289), .b(n_2515), .o(n_2592) );
no02s01 g778669 ( .a(n_2289), .b(n_2858), .o(n_2341) );
in01s01 g778670 ( .a(n_2348), .o(n_2322) );
no02s02 g778671 ( .a(n_2289), .b(n_2292), .o(n_2348) );
no02s01 g778672 ( .a(FE_OCP_RBN6614_n_2289), .b(n_2611), .o(n_2660) );
in01s01 g778673 ( .a(n_2306), .o(n_2274) );
na02s01 g778674 ( .a(FE_OCP_RBN5597_n_45903), .b(n_2255), .o(n_2306) );
na02s01 g778675 ( .a(FE_OCP_RBN4071_n_2289), .b(n_2929), .o(n_2412) );
in01s01 g778676 ( .a(n_2331), .o(n_2350) );
na02s01 g778677 ( .a(n_2277), .b(n_2270), .o(n_2331) );
no02s01 g778678 ( .a(FE_OCP_RBN6606_n_2289), .b(n_2472), .o(n_2661) );
in01s01 g778679 ( .a(n_2449), .o(n_2388) );
no02s01 g778680 ( .a(FE_OCP_RBN4072_n_2289), .b(n_2363), .o(n_2449) );
in01s02 g778681 ( .a(n_2249), .o(n_2230) );
no02s06 g778682 ( .a(n_45903), .b(n_2606), .o(n_2249) );
no02s02 g778683 ( .a(FE_OCP_RBN6606_n_2289), .b(n_2540), .o(n_2634) );
in01s01 g778684 ( .a(n_2651), .o(n_2639) );
no02s01 g778685 ( .a(FE_OCP_RBN6606_n_2289), .b(FE_OFN4807_n_2432), .o(n_2651) );
na02s02 g778687 ( .a(n_2277), .b(n_2276), .o(n_2308) );
in01s01 g778688 ( .a(n_2745), .o(n_2705) );
na02s01 g778689 ( .a(FE_OCP_RBN6616_n_2289), .b(FE_OFN799_n_2644), .o(n_2745) );
na02s02 g778690 ( .a(FE_OCP_RBN6606_n_2289), .b(n_2596), .o(n_2736) );
in01s01 g778691 ( .a(n_2590), .o(n_2591) );
na02s01 g778692 ( .a(FE_OCP_RBN6610_n_2289), .b(n_2577), .o(n_2590) );
no02s06 g778693 ( .a(n_2289), .b(FE_OCP_RBN5567_n_2346), .o(n_2282) );
in01s01 g778694 ( .a(n_2571), .o(n_2635) );
na02s01 g778695 ( .a(FE_OCP_RBN6606_n_2289), .b(n_2540), .o(n_2571) );
no02s01 g778696 ( .a(FE_OCP_RBN5597_n_45903), .b(n_1887), .o(n_2533) );
na02s04 g778698 ( .a(FE_OCP_RBN5595_n_45903), .b(n_2766), .o(n_2233) );
in01s01 g778699 ( .a(n_2652), .o(n_2589) );
no02s01 g778700 ( .a(FE_OCP_RBN6610_n_2289), .b(FE_OFN793_n_2056), .o(n_2652) );
na02s02 g778701 ( .a(FE_OCP_RBN4072_n_2289), .b(n_2364), .o(n_2423) );
in01s01 g778702 ( .a(n_2258), .o(n_2259) );
no02s02 g778703 ( .a(FE_OCP_RBN5594_n_45903), .b(n_2234), .o(n_2258) );
na02s01 g778704 ( .a(FE_OCP_RBN6611_n_2289), .b(n_2562), .o(n_2701) );
in01s01 g778705 ( .a(n_2383), .o(n_2384) );
no02s01 g778706 ( .a(FE_OCP_RBN4072_n_2289), .b(n_2364), .o(n_2383) );
no02s02 g778707 ( .a(FE_OCP_RBN6610_n_2289), .b(n_3039), .o(n_2498) );
na02s01 g778708 ( .a(FE_OCP_RBN4074_n_2289), .b(FE_OFN4807_n_2432), .o(n_2710) );
na02m06 TIMEBOOST_cell_4106 ( .a(TIMEBOOST_net_1143), .b(n_39744), .o(n_39749) );
in01s01 g778710 ( .a(n_2389), .o(n_2448) );
na02s02 g778711 ( .a(FE_OCP_RBN4072_n_2289), .b(n_2363), .o(n_2389) );
no02s02 g778712 ( .a(FE_OCP_RBN6606_n_2289), .b(n_2057), .o(n_3108) );
in01s01 g778713 ( .a(n_2452), .o(n_2404) );
na02s01 g778714 ( .a(FE_OCP_RBN4072_n_2289), .b(n_2357), .o(n_2452) );
in01s01 g778715 ( .a(n_2491), .o(n_2654) );
na02s01 g778716 ( .a(FE_OCP_RBN6606_n_2289), .b(n_2472), .o(n_2491) );
in01s04 g778717 ( .a(n_2245), .o(n_2293) );
na02s08 g778718 ( .a(FE_OCP_RBN5596_n_45903), .b(n_2494), .o(n_2245) );
no02s02 g778719 ( .a(n_2277), .b(n_2276), .o(n_2366) );
in01s01 g778720 ( .a(n_2390), .o(n_2391) );
no02s01 g778721 ( .a(FE_OCP_RBN4072_n_2289), .b(n_2357), .o(n_2390) );
na02s03 g778722 ( .a(FE_OCP_RBN4071_n_2289), .b(n_2898), .o(n_2436) );
no02s02 g778723 ( .a(n_2289), .b(n_2288), .o(n_2290) );
no02s02 g778724 ( .a(n_1888), .b(FE_OCP_RBN6606_n_2289), .o(n_2534) );
no02s02 g778725 ( .a(n_45903), .b(n_2218), .o(n_2219) );
no02s01 g778726 ( .a(FE_OCP_RBN5648_n_2438), .b(FE_OFN799_n_2644), .o(n_2803) );
in01s01 g778727 ( .a(n_2269), .o(n_2326) );
no02s02 g778728 ( .a(n_2215), .b(n_2250), .o(n_2269) );
no02s01 g778729 ( .a(n_2277), .b(n_2270), .o(n_2330) );
in01s01 g778730 ( .a(n_2838), .o(n_2825) );
no02s01 g778731 ( .a(FE_OCP_RBN5654_n_2438), .b(n_2738), .o(n_2838) );
na02s02 g778733 ( .a(FE_OCP_RBN5595_n_45903), .b(n_2234), .o(n_2261) );
in01s01 g778734 ( .a(n_2612), .o(n_2613) );
no02s01 g778735 ( .a(FE_OCP_RBN6606_n_2289), .b(n_2596), .o(n_2612) );
no02s04 g778736 ( .a(n_45903), .b(n_2702), .o(n_2211) );
in01s01 g778737 ( .a(n_2609), .o(n_2643) );
no02s01 g778738 ( .a(FE_OCP_RBN6610_n_2289), .b(n_2562), .o(n_2609) );
in01s01 g778739 ( .a(n_2758), .o(n_2834) );
na02s01 g778740 ( .a(FE_OCP_RBN5654_n_2438), .b(n_2738), .o(n_2758) );
in01s01 g778741 ( .a(n_2402), .o(n_2378) );
na02s01 g778742 ( .a(n_2289), .b(n_2292), .o(n_2402) );
no02m08 TIMEBOOST_cell_8729 ( .a(TIMEBOOST_net_2851), .b(n_40913), .o(n_40926) );
in01s01 g778744 ( .a(n_2251), .o(n_2252) );
ao12s01 g778745 ( .a(n_1415), .b(n_2225), .c(n_1479), .o(n_2251) );
in01s01 g778746 ( .a(n_2212), .o(n_2213) );
ao12s01 g778747 ( .a(n_1470), .b(n_2200), .c(n_1423), .o(n_2212) );
oa22s01 g778748 ( .a(n_2338), .b(n_2029), .c(n_2381), .d(n_2028), .o(n_2476) );
oa22s01 g778749 ( .a(n_2191), .b(n_1499), .c(n_2225), .d(n_1500), .o(n_2807) );
in01s01 g778750 ( .a(n_2420), .o(n_2421) );
ao12s01 g778751 ( .a(n_2355), .b(n_2354), .c(n_2353), .o(n_2420) );
in01s01 g778752 ( .a(n_2473), .o(n_3023) );
oa12s01 g778753 ( .a(n_2223), .b(n_2222), .c(n_2221), .o(n_2473) );
ao12s01 g778754 ( .a(n_2185), .b(n_2184), .c(n_2183), .o(n_2719) );
oa22s01 g778755 ( .a(n_2169), .b(n_1505), .c(n_2200), .d(n_1504), .o(n_2752) );
oa22s01 g778756 ( .a(n_2170), .b(n_1772), .c(n_2171), .d(n_1771), .o(n_2620) );
ao22s01 g778757 ( .a(n_2167), .b(n_1798), .c(n_2166), .d(n_1799), .o(n_2744) );
no02s01 g778758 ( .a(n_2354), .b(n_2353), .o(n_2355) );
na02s01 g778759 ( .a(n_2298), .b(n_1177), .o(n_2385) );
na02s02 g778760 ( .a(n_2327), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_21_), .o(n_2413) );
in01s01 g778761 ( .a(n_2455), .o(n_2434) );
no02s03 g778762 ( .a(n_2381), .b(n_2021), .o(n_2455) );
in01s01 g778763 ( .a(n_2382), .o(n_2370) );
no02s02 g778764 ( .a(n_2354), .b(n_2030), .o(n_2382) );
na02s01 TIMEBOOST_cell_4413 ( .a(FE_OFN4776_n_44463), .b(n_44492), .o(TIMEBOOST_net_1297) );
na02s01 g778767 ( .a(n_45317), .b(n_2358), .o(n_2408) );
in01s01 g778768 ( .a(n_2328), .o(n_2329) );
no02s01 g778769 ( .a(n_2272), .b(n_2313), .o(n_2328) );
no02s01 g778770 ( .a(n_2184), .b(n_2183), .o(n_2185) );
na02s01 g778771 ( .a(n_2297), .b(delay_add_ln22_unr2_stage2_stallmux_q_21_), .o(n_2386) );
in01s01 g778772 ( .a(n_2367), .o(n_2368) );
no02s02 g778773 ( .a(n_2327), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_21_), .o(n_2367) );
na02s01 g778774 ( .a(n_2222), .b(n_2221), .o(n_2223) );
oa12f08 g778776 ( .a(n_1935), .b(n_2189), .c(n_1903), .o(n_2240) );
in01s01 g778777 ( .a(FE_OCP_RBN5596_n_45903), .o(n_2215) );
in01s02 g778808 ( .a(n_3106), .o(n_4093) );
in01s02 g778811 ( .a(n_3106), .o(n_3862) );
in01s06 g778812 ( .a(n_3615), .o(n_3106) );
in01s06 g778815 ( .a(FE_OFN4763_n_3029), .o(n_3615) );
in01s01 g778826 ( .a(FE_OFN4764_n_3029), .o(n_3297) );
in01s03 g778841 ( .a(FE_OFN4764_n_3029), .o(n_3082) );
in01s01 g778851 ( .a(n_2913), .o(n_3029) );
in01s10 g778862 ( .a(FE_OCP_RBN2630_n_2737), .o(n_2913) );
in01m10 g778890 ( .a(n_2277), .o(n_2289) );
in01m10 g778897 ( .a(FE_OCP_RBN5597_n_45903), .o(n_2277) );
oa12s01 g778901 ( .a(n_2178), .b(n_2177), .c(n_2176), .o(n_2644) );
no02s02 g778903 ( .a(n_2190), .b(n_2179), .o(n_3039) );
ao22s01 g778904 ( .a(n_2305), .b(n_2020), .c(n_2279), .d(n_2019), .o(n_2387) );
ao22s01 g778905 ( .a(n_2311), .b(n_2001), .c(n_2268), .d(n_2002), .o(n_2380) );
no02s01 g778906 ( .a(n_2160), .b(n_1956), .o(n_2179) );
na02s01 g778907 ( .a(n_2177), .b(n_2176), .o(n_2178) );
in01m04 g778908 ( .a(n_2338), .o(n_2381) );
no02f06 g778909 ( .a(n_2311), .b(n_1998), .o(n_2338) );
na02s01 g778911 ( .a(n_2324), .b(n_2300), .o(n_2333) );
na02s02 g778912 ( .a(n_2305), .b(n_1973), .o(n_2354) );
no02s02 g778914 ( .a(n_2284), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_20_), .o(n_2314) );
in01s01 g778915 ( .a(n_2271), .o(n_2272) );
na02s02 g778916 ( .a(n_2246), .b(delay_add_ln22_unr2_stage2_stallmux_q_20_), .o(n_2271) );
na02s01 g778918 ( .a(n_2243), .b(n_2265), .o(n_2286) );
na02s02 g778919 ( .a(n_2284), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_20_), .o(n_2358) );
no02s01 g778920 ( .a(n_2189), .b(n_1957), .o(n_2190) );
no02s02 g778921 ( .a(n_2246), .b(delay_add_ln22_unr2_stage2_stallmux_q_20_), .o(n_2313) );
in01s01 g778922 ( .a(n_2191), .o(n_2225) );
na02s01 g778923 ( .a(n_2152), .b(n_1840), .o(n_2191) );
in01s01 g778924 ( .a(n_2166), .o(n_2167) );
ao12s01 g778925 ( .a(n_1749), .b(n_2144), .c(n_1743), .o(n_2166) );
in01s01 g778926 ( .a(n_2169), .o(n_2200) );
oa12s01 g778927 ( .a(n_1781), .b(n_2148), .c(n_1722), .o(n_2169) );
oa12s01 g778928 ( .a(n_1663), .b(n_2148), .c(n_1783), .o(n_2184) );
in01s01 g778929 ( .a(n_2170), .o(n_2171) );
oa12s01 g778930 ( .a(n_1751), .b(n_2143), .c(n_1801), .o(n_2170) );
na03f04 TIMEBOOST_cell_6565 ( .a(n_31233), .b(n_31100), .c(TIMEBOOST_net_955), .o(n_31379) );
oa12s01 g778933 ( .a(n_2121), .b(n_2148), .c(n_2120), .o(n_2738) );
ao12s01 g778934 ( .a(n_2135), .b(n_2143), .c(n_2134), .o(n_2562) );
in01s01 g778935 ( .a(n_2297), .o(n_2298) );
oa22s01 g778936 ( .a(n_2214), .b(n_1984), .c(n_2257), .d(n_1983), .o(n_2297) );
in01s01 g778937 ( .a(n_2898), .o(n_2206) );
oa12s02 g778938 ( .a(n_2157), .b(n_2158), .c(n_2156), .o(n_2898) );
oa12s01 g778939 ( .a(n_2130), .b(n_2129), .c(n_2128), .o(n_2472) );
ao12s01 g778940 ( .a(n_2254), .b(n_2260), .c(n_2253), .o(n_2327) );
no02s01 g778941 ( .a(n_2260), .b(n_2253), .o(n_2254) );
na02s01 g778942 ( .a(n_2158), .b(n_2156), .o(n_2157) );
in01s03 g778943 ( .a(n_2268), .o(n_2311) );
no02s06 g778944 ( .a(n_1971), .b(n_2257), .o(n_2268) );
in01s01 g778945 ( .a(n_2300), .o(n_2301) );
na02s01 g778946 ( .a(n_2229), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_19_), .o(n_2300) );
na02s01 g778948 ( .a(n_2264), .b(n_2263), .o(n_2280) );
no02s01 g778949 ( .a(n_2143), .b(n_2134), .o(n_2135) );
in01s01 g778950 ( .a(n_2305), .o(n_2279) );
no02s04 g778951 ( .a(n_1990), .b(n_2260), .o(n_2305) );
no02f08 TIMEBOOST_cell_5485 ( .a(n_35365), .b(TIMEBOOST_net_1690), .o(n_35401) );
in01s01 g778953 ( .a(n_2243), .o(n_2244) );
na02s01 g778954 ( .a(n_2198), .b(delay_add_ln22_unr2_stage2_stallmux_q_19_), .o(n_2243) );
na02s02 g778955 ( .a(n_2197), .b(n_1101), .o(n_2265) );
na02s02 g778956 ( .a(n_2228), .b(n_1141), .o(n_2324) );
in01s01 g778957 ( .a(n_2247), .o(n_2248) );
na02s01 g778958 ( .a(n_2232), .b(n_2231), .o(n_2247) );
na02s01 g778959 ( .a(n_2129), .b(n_2128), .o(n_2130) );
no02m08 TIMEBOOST_cell_1792 ( .a(TIMEBOOST_net_510), .b(n_6013), .o(n_6059) );
na02s01 g778961 ( .a(n_2148), .b(n_2120), .o(n_2121) );
in01f06 g778962 ( .a(n_2160), .o(n_2189) );
oa12f08 g778963 ( .a(n_1890), .b(FE_OCP_RBN5568_n_2103), .c(n_1856), .o(n_2160) );
in01s01 g778964 ( .a(n_2140), .o(n_2611) );
ao12s01 g778965 ( .a(n_2094), .b(n_2093), .c(n_2092), .o(n_2140) );
oa22s01 g778967 ( .a(n_2103), .b(n_1901), .c(FE_OCP_RBN5569_n_2103), .d(n_1902), .o(n_2929) );
in01s01 g778968 ( .a(n_2151), .o(n_2152) );
ao12s01 g778970 ( .a(n_2133), .b(n_2132), .c(n_2131), .o(n_2577) );
oa22s01 g778971 ( .a(n_2186), .b(n_1961), .c(n_2201), .d(n_1960), .o(n_2246) );
ao22s01 g778972 ( .a(n_2199), .b(n_1996), .c(n_2224), .d(n_1997), .o(n_2284) );
no02s01 g778973 ( .a(n_2101), .b(n_1787), .o(n_2143) );
na02s01 g778974 ( .a(n_2101), .b(n_1741), .o(n_2144) );
na02s02 g778975 ( .a(n_2204), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_18_), .o(n_2263) );
in01s01 g778976 ( .a(n_2216), .o(n_2217) );
na02s02 g778977 ( .a(n_2202), .b(n_2182), .o(n_2216) );
na02s02 g778978 ( .a(n_2205), .b(n_1126), .o(n_2264) );
na02s04 g778979 ( .a(n_2224), .b(n_1946), .o(n_2260) );
na02s01 g778980 ( .a(n_2188), .b(n_1037), .o(n_2231) );
na02s02 g778981 ( .a(n_2187), .b(delay_add_ln22_unr2_stage2_stallmux_q_18_), .o(n_2232) );
in01s01 g778982 ( .a(n_2226), .o(n_2227) );
no02s02 g778983 ( .a(n_2209), .b(n_2208), .o(n_2226) );
in01s02 g778984 ( .a(n_2214), .o(n_2257) );
no02s04 g778985 ( .a(n_2201), .b(n_1947), .o(n_2214) );
no02s01 g778986 ( .a(n_2132), .b(n_2131), .o(n_2133) );
no02s01 g778987 ( .a(n_2093), .b(n_2092), .o(n_2094) );
na02f02 TIMEBOOST_cell_8025 ( .a(TIMEBOOST_net_2643), .b(n_16557), .o(TIMEBOOST_net_1762) );
ao12s01 g778989 ( .a(n_1561), .b(n_2074), .c(n_1516), .o(n_2129) );
in01s01 g778991 ( .a(n_2197), .o(n_2198) );
ao12s01 g778992 ( .a(n_2165), .b(n_2172), .c(n_2164), .o(n_2197) );
in01s01 g778993 ( .a(n_2228), .o(n_2229) );
oa12s01 g778994 ( .a(n_2196), .b(n_2195), .c(n_2194), .o(n_2228) );
in01s01 g778995 ( .a(n_2394), .o(n_2863) );
oa12s02 g778996 ( .a(n_2096), .b(n_2106), .c(n_2095), .o(n_2394) );
na02s01 g778997 ( .a(n_2195), .b(n_2194), .o(n_2196) );
no02s01 g778998 ( .a(n_2077), .b(n_1629), .o(n_2101) );
no02s01 g778999 ( .a(n_2172), .b(n_2164), .o(n_2165) );
na02s02 g779000 ( .a(n_2161), .b(delay_add_ln22_unr2_stage2_stallmux_q_17_), .o(n_2202) );
in01s01 g779001 ( .a(n_2181), .o(n_2182) );
no02s02 g779002 ( .a(n_2161), .b(delay_add_ln22_unr2_stage2_stallmux_q_17_), .o(n_2181) );
in01s02 g779003 ( .a(n_2186), .o(n_2201) );
no02s02 g779004 ( .a(n_2172), .b(n_1930), .o(n_2186) );
in01s01 g779005 ( .a(n_2192), .o(n_2193) );
na02s01 g779006 ( .a(n_2180), .b(n_2142), .o(n_2192) );
no02s02 g779007 ( .a(n_2173), .b(n_1083), .o(n_2208) );
na02s02 TIMEBOOST_cell_8019 ( .a(TIMEBOOST_net_2640), .b(n_11362), .o(TIMEBOOST_net_1756) );
na02s01 g779009 ( .a(n_2077), .b(n_1628), .o(n_2093) );
na02s01 g779010 ( .a(n_2106), .b(n_2095), .o(n_2096) );
no02s02 g779011 ( .a(n_2174), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_17_), .o(n_2209) );
in01s01 g779012 ( .a(n_2224), .o(n_2199) );
no02s04 g779013 ( .a(n_2195), .b(n_1913), .o(n_2224) );
na02s01 g779015 ( .a(FE_RN_824_0), .b(n_2175), .o(n_2698) );
na02s01 g779016 ( .a(n_2075), .b(n_1506), .o(n_2132) );
na02f08 TIMEBOOST_cell_6030 ( .a(TIMEBOOST_net_1866), .b(n_2063), .o(n_2103) );
in01s01 g779019 ( .a(n_2858), .o(n_2102) );
ao12s02 g779020 ( .a(n_2064), .b(n_2063), .c(n_2062), .o(n_2858) );
oa22s01 g779021 ( .a(n_45717), .b(n_1498), .c(n_45716), .d(n_1497), .o(n_2432) );
ao12s01 g779022 ( .a(n_2055), .b(n_2054), .c(n_2053), .o(n_2596) );
in01s01 g779023 ( .a(n_2204), .o(n_2205) );
ao22s01 g779024 ( .a(n_2163), .b(n_1932), .c(n_2147), .d(n_1931), .o(n_2204) );
in01s01 g779025 ( .a(n_2187), .o(n_2188) );
oa22s02 g779026 ( .a(n_2110), .b(n_1917), .c(n_2118), .d(n_1918), .o(n_2187) );
na02s01 g779027 ( .a(n_45717), .b(n_1597), .o(n_2077) );
no02s01 g779028 ( .a(n_2054), .b(n_2053), .o(n_2055) );
in01s01 g779029 ( .a(n_2141), .o(n_2142) );
no02s02 g779030 ( .a(n_2127), .b(delay_add_ln22_unr2_stage2_stallmux_q_16_), .o(n_2141) );
na02s01 g779031 ( .a(n_2119), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_16_), .o(n_2175) );
na02s02 g779032 ( .a(n_2127), .b(delay_add_ln22_unr2_stage2_stallmux_q_16_), .o(n_2180) );
na02s04 g779033 ( .a(n_2163), .b(n_1883), .o(n_2195) );
no02m08 TIMEBOOST_cell_8865 ( .a(TIMEBOOST_net_2919), .b(n_11560), .o(n_11776) );
no02s01 g779035 ( .a(n_2063), .b(n_2062), .o(n_2064) );
in01s01 g779036 ( .a(n_2154), .o(n_2155) );
na02s02 g779037 ( .a(n_2123), .b(FE_OCP_RBN2528_n_2097), .o(n_2154) );
no02s01 g779038 ( .a(n_2153), .b(n_2112), .o(n_2587) );
no02s01 g779040 ( .a(n_2119), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_16_), .o(n_2149) );
na02s02 g779041 ( .a(n_2118), .b(n_1879), .o(n_2172) );
in01s01 g779042 ( .a(n_2074), .o(n_2075) );
no02s01 g779043 ( .a(n_45716), .b(n_1512), .o(n_2074) );
na02m08 g779044 ( .a(n_2044), .b(n_1899), .o(n_2106) );
in01s02 g779045 ( .a(FE_OCP_RBN5566_n_2346), .o(n_2870) );
ao12m01 g779046 ( .a(n_2041), .b(n_2043), .c(n_2040), .o(n_2346) );
in01s01 g779047 ( .a(n_2173), .o(n_2174) );
oa22s02 g779048 ( .a(FE_OCP_RBN5598_n_2100), .b(n_1876), .c(n_2100), .d(n_1877), .o(n_2173) );
oa12s01 g779049 ( .a(n_2089), .b(n_2105), .c(n_2088), .o(n_2161) );
na02s01 g779050 ( .a(n_2105), .b(n_2088), .o(n_2089) );
no02s04 g779052 ( .a(FE_OCP_RBN4053_n_2086), .b(delay_add_ln22_unr2_stage2_stallmux_q_15_), .o(n_2097) );
no02s02 g779053 ( .a(n_2104), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_15_), .o(n_2153) );
na02s08 g779054 ( .a(n_2043), .b(n_1900), .o(n_2044) );
in01s01 g779055 ( .a(n_2163), .o(n_2147) );
no02s04 g779056 ( .a(FE_OCP_RBN5599_n_2100), .b(n_1861), .o(n_2163) );
in01s01 g779057 ( .a(n_2118), .o(n_2110) );
no02s02 g779058 ( .a(n_2105), .b(n_1881), .o(n_2118) );
no02s01 g779059 ( .a(n_2043), .b(n_2040), .o(n_2041) );
na02s02 g779060 ( .a(FE_OCP_RBN4052_n_2086), .b(delay_add_ln22_unr2_stage2_stallmux_q_15_), .o(n_2123) );
na02s01 g779061 ( .a(n_2085), .b(n_2084), .o(n_2518) );
in01s01 g779062 ( .a(n_2111), .o(n_2112) );
na02s02 g779063 ( .a(n_2104), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_15_), .o(n_2111) );
ao12s01 g779064 ( .a(n_1484), .b(n_2023), .c(n_1682), .o(n_2054) );
in01s01 g779066 ( .a(n_2288), .o(n_2794) );
ao12m01 g779067 ( .a(n_2010), .b(n_2009), .c(n_2008), .o(n_2288) );
in01s01 g779068 ( .a(FE_OFN793_n_2056), .o(n_2057) );
ao12s01 g779069 ( .a(n_2014), .b(n_2023), .c(n_2013), .o(n_2056) );
oa22s01 g779072 ( .a(n_1974), .b(n_1779), .c(n_1975), .d(n_1778), .o(n_2515) );
oa22s01 g779073 ( .a(n_2076), .b(n_1830), .c(n_2065), .d(n_1829), .o(n_2127) );
ao22s02 g779074 ( .a(n_2087), .b(n_1854), .c(n_2067), .d(n_1855), .o(n_2119) );
na02s01 g779076 ( .a(FE_OCP_RBN4038_n_2059), .b(n_2081), .o(n_2427) );
na02s04 g779077 ( .a(n_1765), .b(n_2076), .o(n_2105) );
in01s01 g779078 ( .a(n_2068), .o(n_2069) );
na02s02 g779079 ( .a(n_2049), .b(n_2018), .o(n_2068) );
no02s04 g779081 ( .a(n_2087), .b(n_1832), .o(n_2100) );
na02s02 g779082 ( .a(n_2035), .b(delay_add_ln22_unr2_stage2_stallmux_q_14_), .o(n_2085) );
na02s01 g779083 ( .a(n_2034), .b(n_1173), .o(n_2084) );
no02s01 g779084 ( .a(n_2009), .b(n_2008), .o(n_2010) );
no02s01 g779085 ( .a(n_2023), .b(n_2013), .o(n_2014) );
na02s06 g779086 ( .a(n_1988), .b(n_1833), .o(n_2043) );
in01s01 g779087 ( .a(n_2766), .o(n_2031) );
oa12s02 g779088 ( .a(n_1982), .b(n_1987), .c(n_1981), .o(n_2766) );
oa22s01 g779089 ( .a(n_2042), .b(n_1804), .c(n_2024), .d(n_1805), .o(n_2086) );
ao12s02 g779090 ( .a(n_2052), .b(n_2051), .c(n_2050), .o(n_2104) );
no02s02 g779091 ( .a(n_2051), .b(n_2050), .o(n_2052) );
no02s02 g779092 ( .a(n_2061), .b(n_2033), .o(n_2351) );
na02s01 g779093 ( .a(n_2038), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_13_), .o(n_2081) );
na02s02 g779094 ( .a(n_2004), .b(delay_add_ln22_unr2_stage2_stallmux_q_13_), .o(n_2049) );
in01s04 g779095 ( .a(n_2067), .o(n_2087) );
no02s06 g779096 ( .a(n_1797), .b(n_2051), .o(n_2067) );
na02s01 g779097 ( .a(n_1987), .b(n_1981), .o(n_1982) );
na02s01 g779098 ( .a(n_2005), .b(n_1977), .o(n_2317) );
in01s01 g779099 ( .a(n_2017), .o(n_2018) );
no02s02 g779100 ( .a(n_2004), .b(delay_add_ln22_unr2_stage2_stallmux_q_13_), .o(n_2017) );
no02s01 g779102 ( .a(n_2038), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_13_), .o(n_2059) );
in01s01 g779103 ( .a(n_2076), .o(n_2065) );
no02s04 g779104 ( .a(n_2042), .b(n_1770), .o(n_2076) );
na02s06 g779105 ( .a(n_1987), .b(n_1834), .o(n_1988) );
in01s01 g779106 ( .a(n_1974), .o(n_1975) );
oa12s01 g779107 ( .a(n_1794), .b(n_1958), .c(n_1619), .o(n_1974) );
ao12s01 g779109 ( .a(n_1669), .b(n_1964), .c(n_1646), .o(n_2023) );
na02f06 g779110 ( .a(n_1943), .b(n_1815), .o(n_2009) );
oa22s01 g779111 ( .a(n_1958), .b(n_1803), .c(n_1964), .d(n_1802), .o(n_2540) );
in01s01 g779112 ( .a(n_2237), .o(n_2717) );
oa12s01 g779113 ( .a(n_1951), .b(n_1950), .c(n_1949), .o(n_2237) );
in01s01 g779114 ( .a(n_2066), .o(n_2523) );
ao22s02 g779115 ( .a(n_2003), .b(n_1824), .c(n_2025), .d(n_1825), .o(n_2066) );
in01s01 g779116 ( .a(n_2034), .o(n_2035) );
ao22s01 g779117 ( .a(n_1967), .b(n_1774), .c(n_1999), .d(n_1773), .o(n_2034) );
in01s01 g779118 ( .a(n_1976), .o(n_1977) );
no02s01 g779119 ( .a(n_1955), .b(delay_add_ln22_unr2_stage2_stallmux_q_12_), .o(n_1976) );
in01s02 g779120 ( .a(n_2024), .o(n_2042) );
no02s04 g779121 ( .a(n_1759), .b(n_1999), .o(n_2024) );
na02s01 g779122 ( .a(n_1950), .b(n_1949), .o(n_1951) );
na02s01 g779123 ( .a(n_1979), .b(FE_RN_773_0), .o(n_2239) );
na02s06 TIMEBOOST_cell_7949 ( .a(TIMEBOOST_net_2605), .b(n_10877), .o(n_10992) );
na02m06 TIMEBOOST_cell_7090 ( .a(TIMEBOOST_net_2303), .b(n_36593), .o(n_36673) );
in01s01 g779126 ( .a(n_2032), .o(n_2033) );
na02s02 g779127 ( .a(n_2015), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_12_), .o(n_2032) );
na02s01 g779128 ( .a(n_1955), .b(delay_add_ln22_unr2_stage2_stallmux_q_12_), .o(n_2005) );
na02m06 g779129 ( .a(n_1950), .b(n_1814), .o(n_1943) );
no02s02 g779130 ( .a(n_2015), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_12_), .o(n_2061) );
na02s06 g779131 ( .a(n_1704), .b(n_2025), .o(n_2051) );
na02f08 TIMEBOOST_cell_8139 ( .a(TIMEBOOST_net_2700), .b(n_23350), .o(n_23424) );
ao12s01 g779134 ( .a(n_1929), .b(n_1928), .c(n_1927), .o(n_2357) );
in01s01 g779135 ( .a(n_2702), .o(n_1978) );
ao12m01 g779136 ( .a(n_1920), .b(n_1921), .c(n_1919), .o(n_2702) );
oa12s01 g779137 ( .a(n_1942), .b(n_2606), .c(n_1941), .o(n_4117) );
ao12s02 g779138 ( .a(n_1994), .b(n_1993), .c(n_1992), .o(n_2038) );
oa22s02 g779139 ( .a(n_1916), .b(n_1720), .c(n_1962), .d(n_1719), .o(n_2004) );
oa12s01 g779140 ( .a(n_1886), .b(n_1885), .c(n_1884), .o(n_2363) );
ao22s01 g779141 ( .a(n_1895), .b(n_1790), .c(n_1894), .d(n_1791), .o(n_2270) );
no02s02 g779142 ( .a(n_1993), .b(n_1992), .o(n_1994) );
in01s01 g779143 ( .a(n_1958), .o(n_1964) );
in01s01 g779145 ( .a(n_1956), .o(n_1957) );
na02s01 g779146 ( .a(n_1935), .b(n_1904), .o(n_1956) );
no02s01 g779147 ( .a(n_1928), .b(n_1927), .o(n_1929) );
no02m02 TIMEBOOST_cell_4955 ( .a(TIMEBOOST_net_1425), .b(n_33258), .o(n_33297) );
in01s01 g779149 ( .a(n_2025), .o(n_2003) );
no02s08 g779150 ( .a(n_1706), .b(n_1993), .o(n_2025) );
no02s01 g779152 ( .a(n_1915), .b(delay_add_ln22_unr2_stage2_stallmux_q_11_), .o(n_1936) );
in01s04 g779153 ( .a(n_1967), .o(n_1999) );
no02s06 g779154 ( .a(n_1962), .b(n_1685), .o(n_1967) );
na02s01 g779155 ( .a(n_1915), .b(delay_add_ln22_unr2_stage2_stallmux_q_11_), .o(n_1979) );
no02s01 g779156 ( .a(n_1921), .b(n_1919), .o(n_1920) );
na02s01 g779157 ( .a(n_2007), .b(n_2006), .o(n_2221) );
na02s01 g779158 ( .a(n_1885), .b(n_1884), .o(n_1886) );
na02s01 g779159 ( .a(n_2606), .b(n_1941), .o(n_1942) );
na02s02 g779160 ( .a(n_2487), .b(n_2405), .o(n_1933) );
in01s01 g779161 ( .a(n_1940), .o(n_2445) );
na02s01 g779162 ( .a(n_1908), .b(n_1941), .o(n_1940) );
na02s02 TIMEBOOST_cell_8676 ( .a(n_36613), .b(n_36750), .o(TIMEBOOST_net_2825) );
in01s01 g779165 ( .a(n_2218), .o(n_2622) );
ao12s01 g779166 ( .a(n_1875), .b(n_1874), .c(n_1873), .o(n_2218) );
oa12s01 g779167 ( .a(n_1910), .b(n_2494), .c(FE_OFN792_n_1909), .o(n_3944) );
oa22s01 g779168 ( .a(n_1864), .b(n_1689), .c(FE_OCP_RBN4011_n_1864), .d(n_1688), .o(n_1955) );
ao22s02 g779169 ( .a(n_1934), .b(n_1717), .c(n_1959), .d(n_1718), .o(n_2015) );
in01s01 g779170 ( .a(n_1901), .o(n_1902) );
na02s02 g779171 ( .a(n_1890), .b(n_1857), .o(n_1901) );
no02s01 g779172 ( .a(n_1874), .b(n_1873), .o(n_1875) );
na02s01 g779173 ( .a(n_1969), .b(n_1968), .o(n_2156) );
na02s10 g779174 ( .a(n_1959), .b(n_1665), .o(n_1993) );
in01s01 g779176 ( .a(n_1903), .o(n_1904) );
no02s02 g779177 ( .a(n_1898), .b(delay_add_ln22_unr2_stage2_stallmux_q_10_), .o(n_1903) );
na02s02 g779178 ( .a(n_1898), .b(delay_add_ln22_unr2_stage2_stallmux_q_10_), .o(n_1935) );
in01s06 g779179 ( .a(n_1916), .o(n_1962) );
no02s06 g779180 ( .a(n_1668), .b(FE_OCP_RBN4012_n_1864), .o(n_1916) );
na02s02 g779181 ( .a(n_1939), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_10_), .o(n_2006) );
na02s02 g779182 ( .a(n_1938), .b(n_1011), .o(n_2007) );
no02s04 TIMEBOOST_cell_1669 ( .a(n_31107), .b(TIMEBOOST_net_1793), .o(TIMEBOOST_net_449) );
in01s01 g779184 ( .a(n_2487), .o(n_1911) );
no02s01 g779185 ( .a(n_1880), .b(FE_OFN792_n_1909), .o(n_2487) );
na02s01 g779186 ( .a(n_2494), .b(FE_OFN792_n_1909), .o(n_1910) );
ao12s01 g779187 ( .a(n_1630), .b(n_44811), .c(n_1586), .o(n_1885) );
in01s01 g779189 ( .a(n_1894), .o(n_1895) );
oa12s01 g779190 ( .a(n_1792), .b(n_44812), .c(n_1569), .o(n_1894) );
na02m06 TIMEBOOST_cell_4017 ( .a(n_25412), .b(n_25511), .o(TIMEBOOST_net_1099) );
in01s01 g779192 ( .a(n_1908), .o(n_2606) );
oa12s01 g779193 ( .a(n_1848), .b(n_1847), .c(n_1846), .o(n_1908) );
in01s01 g779195 ( .a(n_1965), .o(n_2302) );
ao12s02 g779196 ( .a(n_1925), .b(n_1924), .c(n_1923), .o(n_1965) );
in01s01 g779197 ( .a(n_1887), .o(n_1888) );
ao22s01 g779198 ( .a(n_44811), .b(n_1809), .c(n_44812), .d(n_1810), .o(n_1887) );
oa12s01 g779199 ( .a(n_1860), .b(n_1859), .c(n_1858), .o(n_2292) );
no02s01 g779200 ( .a(n_1924), .b(n_1923), .o(n_1925) );
na02s01 g779201 ( .a(n_1862), .b(n_1850), .o(n_1851) );
na02s01 g779202 ( .a(n_1892), .b(n_1891), .o(n_2062) );
na02s01 g779203 ( .a(n_1847), .b(n_1846), .o(n_1848) );
na02s02 g779204 ( .a(n_1837), .b(delay_add_ln22_unr2_stage2_stallmux_q_9_), .o(n_1890) );
na02s01 g779205 ( .a(n_1953), .b(n_1952), .o(n_2095) );
na02m04 TIMEBOOST_cell_8833 ( .a(TIMEBOOST_net_2903), .b(n_5049), .o(TIMEBOOST_net_2155) );
na02s02 g779207 ( .a(n_1905), .b(n_944), .o(n_1969) );
in01s01 g779208 ( .a(n_1856), .o(n_1857) );
no02s02 g779209 ( .a(n_1837), .b(delay_add_ln22_unr2_stage2_stallmux_q_9_), .o(n_1856) );
in01s01 g779210 ( .a(n_1959), .o(n_1934) );
no02s10 g779211 ( .a(n_1924), .b(n_1695), .o(n_1959) );
no02s06 g779213 ( .a(n_1862), .b(n_1632), .o(n_1864) );
na02s02 g779214 ( .a(FE_OCP_RBN6551_n_1905), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_9_), .o(n_1968) );
na02s01 g779215 ( .a(n_1859), .b(n_1858), .o(n_1860) );
oa12f06 g779216 ( .a(n_1724), .b(n_1838), .c(n_1678), .o(n_1874) );
na02f06 g779217 ( .a(n_1863), .b(n_1624), .o(n_1869) );
in01s01 g779218 ( .a(n_2255), .o(n_1871) );
ao12s01 g779219 ( .a(n_1819), .b(n_1818), .c(n_1817), .o(n_2255) );
in01s02 g779220 ( .a(n_1880), .o(n_2494) );
ao22s01 g779221 ( .a(n_1761), .b(n_1838), .c(n_1760), .d(n_1811), .o(n_1880) );
oa22s01 g779222 ( .a(n_1820), .b(n_1483), .c(n_1821), .d(n_1482), .o(n_2364) );
oa22s02 g779223 ( .a(n_1812), .b(n_1610), .c(FE_OCP_RBN5553_n_1812), .d(n_1609), .o(n_1898) );
in01s01 g779224 ( .a(n_1938), .o(n_1939) );
oa22s02 g779225 ( .a(n_1889), .b(n_1650), .c(FE_OCP_RBN5560_n_1889), .d(n_1649), .o(n_1938) );
no02s01 g779226 ( .a(n_1818), .b(n_1817), .o(n_1819) );
na02s01 g779227 ( .a(n_1822), .b(n_1047), .o(n_1891) );
na02s02 g779228 ( .a(n_1845), .b(n_1844), .o(n_2008) );
na02s01 g779229 ( .a(FE_OCP_RBN5554_n_1822), .b(delay_add_ln22_unr2_stage2_stallmux_q_8_), .o(n_1892) );
na02s06 g779230 ( .a(n_1812), .b(n_1555), .o(n_1862) );
na02s02 g779231 ( .a(n_1900), .b(n_1899), .o(n_2040) );
na02s02 g779232 ( .a(n_1865), .b(n_946), .o(n_1953) );
na02s10 g779233 ( .a(n_1889), .b(n_1600), .o(n_1924) );
na02s02 g779234 ( .a(n_1866), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_8_), .o(n_1952) );
ao12f06 g779236 ( .a(n_1451), .b(n_1806), .c(n_1591), .o(n_1863) );
ao12s01 g779238 ( .a(n_1590), .b(n_1756), .c(n_1463), .o(n_1859) );
in01s01 g779241 ( .a(n_1835), .o(n_1836) );
oa12s01 g779242 ( .a(n_1769), .b(n_1795), .c(n_1768), .o(n_1835) );
oa22s01 g779243 ( .a(n_1725), .b(n_1564), .c(FE_OCP_RBN6548_n_1725), .d(n_1563), .o(n_1837) );
na02s01 g779244 ( .a(n_1853), .b(n_1842), .o(n_1843) );
na02s02 g779245 ( .a(n_1766), .b(n_1038), .o(n_1844) );
na02s03 g779246 ( .a(FE_OCP_RBN5555_n_1827), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_7_), .o(n_1899) );
na02s02 g779247 ( .a(n_1827), .b(n_1033), .o(n_1900) );
no02s10 g779249 ( .a(n_1595), .b(n_1853), .o(n_1889) );
na02s02 g779250 ( .a(n_1834), .b(n_1833), .o(n_1981) );
na02s01 g779251 ( .a(n_1795), .b(n_1768), .o(n_1769) );
no02s06 g779254 ( .a(FE_OCP_RBN6547_n_1725), .b(n_1544), .o(n_1812) );
na02s01 g779255 ( .a(n_1755), .b(n_1558), .o(n_1818) );
na02s04 g779256 ( .a(n_1767), .b(delay_add_ln22_unr2_stage2_stallmux_q_7_), .o(n_1845) );
na02s01 g779257 ( .a(n_1815), .b(n_1814), .o(n_1949) );
in01s01 g779258 ( .a(n_1838), .o(n_1811) );
ao12f06 g779259 ( .a(n_1653), .b(n_1789), .c(n_1694), .o(n_1838) );
in01s01 g779260 ( .a(n_1820), .o(n_1821) );
no02s04 TIMEBOOST_cell_1657 ( .a(FE_OCP_RBN4224_n_8799), .b(FE_OCP_RBN2782_n_8664), .o(TIMEBOOST_net_443) );
oa12s01 g779262 ( .a(n_1763), .b(n_1762), .c(n_1789), .o(n_2466) );
ao12s01 g779263 ( .a(n_1737), .b(n_1736), .c(n_1735), .o(n_2250) );
in01s01 g779264 ( .a(n_1865), .o(n_1866) );
na02s10 g779268 ( .a(n_1520), .b(n_1813), .o(n_1853) );
na02s01 g779269 ( .a(n_1745), .b(n_1744), .o(n_1873) );
in01s01 g779272 ( .a(n_1755), .o(n_1756) );
na02s01 g779273 ( .a(n_1736), .b(n_1559), .o(n_1755) );
na02s06 g779274 ( .a(n_1754), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_6_), .o(n_1833) );
na02s02 g779275 ( .a(n_1727), .b(n_912), .o(n_1814) );
na02s03 g779276 ( .a(n_1728), .b(delay_add_ln22_unr2_stage2_stallmux_q_6_), .o(n_1815) );
na02s02 g779277 ( .a(n_1753), .b(n_959), .o(n_1834) );
na02s01 g779278 ( .a(n_1785), .b(n_1784), .o(n_1919) );
no02s01 g779279 ( .a(n_1736), .b(n_1735), .o(n_1737) );
na02f08 g779280 ( .a(n_1736), .b(n_1557), .o(n_1806) );
na02s01 g779281 ( .a(n_1762), .b(n_1789), .o(n_1763) );
na02m04 TIMEBOOST_cell_8849 ( .a(TIMEBOOST_net_2911), .b(n_16513), .o(n_16601) );
oa22s02 g779284 ( .a(n_1776), .b(n_1534), .c(n_1732), .d(n_1535), .o(n_1827) );
in01s01 g779285 ( .a(n_2463), .o(n_2492) );
oa12s01 g779286 ( .a(n_1700), .b(n_1699), .c(n_1698), .o(n_2463) );
in01s01 g779288 ( .a(n_1766), .o(n_1767) );
na02s01 g779290 ( .a(n_1742), .b(n_1741), .o(n_1743) );
no02s01 g779291 ( .a(n_1712), .b(n_1711), .o(n_1713) );
na02s06 g779292 ( .a(n_1659), .b(delay_add_ln22_unr2_stage2_stallmux_q_5_), .o(n_1745) );
in01s01 g779293 ( .a(n_1760), .o(n_1761) );
na02s02 g779294 ( .a(n_1724), .b(n_1679), .o(n_1760) );
na02s02 g779295 ( .a(n_1658), .b(n_1039), .o(n_1744) );
na02s06 g779296 ( .a(n_1702), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_5_), .o(n_1784) );
in01s01 g779297 ( .a(n_1813), .o(n_1808) );
no02s10 g779298 ( .a(n_1503), .b(n_1776), .o(n_1813) );
na02s02 g779299 ( .a(n_1701), .b(n_1032), .o(n_1785) );
no02s06 g779301 ( .a(n_1712), .b(FE_OCPN3546_n_1705), .o(n_1733) );
na02s01 g779302 ( .a(n_1730), .b(n_1729), .o(n_1846) );
na02s01 g779303 ( .a(n_1699), .b(n_1698), .o(n_1700) );
na02s02 TIMEBOOST_cell_7098 ( .a(TIMEBOOST_net_2307), .b(n_22259), .o(n_22377) );
na02f08 g779305 ( .a(n_1636), .b(n_47027), .o(n_1736) );
na02s06 g779306 ( .a(n_1671), .b(n_1652), .o(n_1789) );
in01s01 g779307 ( .a(n_2442), .o(n_2461) );
ao12s01 g779308 ( .a(n_1709), .b(n_1708), .c(n_1707), .o(n_2442) );
in01s01 g779309 ( .a(n_2405), .o(n_1758) );
ao12s01 g779310 ( .a(n_1692), .b(n_1691), .c(n_1690), .o(n_2405) );
in01s01 g779311 ( .a(n_1727), .o(n_1728) );
in01s01 g779313 ( .a(n_1753), .o(n_1754) );
oa22s02 g779314 ( .a(FE_OCP_RBN6546_n_1672), .b(n_1476), .c(n_1672), .d(n_1477), .o(n_1753) );
in01s01 TIMEBOOST_cell_7384 ( .a(FE_OCPN1951_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(TIMEBOOST_net_2320) );
na02s01 g779316 ( .a(n_1667), .b(n_1666), .o(n_1768) );
no02s01 g779317 ( .a(n_1691), .b(n_1690), .o(n_1692) );
na02s06 g779318 ( .a(n_1675), .b(n_1402), .o(n_1712) );
na02s01 g779319 ( .a(n_1654), .b(n_1694), .o(n_1762) );
na02s02 g779320 ( .a(n_1639), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_4_), .o(n_1729) );
na02s02 g779321 ( .a(n_1660), .b(delay_add_ln22_unr2_stage2_stallmux_q_4_), .o(n_1724) );
na02s01 g779322 ( .a(n_1638), .b(n_892), .o(n_1730) );
in01m08 g779323 ( .a(n_1732), .o(n_1776) );
no02s10 g779324 ( .a(FE_OCP_RBN6545_n_1672), .b(n_1450), .o(n_1732) );
in01s01 g779325 ( .a(n_1678), .o(n_1679) );
no02s03 g779326 ( .a(n_1660), .b(delay_add_ln22_unr2_stage2_stallmux_q_4_), .o(n_1678) );
no02s01 g779327 ( .a(n_1708), .b(n_1707), .o(n_1709) );
oa12s04 g779328 ( .a(n_1616), .b(n_1644), .c(n_1690), .o(n_1699) );
no02s40 TIMEBOOST_cell_4862 ( .a(FE_OCP_RBN7113_n_44365), .b(delay_xor_ln22_unr12_stage5_stallmux_q_1_), .o(TIMEBOOST_net_1379) );
oa12f06 g779330 ( .a(n_1452), .b(n_1635), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_), .o(n_1636) );
no02m08 TIMEBOOST_cell_5056 ( .a(FE_OCP_RBN7036_n_18982), .b(n_18546), .o(TIMEBOOST_net_1476) );
in01s01 g779332 ( .a(n_1658), .o(n_1659) );
in01s01 g779334 ( .a(n_1701), .o(n_1702) );
oa12s01 g779336 ( .a(n_1627), .b(n_1635), .c(n_1626), .o(n_2276) );
na02s06 g779337 ( .a(n_1594), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_3_), .o(n_1666) );
no02s01 g779338 ( .a(n_1644), .b(n_1617), .o(n_1691) );
na02s04 g779339 ( .a(n_1623), .b(n_1622), .o(n_1694) );
na02s01 g779340 ( .a(n_1657), .b(n_1656), .o(n_1698) );
no02m10 g779342 ( .a(FE_OCP_RBN6535_n_1602), .b(n_1385), .o(n_1675) );
na02s40 TIMEBOOST_cell_7404 ( .a(FE_OCP_RBN7109_n_44365), .b(FE_OCP_RBN1120_delay_xor_ln22_unr12_stage5_stallmux_q_2_), .o(TIMEBOOST_net_2333) );
na02s06 g779344 ( .a(n_1625), .b(delay_add_ln22_unr2_stage2_stallmux_q_2_), .o(n_1652) );
na02s03 g779345 ( .a(n_1593), .b(n_1178), .o(n_1667) );
in01s01 g779346 ( .a(n_1653), .o(n_1654) );
no02s03 g779347 ( .a(n_1623), .b(n_1622), .o(n_1653) );
na02s01 g779350 ( .a(n_1635), .b(n_1626), .o(n_1627) );
in01s01 g779351 ( .a(n_2343), .o(n_1687) );
oa12s01 g779352 ( .a(n_1707), .b(n_1585), .c(delay_add_ln22_unr2_stage2_stallmux_q_1_), .o(n_2343) );
in01s02 g779353 ( .a(n_1787), .o(n_1648) );
ao12s04 g779354 ( .a(n_1629), .b(n_1628), .c(n_1613), .o(n_1787) );
ao22s01 g779355 ( .a(n_1604), .b(n_1633), .c(n_1662), .d(delay_add_ln22_unr2_stage2_stallmux_q_2_), .o(n_1708) );
in01s01 g779356 ( .a(n_1638), .o(n_1639) );
no02s06 TIMEBOOST_cell_4269 ( .a(n_33451), .b(n_33406), .o(TIMEBOOST_net_1225) );
no02s02 g779361 ( .a(n_1588), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_1_), .o(n_1644) );
in01s01 g779362 ( .a(n_1616), .o(n_1617) );
na02s02 g779363 ( .a(n_1588), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_1_), .o(n_1616) );
na02s02 g779364 ( .a(n_1541), .b(n_1447), .o(n_1560) );
no03m04 TIMEBOOST_cell_7325 ( .a(TIMEBOOST_net_1743), .b(n_26069), .c(n_26029), .o(n_26173) );
na02s02 g779367 ( .a(n_1571), .b(n_1107), .o(n_1656) );
na02s04 TIMEBOOST_cell_3887 ( .a(n_1785), .b(n_1784), .o(TIMEBOOST_net_1034) );
na02s02 g779370 ( .a(n_1572), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_2_), .o(n_1657) );
in01s01 g779371 ( .a(n_1625), .o(n_1707) );
in01s02 g779372 ( .a(n_1608), .o(n_1625) );
na02s06 g779373 ( .a(n_1585), .b(delay_add_ln22_unr2_stage2_stallmux_q_1_), .o(n_1608) );
in01s02 g779376 ( .a(n_1593), .o(n_1594) );
oa12m02 g779377 ( .a(n_1530), .b(n_1533), .c(n_1529), .o(n_1593) );
no02s04 g779378 ( .a(n_1548), .b(n_1524), .o(n_1623) );
ao12s01 g779379 ( .a(n_1546), .b(n_1551), .c(FE_OFN5064_n_1545), .o(n_2234) );
na02s02 g779380 ( .a(n_1533), .b(n_1529), .o(n_1530) );
no02s02 g779381 ( .a(n_1547), .b(n_1436), .o(n_1548) );
no02s02 g779382 ( .a(n_1513), .b(n_1437), .o(n_1524) );
no02s01 g779383 ( .a(n_1551), .b(FE_OFN5064_n_1545), .o(n_1546) );
no02m10 g779385 ( .a(n_1440), .b(n_1533), .o(n_1541) );
no02s06 g779387 ( .a(n_1547), .b(n_1542), .o(n_1577) );
na02s02 g779388 ( .a(n_1782), .b(n_1746), .o(n_1840) );
ao12s02 g779392 ( .a(FE_OCPN6911_n_1444), .b(n_1561), .c(n_1396), .o(n_1628) );
ao12s01 g779394 ( .a(n_1538), .b(n_1537), .c(delay_sub_ln21_0_unr2_stage2_stallmux_q_0_), .o(n_1909) );
in01s02 g779396 ( .a(n_1571), .o(n_1572) );
in01s01 g779398 ( .a(n_1662), .o(n_1604) );
na02s02 g779399 ( .a(n_1525), .b(n_1556), .o(n_1662) );
na02s01 g779401 ( .a(n_1590), .b(n_1549), .o(n_1550) );
no02s02 g779402 ( .a(n_1478), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_0_), .o(n_1690) );
na02s02 g779403 ( .a(n_1509), .b(n_1486), .o(n_1525) );
na02s02 g779404 ( .a(n_1485), .b(n_1510), .o(n_1556) );
in01s06 g779405 ( .a(n_1513), .o(n_1547) );
no02s01 g779407 ( .a(n_1537), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_0_), .o(n_1538) );
oa12s01 g779409 ( .a(n_1781), .b(n_1493), .c(n_1780), .o(n_1782) );
oa12m08 g779411 ( .a(n_1407), .b(n_1515), .c(n_1456), .o(n_1551) );
ao12s01 g779413 ( .a(n_1502), .b(n_1501), .c(n_1515), .o(n_1565) );
in01s01 g779414 ( .a(n_1509), .o(n_1510) );
no02m01 g779415 ( .a(n_1494), .b(n_1427), .o(n_1509) );
in01s01 g779416 ( .a(n_1495), .o(n_1496) );
na02s02 g779417 ( .a(n_1467), .b(n_1455), .o(n_1495) );
no02s02 g779418 ( .a(n_1587), .b(n_1603), .o(n_1624) );
no02s01 g779421 ( .a(n_1501), .b(n_1515), .o(n_1502) );
ao12s01 g779422 ( .a(n_2030), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_23_), .o(n_2353) );
ao12s02 g779423 ( .a(n_1508), .b(n_1507), .c(n_1506), .o(n_1561) );
ao12s01 g779424 ( .a(FE_OCPN3546_n_1705), .b(FE_OCP_RBN3976_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_7_), .o(n_1711) );
ao12s01 g779425 ( .a(n_2082), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_25_), .o(n_2439) );
in01s01 g779426 ( .a(n_1688), .o(n_1689) );
ao12s01 g779427 ( .a(n_1668), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_12_), .o(n_1688) );
in01s01 g779428 ( .a(n_1460), .o(n_1461) );
no02s02 g779429 ( .a(n_1397), .b(n_1399), .o(n_1460) );
ao12s02 g779430 ( .a(n_1595), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_9_), .o(n_1842) );
in01s01 g779431 ( .a(n_2116), .o(n_2117) );
ao12s01 g779432 ( .a(n_2108), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_26_), .o(n_2116) );
in01s01 g779433 ( .a(n_1534), .o(n_1535) );
ao12s02 g779434 ( .a(n_1503), .b(FE_OCP_RBN2378_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_7_), .o(n_1534) );
na02s01 TIMEBOOST_cell_8028 ( .a(FE_OCP_RBN6791_n_20242), .b(FE_OCPN1923_n_20430), .o(TIMEBOOST_net_2645) );
in01s01 g779436 ( .a(n_1829), .o(n_1830) );
ao12s01 g779437 ( .a(n_1764), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_16_), .o(n_1829) );
in01s01 g779438 ( .a(n_1563), .o(n_1564) );
ao12s01 g779439 ( .a(n_1544), .b(FE_OCP_RBN2377_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_9_), .o(n_1563) );
in01s01 g779440 ( .a(n_1960), .o(n_1961) );
ao12s01 g779441 ( .a(n_1947), .b(n_1852), .c(delay_xor_ln22_unr3_stage2_stallmux_q_20_), .o(n_1960) );
in01s01 g779442 ( .a(n_1917), .o(n_1918) );
ao12s01 g779443 ( .a(n_1878), .b(n_1852), .c(delay_xor_ln22_unr3_stage2_stallmux_q_18_), .o(n_1917) );
in01s01 g779444 ( .a(n_1474), .o(n_1475) );
no02s02 g779445 ( .a(n_1434), .b(n_1400), .o(n_1474) );
in01s01 g779446 ( .a(n_1649), .o(n_1650) );
ao12s01 g779447 ( .a(n_1599), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_10_), .o(n_1649) );
in01s01 g779448 ( .a(n_2070), .o(n_2071) );
ao12s01 g779449 ( .a(n_2026), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_24_), .o(n_2070) );
ao22s01 g779451 ( .a(n_1373), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(FE_OCP_RBN6517_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .d(delay_xor_ln21_unr3_stage2_stallmux_q_5_), .o(n_1438) );
in01s01 g779452 ( .a(n_2001), .o(n_2002) );
ao12s01 g779453 ( .a(n_1998), .b(n_1852), .c(delay_xor_ln22_unr3_stage2_stallmux_q_22_), .o(n_2001) );
ao12s01 g779454 ( .a(n_1797), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_15_), .o(n_2050) );
ao12s01 g779455 ( .a(n_1706), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_13_), .o(n_1992) );
in01s01 g779456 ( .a(n_2145), .o(n_2146) );
ao12s01 g779457 ( .a(n_2126), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_27_), .o(n_2145) );
in01s01 TIMEBOOST_cell_7385 ( .a(TIMEBOOST_net_2320), .o(TIMEBOOST_net_2321) );
oa12s01 g779460 ( .a(n_2113), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_28_), .o(n_2683) );
in01s01 g779461 ( .a(n_2019), .o(n_2020) );
ao12s01 g779462 ( .a(n_1972), .b(n_1852), .c(delay_xor_ln21_unr3_stage2_stallmux_q_22_), .o(n_2019) );
in01s01 g779463 ( .a(n_1773), .o(n_1774) );
ao12s01 g779464 ( .a(n_1759), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_14_), .o(n_1773) );
in01s01 g779465 ( .a(n_1854), .o(n_1855) );
ao12s01 g779466 ( .a(n_1832), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_16_), .o(n_1854) );
in01s01 g779467 ( .a(n_1476), .o(n_1477) );
ao12s02 g779468 ( .a(n_1450), .b(FE_OCP_RBN6517_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_6_), .o(n_1476) );
in01s01 g779469 ( .a(n_1804), .o(n_1805) );
ao12s01 g779470 ( .a(n_1770), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_15_), .o(n_1804) );
in01s01 g779471 ( .a(n_1931), .o(n_1932) );
ao12s01 g779472 ( .a(n_1882), .b(n_1852), .c(delay_xor_ln21_unr3_stage2_stallmux_q_18_), .o(n_1931) );
ao12s01 g779473 ( .a(n_1881), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_17_), .o(n_2088) );
ao12s01 g779474 ( .a(n_2073), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_25_), .o(n_2496) );
in01s01 g779475 ( .a(n_1824), .o(n_1825) );
ao12s01 g779476 ( .a(n_1703), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_14_), .o(n_1824) );
in01s01 g779478 ( .a(n_2028), .o(n_2029) );
ao12s01 g779479 ( .a(n_2021), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_23_), .o(n_2028) );
in01s01 g779480 ( .a(n_1996), .o(n_1997) );
ao12s01 g779481 ( .a(n_1945), .b(n_1852), .c(delay_xor_ln21_unr3_stage2_stallmux_q_20_), .o(n_1996) );
in01s01 g779482 ( .a(n_1717), .o(n_1718) );
ao12s01 g779483 ( .a(n_1664), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_12_), .o(n_1717) );
ao12s01 g779484 ( .a(n_1695), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_11_), .o(n_1923) );
ao12s01 g779485 ( .a(n_1990), .b(n_1852), .c(delay_xor_ln21_unr3_stage2_stallmux_q_21_), .o(n_2253) );
in01s01 g779487 ( .a(n_2090), .o(n_2091) );
ao12s01 g779488 ( .a(n_2083), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_26_), .o(n_2090) );
na02s04 g779490 ( .a(n_1376), .b(n_1455), .o(n_1472) );
in01s01 g779491 ( .a(n_1876), .o(n_1877) );
ao12s01 g779492 ( .a(n_1861), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_17_), .o(n_1876) );
in01s02 g779494 ( .a(n_1436), .o(n_1437) );
in01s01 g779496 ( .a(n_2046), .o(n_2047) );
ao12s01 g779497 ( .a(n_2011), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_24_), .o(n_2046) );
ao22s01 g779499 ( .a(n_1370), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(FE_OCP_RBN6410_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .d(delay_xor_ln22_unr3_stage2_stallmux_q_4_), .o(n_1448) );
ao12s01 g779500 ( .a(n_1930), .b(n_1852), .c(delay_xor_ln22_unr3_stage2_stallmux_q_19_), .o(n_2164) );
no02m02 g779501 ( .a(n_1440), .b(n_1406), .o(n_1529) );
in01s01 g779502 ( .a(n_1485), .o(n_1486) );
no02s01 TIMEBOOST_cell_1551 ( .a(n_30001), .b(n_29877), .o(TIMEBOOST_net_390) );
ao12s01 g779504 ( .a(n_1913), .b(n_1852), .c(delay_xor_ln21_unr3_stage2_stallmux_q_19_), .o(n_2194) );
in01s01 g779506 ( .a(n_1609), .o(n_1610) );
ao12s01 g779507 ( .a(n_1554), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_10_), .o(n_1609) );
in01s01 g779508 ( .a(n_1446), .o(n_1447) );
ao22s01 g779509 ( .a(n_1368), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(FE_OCP_RBN6410_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .d(delay_xor_ln21_unr3_stage2_stallmux_q_4_), .o(n_1446) );
in01s01 g779510 ( .a(n_1983), .o(n_1984) );
ao12s01 g779511 ( .a(n_1971), .b(n_1852), .c(delay_xor_ln22_unr3_stage2_stallmux_q_21_), .o(n_1983) );
in01s01 g779512 ( .a(n_1453), .o(n_1454) );
ao22m01 g779513 ( .a(n_1372), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(FE_OCP_RBN6516_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .d(delay_xor_ln22_unr3_stage2_stallmux_q_5_), .o(n_1453) );
in01s01 g779514 ( .a(n_1719), .o(n_1720) );
ao12s01 g779515 ( .a(n_1685), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_13_), .o(n_1719) );
in01s01 g779516 ( .a(n_1567), .o(n_1568) );
ao12s01 g779517 ( .a(n_1519), .b(FE_OCP_RBN2378_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_8_), .o(n_1567) );
oa12s02 g779519 ( .a(n_1686), .b(n_1739), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_), .o(n_1781) );
ao22s01 g779520 ( .a(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(n_1371), .c(FE_OCP_RBN3762_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .d(delay_xor_ln22_unr3_stage2_stallmux_q_0_), .o(n_1941) );
in01s01 g779521 ( .a(n_1478), .o(n_1537) );
na02m06 TIMEBOOST_cell_5026 ( .a(FE_OCP_RBN1827_n_19538), .b(FE_OCPN4528_n_18117), .o(TIMEBOOST_net_1461) );
in01s01 g779523 ( .a(n_2359), .o(n_2360) );
oa22s01 g779524 ( .a(n_1433), .b(n_607), .c(n_1403), .d(delay_sub_ln23_0_unr1_stage2_stallmux_q_1_), .o(n_2359) );
in01s01 g779525 ( .a(n_1586), .o(n_1587) );
no02s02 g779526 ( .a(n_1569), .b(n_1570), .o(n_1586) );
no02s08 g779527 ( .a(n_1433), .b(delay_sub_ln23_0_unr1_stage2_stallmux_q_1_), .o(n_1515) );
na02s04 TIMEBOOST_cell_5025 ( .a(TIMEBOOST_net_1460), .b(n_41608), .o(n_41740) );
no02s01 g779530 ( .a(n_1619), .b(n_1620), .o(n_1646) );
no02s01 g779531 ( .a(n_1470), .b(n_1445), .o(n_1746) );
no02s02 g779533 ( .a(n_1643), .b(n_1801), .o(n_1741) );
na02s02 g779535 ( .a(n_1527), .b(n_1780), .o(n_1528) );
na02m08 TIMEBOOST_cell_6671 ( .a(n_24488), .b(n_24457), .o(TIMEBOOST_net_2093) );
no02s01 g779538 ( .a(n_1553), .b(n_1603), .o(n_1884) );
in01s02 g779539 ( .a(n_1397), .o(n_1398) );
no02s06 g779540 ( .a(FE_OCP_RBN6408_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_2_), .o(n_1397) );
in01s02 g779541 ( .a(n_1519), .o(n_1520) );
no02s02 g779542 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_8_), .b(FE_OCP_RBN2378_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1519) );
no02s02 g779543 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_13_), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1706) );
in01s01 g779544 ( .a(n_1878), .o(n_1879) );
no02s01 g779545 ( .a(n_1852), .b(delay_xor_ln22_unr3_stage2_stallmux_q_18_), .o(n_1878) );
no02s01 g779546 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_26_), .o(n_2108) );
no02s01 g779547 ( .a(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_15_), .o(n_1770) );
in01s06 g779548 ( .a(n_1426), .o(n_1427) );
na02m03 g779550 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(n_1365), .o(n_1426) );
no02s03 g779551 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_7_), .b(FE_OCP_RBN6517_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1503) );
no02s02 g779552 ( .a(FE_OCP_RBN3976_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_9_), .o(n_1544) );
no02s03 g779553 ( .a(FE_OCP_RBN6408_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_2_), .o(n_1435) );
na02s10 g779554 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(n_1366), .o(n_1455) );
in01s01 g779555 ( .a(n_1664), .o(n_1665) );
no02s01 g779556 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_12_), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1664) );
in01s01 g779557 ( .a(n_2113), .o(n_2114) );
na02s01 g779558 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_28_), .o(n_2113) );
no02s01 g779559 ( .a(n_1456), .b(n_1408), .o(n_1501) );
na02s06 g779560 ( .a(FE_OCP_RBN6407_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_1_), .o(n_1376) );
no02s01 g779561 ( .a(n_1800), .b(delay_xor_ln22_unr3_stage2_stallmux_q_17_), .o(n_1881) );
no02s01 g779562 ( .a(n_1852), .b(delay_xor_ln22_unr3_stage2_stallmux_q_20_), .o(n_1947) );
in01s01 g779563 ( .a(n_1554), .o(n_1555) );
no02s01 g779564 ( .a(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_10_), .o(n_1554) );
no02s01 g779565 ( .a(n_1471), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_26_), .o(n_1493) );
in01s01 g779566 ( .a(n_1599), .o(n_1600) );
no02s01 g779567 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_10_), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1599) );
no02s06 g779568 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_5_), .b(FE_OCP_RBN6516_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1385) );
no02s20 g779569 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_3_), .b(FE_OCP_RBN6407_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1440) );
in01s01 g779570 ( .a(n_1809), .o(n_1810) );
na02s01 g779571 ( .a(n_1792), .b(n_1514), .o(n_1809) );
no02s03 g779573 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_11_), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1695) );
no02s01 g779574 ( .a(n_1852), .b(delay_xor_ln22_unr3_stage2_stallmux_q_21_), .o(n_1971) );
in01s01 g779575 ( .a(n_1467), .o(n_1421) );
na02s10 g779576 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(n_1362), .o(n_1467) );
no02s01 g779577 ( .a(n_1783), .b(n_1739), .o(n_2120) );
no02s02 g779578 ( .a(n_1374), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1399) );
in01s06 g779579 ( .a(n_1434), .o(n_1402) );
no02s06 g779580 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_6_), .b(FE_OCP_RBN6516_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1434) );
no02s01 g779581 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_12_), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1668) );
no02s06 g779582 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_9_), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1595) );
no02s01 g779583 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_27_), .o(n_2126) );
in01s01 g779584 ( .a(n_2026), .o(n_2027) );
no02s01 g779585 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_24_), .o(n_2026) );
no02s20 g779586 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_3_), .b(FE_OCP_RBN6407_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1542) );
no02s01 g779587 ( .a(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_14_), .o(n_1759) );
no02s01 g779588 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_17_), .b(n_1800), .o(n_1861) );
in01s01 g779589 ( .a(n_1972), .o(n_1973) );
no02s01 g779590 ( .a(n_1852), .b(delay_xor_ln21_unr3_stage2_stallmux_q_22_), .o(n_1972) );
no02s02 g779592 ( .a(n_1364), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1406) );
no02s02 g779593 ( .a(n_1363), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1400) );
no02s06 g779595 ( .a(FE_OCP_RBN6408_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_0_), .o(n_1494) );
in01s01 g779596 ( .a(n_2011), .o(n_2012) );
no02s01 g779597 ( .a(n_1800), .b(delay_xor_ln22_unr3_stage2_stallmux_q_24_), .o(n_2011) );
in01s01 g779598 ( .a(n_1882), .o(n_1883) );
no02s01 g779599 ( .a(n_1852), .b(delay_xor_ln21_unr3_stage2_stallmux_q_18_), .o(n_1882) );
na02s01 g779600 ( .a(n_1721), .b(n_1715), .o(n_2176) );
no02s08 g779601 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_6_), .b(FE_OCP_RBN6517_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1450) );
in01s01 g779602 ( .a(n_1703), .o(n_1704) );
no02s01 g779603 ( .a(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_14_), .o(n_1703) );
no02s04 TIMEBOOST_cell_2932 ( .a(n_19255), .b(n_18507), .o(TIMEBOOST_net_757) );
no02s02 g779605 ( .a(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_13_), .o(n_1685) );
no02s01 g779606 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_16_), .o(n_1832) );
no02s01 g779607 ( .a(n_1800), .b(delay_xor_ln22_unr3_stage2_stallmux_q_25_), .o(n_2073) );
no02s01 g779608 ( .a(n_1518), .b(n_1543), .o(n_1858) );
in01s01 g779609 ( .a(n_1802), .o(n_1803) );
na02s01 g779610 ( .a(n_1794), .b(n_1584), .o(n_1802) );
na02m08 TIMEBOOST_cell_5027 ( .a(TIMEBOOST_net_1461), .b(n_19568), .o(n_19730) );
na02s01 g779612 ( .a(n_1559), .b(n_1558), .o(n_1735) );
na02s01 g779613 ( .a(n_1516), .b(n_1507), .o(n_2131) );
no02s02 g779614 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_15_), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1797) );
na02s01 g779615 ( .a(n_1596), .b(n_1613), .o(n_2092) );
no02s01 g779616 ( .a(n_1800), .b(delay_xor_ln22_unr3_stage2_stallmux_q_26_), .o(n_2083) );
in01s01 g779617 ( .a(n_1945), .o(n_1946) );
no02s01 g779618 ( .a(n_1852), .b(delay_xor_ln21_unr3_stage2_stallmux_q_20_), .o(n_1945) );
na03m10 TIMEBOOST_cell_8284 ( .a(n_18119), .b(n_19454), .c(n_19427), .o(n_19585) );
no02s01 g779620 ( .a(n_1852), .b(delay_xor_ln21_unr3_stage2_stallmux_q_21_), .o(n_1990) );
no02s01 g779621 ( .a(n_1852), .b(delay_xor_ln22_unr3_stage2_stallmux_q_19_), .o(n_1930) );
no02s01 g779622 ( .a(n_1852), .b(delay_xor_ln22_unr3_stage2_stallmux_q_23_), .o(n_2021) );
no02s06 g779623 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_7_), .b(FE_OCP_RBN6516_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1705) );
no02s01 g779624 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_25_), .o(n_2082) );
na02s01 g779625 ( .a(n_1674), .b(n_1681), .o(n_2053) );
no02s01 g779626 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_22_), .b(n_1852), .o(n_1998) );
no02s01 g779627 ( .a(n_1852), .b(delay_xor_ln21_unr3_stage2_stallmux_q_19_), .o(n_1913) );
na02f02 TIMEBOOST_cell_6827 ( .a(n_16661), .b(n_16662), .o(TIMEBOOST_net_2171) );
no02s01 g779629 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_23_), .o(n_2030) );
in01s01 g779630 ( .a(n_1764), .o(n_1765) );
no02s01 g779631 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_16_), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1764) );
no02s01 g779632 ( .a(n_1752), .b(n_1801), .o(n_2134) );
in01s01 g779633 ( .a(n_1504), .o(n_1505) );
no02s01 g779634 ( .a(n_1471), .b(n_1470), .o(n_1504) );
na02s01 g779635 ( .a(n_1463), .b(n_1462), .o(n_1817) );
no02s01 g779636 ( .a(n_1444), .b(n_1443), .o(n_2128) );
no02s01 g779637 ( .a(n_1409), .b(n_1484), .o(n_2013) );
in01s01 g779638 ( .a(n_1497), .o(n_1498) );
no02s01 g779639 ( .a(n_1512), .b(n_1420), .o(n_1497) );
na02s01 g779640 ( .a(n_1442), .b(n_1441), .o(n_1927) );
in01s01 g779641 ( .a(n_1499), .o(n_1500) );
na02s01 g779642 ( .a(n_1480), .b(n_1479), .o(n_1499) );
in01s01 g779643 ( .a(n_1487), .o(n_1488) );
ao12s01 g779644 ( .a(n_1431), .b(FE_OCPN4927_n_1452), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_28_), .o(n_1487) );
in01s01 g779645 ( .a(n_1790), .o(n_1791) );
ao12s01 g779646 ( .a(n_1570), .b(n_1686), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_8_), .o(n_1790) );
in01s01 g779647 ( .a(n_1482), .o(n_1483) );
ao12s01 g779648 ( .a(n_1451), .b(n_1452), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_6_), .o(n_1482) );
in01s01 g779649 ( .a(n_1489), .o(n_1490) );
ao12s01 g779650 ( .a(n_1445), .b(FE_OCPN4927_n_1452), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_26_), .o(n_1489) );
in01s01 g779651 ( .a(n_1771), .o(n_1772) );
ao12s01 g779652 ( .a(n_1643), .b(n_1686), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_20_), .o(n_1771) );
in01s01 g779653 ( .a(n_1798), .o(n_1799) );
ao12s01 g779654 ( .a(n_1748), .b(n_1686), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_22_), .o(n_1798) );
in01s01 g779655 ( .a(n_1778), .o(n_1779) );
ao12s01 g779656 ( .a(n_1620), .b(n_1686), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_12_), .o(n_1778) );
oa12s01 g779657 ( .a(n_1731), .b(n_1686), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_), .o(n_2183) );
oa22s01 g779658 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_1_), .c(n_1780), .d(n_1392), .o(n_1545) );
oa22s01 g779659 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_), .c(n_1780), .d(n_756), .o(n_1626) );
in01s01 g779663 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_0_), .o(n_1369) );
in01s10 g779664 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_0_), .o(n_1362) );
in01s01 g779675 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_0_), .o(n_1371) );
in01s01 g779678 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_2_), .o(n_1374) );
in01s10 g779681 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_1_), .o(n_1366) );
in01m03 g779684 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_1_), .o(n_1365) );
in01s01 g779690 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_4_), .o(n_1370) );
in01s02 g779693 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_3_), .o(n_1364) );
in01s01 g779696 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_2_), .o(n_1367) );
in01s01 g779699 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_5_), .o(n_1373) );
in01s01 g779701 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_6_), .o(n_1363) );
in01s01 g779712 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_4_), .o(n_1368) );
in01s06 g779714 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_5_), .o(n_1372) );
na02s01 g779727 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_11_), .o(n_1794) );
no02s01 g779728 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_12_), .o(n_1620) );
no02s01 g779729 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_19_), .o(n_1801) );
no02s01 g779730 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_8_), .o(n_1570) );
no02s02 g779731 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_22_), .o(n_1748) );
in01s01 g779732 ( .a(n_1521), .o(n_1559) );
no02s01 g779733 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_3_), .o(n_1521) );
in01s01 g779734 ( .a(n_1407), .o(n_1408) );
na02s10 g779735 ( .a(n_1379), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_0_), .o(n_1407) );
na02s01 g779736 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_7_), .o(n_1792) );
na02s01 g779737 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_18_), .o(n_1613) );
no02s08 g779738 ( .a(n_1379), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_0_), .o(n_1456) );
no02s01 g779739 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_20_), .o(n_1643) );
no02s01 g779740 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_23_), .o(n_1783) );
in01s01 g779741 ( .a(n_1629), .o(n_1596) );
no02s01 g779742 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_18_), .o(n_1629) );
in01s01 g779743 ( .a(n_1751), .o(n_1752) );
na02s01 g779744 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_19_), .o(n_1751) );
in01s01 g779745 ( .a(n_1580), .o(n_1553) );
na02s01 g779746 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_9_), .o(n_1580) );
in01s01 g779747 ( .a(n_1527), .o(n_1518) );
na02s02 g779748 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_5_), .o(n_1527) );
in01s01 g779749 ( .a(n_1673), .o(n_1674) );
no02s01 g779750 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_14_), .b(n_1575), .o(n_1673) );
in01s01 g779751 ( .a(n_1508), .o(n_1516) );
no02s01 g779752 ( .a(n_1379), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_16_), .o(n_1508) );
na02s06 g779753 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_3_), .o(n_1558) );
na02s01 g779754 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_), .o(n_1731) );
na02s01 g779755 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_21_), .o(n_1715) );
na02s01 g779756 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_14_), .b(n_1575), .o(n_1681) );
in01s01 g779757 ( .a(n_1663), .o(n_1739) );
na02s02 g779758 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_23_), .o(n_1663) );
in01s01 g779759 ( .a(n_1569), .o(n_1514) );
no02s01 g779760 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_7_), .o(n_1569) );
in01s01 g779761 ( .a(n_1749), .o(n_1721) );
no02s01 g779762 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_21_), .o(n_1749) );
in01s01 g779763 ( .a(n_1619), .o(n_1584) );
no02s01 g779764 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_11_), .o(n_1619) );
in01s01 g779765 ( .a(n_1543), .o(n_1549) );
no02s06 g779766 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_5_), .o(n_1543) );
no02s01 g779767 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_9_), .o(n_1603) );
na02s02 g779768 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_16_), .o(n_1507) );
na02s01 g779770 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_27_), .b(n_1452), .o(n_1479) );
no02s01 g779771 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_25_), .o(n_1470) );
na02s01 g779773 ( .a(n_1780), .b(n_1392), .o(n_1393) );
no02s01 g779774 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_15_), .o(n_1512) );
no02s01 g779775 ( .a(n_1780), .b(n_1381), .o(n_1444) );
in01s01 g779776 ( .a(n_1396), .o(n_1443) );
na02s01 g779777 ( .a(n_1780), .b(n_1381), .o(n_1396) );
in01s01 g779778 ( .a(n_1423), .o(n_1471) );
na02s01 g779779 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_25_), .o(n_1423) );
in01s01 g779780 ( .a(n_1415), .o(n_1480) );
no02s01 g779781 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_27_), .b(n_1452), .o(n_1415) );
na02s01 g779782 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_10_), .o(n_1441) );
in01s01 g779783 ( .a(n_1422), .o(n_1463) );
no02s01 g779784 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_4_), .o(n_1422) );
na02s01 g779786 ( .a(n_1780), .b(n_1131), .o(n_1442) );
no02s01 g779787 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_26_), .o(n_1445) );
na02s02 g779788 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_4_), .o(n_1462) );
no02s02 g779789 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_6_), .o(n_1451) );
no02s01 g779791 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_28_), .b(n_1452), .o(n_1431) );
in01s01 g779792 ( .a(n_1506), .o(n_1420) );
na02s01 g779793 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_15_), .o(n_1506) );
in01s01 g779794 ( .a(n_1484), .o(n_1645) );
no02s01 g779795 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_13_), .b(n_1452), .o(n_1484) );
in01s01 g779796 ( .a(n_1682), .o(n_1409) );
na02s01 g779797 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_13_), .o(n_1682) );
oa12s01 g779799 ( .a(n_2115), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_28_), .o(n_2137) );
ao12s01 g779801 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_23_), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_), .o(n_1722) );
in01s01 g779802 ( .a(n_1433), .o(n_1403) );
na02m02 TIMEBOOST_cell_1544 ( .a(TIMEBOOST_net_386), .b(n_14478), .o(FE_RN_1466_0) );
in01s01 g779805 ( .a(n_1601), .o(n_1630) );
in01s01 g779807 ( .a(n_1539), .o(n_1540) );
ao12s01 g779808 ( .a(n_1517), .b(FE_OCP_RBN2377_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_8_), .o(n_1539) );
in01s01 g779809 ( .a(n_2124), .o(n_2125) );
ao12s01 g779810 ( .a(n_2109), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_27_), .o(n_2124) );
ao12s01 g779811 ( .a(n_1632), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_11_), .o(n_1850) );
oa12s01 g779812 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_20_), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_19_), .o(n_1714) );
na02m03 g779815 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln23_unr3_stage2_stallmux_q), .o(n_1387) );
no02s02 g779816 ( .a(FE_OCP_RBN3976_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_8_), .o(n_1517) );
in01s06 g779817 ( .a(n_1780), .o(n_1452) );
no02s40 g779818 ( .a(delay_xor_ln23_unr3_stage2_stallmux_q), .b(FE_OCP_RBN6408_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1780) );
na02s01 g779819 ( .a(n_1800), .b(delay_xor_ln22_unr3_stage2_stallmux_q_28_), .o(n_2115) );
no02s01 g779820 ( .a(n_1800), .b(delay_xor_ln22_unr3_stage2_stallmux_q_27_), .o(n_2109) );
in01s02 g779825 ( .a(n_1377), .o(n_1686) );
in01s02 g779835 ( .a(n_1377), .o(n_1575) );
in01s10 g779842 ( .a(n_1377), .o(n_1416) );
in01s10 g779844 ( .a(n_1379), .o(n_1377) );
na02s40 g779845 ( .a(FE_OCP_RBN6409_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln23_unr3_stage2_stallmux_q), .o(n_1379) );
no02s01 g779846 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_11_), .b(FE_OCP_RBN3763_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1632) );
oa22s01 g779847 ( .a(n_44652), .b(n_1190), .c(n_44623), .d(n_1183), .o(n_1302) );
oa22s01 g779849 ( .a(n_44652), .b(n_1022), .c(n_44623), .d(n_957), .o(n_1355) );
oa22s01 g779852 ( .a(n_44652), .b(n_1025), .c(n_44623), .d(n_989), .o(n_1300) );
oa22s01 g779856 ( .a(n_44659), .b(n_973), .c(n_44623), .d(n_899), .o(n_1288) );
oa22s01 g779859 ( .a(n_44652), .b(n_1163), .c(n_44623), .d(n_1151), .o(n_1315) );
oa22s02 g779861 ( .a(n_44652), .b(n_1018), .c(n_44637), .d(n_975), .o(n_1345) );
oa22s01 g779862 ( .a(FE_OCPN838_n_44672), .b(n_1001), .c(n_44637), .d(n_954), .o(n_1332) );
oa22s01 g779865 ( .a(n_44659), .b(n_1169), .c(n_44623), .d(n_1158), .o(n_1322) );
oa22s01 g779871 ( .a(n_44659), .b(n_981), .c(n_44623), .d(n_924), .o(n_1357) );
in01s01 g779872 ( .a(n_1285), .o(n_1286) );
oa22s01 g779873 ( .a(n_44636), .b(n_990), .c(FE_OCPN5099_n_1282), .d(n_1014), .o(n_1285) );
oa22s01 g779874 ( .a(n_44659), .b(n_886), .c(n_44661), .d(n_822), .o(n_1291) );
oa22s01 g779876 ( .a(FE_OCPN838_n_44672), .b(n_1118), .c(n_44637), .d(n_1068), .o(n_1289) );
in01s01 g779877 ( .a(n_1356), .o(n_1360) );
ao22s01 g779878 ( .a(FE_OCPN5099_n_1282), .b(n_902), .c(n_44650), .d(n_934), .o(n_1356) );
oa22s01 g779880 ( .a(n_44652), .b(n_1129), .c(n_44637), .d(n_1087), .o(n_1287) );
oa22s01 g779881 ( .a(FE_OCPN838_n_44672), .b(n_1040), .c(n_44637), .d(n_984), .o(n_1348) );
oa22s01 g779883 ( .a(n_44659), .b(n_1066), .c(n_44623), .d(n_1028), .o(n_1346) );
oa22s01 g779884 ( .a(n_44652), .b(n_1144), .c(n_44623), .d(n_1125), .o(n_1351) );
oa22s01 g779886 ( .a(FE_OCPN839_n_44672), .b(n_1137), .c(n_44623), .d(n_1121), .o(n_1306) );
oa22s01 g779888 ( .a(n_44652), .b(n_1009), .c(n_44623), .d(n_962), .o(n_1308) );
oa22s01 g779890 ( .a(n_44652), .b(n_1134), .c(n_44623), .d(n_1120), .o(n_1324) );
oa22s01 g779891 ( .a(FE_OCPN838_n_44672), .b(n_1005), .c(n_44623), .d(n_949), .o(n_1297) );
oa22s01 g779892 ( .a(n_44659), .b(FE_OFN4817_n_920), .c(n_44623), .d(n_920), .o(n_1340) );
oa22s01 g779894 ( .a(n_44659), .b(n_1092), .c(n_44623), .d(n_1050), .o(n_1292) );
oa22s01 g779895 ( .a(n_44652), .b(n_1019), .c(n_44623), .d(n_947), .o(n_1320) );
oa22s02 g779896 ( .a(n_44652), .b(n_1017), .c(n_44661), .d(n_972), .o(n_1335) );
oa22s01 g779899 ( .a(n_44652), .b(FE_OFN4785_n_45813), .c(n_44623), .d(n_1203), .o(n_1325) );
in01s02 g779929 ( .a(FE_OCP_RBN3762_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1852) );
in01s03 g779940 ( .a(FE_OCP_RBN3762_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1800) );
oa22s01 g779978 ( .a(n_1268), .b(n_999), .c(n_1267), .d(n_1000), .o(n_1274) );
no02f10 g780009 ( .a(n_1026), .b(n_1269), .o(n_1282) );
oa22s01 g780010 ( .a(n_1270), .b(n_1044), .c(n_1271), .d(n_1043), .o(n_1275) );
no02f08 g780012 ( .a(n_1266), .b(n_1027), .o(n_1269) );
in01s01 g780013 ( .a(n_1267), .o(n_1268) );
oa12s01 g780014 ( .a(n_977), .b(n_1259), .c(n_925), .o(n_1267) );
oa22s01 g780015 ( .a(n_1259), .b(n_982), .c(n_1264), .d(n_983), .o(n_1272) );
oa22s01 g780016 ( .a(n_1263), .b(n_1072), .c(n_1262), .d(n_1073), .o(n_1273) );
in01s01 g780018 ( .a(n_1270), .o(n_1271) );
in01s01 g780019 ( .a(n_1266), .o(n_1270) );
no02s01 TIMEBOOST_cell_1032 ( .a(n_33005), .b(TIMEBOOST_net_130), .o(n_33122) );
oa22s01 g780021 ( .a(n_1253), .b(n_988), .c(n_1254), .d(n_987), .o(n_1261) );
in01s01 g780024 ( .a(n_1262), .o(n_1263) );
no02s01 g780025 ( .a(n_1256), .b(n_985), .o(n_1262) );
no02s01 TIMEBOOST_cell_1031 ( .a(n_33028), .b(n_32488), .o(TIMEBOOST_net_130) );
in01s01 g780028 ( .a(n_1259), .o(n_1264) );
oa12s01 g780029 ( .a(n_866), .b(n_1250), .c(n_929), .o(n_1259) );
oa22s01 g780030 ( .a(n_1251), .b(n_1070), .c(n_1250), .d(n_1071), .o(n_1260) );
in01s01 g780032 ( .a(n_1255), .o(n_1256) );
na02f06 g780033 ( .a(n_1248), .b(n_1053), .o(n_1255) );
in01s01 g780034 ( .a(n_1253), .o(n_1254) );
oa12s01 g780035 ( .a(n_891), .b(n_1245), .c(n_844), .o(n_1253) );
oa22s01 g780036 ( .a(n_1245), .b(n_930), .c(n_1246), .d(n_931), .o(n_1257) );
oa22s01 g780037 ( .a(n_1243), .b(n_1059), .c(n_1242), .d(n_1060), .o(n_1249) );
in01s01 g780040 ( .a(n_1250), .o(n_1251) );
in01s01 g780041 ( .a(n_1248), .o(n_1250) );
no02s02 TIMEBOOST_cell_996 ( .a(TIMEBOOST_net_112), .b(n_23195), .o(n_23312) );
oa22s01 g780043 ( .a(n_1233), .b(n_896), .c(n_1232), .d(n_895), .o(n_1241) );
in01s01 g780044 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_17_), .o(n_1381) );
in01s01 g780048 ( .a(n_1245), .o(n_1246) );
na02s01 g780049 ( .a(n_1239), .b(n_888), .o(n_1245) );
in01s01 g780050 ( .a(n_1242), .o(n_1243) );
ao12s01 g780051 ( .a(n_816), .b(n_1231), .c(n_1052), .o(n_1242) );
no02s04 TIMEBOOST_cell_8737 ( .a(TIMEBOOST_net_2855), .b(n_13807), .o(TIMEBOOST_net_2703) );
oa22s01 g780053 ( .a(n_1231), .b(n_1054), .c(n_1235), .d(n_1055), .o(n_1244) );
in01s01 g780054 ( .a(n_1238), .o(n_1239) );
no02f06 g780055 ( .a(n_1230), .b(n_894), .o(n_1238) );
in01s01 g780056 ( .a(n_1232), .o(n_1233) );
ao12s01 g780057 ( .a(n_818), .b(n_1225), .c(n_842), .o(n_1232) );
oa22s01 g780058 ( .a(n_1229), .b(n_1062), .c(n_1228), .d(n_1063), .o(n_1237) );
oa22s01 g780059 ( .a(n_1225), .b(n_825), .c(n_1226), .d(n_826), .o(n_1234) );
in01s01 g780062 ( .a(n_1231), .o(n_1235) );
in01s01 g780063 ( .a(n_1230), .o(n_1231) );
na02s04 TIMEBOOST_cell_8804 ( .a(n_14524), .b(n_15598), .o(TIMEBOOST_net_2889) );
in01s01 g780066 ( .a(n_1225), .o(n_1226) );
na02s01 g780067 ( .a(n_1222), .b(n_769), .o(n_1225) );
no02s01 TIMEBOOST_cell_957 ( .a(n_18052), .b(n_18051), .o(TIMEBOOST_net_93) );
in01s01 g780069 ( .a(n_1228), .o(n_1229) );
ao12s01 g780070 ( .a(n_1016), .b(n_1215), .c(n_1051), .o(n_1228) );
oa22s01 g780071 ( .a(n_1218), .b(n_1057), .c(n_1220), .d(n_1058), .o(n_1224) );
na02f06 g780073 ( .a(n_1215), .b(n_811), .o(n_1222) );
in01s01 g780074 ( .a(n_1220), .o(n_1218) );
in01s01 g780076 ( .a(n_1215), .o(n_1220) );
oa12m06 g780077 ( .a(n_841), .b(n_1199), .c(n_793), .o(n_1215) );
oa12s01 g780078 ( .a(n_1214), .b(n_1213), .c(n_1212), .o(n_1219) );
na02s01 g780080 ( .a(n_1213), .b(n_1212), .o(n_1214) );
ao12m06 g780081 ( .a(n_1191), .b(n_1198), .c(n_814), .o(n_1199) );
no02s01 g780082 ( .a(n_1192), .b(n_790), .o(n_1213) );
oa12s01 g780083 ( .a(n_1196), .b(n_1198), .c(n_1195), .o(n_1207) );
na02s01 g780085 ( .a(n_1198), .b(n_1195), .o(n_1196) );
no02s01 g780086 ( .a(n_1198), .b(n_1191), .o(n_1192) );
no02s01 TIMEBOOST_cell_1552 ( .a(TIMEBOOST_net_390), .b(n_30442), .o(n_30549) );
oa12m08 g780088 ( .a(n_742), .b(n_1184), .c(n_781), .o(n_1198) );
oa12s01 g780089 ( .a(n_1172), .b(n_1184), .c(n_1171), .o(n_1187) );
na02s01 g780091 ( .a(n_1184), .b(n_1171), .o(n_1172) );
ao12m08 g780092 ( .a(n_746), .b(n_1153), .c(n_771), .o(n_1184) );
oa12s01 g780093 ( .a(n_1146), .b(n_1153), .c(n_1145), .o(n_1166) );
na02s01 g780095 ( .a(n_1153), .b(n_1145), .o(n_1146) );
oa12m08 g780097 ( .a(n_725), .b(n_1119), .c(n_751), .o(n_1153) );
oa12s01 g780098 ( .a(n_1097), .b(n_1119), .c(n_1096), .o(n_1136) );
in01s01 g780099 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_10_), .o(n_1131) );
na02s01 g780101 ( .a(n_1119), .b(n_1096), .o(n_1097) );
in01s01 g780102 ( .a(n_1217), .o(n_1216) );
oa12s01 g780103 ( .a(n_1210), .b(n_45818), .c(n_1208), .o(n_1217) );
na02s01 g780109 ( .a(n_45818), .b(n_1208), .o(n_1210) );
ao12m08 g780110 ( .a(n_732), .b(n_1029), .c(n_753), .o(n_1119) );
oa12s01 g780111 ( .a(n_1013), .b(n_1029), .c(n_1012), .o(n_1082) );
na02s01 g780112 ( .a(n_1029), .b(n_1012), .o(n_1013) );
in01s01 g780114 ( .a(n_1206), .o(n_1201) );
oa12s01 g780115 ( .a(n_1182), .b(n_1181), .c(n_1180), .o(n_1206) );
oa12s01 g780116 ( .a(n_1086), .b(n_1085), .c(n_1084), .o(n_1135) );
in01s01 g780117 ( .a(n_1205), .o(n_1200) );
oa22s01 g780118 ( .a(n_1175), .b(FE_OFN759_n_45813), .c(n_1176), .d(n_1203), .o(n_1205) );
in01s01 g780119 ( .a(n_1211), .o(n_1204) );
oa22s01 g780120 ( .a(n_1194), .b(n_1203), .c(n_1185), .d(FE_OFN759_n_45813), .o(n_1211) );
in01s01 g780121 ( .a(n_1188), .o(n_1186) );
oa12s01 g780122 ( .a(n_1161), .b(n_1160), .c(n_1159), .o(n_1188) );
in01s01 g780123 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_24_), .o(n_1197) );
in01s01 g780126 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_22_), .o(n_2379) );
in01s01 g780128 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_14_), .o(n_1173) );
na02s01 g780131 ( .a(n_1160), .b(n_1159), .o(n_1161) );
na02s01 g780132 ( .a(n_1181), .b(n_1180), .o(n_1182) );
na02s01 g780133 ( .a(n_1085), .b(n_1084), .o(n_1086) );
ao12m08 g780134 ( .a(n_711), .b(n_948), .c(n_727), .o(n_1029) );
in01s01 g780138 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_21_), .o(n_1177) );
in01s01 g780140 ( .a(n_1194), .o(n_1185) );
na02s01 g780141 ( .a(n_1147), .b(n_832), .o(n_1194) );
na02s01 g780142 ( .a(n_948), .b(n_1006), .o(n_1085) );
oa12s01 g780143 ( .a(n_881), .b(n_1139), .c(n_802), .o(n_1160) );
oa12s01 g780144 ( .a(n_1111), .b(n_1170), .c(n_936), .o(n_1181) );
in01s01 g780145 ( .a(n_1175), .o(n_1176) );
oa12s01 g780146 ( .a(n_935), .b(n_1162), .c(n_1061), .o(n_1175) );
in01s01 g780147 ( .a(n_1189), .o(n_1179) );
oa12s01 g780148 ( .a(n_1156), .b(n_1162), .c(n_1155), .o(n_1189) );
in01s01 g780149 ( .a(n_1169), .o(n_1158) );
oa22s01 g780150 ( .a(n_1091), .b(FE_OFN4781_n_45813), .c(n_1090), .d(n_1203), .o(n_1169) );
oa12s01 g780151 ( .a(n_1076), .b(n_1075), .c(n_1074), .o(n_1112) );
in01s01 g780152 ( .a(n_1190), .o(n_1183) );
oa12s01 g780153 ( .a(n_1149), .b(n_1170), .c(n_1148), .o(n_1190) );
in01s01 g780154 ( .a(n_1164), .o(n_1157) );
oa12s01 g780155 ( .a(n_1123), .b(n_1139), .c(n_1122), .o(n_1164) );
in01s01 g780156 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_3_), .o(n_1178) );
in01s01 g780159 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_23_), .o(n_1174) );
na02s01 g780162 ( .a(n_1170), .b(n_1148), .o(n_1149) );
na02s01 g780163 ( .a(n_1139), .b(n_1122), .o(n_1123) );
na02s01 g780164 ( .a(n_1162), .b(n_1155), .o(n_1156) );
na02m08 g780165 ( .a(n_1075), .b(n_882), .o(n_948) );
na02s01 g780166 ( .a(n_1075), .b(n_1074), .o(n_1076) );
na02s02 g780167 ( .a(n_1170), .b(n_797), .o(n_1147) );
in01s01 g780168 ( .a(n_1124), .o(n_1100) );
oa22s01 g780169 ( .a(n_997), .b(n_1098), .c(n_45819), .d(n_1099), .o(n_1124) );
in01s01 g780170 ( .a(n_1142), .o(n_1130) );
oa12s01 g780171 ( .a(n_1078), .b(n_1077), .c(n_1159), .o(n_1142) );
in01s01 g780172 ( .a(n_1163), .o(n_1151) );
oa22s01 g780173 ( .a(n_1093), .b(n_1203), .c(n_1094), .d(FE_OFN4786_n_45813), .o(n_1163) );
in01s01 g780174 ( .a(n_1168), .o(n_1150) );
oa12s01 g780175 ( .a(n_1117), .b(n_1116), .c(n_1148), .o(n_1168) );
in01s01 g780180 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_19_), .o(n_1101) );
in01s01 g780182 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_28_), .o(n_1095) );
na02s01 g780184 ( .a(n_848), .b(n_1128), .o(n_1170) );
na02s01 g780185 ( .a(n_1116), .b(n_1148), .o(n_1117) );
na02s01 g780186 ( .a(n_1128), .b(n_45814), .o(n_1162) );
na02s01 g780187 ( .a(n_1077), .b(n_1159), .o(n_1078) );
in01s01 g780188 ( .a(n_1090), .o(n_1091) );
ao12s01 g780189 ( .a(n_796), .b(n_1069), .c(n_762), .o(n_1090) );
oa22s01 g780190 ( .a(n_1069), .b(n_817), .c(n_1061), .d(n_779), .o(n_1139) );
oa12m08 g780191 ( .a(n_703), .b(n_837), .c(n_730), .o(n_1075) );
in01s01 g780192 ( .a(n_1143), .o(n_1165) );
ao22s01 g780193 ( .a(n_1067), .b(FE_OFN759_n_45813), .c(n_1089), .d(n_1203), .o(n_1143) );
oa12s01 g780194 ( .a(n_813), .b(n_837), .c(n_812), .o(n_854) );
in01s01 g780195 ( .a(n_1137), .o(n_1121) );
oa12s01 g780196 ( .a(n_1030), .b(n_1069), .c(n_1180), .o(n_1137) );
in01s01 g780197 ( .a(n_1167), .o(n_1154) );
oa12s02 g780198 ( .a(n_1115), .b(n_1114), .c(n_1113), .o(n_1167) );
in01s01 g780201 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_19_), .o(n_1141) );
in01s01 g780204 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_5_), .o(n_1039) );
in01s01 g780208 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_7_), .o(n_1038) );
na02s01 g780210 ( .a(n_1069), .b(n_1180), .o(n_1030) );
na02s01 g780211 ( .a(n_45809), .b(n_1041), .o(n_1116) );
na02s02 g780212 ( .a(n_1111), .b(n_1042), .o(n_1128) );
in01s01 g780213 ( .a(n_1125), .o(n_1144) );
no02s01 g780214 ( .a(n_1089), .b(n_883), .o(n_1125) );
na02s01 g780215 ( .a(n_837), .b(n_812), .o(n_813) );
na02s01 g780216 ( .a(n_1114), .b(n_1113), .o(n_1115) );
in01s01 g780217 ( .a(n_1093), .o(n_1094) );
oa12s01 g780218 ( .a(n_749), .b(n_1056), .c(n_845), .o(n_1093) );
no02s01 g780219 ( .a(n_45817), .b(n_763), .o(n_1077) );
in01s01 g780220 ( .a(n_45819), .o(n_997) );
in01s01 g780222 ( .a(n_1134), .o(n_1120) );
oa22s01 g780223 ( .a(n_1008), .b(n_1099), .c(n_1056), .d(n_1098), .o(n_1134) );
in01s01 g780224 ( .a(n_1102), .o(n_1064) );
oa22s01 g780225 ( .a(n_1003), .b(n_1203), .c(n_969), .d(FE_OFN4780_n_45813), .o(n_1102) );
in01s01 g780226 ( .a(n_1065), .o(n_1049) );
oa12s01 g780227 ( .a(n_961), .b(n_960), .c(n_1155), .o(n_1065) );
in01s01 g780228 ( .a(n_1028), .o(n_1066) );
ao22s01 g780229 ( .a(n_970), .b(FE_OFN759_n_45813), .c(n_904), .d(n_1203), .o(n_1028) );
in01s01 g780230 ( .a(n_1138), .o(n_1152) );
ao12s01 g780231 ( .a(n_1081), .b(n_1080), .c(n_1079), .o(n_1138) );
in01s01 g780232 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_2_), .o(n_1107) );
in01s01 g780234 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_18_), .o(n_1126) );
in01s01 g780236 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_18_), .o(n_1037) );
in01s01 g780240 ( .a(n_1041), .o(n_1042) );
na02s01 g780241 ( .a(n_1002), .b(n_1003), .o(n_1041) );
no02s01 g780242 ( .a(n_1080), .b(n_1079), .o(n_1081) );
na02s01 g780243 ( .a(n_960), .b(n_1155), .o(n_961) );
ao22s01 g780244 ( .a(n_995), .b(n_798), .c(n_849), .d(n_45809), .o(n_1069) );
in01s01 g780246 ( .a(n_1089), .o(n_1067) );
ao12s01 g780247 ( .a(n_1098), .b(n_1046), .c(FE_OFN824_n_1045), .o(n_1089) );
ao12m08 g780248 ( .a(n_684), .b(n_786), .c(n_698), .o(n_837) );
in01s01 g780249 ( .a(n_1106), .o(n_1132) );
ao22s01 g780250 ( .a(n_980), .b(n_1099), .c(n_979), .d(n_1098), .o(n_1106) );
in01s01 g780251 ( .a(n_1088), .o(n_1127) );
ao22s01 g780252 ( .a(n_974), .b(n_1203), .c(n_1046), .d(FE_OFN759_n_45813), .o(n_1088) );
oa12s01 g780253 ( .a(n_1105), .b(n_1104), .c(n_1103), .o(n_1133) );
in01s01 g780254 ( .a(n_1025), .o(n_989) );
oa12s01 g780255 ( .a(n_911), .b(n_910), .c(n_1159), .o(n_1025) );
oa12s01 g780256 ( .a(n_1024), .b(n_1023), .c(FE_OFN824_n_1045), .o(n_1114) );
in01s01 g780257 ( .a(n_1087), .o(n_1129) );
ao22s01 g780258 ( .a(n_991), .b(FE_OFN4784_n_45813), .c(n_992), .d(n_1203), .o(n_1087) );
in01s01 g780259 ( .a(n_1010), .o(n_993) );
oa22s01 g780260 ( .a(n_45816), .b(n_1122), .c(n_863), .d(n_1208), .o(n_1010) );
in01s01 g780261 ( .a(n_1018), .o(n_975) );
oa12s01 g780262 ( .a(n_909), .b(n_908), .c(n_1148), .o(n_1018) );
oa12s01 g780263 ( .a(n_766), .b(n_786), .c(n_765), .o(n_791) );
in01s01 g780264 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_17_), .o(n_1083) );
in01s01 g780267 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_5_), .o(n_1032) );
in01s01 g780270 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_8_), .o(n_1047) );
in01s01 g780276 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_10_), .o(n_1011) );
in01s01 g780278 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_27_), .o(n_1031) );
in01s01 g780280 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_7_), .o(n_1033) );
in01s01 g780282 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_4_), .o(n_792) );
in01s01 g780284 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_3_), .o(n_1622) );
in01s01 g780286 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_24_), .o(n_2483) );
na02s01 g780288 ( .a(n_910), .b(n_1159), .o(n_911) );
na02s01 g780289 ( .a(n_908), .b(n_1148), .o(n_909) );
in01s01 g780290 ( .a(n_970), .o(n_904) );
na02s01 g780291 ( .a(n_833), .b(n_881), .o(n_970) );
na02s01 g780292 ( .a(n_1046), .b(n_1203), .o(n_1080) );
na02s01 g780293 ( .a(n_1104), .b(n_1103), .o(n_1105) );
na02s01 g780294 ( .a(n_1023), .b(FE_OFN824_n_1045), .o(n_1024) );
na02s01 g780295 ( .a(n_1113), .b(n_956), .o(n_1021) );
na02s01 g780296 ( .a(n_786), .b(n_765), .o(n_766) );
in01s01 g780297 ( .a(n_1056), .o(n_1008) );
ao12s01 g780298 ( .a(n_827), .b(n_995), .c(n_1002), .o(n_1056) );
oa12s01 g780299 ( .a(n_750), .b(n_903), .c(n_795), .o(n_960) );
in01s01 g780300 ( .a(n_998), .o(n_1048) );
ao22s01 g780301 ( .a(n_950), .b(n_1098), .c(n_864), .d(n_1099), .o(n_998) );
oa12s01 g780302 ( .a(n_1113), .b(n_941), .c(FE_OFN824_n_1045), .o(n_1007) );
in01s01 g780303 ( .a(n_1050), .o(n_1092) );
ao12s01 g780304 ( .a(n_965), .b(n_964), .c(n_1079), .o(n_1050) );
in01s01 g780305 ( .a(n_954), .o(n_1001) );
ao22s01 g780306 ( .a(n_922), .b(n_1148), .c(n_903), .d(n_770), .o(n_954) );
in01s01 g780307 ( .a(n_969), .o(n_1003) );
ao22s01 g780308 ( .a(n_855), .b(n_936), .c(n_922), .d(n_935), .o(n_969) );
in01s01 g780309 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_2_), .o(n_1633) );
in01s01 g780311 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_8_), .o(n_946) );
in01s01 g780314 ( .a(n_991), .o(n_992) );
no02s01 g780315 ( .a(n_995), .b(n_1061), .o(n_991) );
no02s01 g780316 ( .a(n_964), .b(n_1079), .o(n_965) );
in01s01 g780317 ( .a(n_979), .o(n_980) );
na02s01 g780318 ( .a(n_950), .b(n_942), .o(n_979) );
oa12s01 g780319 ( .a(n_945), .b(n_889), .c(n_870), .o(n_963) );
na02s01 g780320 ( .a(n_941), .b(FE_OFN824_n_1045), .o(n_1113) );
na02s01 g780321 ( .a(n_848), .b(n_755), .o(n_849) );
ao12s01 g780322 ( .a(n_831), .b(n_851), .c(n_45809), .o(n_908) );
in01s01 g780323 ( .a(n_45816), .o(n_863) );
in01s01 g780325 ( .a(n_984), .o(n_1040) );
ao12s01 g780326 ( .a(n_964), .b(n_907), .c(n_1203), .o(n_984) );
in01s01 g780327 ( .a(n_1046), .o(n_974) );
na02s01 g780328 ( .a(n_850), .b(n_942), .o(n_1046) );
oa12s01 g780329 ( .a(n_690), .b(n_739), .c(n_706), .o(n_1104) );
oa12m08 g780330 ( .a(n_686), .b(n_739), .c(n_689), .o(n_786) );
in01s01 g780331 ( .a(n_957), .o(n_1022) );
ao12s01 g780332 ( .a(n_879), .b(n_937), .c(n_878), .o(n_957) );
in01s01 g780333 ( .a(n_962), .o(n_1009) );
ao12s01 g780334 ( .a(n_861), .b(n_937), .c(n_860), .o(n_962) );
oa12s01 g780335 ( .a(n_716), .b(n_715), .c(n_714), .o(n_738) );
in01s01 g780336 ( .a(n_897), .o(n_966) );
ao22s01 g780337 ( .a(n_1208), .b(n_801), .c(n_1122), .d(n_800), .o(n_897) );
in01s01 g780338 ( .a(n_967), .o(n_1004) );
ao12s01 g780339 ( .a(n_874), .b(n_1079), .c(n_919), .o(n_967) );
oa12s01 g780340 ( .a(n_915), .b(n_955), .c(n_580), .o(n_1023) );
oa12s01 g780341 ( .a(n_718), .b(n_739), .c(n_717), .o(n_740) );
in01s01 g780342 ( .a(n_924), .o(n_981) );
ao22s01 g780343 ( .a(n_824), .b(n_1203), .c(n_823), .d(FE_OFN759_n_45813), .o(n_924) );
in01s01 g780344 ( .a(n_918), .o(n_958) );
ao22s01 g780345 ( .a(n_807), .b(n_1203), .c(n_851), .d(FE_OFN4782_n_45813), .o(n_918) );
oa12s01 g780346 ( .a(n_45815), .b(n_832), .c(n_831), .o(n_833) );
in01s01 g780347 ( .a(n_990), .o(n_1014) );
oa22s01 g780348 ( .a(n_921), .b(n_840), .c(n_920), .d(n_919), .o(n_990) );
in01s01 g780349 ( .a(n_899), .o(n_973) );
ao22s01 g780350 ( .a(n_1122), .b(n_789), .c(n_1208), .d(n_856), .o(n_899) );
in01s01 g780351 ( .a(n_972), .o(n_1017) );
ao12s01 g780352 ( .a(n_873), .b(n_937), .c(n_872), .o(n_972) );
ao12s01 g780353 ( .a(n_901), .b(n_955), .c(n_46055), .o(n_956) );
in01s01 g780354 ( .a(n_947), .o(n_1019) );
ao12s01 g780355 ( .a(n_877), .b(n_1155), .c(n_876), .o(n_947) );
in01s01 g780356 ( .a(n_949), .o(n_1005) );
ao22s01 g780357 ( .a(n_1079), .b(FE_OFN759_n_45813), .c(n_853), .d(n_1203), .o(n_949) );
ao22s01 g780358 ( .a(n_806), .b(n_856), .c(n_855), .d(n_420), .o(n_910) );
in01s01 g780360 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_9_), .o(n_944) );
in01s01 g780362 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_6_), .o(n_959) );
in01s01 g780364 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_1_), .o(n_1392) );
in01s01 g780368 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_), .o(n_756) );
in01s01 g780370 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_4_), .o(n_892) );
in01s01 g780372 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_6_), .o(n_912) );
in01s01 g780374 ( .a(n_903), .o(n_922) );
na02s01 g780375 ( .a(n_856), .b(n_778), .o(n_903) );
no02s01 g780376 ( .a(n_858), .b(n_782), .o(n_995) );
no02s01 g780377 ( .a(n_1155), .b(n_876), .o(n_877) );
no02s01 g780378 ( .a(n_955), .b(n_46055), .o(n_901) );
na02s01 g780379 ( .a(n_955), .b(n_580), .o(n_915) );
no02s01 g780380 ( .a(n_907), .b(n_1203), .o(n_964) );
na02s01 g780381 ( .a(n_907), .b(n_805), .o(n_942) );
na02s01 g780382 ( .a(n_715), .b(n_714), .o(n_716) );
no02s01 g780383 ( .a(n_860), .b(n_1098), .o(n_850) );
no02s01 g780384 ( .a(n_937), .b(n_878), .o(n_879) );
no02s01 g780385 ( .a(n_937), .b(n_860), .o(n_861) );
no02s01 g780386 ( .a(n_1079), .b(n_919), .o(n_874) );
no02s01 g780387 ( .a(n_937), .b(n_872), .o(n_873) );
in01s01 g780388 ( .a(n_950), .o(n_864) );
no02s01 g780389 ( .a(n_860), .b(n_847), .o(n_950) );
na02s01 g780390 ( .a(n_739), .b(n_717), .o(n_718) );
in01s01 g780391 ( .a(n_848), .o(n_827) );
no02f08 TIMEBOOST_cell_6836 ( .a(n_35923), .b(TIMEBOOST_net_2175), .o(n_36015) );
in01s01 g780393 ( .a(n_875), .o(n_928) );
ao22s01 g780394 ( .a(n_847), .b(n_1098), .c(n_815), .d(n_1099), .o(n_875) );
oa22s01 g780395 ( .a(n_836), .b(n_420), .c(n_846), .d(n_580), .o(n_941) );
in01s01 g780396 ( .a(FE_OFN1178_n_916), .o(n_938) );
ao22s01 g780397 ( .a(n_883), .b(FE_OFN759_n_45813), .c(n_834), .d(n_1203), .o(n_916) );
oa22s01 g780398 ( .a(n_881), .b(n_780), .c(n_803), .d(n_1159), .o(n_835) );
in01s01 g780399 ( .a(n_789), .o(n_856) );
no02s01 g780400 ( .a(n_802), .b(n_767), .o(n_789) );
in01s01 g780401 ( .a(n_876), .o(n_858) );
na02s01 g780402 ( .a(n_804), .b(n_45814), .o(n_876) );
no02s06 TIMEBOOST_cell_6835 ( .a(n_35878), .b(n_34918), .o(TIMEBOOST_net_2175) );
in01s01 g780404 ( .a(n_800), .o(n_801) );
na02s01 g780405 ( .a(n_881), .b(n_778), .o(n_800) );
in01s01 g780406 ( .a(n_851), .o(n_807) );
na02s01 g780407 ( .a(n_806), .b(n_881), .o(n_851) );
na02s01 g780408 ( .a(n_787), .b(n_1002), .o(n_817) );
na02s01 g780409 ( .a(n_935), .b(n_784), .o(n_1155) );
no02s01 g780410 ( .a(n_796), .b(n_795), .o(n_797) );
no02s01 g780411 ( .a(n_796), .b(n_788), .o(n_1180) );
no02s01 g780412 ( .a(n_788), .b(n_936), .o(n_832) );
in01s01 g780414 ( .a(n_1208), .o(n_1122) );
no02s01 g780415 ( .a(n_802), .b(n_803), .o(n_1208) );
no02s02 g780416 ( .a(n_846), .b(n_845), .o(n_955) );
no02s01 g780417 ( .a(n_888), .b(n_887), .o(n_889) );
in01s01 g780418 ( .a(n_823), .o(n_824) );
na02s01 g780419 ( .a(n_815), .b(n_1098), .o(n_823) );
ao12s01 g780420 ( .a(n_884), .b(n_820), .c(n_799), .o(n_885) );
no02s01 g780421 ( .a(n_821), .b(FE_OFN759_n_45813), .o(n_860) );
in01s01 g780422 ( .a(n_1079), .o(n_853) );
no02s02 g780423 ( .a(n_847), .b(n_821), .o(n_1079) );
in01s01 g780424 ( .a(n_902), .o(n_934) );
ao12s01 g780425 ( .a(n_878), .b(n_1203), .c(n_1099), .o(n_902) );
ao12s01 g780426 ( .a(n_878), .b(n_1099), .c(FE_OFN824_n_1045), .o(n_907) );
oa12s01 g780427 ( .a(n_834), .b(n_1098), .c(FE_OFN824_n_1045), .o(n_937) );
oa12s01 g780428 ( .a(n_675), .b(n_707), .c(n_687), .o(n_715) );
na02s01 g780429 ( .a(n_943), .b(n_926), .o(n_1020) );
no02m08 g780430 ( .a(n_688), .b(n_676), .o(n_739) );
in01s01 g780431 ( .a(n_921), .o(n_920) );
oa12s01 g780432 ( .a(n_872), .b(n_1203), .c(FE_OFN824_n_1045), .o(n_921) );
oa12s01 g780433 ( .a(n_1110), .b(n_1109), .c(n_1108), .o(n_1140) );
oa12s01 g780434 ( .a(n_709), .b(n_708), .c(n_707), .o(n_729) );
in01s01 g780435 ( .a(n_822), .o(n_886) );
ao22s01 g780436 ( .a(n_1203), .b(n_855), .c(FE_OFN4782_n_45813), .d(n_764), .o(n_822) );
in01s01 g780437 ( .a(n_1068), .o(n_1118) );
ao22s01 g780438 ( .a(FE_OFN4782_n_45813), .b(n_923), .c(n_1203), .d(n_890), .o(n_1068) );
in01s01 g780441 ( .a(n_788), .o(n_762) );
no02s01 g780442 ( .a(n_46055), .b(n_855), .o(n_788) );
in01s01 g780443 ( .a(n_796), .o(n_787) );
no02s01 g780444 ( .a(n_764), .b(n_7), .o(n_796) );
in01s01 g780445 ( .a(n_784), .o(n_1061) );
na02s01 g780446 ( .a(n_7), .b(n_855), .o(n_784) );
in01s01 g780447 ( .a(n_935), .o(n_782) );
na02s01 g780448 ( .a(n_46055), .b(n_764), .o(n_935) );
no02s01 g780449 ( .a(n_855), .b(n_521), .o(n_802) );
na02s01 g780450 ( .a(n_764), .b(n_580), .o(n_806) );
in01s01 g780451 ( .a(n_881), .o(n_803) );
na02s01 g780452 ( .a(n_855), .b(n_580), .o(n_881) );
no02s01 g780453 ( .a(n_1203), .b(n_845), .o(n_798) );
no02s01 g780454 ( .a(n_1203), .b(n_1099), .o(n_878) );
in01s01 g780455 ( .a(n_840), .o(n_919) );
no02s01 g780456 ( .a(FE_OFN4783_n_45813), .b(n_1099), .o(n_840) );
in01s01 g780457 ( .a(n_834), .o(n_883) );
na02s01 g780458 ( .a(n_1098), .b(FE_OFN824_n_1045), .o(n_834) );
in01s01 g780459 ( .a(n_846), .o(n_836) );
no02s02 g780460 ( .a(FE_OFN4782_n_45813), .b(n_745), .o(n_846) );
in01s01 g780461 ( .a(n_815), .o(n_847) );
na02s01 g780462 ( .a(FE_OFN759_n_45813), .b(FE_OFN824_n_1045), .o(n_815) );
na02s01 g780463 ( .a(n_1203), .b(FE_OFN824_n_1045), .o(n_872) );
in01s01 g780464 ( .a(n_821), .o(n_805) );
no02s01 g780465 ( .a(FE_OFN759_n_45813), .b(FE_OFN824_n_1045), .o(n_821) );
na02s01 g780466 ( .a(n_1109), .b(n_1108), .o(n_1110) );
na02s01 g780467 ( .a(n_708), .b(n_707), .o(n_709) );
na02s01 g780469 ( .a(n_855), .b(n_759), .o(n_804) );
no02m04 g780470 ( .a(n_671), .b(n_707), .o(n_688) );
oa12s01 g780471 ( .a(n_893), .b(n_816), .c(n_779), .o(n_888) );
na03s01 g780472 ( .a(n_976), .b(n_951), .c(n_977), .o(n_978) );
no02s06 TIMEBOOST_cell_8687 ( .a(TIMEBOOST_net_2830), .b(TIMEBOOST_net_916), .o(n_21571) );
in01s01 g780474 ( .a(n_1159), .o(n_780) );
no02s02 g780475 ( .a(n_767), .b(n_724), .o(n_1159) );
in01s01 g780476 ( .a(n_1098), .o(n_1099) );
no02s02 g780477 ( .a(n_754), .b(n_845), .o(n_1098) );
no02s01 g780478 ( .a(n_831), .b(n_754), .o(n_755) );
na02s01 g780479 ( .a(n_1002), .b(n_736), .o(n_763) );
no02s01 g780480 ( .a(n_831), .b(n_795), .o(n_759) );
in01s01 g780481 ( .a(n_1148), .o(n_770) );
na02s02 g780482 ( .a(n_1111), .b(n_750), .o(n_1148) );
in01s02 g780483 ( .a(FE_OFN759_n_45813), .o(n_1203) );
no02s01 g780485 ( .a(n_887), .b(n_900), .o(n_927) );
na02m02 g780486 ( .a(n_664), .b(n_670), .o(n_671) );
na02m04 g780487 ( .a(n_675), .b(n_674), .o(n_676) );
na02s01 g780488 ( .a(n_869), .b(n_868), .o(n_870) );
no02s01 g780489 ( .a(n_925), .b(n_913), .o(n_926) );
no02s01 g780490 ( .a(n_743), .b(n_781), .o(n_1171) );
in01s01 g780491 ( .a(n_895), .o(n_896) );
no02s01 g780492 ( .a(n_819), .b(n_884), .o(n_895) );
in01s01 g780493 ( .a(n_1057), .o(n_1058) );
na02s01 g780494 ( .a(n_1015), .b(n_1051), .o(n_1057) );
in01s01 g780495 ( .a(n_982), .o(n_983) );
na02s01 g780496 ( .a(n_977), .b(n_898), .o(n_982) );
in01s01 g780497 ( .a(n_1043), .o(n_1044) );
no02s01 g780498 ( .a(n_1027), .b(n_1026), .o(n_1043) );
in01s01 g780499 ( .a(n_930), .o(n_931) );
na02s01 g780500 ( .a(n_869), .b(n_891), .o(n_930) );
no02s01 g780501 ( .a(n_691), .b(n_706), .o(n_717) );
na02s01 g780502 ( .a(n_733), .b(n_753), .o(n_1012) );
na02s01 g780503 ( .a(n_768), .b(n_842), .o(n_799) );
na02s01 g780504 ( .a(n_752), .b(n_814), .o(n_1195) );
no02s01 g780505 ( .a(n_704), .b(n_730), .o(n_812) );
in01s01 g780506 ( .a(n_987), .o(n_988) );
na02s01 g780507 ( .a(n_868), .b(n_945), .o(n_987) );
no02s01 g780508 ( .a(n_667), .b(n_687), .o(n_708) );
na02s01 g780509 ( .a(n_674), .b(n_670), .o(n_714) );
in01s01 g780510 ( .a(n_999), .o(n_1000) );
na02s01 g780511 ( .a(n_951), .b(n_914), .o(n_999) );
na02s01 g780512 ( .a(n_1006), .b(n_882), .o(n_1074) );
no02s01 g780513 ( .a(n_819), .b(n_818), .o(n_820) );
no02s01 g780514 ( .a(n_726), .b(n_751), .o(n_1096) );
in01s01 g780515 ( .a(n_1054), .o(n_1055) );
na02s01 g780516 ( .a(n_1052), .b(n_761), .o(n_1054) );
in01s01 g780517 ( .a(n_1070), .o(n_1071) );
na02s01 g780518 ( .a(n_986), .b(n_1053), .o(n_1070) );
na02s01 g780519 ( .a(n_829), .b(n_842), .o(n_843) );
na02s01 g780520 ( .a(n_794), .b(n_841), .o(n_1212) );
na02s01 g780521 ( .a(n_698), .b(n_685), .o(n_765) );
na02s01 g780522 ( .a(n_771), .b(n_747), .o(n_1145) );
in01s01 g780523 ( .a(n_825), .o(n_826) );
na02s01 g780524 ( .a(n_842), .b(n_776), .o(n_825) );
in01s01 g780525 ( .a(n_1072), .o(n_1073) );
oa12s01 g780526 ( .a(n_976), .b(n_890), .c(n_906), .o(n_1072) );
oa12s01 g780527 ( .a(n_710), .b(n_890), .c(n_701), .o(n_1084) );
na02s06 g780528 ( .a(n_677), .b(n_669), .o(n_689) );
na02m04 TIMEBOOST_cell_2022 ( .a(TIMEBOOST_net_625), .b(n_14025), .o(n_14114) );
no02m04 g780530 ( .a(n_659), .b(n_423), .o(n_707) );
in01s01 g780531 ( .a(n_1062), .o(n_1063) );
oa22s01 g780532 ( .a(n_890), .b(n_809), .c(n_923), .d(n_620), .o(n_1062) );
oa22s01 g780533 ( .a(n_890), .b(n_672), .c(n_923), .d(n_556), .o(n_1103) );
oa22s01 g780534 ( .a(n_890), .b(n_422), .c(n_923), .d(n_412), .o(n_1109) );
in01s01 g780535 ( .a(n_1059), .o(n_1060) );
oa22s01 g780536 ( .a(n_923), .b(n_893), .c(n_890), .d(n_640), .o(n_1059) );
in01s01 g780537 ( .a(n_855), .o(n_764) );
no02s02 g780538 ( .a(n_705), .b(n_692), .o(n_855) );
ao22s01 g780539 ( .a(n_745), .b(n_893), .c(n_779), .d(n_748), .o(n_894) );
na02s02 g780540 ( .a(n_700), .b(n_697), .o(n_727) );
no02s01 g780541 ( .a(n_713), .b(n_46055), .o(n_767) );
in01s01 g780542 ( .a(n_778), .o(n_724) );
na02s01 g780543 ( .a(n_46055), .b(n_713), .o(n_778) );
in01s01 g780544 ( .a(n_831), .o(n_1002) );
no02s02 g780545 ( .a(n_46055), .b(FE_OCPN5097_n_694), .o(n_831) );
in01s01 g780548 ( .a(n_1111), .o(n_795) );
na02s01 g780549 ( .a(n_420), .b(FE_OCPN5097_n_694), .o(n_1111) );
in01s01 g780550 ( .a(n_936), .o(n_750) );
no02s01 g780551 ( .a(FE_OCPN5097_n_694), .b(n_420), .o(n_936) );
in01s01 g780552 ( .a(n_754), .o(n_749) );
no02s01 g780553 ( .a(n_420), .b(n_713), .o(n_754) );
in01s01 g780554 ( .a(n_845), .o(n_736) );
no02s01 g780555 ( .a(FE_OCPN5097_n_694), .b(n_521), .o(n_845) );
in01s01 g780556 ( .a(n_761), .o(n_816) );
na02s01 g780557 ( .a(n_745), .b(n_748), .o(n_761) );
na02m02 g780558 ( .a(n_662), .b(n_545), .o(n_670) );
na02s06 g780559 ( .a(n_679), .b(n_678), .o(n_698) );
in01s01 g780560 ( .a(n_869), .o(n_844) );
na02s01 g780561 ( .a(n_779), .b(n_828), .o(n_869) );
no02s03 g780562 ( .a(n_660), .b(n_923), .o(n_1026) );
no02s02 g780563 ( .a(n_713), .b(n_712), .o(n_751) );
no02s02 g780564 ( .a(n_890), .b(n_661), .o(n_1027) );
na02s01 g780565 ( .a(n_666), .b(n_695), .o(n_700) );
na02s02 g780566 ( .a(n_679), .b(n_695), .o(n_882) );
no02s01 TIMEBOOST_cell_1977 ( .a(n_420), .b(n_46055), .o(TIMEBOOST_net_603) );
in01s01 g780568 ( .a(n_742), .o(n_743) );
na02s02 g780569 ( .a(n_713), .b(n_734), .o(n_742) );
in01s01 g780570 ( .a(n_818), .o(n_776) );
no02s01 g780571 ( .a(n_713), .b(n_757), .o(n_818) );
no02s01 g780572 ( .a(n_745), .b(n_783), .o(n_819) );
in01s01 g780573 ( .a(n_1015), .o(n_1016) );
na02s01 g780574 ( .a(n_923), .b(n_610), .o(n_1015) );
na02s01 g780575 ( .a(n_906), .b(n_745), .o(n_976) );
in01s01 g780576 ( .a(n_1191), .o(n_752) );
no02s02 g780577 ( .a(n_745), .b(n_744), .o(n_1191) );
na02s02 g780578 ( .a(n_663), .b(n_546), .o(n_674) );
no02s01 g780579 ( .a(n_666), .b(n_563), .o(n_705) );
in01s01 g780580 ( .a(n_814), .o(n_790) );
na02s02 g780581 ( .a(n_745), .b(n_744), .o(n_814) );
na02s01 g780582 ( .a(n_923), .b(n_633), .o(n_1052) );
na02s02 g780583 ( .a(n_666), .b(n_672), .o(n_669) );
in01s01 g780584 ( .a(n_829), .o(n_884) );
na02s01 g780585 ( .a(n_745), .b(n_783), .o(n_829) );
in01s01 g780586 ( .a(n_675), .o(n_667) );
na02s03 g780587 ( .a(n_663), .b(n_554), .o(n_675) );
in01s01 g780588 ( .a(n_677), .o(n_706) );
na02s03 g780589 ( .a(n_666), .b(n_665), .o(n_677) );
na02s01 g780590 ( .a(n_890), .b(n_550), .o(n_1006) );
in01s01 g780591 ( .a(n_925), .o(n_898) );
no02s01 g780592 ( .a(n_867), .b(n_779), .o(n_925) );
in01s01 g780593 ( .a(n_793), .o(n_794) );
no02s02 g780594 ( .a(n_745), .b(n_773), .o(n_793) );
in01s01 g780595 ( .a(n_732), .o(n_733) );
no02s02 g780596 ( .a(n_694), .b(n_719), .o(n_732) );
na02s02 g780597 ( .a(n_713), .b(n_731), .o(n_771) );
na02s01 g780598 ( .a(n_867), .b(n_779), .o(n_977) );
na02s02 g780599 ( .a(n_745), .b(n_773), .o(n_841) );
na02s02 g780600 ( .a(n_694), .b(n_719), .o(n_753) );
in01s01 g780601 ( .a(n_690), .o(n_691) );
in01s01 g780602 ( .a(n_682), .o(n_690) );
no02s03 g780603 ( .a(n_666), .b(n_665), .o(n_682) );
in01s01 g780604 ( .a(n_710), .o(n_711) );
na02s01 g780605 ( .a(n_694), .b(n_701), .o(n_710) );
na02s01 g780606 ( .a(n_890), .b(n_905), .o(n_1053) );
in01s01 g780607 ( .a(n_725), .o(n_726) );
na02s02 g780608 ( .a(n_713), .b(n_712), .o(n_725) );
in01s01 g780609 ( .a(n_746), .o(n_747) );
no02s02 g780610 ( .a(n_713), .b(n_731), .o(n_746) );
na02s01 g780611 ( .a(n_779), .b(n_839), .o(n_868) );
in01s01 g780612 ( .a(n_664), .o(n_687) );
na02m02 g780613 ( .a(n_662), .b(n_553), .o(n_664) );
na02s01 g780614 ( .a(n_713), .b(n_757), .o(n_842) );
in01s01 g780615 ( .a(n_913), .o(n_914) );
no02s01 g780616 ( .a(n_779), .b(n_859), .o(n_913) );
na02s01 g780617 ( .a(n_679), .b(n_701), .o(n_697) );
no02s02 g780618 ( .a(n_679), .b(n_693), .o(n_730) );
in01s01 g780619 ( .a(n_985), .o(n_986) );
no02s01 g780620 ( .a(n_890), .b(n_905), .o(n_985) );
no02s01 g780621 ( .a(FE_OCPN5095_n_679), .b(FE_OFN823_n_1045), .o(n_692) );
no02s02 g780622 ( .a(n_713), .b(n_734), .o(n_781) );
in01s01 g780623 ( .a(n_684), .o(n_685) );
no02s06 g780624 ( .a(n_679), .b(n_678), .o(n_684) );
in01s01 g780625 ( .a(n_703), .o(n_704) );
na02s02 g780626 ( .a(n_679), .b(n_693), .o(n_703) );
na02s01 g780627 ( .a(n_890), .b(n_808), .o(n_1051) );
in01s01 g780628 ( .a(n_900), .o(n_945) );
no02s01 g780629 ( .a(n_779), .b(n_839), .o(n_900) );
na02s01 g780630 ( .a(n_859), .b(n_779), .o(n_951) );
in01s01 g780631 ( .a(n_887), .o(n_891) );
no02s01 g780632 ( .a(n_779), .b(n_828), .o(n_887) );
no02m02 g780633 ( .a(n_662), .b(n_413), .o(n_659) );
no02s01 g780634 ( .a(n_923), .b(n_658), .o(n_929) );
oa12s01 g780635 ( .a(n_745), .b(n_809), .c(n_808), .o(n_811) );
in01s01 g780636 ( .a(n_768), .o(n_769) );
ao12s01 g780637 ( .a(n_745), .b(n_809), .c(n_808), .o(n_768) );
in01s01 g780638 ( .a(n_865), .o(n_866) );
ao12s01 g780639 ( .a(n_745), .b(n_906), .c(n_905), .o(n_865) );
in01s01 g780655 ( .a(n_890), .o(n_923) );
in01s02 g780656 ( .a(n_779), .o(n_890) );
in01s02 g780663 ( .a(n_745), .o(n_779) );
in01s02 g780667 ( .a(n_713), .o(n_745) );
in01s02 g780672 ( .a(n_694), .o(n_713) );
in01s02 g780673 ( .a(n_679), .o(n_694) );
in01m06 g780679 ( .a(n_666), .o(n_679) );
in01m08 g780680 ( .a(n_663), .o(n_666) );
in01m06 g780681 ( .a(n_662), .o(n_663) );
oa12f08 g780682 ( .a(n_513), .b(n_657), .c(n_536), .o(n_662) );
in01s01 g780683 ( .a(n_660), .o(n_661) );
ao12s01 g780684 ( .a(n_656), .b(n_657), .c(n_655), .o(n_660) );
no02s01 g780685 ( .a(n_657), .b(n_655), .o(n_656) );
no02s01 g780686 ( .a(n_906), .b(n_905), .o(n_658) );
ao12s01 g780687 ( .a(n_651), .b(n_650), .c(n_649), .o(n_859) );
no02s01 g780688 ( .a(n_650), .b(n_649), .o(n_651) );
na02f08 g780689 ( .a(n_648), .b(n_515), .o(n_657) );
ao12s01 g780690 ( .a(n_654), .b(n_653), .c(n_652), .o(n_906) );
no02s01 g780691 ( .a(n_653), .b(n_652), .o(n_654) );
ao12s01 g780692 ( .a(n_645), .b(n_647), .c(n_497), .o(n_650) );
oa12f06 g780693 ( .a(n_511), .b(n_647), .c(n_645), .o(n_648) );
ao12s01 g780694 ( .a(n_644), .b(n_647), .c(n_643), .o(n_867) );
no02s01 g780695 ( .a(n_647), .b(n_643), .o(n_644) );
oa12s01 g780696 ( .a(n_488), .b(n_646), .c(n_480), .o(n_653) );
ao12s01 g780697 ( .a(n_642), .b(n_646), .c(n_641), .o(n_905) );
no02s01 g780698 ( .a(n_641), .b(n_646), .o(n_642) );
oa12s01 g780699 ( .a(n_639), .b(n_638), .c(n_637), .o(n_839) );
ao12f08 g780700 ( .a(n_510), .b(n_635), .c(n_492), .o(n_647) );
na02s01 g780701 ( .a(n_637), .b(n_638), .o(n_639) );
na02s01 g780702 ( .a(n_509), .b(n_636), .o(n_646) );
in01s01 g780703 ( .a(n_893), .o(n_640) );
oa12s01 g780704 ( .a(n_632), .b(n_631), .c(n_630), .o(n_893) );
na02s01 g780705 ( .a(n_631), .b(n_630), .o(n_632) );
in01s01 g780706 ( .a(n_635), .o(n_636) );
no02f08 g780707 ( .a(n_634), .b(n_475), .o(n_635) );
na02s01 g780708 ( .a(n_634), .b(n_582), .o(n_638) );
oa12s01 g780709 ( .a(n_629), .b(n_628), .c(n_627), .o(n_828) );
na02f08 g780710 ( .a(n_628), .b(n_581), .o(n_634) );
na02s01 g780711 ( .a(n_628), .b(n_627), .o(n_629) );
oa12s01 g780712 ( .a(n_482), .b(n_626), .c(n_451), .o(n_631) );
ao12s01 g780713 ( .a(n_623), .b(n_622), .c(n_621), .o(n_783) );
in01s01 g780714 ( .a(n_748), .o(n_633) );
oa12s01 g780715 ( .a(n_625), .b(n_626), .c(n_624), .o(n_748) );
no02s01 g780716 ( .a(n_622), .b(n_621), .o(n_623) );
na02s01 g780717 ( .a(n_626), .b(n_624), .o(n_625) );
na02f04 TIMEBOOST_cell_1982 ( .a(TIMEBOOST_net_605), .b(n_44428), .o(n_41362) );
na02s01 g780719 ( .a(n_468), .b(n_617), .o(n_626) );
ao12s01 g780720 ( .a(n_441), .b(n_619), .c(n_567), .o(n_622) );
no02s06 TIMEBOOST_cell_1971 ( .a(n_37608), .b(n_37116), .o(TIMEBOOST_net_600) );
in01s01 g780722 ( .a(n_809), .o(n_620) );
ao12s01 g780723 ( .a(n_613), .b(n_612), .c(n_611), .o(n_809) );
ao12s01 g780724 ( .a(n_615), .b(n_619), .c(n_614), .o(n_757) );
no02s01 g780725 ( .a(n_612), .b(n_611), .o(n_613) );
no02s01 g780726 ( .a(n_614), .b(n_619), .o(n_615) );
in01s01 g780727 ( .a(n_616), .o(n_617) );
no02f06 g780728 ( .a(n_609), .b(n_477), .o(n_616) );
ao12s01 g780729 ( .a(n_448), .b(n_608), .c(n_460), .o(n_612) );
in01s01 g780730 ( .a(n_609), .o(n_619) );
oa12f06 g780731 ( .a(n_453), .b(n_608), .c(n_466), .o(n_609) );
in01s01 g780732 ( .a(n_808), .o(n_610) );
ao12s01 g780733 ( .a(n_603), .b(n_608), .c(n_602), .o(n_808) );
oa12s01 g780734 ( .a(n_606), .b(n_605), .c(n_604), .o(n_773) );
na02s01 g780735 ( .a(n_605), .b(n_604), .o(n_606) );
no02s01 g780736 ( .a(n_608), .b(n_602), .o(n_603) );
ao12s01 g780737 ( .a(n_560), .b(n_601), .c(n_570), .o(n_605) );
oa12f08 g780738 ( .a(n_446), .b(n_596), .c(n_433), .o(n_608) );
ao22s01 g780739 ( .a(n_601), .b(n_571), .c(n_599), .d(n_572), .o(n_744) );
oa12s01 g780740 ( .a(n_595), .b(n_594), .c(n_593), .o(n_734) );
in01s01 g780741 ( .a(n_601), .o(n_599) );
in01s01 g780742 ( .a(n_596), .o(n_601) );
na02f08 g780743 ( .a(n_591), .b(n_438), .o(n_596) );
na02s01 g780744 ( .a(n_594), .b(n_593), .o(n_595) );
ao12s01 g780745 ( .a(n_589), .b(n_590), .c(n_411), .o(n_594) );
ao12s01 g780746 ( .a(n_588), .b(n_590), .c(n_587), .o(n_731) );
oa12f06 g780747 ( .a(n_435), .b(n_590), .c(n_589), .o(n_591) );
no02s01 g780748 ( .a(n_590), .b(n_587), .o(n_588) );
oa12f08 g780749 ( .a(n_426), .b(n_584), .c(n_404), .o(n_590) );
oa12s01 g780750 ( .a(n_579), .b(n_584), .c(n_578), .o(n_712) );
na02s01 g780751 ( .a(n_584), .b(n_578), .o(n_579) );
oa12f08 g780752 ( .a(n_400), .b(n_576), .c(n_416), .o(n_584) );
ao12s01 g780753 ( .a(n_569), .b(n_576), .c(n_568), .o(n_719) );
no02s01 g780754 ( .a(n_576), .b(n_568), .o(n_569) );
na02f08 g780755 ( .a(n_548), .b(n_389), .o(n_576) );
ao12s01 g780756 ( .a(n_544), .b(n_547), .c(n_543), .o(n_701) );
na02f06 g780757 ( .a(n_547), .b(n_396), .o(n_548) );
no02s01 g780758 ( .a(n_547), .b(n_543), .o(n_544) );
oa12s01 g780759 ( .a(n_566), .b(n_565), .c(n_564), .o(n_693) );
in01s01 g780760 ( .a(n_695), .o(n_550) );
ao12s01 g780761 ( .a(n_524), .b(n_523), .c(n_522), .o(n_695) );
na02s01 g780762 ( .a(n_565), .b(n_564), .o(n_566) );
no02s01 g780763 ( .a(n_523), .b(n_522), .o(n_524) );
no02f06 g780764 ( .a(n_506), .b(n_410), .o(n_547) );
no02f04 g780765 ( .a(n_505), .b(n_391), .o(n_506) );
na02s01 g780766 ( .a(n_505), .b(n_408), .o(n_523) );
oa12s01 g780767 ( .a(n_530), .b(n_558), .c(n_542), .o(n_565) );
ao12s02 g780768 ( .a(n_559), .b(n_558), .c(n_557), .o(n_678) );
na02f04 g780769 ( .a(n_490), .b(n_378), .o(n_505) );
no02s01 g780770 ( .a(n_558), .b(n_557), .o(n_559) );
in01s01 g780771 ( .a(n_490), .o(n_558) );
na02f04 g780772 ( .a(n_471), .b(n_456), .o(n_490) );
in01s01 g780773 ( .a(n_672), .o(n_556) );
ao12s01 g780774 ( .a(n_541), .b(n_540), .c(n_539), .o(n_672) );
no02s01 g780775 ( .a(n_540), .b(n_539), .o(n_541) );
oa12f02 g780776 ( .a(n_377), .b(n_455), .c(n_470), .o(n_471) );
ao12s01 g780777 ( .a(n_535), .b(n_534), .c(n_533), .o(n_665) );
no02s01 g780778 ( .a(n_455), .b(n_454), .o(n_540) );
no02s01 g780779 ( .a(n_534), .b(n_533), .o(n_535) );
ao12m02 g780780 ( .a(n_454), .b(n_430), .c(n_470), .o(n_456) );
in01s01 g780781 ( .a(n_545), .o(n_546) );
ao12s01 g780782 ( .a(n_520), .b(n_519), .c(n_518), .o(n_545) );
no02s01 g780783 ( .a(n_519), .b(n_518), .o(n_520) );
ao12s01 g780784 ( .a(n_454), .b(n_425), .c(n_365), .o(n_534) );
na02f04 g780785 ( .a(n_429), .b(n_373), .o(n_455) );
in01s02 g780786 ( .a(n_429), .o(n_430) );
na02f06 g780787 ( .a(n_425), .b(n_370), .o(n_429) );
ao12s01 g780788 ( .a(n_425), .b(n_420), .c(n_501), .o(n_519) );
in01s01 g780789 ( .a(n_553), .o(n_554) );
ao12s01 g780790 ( .a(n_529), .b(n_528), .c(n_527), .o(n_553) );
no02s01 g780791 ( .a(n_528), .b(n_527), .o(n_529) );
no02s01 g780792 ( .a(n_412), .b(n_1108), .o(n_413) );
no02s01 g780793 ( .a(n_422), .b(n_419), .o(n_423) );
no02f08 g780794 ( .a(n_528), .b(n_358), .o(n_425) );
oa12s01 g780795 ( .a(n_472), .b(n_469), .c(n_462), .o(n_496) );
ao12f08 g780796 ( .a(n_360), .b(n_367), .c(n_386), .o(n_528) );
in01s01 g780797 ( .a(n_412), .o(n_422) );
oa12s01 g780798 ( .a(n_383), .b(n_386), .c(n_382), .o(n_412) );
in01s01 g780799 ( .a(delay_sub_ln23_0_unr1_stage2_stallmux_q_1_), .o(n_607) );
na02s01 g780802 ( .a(n_386), .b(n_382), .o(n_383) );
ao12s02 g780803 ( .a(n_491), .b(n_481), .c(n_509), .o(n_510) );
no02s01 g780804 ( .a(n_468), .b(n_467), .o(n_469) );
no02s01 g780805 ( .a(n_514), .b(n_536), .o(n_655) );
in01s01 g780807 ( .a(n_1108), .o(n_419) );
oa12s01 g780808 ( .a(n_381), .b(n_380), .c(n_379), .o(n_1108) );
oa12s01 g780809 ( .a(n_598), .b(n_597), .c(beta_0), .o(n_600) );
na02s01 g780810 ( .a(n_597), .b(beta_0), .o(n_598) );
no02s02 g780811 ( .a(n_504), .b(n_420), .o(n_536) );
in01s01 g780812 ( .a(n_513), .o(n_514) );
na02s02 g780813 ( .a(n_504), .b(n_420), .o(n_513) );
na02s01 g780815 ( .a(n_380), .b(n_379), .o(n_381) );
oa12s01 g780816 ( .a(n_476), .b(n_441), .c(n_403), .o(n_468) );
no02f04 TIMEBOOST_cell_8871 ( .a(TIMEBOOST_net_2922), .b(n_39664), .o(n_39704) );
oa12s01 g780818 ( .a(n_457), .b(n_480), .c(n_479), .o(n_481) );
no02s01 g780819 ( .a(FE_RN_69_0), .b(n_371), .o(n_380) );
na02s01 g780820 ( .a(n_361), .b(n_367), .o(n_382) );
in01s01 g780821 ( .a(n_491), .o(n_492) );
na02s01 g780822 ( .a(n_488), .b(n_464), .o(n_491) );
na02s01 g780823 ( .a(n_408), .b(n_409), .o(n_410) );
no02s01 g780824 ( .a(n_452), .b(n_442), .o(n_453) );
na02s01 g780825 ( .a(n_460), .b(n_432), .o(n_602) );
no02s01 g780826 ( .a(n_434), .b(n_414), .o(n_435) );
na02s01 g780827 ( .a(n_458), .b(n_488), .o(n_641) );
na02s01 g780828 ( .a(n_567), .b(n_427), .o(n_614) );
na02s01 g780829 ( .a(n_582), .b(n_581), .o(n_627) );
no02s01 g780830 ( .a(n_467), .b(n_478), .o(n_484) );
no02s01 g780831 ( .a(n_542), .b(n_531), .o(n_557) );
na02s01 g780832 ( .a(n_415), .b(n_438), .o(n_593) );
no02s01 g780833 ( .a(n_508), .b(n_498), .o(n_511) );
na02s01 g780834 ( .a(n_499), .b(n_515), .o(n_649) );
no02s01 g780835 ( .a(n_645), .b(n_508), .o(n_643) );
no02s01 g780836 ( .a(n_395), .b(n_390), .o(n_543) );
na02s01 g780837 ( .a(n_392), .b(n_409), .o(n_522) );
na02s01 g780838 ( .a(n_426), .b(n_405), .o(n_578) );
na02s01 g780839 ( .a(n_461), .b(n_444), .o(n_462) );
no02s01 g780840 ( .a(n_589), .b(n_434), .o(n_587) );
na02s01 g780841 ( .a(n_461), .b(n_482), .o(n_624) );
in01s01 g780842 ( .a(n_571), .o(n_572) );
na02s01 g780843 ( .a(n_561), .b(n_570), .o(n_571) );
no02s01 g780844 ( .a(n_478), .b(n_445), .o(n_630) );
no02s01 g780845 ( .a(n_401), .b(n_416), .o(n_568) );
no03m10 TIMEBOOST_cell_3614 ( .a(TIMEBOOST_net_829), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .c(n_39092), .o(n_38680) );
ao12s01 g780848 ( .a(n_452), .b(n_521), .c(n_447), .o(n_611) );
ao12s01 g780849 ( .a(n_463), .b(n_521), .c(n_479), .o(n_652) );
ao12s01 g780850 ( .a(n_369), .b(n_420), .c(n_362), .o(n_518) );
oa12s01 g780851 ( .a(n_489), .b(n_521), .c(n_485), .o(n_637) );
ao12s02 g780852 ( .a(n_369), .b(n_354), .c(n_368), .o(n_370) );
ao22s01 g780853 ( .a(n_521), .b(n_476), .c(n_420), .d(n_261), .o(n_621) );
ao22s01 g780854 ( .a(n_521), .b(n_241), .c(n_420), .d(n_235), .o(n_604) );
ao22s01 g780855 ( .a(n_457), .b(n_375), .c(n_420), .d(n_501), .o(n_527) );
ao22s01 g780856 ( .a(n_457), .b(n_193), .c(n_420), .d(n_470), .o(n_539) );
ao22s01 g780857 ( .a(n_457), .b(n_368), .c(n_420), .d(n_372), .o(n_533) );
oa22s01 g780858 ( .a(n_420), .b(n_376), .c(n_457), .d(n_384), .o(n_564) );
oa22s01 g780859 ( .a(n_420), .b(beta_1), .c(n_580), .d(n_353), .o(n_597) );
ao22s01 g780860 ( .a(n_420), .b(n_476), .c(n_403), .d(n_260), .o(n_477) );
in01s01 g780862 ( .a(FE_OFN823_n_1045), .o(n_563) );
na02s01 TIMEBOOST_cell_3338 ( .a(n_35831), .b(n_35955), .o(TIMEBOOST_net_960) );
oa22s01 g780864 ( .a(n_286), .b(n_145), .c(n_285), .d(n_144), .o(n_504) );
no02s06 g780865 ( .a(n_354), .b(beta_2), .o(n_371) );
na02s04 g780867 ( .a(n_354), .b(beta_2), .o(n_363) );
na02s02 g780868 ( .a(n_354), .b(beta_3), .o(n_367) );
in01s01 g780869 ( .a(n_360), .o(n_361) );
no02s02 g780870 ( .a(n_354), .b(beta_3), .o(n_360) );
na03f10 TIMEBOOST_cell_7261 ( .a(n_35184), .b(n_35119), .c(n_35083), .o(n_35275) );
no02s02 TIMEBOOST_cell_4024 ( .a(TIMEBOOST_net_1102), .b(n_20778), .o(n_20784) );
na02s02 g780873 ( .a(n_495), .b(n_457), .o(n_515) );
in01s01 g780874 ( .a(n_414), .o(n_415) );
no02s01 g780875 ( .a(n_403), .b(n_399), .o(n_414) );
no02s02 g780876 ( .a(n_377), .b(n_393), .o(n_416) );
no02s02 g780877 ( .a(n_493), .b(n_457), .o(n_645) );
na02s01 g780878 ( .a(n_521), .b(n_424), .o(n_567) );
in01s01 g780879 ( .a(n_441), .o(n_427) );
no02s01 g780880 ( .a(n_403), .b(n_424), .o(n_441) );
na02s01 g780881 ( .a(n_439), .b(n_420), .o(n_488) );
in01s01 g780882 ( .a(n_497), .o(n_508) );
na02s01 g780883 ( .a(n_457), .b(n_493), .o(n_497) );
na02s02 g780884 ( .a(n_377), .b(n_398), .o(n_426) );
in01s01 g780885 ( .a(n_400), .o(n_401) );
na02s02 g780886 ( .a(n_377), .b(n_393), .o(n_400) );
in01s01 g780887 ( .a(n_391), .o(n_392) );
no02s01 g780888 ( .a(n_374), .b(n_385), .o(n_391) );
na02s02 g780889 ( .a(n_403), .b(n_399), .o(n_438) );
in01s01 g780890 ( .a(n_444), .o(n_445) );
na02s01 g780891 ( .a(n_403), .b(n_437), .o(n_444) );
na02s01 g780892 ( .a(n_521), .b(n_549), .o(n_570) );
na02s01 g780893 ( .a(n_374), .b(n_385), .o(n_409) );
in01s01 g780894 ( .a(n_389), .o(n_390) );
na02s02 g780895 ( .a(n_374), .b(n_387), .o(n_389) );
no02s02 g780896 ( .a(n_403), .b(n_402), .o(n_589) );
in01s01 g780897 ( .a(n_442), .o(n_460) );
no02s01 g780898 ( .a(n_403), .b(n_417), .o(n_442) );
in01s01 g780899 ( .a(n_395), .o(n_396) );
no02s01 g780900 ( .a(n_374), .b(n_387), .o(n_395) );
no02s02 g780901 ( .a(n_357), .b(n_501), .o(n_358) );
in01s01 g780902 ( .a(n_461), .o(n_451) );
na02s01 g780903 ( .a(n_443), .b(n_420), .o(n_461) );
na02s02 g780904 ( .a(n_420), .b(n_465), .o(n_581) );
in01s01 g780905 ( .a(n_432), .o(n_448) );
na02s01 g780906 ( .a(n_403), .b(n_417), .o(n_432) );
in01s01 g780907 ( .a(n_478), .o(n_472) );
no02s01 g780908 ( .a(n_403), .b(n_437), .o(n_478) );
in01s01 g780909 ( .a(n_404), .o(n_405) );
no02s02 g780910 ( .a(n_377), .b(n_398), .o(n_404) );
in01s01 g780911 ( .a(n_480), .o(n_458) );
no02s01 g780912 ( .a(n_420), .b(n_439), .o(n_480) );
in01s01 g780913 ( .a(n_467), .o(n_482) );
no02s01 g780914 ( .a(n_420), .b(n_443), .o(n_467) );
in01s01 g780915 ( .a(n_411), .o(n_434) );
na02s01 g780916 ( .a(n_403), .b(n_402), .o(n_411) );
na02s01 g780917 ( .a(n_521), .b(n_274), .o(n_582) );
in01s01 g780918 ( .a(n_560), .o(n_561) );
no02s01 g780919 ( .a(n_521), .b(n_549), .o(n_560) );
in01s01 g780920 ( .a(n_369), .o(n_365) );
no02s02 g780921 ( .a(n_357), .b(n_362), .o(n_369) );
no02s01 g780922 ( .a(n_457), .b(n_516), .o(n_542) );
in01s01 g780923 ( .a(n_530), .o(n_531) );
na02s01 g780924 ( .a(n_457), .b(n_516), .o(n_530) );
in01s01 g780925 ( .a(n_498), .o(n_499) );
no02s01 g780926 ( .a(n_457), .b(n_495), .o(n_498) );
no02s01 g780927 ( .a(n_403), .b(n_447), .o(n_452) );
in01s01 g780928 ( .a(n_463), .o(n_464) );
no02s01 g780929 ( .a(n_457), .b(n_479), .o(n_463) );
na02s01 g780930 ( .a(n_357), .b(n_372), .o(n_373) );
in01s01 g780931 ( .a(n_489), .o(n_475) );
na02s01 g780932 ( .a(n_457), .b(n_485), .o(n_489) );
no02s01 TIMEBOOST_cell_8540 ( .a(n_14454), .b(n_14456), .o(TIMEBOOST_net_2757) );
no02s02 g780935 ( .a(n_420), .b(n_240), .o(n_433) );
oa12s01 g780936 ( .a(n_377), .b(n_376), .c(n_200), .o(n_378) );
ao12s01 g780937 ( .a(n_374), .b(n_176), .c(n_375), .o(n_454) );
oa12s01 g780938 ( .a(n_374), .b(n_384), .c(n_516), .o(n_408) );
in01s01 g780939 ( .a(n_285), .o(n_286) );
ao12s01 g780940 ( .a(n_56), .b(n_284), .c(n_128), .o(n_285) );
in01s01 g780949 ( .a(n_420), .o(n_580) );
in01s01 g780960 ( .a(n_420), .o(n_521) );
in01s02 g780972 ( .a(n_420), .o(n_457) );
in01s06 g780980 ( .a(n_403), .o(n_420) );
in01s02 g780985 ( .a(n_377), .o(n_403) );
in01s02 g780988 ( .a(n_374), .o(n_377) );
in01s02 g780989 ( .a(n_357), .o(n_374) );
in01s02 g780992 ( .a(n_354), .o(n_357) );
no02f10 g780996 ( .a(n_283), .b(n_129), .o(n_354) );
ao22s01 g780997 ( .a(n_284), .b(n_139), .c(n_281), .d(n_138), .o(n_495) );
no02f10 g780998 ( .a(n_284), .b(n_108), .o(n_283) );
oa12s01 g780999 ( .a(n_280), .b(n_279), .c(n_278), .o(n_493) );
ao22s01 g781000 ( .a(n_276), .b(n_154), .c(n_277), .d(n_153), .o(n_439) );
na02s01 g781001 ( .a(n_279), .b(n_278), .o(n_280) );
in01f08 g781002 ( .a(n_281), .o(n_284) );
oa12f08 g781003 ( .a(n_269), .b(n_263), .c(n_88), .o(n_281) );
oa12s01 g781004 ( .a(n_87), .b(n_273), .c(n_100), .o(n_279) );
in01s01 g781005 ( .a(n_276), .o(n_277) );
ao12s01 g781006 ( .a(n_52), .b(n_272), .c(n_103), .o(n_276) );
ao22s01 g781007 ( .a(n_272), .b(n_142), .c(n_259), .d(n_141), .o(n_485) );
oa12s01 g781008 ( .a(n_271), .b(n_273), .c(n_270), .o(n_479) );
in01s01 g781009 ( .a(n_465), .o(n_274) );
ao12s01 g781010 ( .a(n_268), .b(n_267), .c(n_266), .o(n_465) );
na02s01 g781011 ( .a(cos_out_0), .b(FE_OFN4653_n_43918), .o(n_317) );
na02s01 g781012 ( .a(cos_out_7), .b(FE_OFN4_n_43918), .o(n_287) );
na02s01 g781013 ( .a(sin_out_19), .b(FE_OFN5_n_43918), .o(n_328) );
na02s01 g781014 ( .a(sin_out_12), .b(FE_OFN4651_n_43918), .o(n_325) );
na02s01 g781015 ( .a(cos_out_1), .b(FE_OFN1_n_43918), .o(n_321) );
na02s01 g781016 ( .a(cos_out_25), .b(FE_OFN2_n_43918), .o(n_339) );
na02s01 g781017 ( .a(sin_out_21), .b(FE_OFN5_n_43918), .o(n_290) );
na02s01 g781018 ( .a(sin_out_6), .b(FE_OFN5_n_43918), .o(n_326) );
na02s01 g781019 ( .a(cos_out_4), .b(FE_OFN1_n_43918), .o(n_345) );
na02s01 g781020 ( .a(cos_out_9), .b(FE_OFN4_n_43918), .o(n_314) );
na02s01 g781021 ( .a(sin_out_22), .b(FE_OFN5_n_43918), .o(n_310) );
na02s01 g781022 ( .a(cos_out_2), .b(FE_OFN4_n_43918), .o(n_343) );
na02s01 g781023 ( .a(cos_out_11), .b(FE_OFN4_n_43918), .o(n_303) );
na02s01 g781024 ( .a(cos_out_27), .b(FE_OFN2_n_43918), .o(n_297) );
na02s01 g781025 ( .a(sin_out_5), .b(FE_OFN5_n_43918), .o(n_311) );
na02s01 g781026 ( .a(sin_out_18), .b(FE_OFN5_n_43918), .o(n_288) );
na02s01 g781027 ( .a(sin_out_2), .b(FE_OFN4653_n_43918), .o(n_306) );
na02s01 g781028 ( .a(cos_out_3), .b(FE_OFN4_n_43918), .o(n_301) );
na02s01 g781029 ( .a(cos_out_21), .b(FE_OFN2_n_43918), .o(n_342) );
na02s01 g781030 ( .a(sin_out_28), .b(FE_OFN1_n_43918), .o(n_322) );
na02s01 g781031 ( .a(cos_out_17), .b(FE_OFN1_n_43918), .o(n_329) );
na02s01 g781032 ( .a(cos_out_31), .b(FE_OFN4_n_43918), .o(n_305) );
na02s01 g781033 ( .a(sin_out_0), .b(FE_OFN4653_n_43918), .o(n_334) );
na02s01 g781034 ( .a(sin_out_3), .b(FE_OFN4653_n_43918), .o(n_304) );
na02s01 g781035 ( .a(sin_out_25), .b(FE_OFN1_n_43918), .o(n_331) );
na02s01 g781036 ( .a(sin_out_13), .b(FE_OFN5_n_43918), .o(n_300) );
na02s01 g781037 ( .a(cos_out_22), .b(FE_OFN2_n_43918), .o(n_347) );
na02s01 g781038 ( .a(sin_out_14), .b(FE_OFN4651_n_43918), .o(n_312) );
na02s01 g781039 ( .a(cos_out_14), .b(FE_OFN4_n_43918), .o(n_344) );
na02s01 g781040 ( .a(sin_out_11), .b(FE_OFN4651_n_43918), .o(n_349) );
na02s01 g781041 ( .a(sin_out_26), .b(FE_OFN1_n_43918), .o(n_302) );
na02s01 g781042 ( .a(cos_out_12), .b(FE_OFN4_n_43918), .o(n_348) );
na02s01 g781043 ( .a(cos_out_30), .b(FE_OFN2_n_43918), .o(n_308) );
na02s01 g781045 ( .a(cos_out_18), .b(FE_OFN1_n_43918), .o(n_315) );
na02s01 g781046 ( .a(cos_out_6), .b(FE_OFN4_n_43918), .o(n_319) );
na02s01 g781047 ( .a(sin_out_10), .b(FE_OFN5_n_43918), .o(n_327) );
na02s01 g781048 ( .a(sin_out_9), .b(FE_OFN4651_n_43918), .o(n_320) );
na02s01 g781049 ( .a(sin_out_30), .b(FE_OFN1_n_43918), .o(n_294) );
na02s01 g781050 ( .a(cos_out_20), .b(FE_OFN2_n_43918), .o(n_338) );
na02s01 g781051 ( .a(cos_out_5), .b(FE_OFN4_n_43918), .o(n_341) );
na02s01 g781052 ( .a(cos_out_28), .b(FE_OFN1_n_43918), .o(n_316) );
na02s01 g781053 ( .a(cos_out_23), .b(FE_OFN2_n_43918), .o(n_298) );
na02s01 g781054 ( .a(sin_out_8), .b(FE_OFN5_n_43918), .o(n_335) );
na02s01 g781055 ( .a(cos_out_16), .b(FE_OFN4_n_43918), .o(n_336) );
na02s01 g781056 ( .a(sin_out_15), .b(FE_OFN4651_n_43918), .o(n_340) );
na02s01 g781057 ( .a(sin_out_17), .b(FE_OFN4651_n_43918), .o(n_324) );
na02s01 g781058 ( .a(cos_out_8), .b(FE_OFN4_n_43918), .o(n_313) );
na02s01 g781059 ( .a(sin_out_4), .b(FE_OFN1_n_43918), .o(n_318) );
na02s01 g781060 ( .a(cos_out_10), .b(FE_OFN4_n_43918), .o(n_330) );
na02s01 g781061 ( .a(sin_out_31), .b(FE_OFN4653_n_43918), .o(n_295) );
na02s01 g781062 ( .a(cos_out_26), .b(FE_OFN2_n_43918), .o(n_337) );
na02s01 g781063 ( .a(sin_out_29), .b(FE_OFN1_n_43918), .o(n_333) );
na02s01 g781064 ( .a(cos_out_15), .b(FE_OFN4_n_43918), .o(n_350) );
na02s01 g781065 ( .a(sin_out_27), .b(FE_OFN1_n_43918), .o(n_293) );
na02s01 g781066 ( .a(sin_out_7), .b(FE_OFN5_n_43918), .o(n_323) );
na02s01 g781067 ( .a(sin_out_16), .b(FE_OFN5_n_43918), .o(n_332) );
na02s01 g781068 ( .a(cos_out_29), .b(FE_OFN1_n_43918), .o(n_292) );
na02s01 g781069 ( .a(cos_out_24), .b(FE_OFN2_n_43918), .o(n_291) );
na02s01 g781070 ( .a(cos_out_19), .b(FE_OFN4_n_43918), .o(n_309) );
na02s01 g781071 ( .a(cos_out_13), .b(FE_OFN4_n_43918), .o(n_346) );
na02s01 g781072 ( .a(sin_out_24), .b(FE_OFN1_n_43918), .o(n_296) );
na02s01 g781073 ( .a(sin_out_1), .b(FE_OFN4653_n_43918), .o(n_299) );
na02s01 g781074 ( .a(sin_out_23), .b(FE_OFN5_n_43918), .o(n_289) );
no02s01 g781075 ( .a(n_267), .b(n_266), .o(n_268) );
na02s01 g781076 ( .a(n_270), .b(n_273), .o(n_271) );
na02m08 g781077 ( .a(n_262), .b(n_48), .o(n_269) );
no02f08 g781078 ( .a(n_262), .b(n_46), .o(n_263) );
oa12s01 g781079 ( .a(n_256), .b(n_255), .c(n_254), .o(n_443) );
in01s01 g781080 ( .a(n_262), .o(n_273) );
oa12f10 g781081 ( .a(n_163), .b(n_258), .c(n_159), .o(n_262) );
na02s01 g781082 ( .a(n_254), .b(n_255), .o(n_256) );
in01s01 g781083 ( .a(n_259), .o(n_272) );
oa12s01 g781084 ( .a(n_89), .b(n_258), .c(n_120), .o(n_259) );
na02s01 g781085 ( .a(state_cordic_1_), .b(n_282), .o(n_43918) );
oa12s01 g781086 ( .a(n_72), .b(n_258), .c(n_140), .o(n_267) );
in01s01 g781087 ( .a(n_476), .o(n_261) );
oa12s01 g781088 ( .a(n_253), .b(n_252), .c(n_251), .o(n_476) );
in01s01 g781089 ( .a(n_424), .o(n_260) );
ao12s01 g781090 ( .a(n_248), .b(n_247), .c(n_246), .o(n_424) );
oa12s01 g781091 ( .a(n_250), .b(n_258), .c(n_249), .o(n_437) );
no02s01 g781092 ( .a(n_275), .b(n_264), .o(n_282) );
no02s01 g781093 ( .a(n_247), .b(n_246), .o(n_248) );
na02s01 g781094 ( .a(n_249), .b(n_258), .o(n_250) );
na02s01 g781095 ( .a(n_251), .b(n_252), .o(n_253) );
ao12s01 g781096 ( .a(n_105), .b(n_245), .c(n_155), .o(n_255) );
in01s01 g781097 ( .a(mux_while_ln12_psv_q_8_), .o(n_275) );
na02s06 TIMEBOOST_cell_8638 ( .a(n_30842), .b(n_27131), .o(TIMEBOOST_net_2806) );
no02s01 g781100 ( .a(n_74), .b(n_245), .o(n_252) );
oa12s01 g781101 ( .a(n_70), .b(n_244), .c(n_135), .o(n_247) );
oa12s01 g781102 ( .a(n_238), .b(n_244), .c(n_237), .o(n_447) );
no02s01 g781103 ( .a(n_244), .b(n_94), .o(n_245) );
na02s01 g781104 ( .a(n_244), .b(n_237), .o(n_238) );
no02s01 g781105 ( .a(n_549), .b(n_241), .o(n_240) );
no03s02 TIMEBOOST_cell_8148 ( .a(n_12768), .b(n_12247), .c(n_12942), .o(TIMEBOOST_net_2705) );
no02s01 g781107 ( .a(n_257), .b(n_264), .o(n_265) );
na02m08 TIMEBOOST_cell_8549 ( .a(TIMEBOOST_net_2761), .b(n_19301), .o(n_19445) );
oa12s01 g781109 ( .a(n_234), .b(n_233), .c(n_232), .o(n_417) );
na02s01 g781110 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_7_), .o(n_257) );
na02s01 g781111 ( .a(n_233), .b(n_232), .o(n_234) );
no02f04 TIMEBOOST_cell_1788 ( .a(TIMEBOOST_net_508), .b(FE_OCP_RBN6831_n_15676), .o(n_15680) );
in01s01 g781113 ( .a(n_241), .o(n_235) );
ao12s01 g781114 ( .a(n_230), .b(n_229), .c(n_228), .o(n_241) );
ao22s01 g781115 ( .a(n_226), .b(n_125), .c(n_225), .d(n_126), .o(n_549) );
no02s01 g781117 ( .a(n_228), .b(n_229), .o(n_230) );
no03s10 TIMEBOOST_cell_2146 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_4_), .o(n_11686) );
oa12s01 g781119 ( .a(n_161), .b(n_224), .c(n_111), .o(n_233) );
na02s01 g781120 ( .a(n_143), .b(n_224), .o(n_229) );
in01s01 g781121 ( .a(n_225), .o(n_226) );
oa12s01 g781122 ( .a(n_42), .b(n_222), .c(n_109), .o(n_225) );
no02s01 g781123 ( .a(n_236), .b(n_264), .o(n_243) );
no02m06 TIMEBOOST_cell_4293 ( .a(n_29371), .b(n_29561), .o(TIMEBOOST_net_1237) );
ao12s01 g781125 ( .a(n_218), .b(n_222), .c(n_217), .o(n_399) );
oa22s01 g781126 ( .a(n_219), .b(n_114), .c(n_220), .d(n_113), .o(n_402) );
na02s01 g781127 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_6_), .o(n_236) );
na02s01 g781128 ( .a(n_222), .b(n_75), .o(n_224) );
no02s01 g781129 ( .a(n_222), .b(n_217), .o(n_218) );
na03f04 TIMEBOOST_cell_3561 ( .a(FE_OCP_RBN5041_n_14201), .b(FE_RN_2260_0), .c(FE_RN_481_0), .o(n_14283) );
in01s01 g781132 ( .a(n_219), .o(n_220) );
oa12s01 g781133 ( .a(n_116), .b(n_215), .c(n_82), .o(n_219) );
oa12f10 g781134 ( .a(n_83), .b(n_214), .c(n_115), .o(n_222) );
ao22s01 g781135 ( .a(n_215), .b(n_134), .c(n_214), .d(n_133), .o(n_398) );
no02s01 g781136 ( .a(n_221), .b(n_264), .o(n_227) );
oa12s01 g781137 ( .a(n_212), .b(n_211), .c(n_210), .o(n_393) );
na02s01 g781138 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_5_), .o(n_221) );
na02s01 g781139 ( .a(n_210), .b(n_211), .o(n_212) );
in01s01 g781140 ( .a(n_214), .o(n_215) );
na02f10 g781141 ( .a(n_205), .b(n_207), .o(n_214) );
oa12f08 g781143 ( .a(beta_12), .b(n_206), .c(n_59), .o(n_205) );
oa12s01 g781144 ( .a(n_127), .b(n_208), .c(n_92), .o(n_211) );
ao22s01 g781145 ( .a(n_206), .b(n_147), .c(n_208), .d(n_148), .o(n_387) );
oa22s01 g781146 ( .a(n_203), .b(n_96), .c(n_202), .d(n_97), .o(n_385) );
no02s01 g781148 ( .a(n_209), .b(n_264), .o(n_213) );
na02s01 g781149 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_4_), .o(n_209) );
in01s01 g781150 ( .a(n_202), .o(n_203) );
ao12s01 g781151 ( .a(n_57), .b(n_199), .c(n_101), .o(n_202) );
in01s01 g781152 ( .a(n_206), .o(n_208) );
ao12f10 g781153 ( .a(n_112), .b(n_199), .c(n_130), .o(n_206) );
in01s01 g781154 ( .a(n_384), .o(n_376) );
oa22s01 g781155 ( .a(n_194), .b(n_149), .c(n_199), .d(n_150), .o(n_384) );
in01s01 g781157 ( .a(n_516), .o(n_200) );
oa12s01 g781158 ( .a(n_190), .b(n_189), .c(n_188), .o(n_516) );
na02s01 g781159 ( .a(n_189), .b(n_188), .o(n_190) );
no02s01 g781160 ( .a(n_198), .b(n_264), .o(n_204) );
in01s01 g781161 ( .a(n_199), .o(n_194) );
no02m10 g781162 ( .a(n_183), .b(n_180), .o(n_199) );
na02s01 g781163 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_3_), .o(n_198) );
ao12m10 g781164 ( .a(n_77), .b(n_182), .c(n_49), .o(n_183) );
oa12s01 g781165 ( .a(n_118), .b(n_182), .c(n_63), .o(n_189) );
in01s01 g781166 ( .a(n_470), .o(n_193) );
oa22s01 g781167 ( .a(n_178), .b(n_131), .c(n_182), .d(n_132), .o(n_470) );
no02s10 g781169 ( .a(n_182), .b(n_58), .o(n_180) );
no02s01 g781171 ( .a(n_177), .b(n_264), .o(n_181) );
in01s01 g781172 ( .a(n_182), .o(n_178) );
no02m20 g781173 ( .a(n_175), .b(n_170), .o(n_182) );
na02s01 g781175 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_2_), .o(n_177) );
ao12m10 g781176 ( .a(n_67), .b(n_174), .c(beta_31), .o(n_175) );
in01s01 g781177 ( .a(n_368), .o(n_372) );
ao22s01 g781178 ( .a(n_174), .b(n_124), .c(n_171), .d(n_123), .o(n_368) );
in01s06 g781191 ( .a(n_186), .o(n_179) );
in01s01 g781193 ( .a(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_24105) );
in01s01 g781195 ( .a(n_174), .o(n_171) );
ao12s10 g781196 ( .a(n_45), .b(n_162), .c(n_117), .o(n_174) );
no02s01 g781198 ( .a(n_168), .b(n_264), .o(n_173) );
ao12s01 g781199 ( .a(n_93), .b(n_157), .c(n_104), .o(n_172) );
in01s01 g781200 ( .a(n_362), .o(n_176) );
oa22s01 g781201 ( .a(n_164), .b(n_136), .c(n_169), .d(n_137), .o(n_362) );
in01s06 g781202 ( .a(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_17427) );
na02s01 g781204 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_1_), .o(n_168) );
na02s01 g781205 ( .a(n_95), .b(n_155), .o(n_156) );
na02s03 g781206 ( .a(n_121), .b(n_158), .o(n_159) );
ao22s03 g781207 ( .a(n_90), .b(n_158), .c(n_85), .d(beta_26), .o(n_163) );
in01s01 g781208 ( .a(n_501), .o(n_375) );
oa12s01 g781209 ( .a(n_166), .b(n_165), .c(beta_3), .o(n_501) );
na02s01 g781213 ( .a(n_104), .b(n_84), .o(n_105) );
no02s01 g781214 ( .a(n_120), .b(n_119), .o(n_121) );
no02s01 g781215 ( .a(n_93), .b(n_94), .o(n_95) );
in01s01 g781216 ( .a(n_160), .o(n_161) );
na02s01 g781217 ( .a(n_143), .b(n_54), .o(n_160) );
na02s01 g781218 ( .a(n_165), .b(beta_3), .o(n_166) );
in01s01 g781219 ( .a(n_169), .o(n_164) );
in01s06 g781220 ( .a(n_162), .o(n_169) );
oa12s20 g781221 ( .a(n_146), .b(n_78), .c(n_12), .o(n_162) );
ao12s02 g781222 ( .a(n_110), .b(n_128), .c(n_46055), .o(n_129) );
ao12s01 g781223 ( .a(n_11), .b(n_62), .c(beta_31), .o(n_99) );
oa12s02 g781224 ( .a(beta_22), .b(n_152), .c(beta_31), .o(n_157) );
ao12s03 g781225 ( .a(n_7), .b(n_116), .c(n_40), .o(n_115) );
na02s06 g781226 ( .a(n_80), .b(beta_31), .o(n_130) );
in01s01 g781227 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_0_), .o(n_167) );
na02s03 g781229 ( .a(n_102), .b(n_61), .o(n_112) );
na02s01 g781230 ( .a(n_103), .b(beta_31), .o(n_85) );
no02s03 g781231 ( .a(n_82), .b(n_81), .o(n_83) );
na02s02 g781232 ( .a(n_107), .b(n_106), .o(n_108) );
no02s01 g781233 ( .a(n_109), .b(n_68), .o(n_143) );
na02s01 g781234 ( .a(n_101), .b(n_38), .o(n_80) );
in01s01 g781235 ( .a(n_131), .o(n_132) );
na02s01 g781236 ( .a(n_64), .b(n_118), .o(n_131) );
in01s01 g781237 ( .a(n_136), .o(n_137) );
na02s01 g781238 ( .a(n_117), .b(n_44), .o(n_136) );
in01s01 g781239 ( .a(n_138), .o(n_139) );
na02s01 g781240 ( .a(n_106), .b(n_128), .o(n_138) );
in01s01 g781241 ( .a(n_141), .o(n_142) );
na02s01 g781242 ( .a(n_158), .b(n_103), .o(n_141) );
in01s01 g781243 ( .a(n_149), .o(n_150) );
na02s01 g781244 ( .a(n_102), .b(n_101), .o(n_149) );
no02s01 g781245 ( .a(n_111), .b(n_53), .o(n_228) );
no02s01 g781246 ( .a(n_43), .b(n_109), .o(n_217) );
in01s01 g781247 ( .a(n_133), .o(n_134) );
na02s01 g781248 ( .a(n_55), .b(n_116), .o(n_133) );
no02s01 g781249 ( .a(n_86), .b(n_100), .o(n_270) );
no02s01 g781250 ( .a(n_140), .b(n_73), .o(n_249) );
na02s01 g781251 ( .a(n_79), .b(n_146), .o(n_165) );
in01s01 g781252 ( .a(n_147), .o(n_148) );
na02s01 g781253 ( .a(n_127), .b(n_91), .o(n_147) );
no02s01 g781254 ( .a(n_69), .b(n_152), .o(n_251) );
no02s01 g781255 ( .a(n_135), .b(n_71), .o(n_237) );
no02s01 g781256 ( .a(n_66), .b(n_264), .o(n_98) );
ao12s01 g781257 ( .a(n_122), .b(n_7), .c(beta_18), .o(n_232) );
ao12s01 g781258 ( .a(n_7), .b(beta_20), .c(beta_19), .o(n_94) );
in01s01 g781259 ( .a(n_144), .o(n_145) );
oa12s01 g781260 ( .a(n_107), .b(n_110), .c(n_46055), .o(n_144) );
in01s01 g781261 ( .a(n_75), .o(n_76) );
oa12s01 g781262 ( .a(beta_31), .b(beta_16), .c(beta_15), .o(n_75) );
in01s01 g781263 ( .a(n_125), .o(n_126) );
ao12s01 g781264 ( .a(n_68), .b(n_46055), .c(beta_16), .o(n_125) );
in01s01 g781265 ( .a(n_96), .o(n_97) );
ao12s01 g781266 ( .a(n_60), .b(n_46055), .c(beta_10), .o(n_96) );
ao12s01 g781267 ( .a(n_7), .b(beta_24), .c(beta_23), .o(n_120) );
in01s01 g781268 ( .a(n_89), .o(n_90) );
oa12s01 g781269 ( .a(n_7), .b(beta_24), .c(beta_23), .o(n_89) );
in01s01 g781270 ( .a(n_113), .o(n_114) );
ao12s01 g781271 ( .a(n_81), .b(n_46055), .c(beta_14), .o(n_113) );
in01s01 g781272 ( .a(n_153), .o(n_154) );
ao12s01 g781273 ( .a(n_119), .b(n_7), .c(beta_26), .o(n_153) );
ao12s01 g781274 ( .a(n_93), .b(n_46055), .c(beta_22), .o(n_254) );
in01s01 g781275 ( .a(n_104), .o(n_74) );
oa12s01 g781276 ( .a(n_7), .b(beta_20), .c(beta_19), .o(n_104) );
oa22s01 g781277 ( .a(n_46055), .b(beta_12), .c(n_7), .d(n_27), .o(n_210) );
oa22s01 g781278 ( .a(n_46055), .b(beta_28), .c(n_7), .d(n_88), .o(n_278) );
oa22s01 g781279 ( .a(n_18), .b(n_46055), .c(n_7), .d(beta_20), .o(n_246) );
oa22s01 g781280 ( .a(n_77), .b(n_46055), .c(n_7), .d(beta_8), .o(n_188) );
in01s01 g781281 ( .a(n_123), .o(n_124) );
oa22s01 g781282 ( .a(n_67), .b(n_46055), .c(n_7), .d(beta_6), .o(n_123) );
oa22s01 g781283 ( .a(n_13), .b(n_46055), .c(n_7), .d(beta_24), .o(n_266) );
in01s01 g781284 ( .a(delay_sub_ln23_0_unr1_stage2_stallmux_q_0_), .o(n_151) );
in01s01 g781287 ( .a(state_cordic_1_), .o(n_66) );
in01s01 g781289 ( .a(n_63), .o(n_64) );
no02s01 g781290 ( .a(n_46055), .b(beta_7), .o(n_63) );
in01s01 g781291 ( .a(n_52), .o(n_158) );
no02s01 g781292 ( .a(beta_31), .b(beta_25), .o(n_52) );
no02s01 g781293 ( .a(beta_22), .b(beta_31), .o(n_93) );
na02s01 g781294 ( .a(beta_31), .b(beta_9), .o(n_101) );
in01s01 g781295 ( .a(n_82), .o(n_55) );
no02s01 g781296 ( .a(beta_31), .b(beta_13), .o(n_82) );
in01s01 g781297 ( .a(n_62), .o(n_111) );
na02s01 g781298 ( .a(beta_31), .b(beta_17), .o(n_62) );
no02s01 g781299 ( .a(beta_31), .b(beta_15), .o(n_109) );
na02s01 g781300 ( .a(n_7), .b(n_47), .o(n_46) );
na02s01 g781301 ( .a(beta_29), .b(beta_31), .o(n_128) );
in01s06 g781302 ( .a(n_44), .o(n_45) );
na02s06 g781303 ( .a(beta_31), .b(beta_5), .o(n_44) );
na02s01 g781304 ( .a(n_46055), .b(beta_7), .o(n_118) );
no02s01 g781305 ( .a(beta_31), .b(beta_16), .o(n_68) );
na02s02 g781306 ( .a(n_1), .b(n_51), .o(n_59) );
no02s01 g781307 ( .a(beta_31), .b(beta_14), .o(n_81) );
in01s01 g781308 ( .a(n_57), .o(n_102) );
no02s01 g781309 ( .a(beta_31), .b(beta_9), .o(n_57) );
no02s01 g781310 ( .a(n_7), .b(n_47), .o(n_48) );
in01s01 g781311 ( .a(n_60), .o(n_61) );
no02s01 g781312 ( .a(beta_31), .b(beta_10), .o(n_60) );
in01s01 g781313 ( .a(n_53), .o(n_54) );
no02s01 g781314 ( .a(beta_31), .b(beta_17), .o(n_53) );
na02s01 g781315 ( .a(beta_31), .b(beta_13), .o(n_116) );
na02s01 g781316 ( .a(beta_31), .b(beta_25), .o(n_103) );
in01s01 g781317 ( .a(n_56), .o(n_106) );
no02s01 g781318 ( .a(beta_29), .b(beta_31), .o(n_56) );
in01s06 g781319 ( .a(n_65), .o(n_117) );
no02s06 g781320 ( .a(beta_31), .b(beta_5), .o(n_65) );
in01s01 g781321 ( .a(n_42), .o(n_43) );
na02s01 g781322 ( .a(n_46055), .b(beta_15), .o(n_42) );
no02s01 g781323 ( .a(n_7), .b(beta_19), .o(n_135) );
no02s01 g781324 ( .a(n_7), .b(beta_26), .o(n_119) );
in01s01 g781325 ( .a(n_78), .o(n_79) );
no02s40 g781326 ( .a(n_1), .b(beta_4), .o(n_78) );
in01s01 g781327 ( .a(n_84), .o(n_152) );
na02s01 g781328 ( .a(n_7), .b(beta_21), .o(n_84) );
in01s01 g781329 ( .a(n_69), .o(n_155) );
no02m01 g781330 ( .a(beta_21), .b(n_7), .o(n_69) );
na02s02 g781331 ( .a(n_1), .b(beta_7), .o(n_58) );
no02s01 g781332 ( .a(n_7), .b(beta_23), .o(n_140) );
no02s03 g781333 ( .a(n_1), .b(beta_7), .o(n_49) );
no02s02 g781334 ( .a(n_7), .b(beta_18), .o(n_122) );
in01s01 g781335 ( .a(n_70), .o(n_71) );
na02s01 g781336 ( .a(beta_19), .b(n_7), .o(n_70) );
in01s01 g781337 ( .a(n_91), .o(n_92) );
na02s01 g781338 ( .a(n_51), .b(n_46055), .o(n_91) );
in01s01 g781339 ( .a(n_72), .o(n_73) );
na02s01 g781340 ( .a(n_7), .b(beta_23), .o(n_72) );
in01s01 g781341 ( .a(n_86), .o(n_87) );
no02s01 g781342 ( .a(n_46055), .b(n_47), .o(n_86) );
na02s40 g781343 ( .a(n_29), .b(beta_4), .o(n_146) );
na02s01 g781344 ( .a(n_110), .b(beta_31), .o(n_107) );
na02s01 g781345 ( .a(n_7), .b(beta_11), .o(n_127) );
no02s01 g781346 ( .a(n_7), .b(beta_27), .o(n_100) );
in01s01 g781347 ( .a(beta_27), .o(n_47) );
in01s01 g781348 ( .a(beta_1), .o(n_353) );
in01s01 g781349 ( .a(beta_0), .o(n_50) );
in01s06 g781350 ( .a(beta_3), .o(n_12) );
in01s01 g781351 ( .a(beta_28), .o(n_88) );
in01s01 g781352 ( .a(beta_18), .o(n_11) );
in01s01 g781353 ( .a(beta_30), .o(n_110) );
in01s01 g781354 ( .a(beta_10), .o(n_38) );
in01s80 g781357 ( .a(beta_31), .o(n_29) );
in01s80 g781366 ( .a(beta_31), .o(n_1) );
in01s01 g781390 ( .a(beta_24), .o(n_13) );
in01s02 g781391 ( .a(beta_8), .o(n_77) );
in01s01 g781392 ( .a(beta_14), .o(n_40) );
in01s02 g781393 ( .a(beta_6), .o(n_67) );
in01s01 g781394 ( .a(rst), .o(n_264) );
in01s01 g781395 ( .a(beta_11), .o(n_51) );
in01s01 g781396 ( .a(beta_12), .o(n_27) );
in01s01 g781397 ( .a(beta_20), .o(n_18) );
in01m01 g782628 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_20_), .o(n_44021) );
in01s01 g782633 ( .a(n_44060), .o(n_509) );
na02f20 g782634 ( .a(n_40654), .b(n_40655), .o(n_44027) );
oa12s06 g782635 ( .a(n_44610), .b(n_40604), .c(n_40611), .o(n_44028) );
oa12f04 g782636 ( .a(n_38028), .b(n_37985), .c(n_37638), .o(n_44029) );
ao12s02 g782637 ( .a(n_44875), .b(n_38270), .c(FE_OCP_RBN4027_n_37577), .o(n_44030) );
in01s01 g782638 ( .a(n_44032), .o(n_44033) );
oa12s02 g782639 ( .a(n_44877), .b(n_37965), .c(n_38290), .o(n_44032) );
in01s02 g782640 ( .a(n_44034), .o(n_44035) );
ao12s06 g782641 ( .a(n_44875), .b(n_37490), .c(n_38268), .o(n_44034) );
oa12f08 g782642 ( .a(n_37916), .b(n_37891), .c(n_37835), .o(n_44036) );
oa12s02 g782643 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_36950), .c(n_36992), .o(n_44037) );
oa12s02 g782644 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_36991), .c(FE_OCP_RBN2338_delay_sub_ln21_0_unr23_stage9_stallmux_q_20_), .o(n_44038) );
no02s03 g782645 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_18_), .b(delay_add_ln22_unr23_stage9_stallmux_q_19_), .o(n_44039) );
oa12s01 g782647 ( .a(FE_OCPN950_n_44180), .b(FE_OCP_RBN4925_n_34980), .c(n_35774), .o(n_44040) );
ao12s02 g782648 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n_32312), .c(n_32492), .o(n_44042) );
ao12s02 g782651 ( .a(n_28836), .b(n_28883), .c(n_28690), .o(n_44045) );
ao12s04 g782652 ( .a(n_27923), .b(n_27931), .c(n_27854), .o(n_44046) );
in01s02 g782657 ( .a(n_44051), .o(n_44052) );
ao12s04 g782658 ( .a(n_15142), .b(n_15228), .c(n_14239), .o(n_44051) );
in01m02 g782659 ( .a(n_44053), .o(n_44054) );
ao12m02 g782660 ( .a(FE_OCP_RBN5911_n_44563), .b(n_10411), .c(n_10270), .o(n_44053) );
oa12f02 g782662 ( .a(FE_OCP_RBN4240_n_44594), .b(n_9035), .c(n_9034), .o(n_44055) );
no02m06 g782663 ( .a(n_8532), .b(n_8634), .o(n_44057) );
oa12m06 g782664 ( .a(n_8493), .b(n_8443), .c(n_8316), .o(n_44058) );
ao12s02 g782665 ( .a(FE_OCP_RBN5662_n_2438), .b(n_3127), .c(n_3217), .o(n_44059) );
ao12s01 g782666 ( .a(n_485), .b(n_457), .c(n_465), .o(n_44060) );
oa12m02 g783677 ( .a(n_15999), .b(n_15856), .c(n_15942), .o(n_45331) );
no02f08 g783678 ( .a(n_15942), .b(n_15856), .o(n_45332) );
in01s02 g783785 ( .a(n_45462), .o(n_45463) );
no02s02 g783786 ( .a(n_47008), .b(FE_OCP_RBN6781_n_4046), .o(n_45462) );
na02f04 g783817 ( .a(n_15392), .b(n_15353), .o(n_45502) );
ao12m06 g783818 ( .a(n_8531), .b(n_8471), .c(n_7594), .o(n_45503) );
ao12m04 g783820 ( .a(n_2424), .b(n_2575), .c(n_2349), .o(n_45505) );
na02s01 g783821 ( .a(n_2575), .b(n_2349), .o(n_45506) );
ao12m40 g783822 ( .a(n_40619), .b(n_45507), .c(n_44610), .o(n_45508) );
na02m80 g783823 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .b(delay_xor_ln22_unr28_stage10_stallmux_q_2_), .o(n_45507) );
na02s20 g783824 ( .a(n_40611), .b(n_44610), .o(n_45511) );
in01s20 g783825 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .o(n_40611) );
na02m10 g783826 ( .a(n_45512), .b(n_44610), .o(n_45513) );
in01s10 g783827 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_2_), .o(n_45512) );
oa12m02 g783828 ( .a(FE_RN_1873_0), .b(n_39596), .c(n_39607), .o(n_45514) );
na02s06 g783830 ( .a(n_32090), .b(n_31880), .o(n_45516) );
in01s04 g783831 ( .a(n_45517), .o(n_45518) );
na02m10 g783832 ( .a(n_32090), .b(n_31880), .o(n_45517) );
na02f06 g783834 ( .a(n_14586), .b(n_14612), .o(n_45520) );
in01s01 g783839 ( .a(n_45528), .o(n_45529) );
no02s01 g783840 ( .a(n_18237), .b(n_45527), .o(n_45528) );
na02s01 g783841 ( .a(n_45525), .b(FE_RN_21_0), .o(n_45527) );
in01s01 g783842 ( .a(n_17533), .o(n_45525) );
oa12m04 g783844 ( .a(FE_RN_1873_0), .b(n_39594), .c(n_39579), .o(n_45530) );
oa12s02 g783846 ( .a(n_25824), .b(n_25678), .c(n_25707), .o(n_45532) );
no02f02 g783847 ( .a(n_25707), .b(n_25678), .o(n_45533) );
no02s02 g784066 ( .a(n_7), .b(FE_OCPN5095_n_679), .o(n_45808) );
no02s02 g784067 ( .a(n_831), .b(n_45812), .o(n_45813) );
oa12s01 g784068 ( .a(n_1111), .b(n_45808), .c(n_936), .o(n_45814) );
no02s01 g784069 ( .a(n_802), .b(n_45812), .o(n_45815) );
oa12s01 g784070 ( .a(n_1002), .b(n_851), .c(n_45808), .o(n_45816) );
no02m04 TIMEBOOST_cell_1926 ( .a(TIMEBOOST_net_577), .b(FE_OCP_RBN6209_n_11486), .o(n_11723) );
oa12s01 g784072 ( .a(n_1002), .b(n_1194), .c(n_45812), .o(n_45818) );
ao12s01 g784073 ( .a(n_45812), .b(n_970), .c(n_1002), .o(n_45819) );
oa12m01 g784077 ( .a(n_7285), .b(n_7284), .c(n_7283), .o(n_45820) );
na02s03 g784078 ( .a(n_7598), .b(n_45824), .o(n_45825) );
na02s01 g784080 ( .a(n_7654), .b(n_45820), .o(n_45826) );
no02m02 g784081 ( .a(n_8199), .b(n_45820), .o(n_45827) );
na02s03 g784082 ( .a(n_8199), .b(n_45824), .o(n_45828) );
ao12m08 g784097 ( .a(n_45845), .b(n_45887), .c(n_7225), .o(n_45846) );
no02s01 g784100 ( .a(n_7156), .b(delay_add_ln22_unr5_stage3_stallmux_q_14_), .o(n_45843) );
no02s01 g784108 ( .a(n_6866), .b(n_45858), .o(n_45861) );
na02s02 g784111 ( .a(n_6851), .b(n_6895), .o(n_45858) );
no02s01 g784112 ( .a(n_45858), .b(n_6819), .o(n_45863) );
na02s02 TIMEBOOST_cell_3198 ( .a(n_25954), .b(n_25748), .o(TIMEBOOST_net_890) );
no02f08 g784115 ( .a(n_47176), .b(n_45858), .o(n_45865) );
na02s02 g784119 ( .a(n_7212), .b(n_7211), .o(n_45866) );
na02s01 g784120 ( .a(n_45873), .b(n_45866), .o(n_45871) );
ao12m08 g784122 ( .a(n_45874), .b(n_45846), .c(n_45866), .o(n_45875) );
no02s01 g784125 ( .a(n_7212), .b(n_7211), .o(n_45872) );
no02s01 g784131 ( .a(n_7136), .b(n_7135), .o(n_45878) );
ao12m08 g784134 ( .a(n_45880), .b(n_7659), .c(n_45884), .o(n_45887) );
na02s02 g784137 ( .a(n_7136), .b(n_7135), .o(n_45884) );
na02s01 g784138 ( .a(n_45879), .b(n_45884), .o(n_45889) );
no02s02 TIMEBOOST_cell_6794 ( .a(TIMEBOOST_net_2154), .b(n_4306), .o(n_4588) );
ao12s01 g784144 ( .a(n_45894), .b(n_37825), .c(n_37790), .o(n_45895) );
oa22s01 g784146 ( .a(n_36898), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_0_), .c(n_45890), .d(n_37023), .o(n_45896) );
ao22s01 g784147 ( .a(n_38193), .b(n_37225), .c(n_38221), .d(n_45894), .o(n_45897) );
oa12s01 g784148 ( .a(n_38525), .b(n_38174), .c(n_45890), .o(n_45898) );
ao12s02 g784149 ( .a(n_38372), .b(n_38371), .c(n_45894), .o(n_45899) );
oa12f08 g784336 ( .a(n_5384), .b(n_6315), .c(n_6304), .o(n_46137) );
oa22s02 g784337 ( .a(FE_OFN4789_n_46137), .b(n_5286), .c(FE_OCP_RBN6200_FE_OFN789_n_46195), .d(n_5379), .o(n_46141) );
oa22m02 g784338 ( .a(FE_OCP_RBN6195_FE_OFN789_n_46195), .b(n_5913), .c(FE_OFN4789_n_46137), .d(n_5906), .o(n_46143) );
oa22s02 g784339 ( .a(FE_OFN4789_n_46137), .b(n_5489), .c(FE_OCP_RBN6195_FE_OFN789_n_46195), .d(n_5527), .o(n_46145) );
oa22s02 g784340 ( .a(FE_OFN4789_n_46137), .b(n_5538), .c(FE_OCP_RBN6195_FE_OFN789_n_46195), .d(n_5569), .o(n_46146) );
oa22s02 g784341 ( .a(FE_OFN768_n_46137), .b(n_6365), .c(FE_OCP_RBN6196_FE_OFN789_n_46195), .d(n_6376), .o(n_46147) );
oa22s02 g784342 ( .a(FE_OCP_RBN6199_FE_OFN789_n_46195), .b(n_5408), .c(FE_OFN4789_n_46137), .d(n_5350), .o(n_46148) );
oa22m02 g784343 ( .a(FE_OFN768_n_46137), .b(n_6318), .c(FE_OCP_RBN6196_FE_OFN789_n_46195), .d(n_46994), .o(n_46149) );
oa22m02 g784344 ( .a(FE_OFN4788_n_46137), .b(n_6137), .c(FE_OCP_RBN6196_FE_OFN789_n_46195), .d(n_6146), .o(n_46150) );
oa22s02 g784345 ( .a(FE_OCP_RBN6196_FE_OFN789_n_46195), .b(n_6248), .c(FE_OFN768_n_46137), .d(n_6206), .o(n_46151) );
oa22s02 g784346 ( .a(FE_OFN4788_n_46137), .b(n_6005), .c(FE_OCP_RBN6195_FE_OFN789_n_46195), .d(n_6047), .o(n_46152) );
oa22s02 g784347 ( .a(FE_OFN4789_n_46137), .b(n_5676), .c(FE_OCP_RBN6195_FE_OFN789_n_46195), .d(n_5748), .o(n_46153) );
oa22m02 g784348 ( .a(FE_OFN768_n_46137), .b(n_6280), .c(FE_OCP_RBN6196_FE_OFN789_n_46195), .d(n_6301), .o(n_46154) );
oa22f02 g784349 ( .a(FE_OCP_RBN6196_FE_OFN789_n_46195), .b(n_6267), .c(FE_OFN768_n_46137), .d(n_6245), .o(n_46155) );
oa22s02 g784350 ( .a(FE_OCP_RBN6195_FE_OFN789_n_46195), .b(n_5483), .c(FE_OFN4789_n_46137), .d(n_5418), .o(n_46156) );
oa22f02 g784351 ( .a(FE_OFN768_n_46137), .b(n_6285), .c(FE_OCP_RBN6196_FE_OFN789_n_46195), .d(n_6313), .o(n_46157) );
oa22m02 g784352 ( .a(FE_OFN4788_n_46137), .b(n_6071), .c(FE_OCP_RBN6195_FE_OFN789_n_46195), .d(n_6105), .o(n_46158) );
oa22s01 g784353 ( .a(FE_OCP_RBN6196_FE_OFN789_n_46195), .b(n_6154), .c(FE_OFN4788_n_46137), .d(n_6124), .o(n_46159) );
oa22s02 g784354 ( .a(FE_OFN4788_n_46137), .b(n_6043), .c(FE_OCP_RBN6195_FE_OFN789_n_46195), .d(n_6063), .o(n_46160) );
oa22s02 g784355 ( .a(FE_OFN768_n_46137), .b(n_6175), .c(FE_OCP_RBN6196_FE_OFN789_n_46195), .d(n_46995), .o(n_46161) );
oa22s02 g784356 ( .a(FE_OFN4789_n_46137), .b(n_5567), .c(FE_OCP_RBN6195_FE_OFN789_n_46195), .d(n_5618), .o(n_46162) );
oa22s02 g784357 ( .a(FE_OCP_RBN6195_FE_OFN789_n_46195), .b(n_5840), .c(FE_OFN4788_n_46137), .d(n_5789), .o(n_46163) );
oa22s02 g784358 ( .a(FE_OFN4789_n_46137), .b(n_5795), .c(FE_OCP_RBN6195_FE_OFN789_n_46195), .d(n_5841), .o(n_46164) );
oa22f02 g784360 ( .a(FE_OFN768_n_46137), .b(n_6254), .c(FE_OCP_RBN6196_FE_OFN789_n_46195), .d(n_6297), .o(n_46166) );
oa22s02 g784361 ( .a(FE_OFN768_n_46137), .b(n_6212), .c(FE_OCP_RBN6196_FE_OFN789_n_46195), .d(n_6233), .o(n_46167) );
oa22s02 g784362 ( .a(FE_OFN4788_n_46137), .b(n_5935), .c(FE_OCP_RBN6195_FE_OFN789_n_46195), .d(n_5971), .o(n_46168) );
oa22s02 g784363 ( .a(FE_OFN771_n_46196), .b(n_5363), .c(FE_OFN4789_n_46137), .d(n_5324), .o(n_46169) );
oa22s02 g784364 ( .a(FE_OFN4789_n_46137), .b(n_5708), .c(FE_OFN771_n_46196), .d(n_5724), .o(n_46170) );
oa22s02 g784365 ( .a(FE_OFN4788_n_46137), .b(n_5937), .c(FE_OFN771_n_46196), .d(n_5972), .o(n_46171) );
oa22s02 g784366 ( .a(FE_OFN4789_n_46137), .b(n_5210), .c(FE_OFN771_n_46196), .d(n_5244), .o(n_46172) );
oa22m02 g784367 ( .a(FE_OFN4788_n_46137), .b(n_6004), .c(FE_OFN771_n_46196), .d(n_46997), .o(n_46173) );
oa22s02 g784368 ( .a(FE_OFN4789_n_46137), .b(n_5285), .c(FE_OFN771_n_46196), .d(n_5323), .o(n_46174) );
oa22s01 g784369 ( .a(FE_OFN768_n_46137), .b(n_6217), .c(FE_OFN771_n_46196), .d(n_6243), .o(n_46175) );
oa22s02 g784370 ( .a(FE_OFN4789_n_46137), .b(n_5613), .c(FE_OFN771_n_46196), .d(n_5645), .o(n_46176) );
oa22s01 g784371 ( .a(FE_OFN768_n_46137), .b(n_6392), .c(FE_OFN770_n_46196), .d(n_6419), .o(n_46177) );
oa22m02 g784372 ( .a(FE_OFN770_n_46196), .b(FE_OCP_RBN3434_n_6379), .c(FE_OFN4787_n_46137), .d(n_6379), .o(n_46178) );
oa22s01 g784373 ( .a(FE_OFN770_n_46196), .b(n_6435), .c(FE_OFN4787_n_46137), .d(n_6407), .o(n_46179) );
oa22s01 g784374 ( .a(FE_OFN768_n_46137), .b(n_6436), .c(n_6476), .d(FE_OFN770_n_46196), .o(n_46180) );
oa22f02 g784376 ( .a(n_6477), .b(FE_OFN4787_n_46137), .c(FE_OCP_RBN6248_n_6477), .d(FE_OFN770_n_46196), .o(n_46182) );
oa22s02 g784377 ( .a(n_6500), .b(FE_OFN770_n_46196), .c(n_6490), .d(FE_OFN4787_n_46137), .o(n_46183) );
oa22s02 g784378 ( .a(n_6519), .b(FE_OFN4787_n_46137), .c(n_6529), .d(FE_OFN770_n_46196), .o(n_46184) );
oa22f02 g784386 ( .a(n_6720), .b(FE_OFN770_n_46196), .c(n_44823), .d(FE_OFN4787_n_46137), .o(n_46192) );
no02f04 TIMEBOOST_cell_8652 ( .a(FE_RN_1179_0), .b(n_16466), .o(TIMEBOOST_net_2813) );
ao12s01 g784390 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_), .o(n_46200) );
in01s03 g784391 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_46197) );
oa12s01 g784392 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_), .o(n_46202) );
oa12s01 g784393 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_), .o(n_46203) );
ao12s01 g784394 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_8_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_7_), .o(n_46205) );
na02s01 g784395 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_), .o(n_46206) );
na02s01 g784396 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_5_), .o(n_46208) );
na02s01 g784397 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_1_), .o(n_46209) );
no02s01 g784398 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_22_), .o(n_46210) );
na02s01 g784399 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_21_), .o(n_46211) );
na02s01 g784400 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_13_), .o(n_46212) );
no02s01 g784401 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_), .o(n_46213) );
na02s01 g784402 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_17_), .o(n_46214) );
na02s01 g784403 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_25_), .o(n_46215) );
no02s01 g784404 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_25_), .o(n_46216) );
no02s01 g784405 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_17_), .o(n_46217) );
no02s01 g784406 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_18_), .o(n_46218) );
na02s01 g784407 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_9_), .o(n_46219) );
no02s01 g784408 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_13_), .o(n_46220) );
no02s01 g784409 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_9_), .o(n_46221) );
no02s01 g784410 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_0_), .o(n_46222) );
na02s01 g784411 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_0_), .o(n_46223) );
no02s01 g784412 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_10_), .o(n_46224) );
no02s01 g784413 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_21_), .o(n_46225) );
no02s01 g784414 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_26_), .o(n_46226) );
no02s01 g784415 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_27_), .o(n_46227) );
na02s01 g784416 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_27_), .o(n_46228) );
ao22s01 g784417 ( .a(n_36355), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46197), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_), .o(n_46229) );
oa22s01 g784418 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_7_), .c(n_36784), .d(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_46230) );
oa22s01 g784419 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_6_), .c(n_36358), .d(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_46231) );
ao22s01 g784420 ( .a(n_36762), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46204), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_), .o(n_46232) );
ao22s01 g784421 ( .a(n_36541), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46197), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_), .o(n_46233) );
oa22s01 g784422 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_8_), .c(n_36785), .d(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_46234) );
ao22s01 g784423 ( .a(n_36497), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46197), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_), .o(n_46235) );
ao22s01 g784424 ( .a(n_36354), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46204), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_), .o(n_46236) );
oa22s01 g784425 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_2_), .c(n_36353), .d(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_46237) );
ao22s01 g784426 ( .a(n_36745), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46204), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_19_), .o(n_46238) );
ao22s01 g784427 ( .a(n_36578), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46197), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_), .o(n_46239) );
oa22s01 g784428 ( .a(n_36637), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46204), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_), .o(n_46240) );
ao22s01 g784429 ( .a(n_36744), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46197), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_20_), .o(n_46241) );
ao22s01 g784430 ( .a(n_36773), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46204), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_), .o(n_46242) );
ao22s01 g784431 ( .a(n_36713), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46197), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_), .o(n_46243) );
ao12s01 g784432 ( .a(n_46218), .b(n_46204), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_18_), .o(n_46244) );
ao12s01 g784433 ( .a(n_46224), .b(n_46197), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_10_), .o(n_46245) );
oa12s01 g784434 ( .a(n_46208), .b(n_46204), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_5_), .o(n_46246) );
ao12s01 g784435 ( .a(n_46226), .b(n_46197), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_26_), .o(n_46247) );
ao12s01 g784436 ( .a(n_46210), .b(n_46204), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_22_), .o(n_46248) );
ao12s01 g784437 ( .a(n_37631), .b(n_36746), .c(n_46197), .o(n_46249) );
ao22s02 g784438 ( .a(n_36902), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_2_), .c(n_36942), .d(n_46204), .o(n_46250) );
oa12s01 g784439 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_6_), .b(n_37138), .c(n_46197), .o(n_46251) );
oa12s01 g784440 ( .a(n_46204), .b(n_37992), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_), .o(n_46252) );
ao12s01 g784441 ( .a(n_37202), .b(n_37169), .c(n_46204), .o(n_46253) );
na02s04 g784469 ( .a(n_11364), .b(n_10385), .o(n_46285) );
no02s10 g784519 ( .a(FE_OCP_RBN6137_n_11364), .b(n_10386), .o(n_46337) );
oa22s02 g784539 ( .a(n_11856), .b(FE_OCP_RBN6862_n_46285), .c(n_11805), .d(FE_OCP_RBN4448_FE_OFN760_n_46337), .o(n_46360) );
oa22f02 g784541 ( .a(n_11759), .b(FE_OCP_RBN6862_n_46285), .c(n_11669), .d(FE_OCP_RBN4447_FE_OFN760_n_46337), .o(n_46362) );
oa22m02 g784543 ( .a(n_11655), .b(FE_OCP_RBN6865_n_46285), .c(n_11527), .d(FE_OCP_RBN4448_FE_OFN760_n_46337), .o(n_46364) );
oa22f02 g784544 ( .a(n_11605), .b(FE_OCP_RBN6862_n_46285), .c(n_11495), .d(FE_OCP_RBN6167_n_46337), .o(n_46365) );
oa22s02 g784545 ( .a(n_11494), .b(FE_OCP_RBN6862_n_46285), .c(n_11463), .d(FE_OCP_RBN6167_n_46337), .o(n_46366) );
oa22m02 g784546 ( .a(n_11453), .b(FE_OCP_RBN6862_n_46285), .c(n_11422), .d(FE_OCP_RBN6167_n_46337), .o(n_46367) );
oa22f02 g784547 ( .a(FE_OCP_RBN6864_n_46285), .b(n_46986), .c(FE_OCP_RBN6168_n_46337), .d(n_11412), .o(n_46368) );
oa22s02 g784548 ( .a(n_11490), .b(FE_OCP_RBN6865_n_46285), .c(n_11409), .d(FE_OCP_RBN4448_FE_OFN760_n_46337), .o(n_46369) );
oa22m02 g784549 ( .a(FE_OCP_RBN6864_n_46285), .b(n_11212), .c(FE_OCP_RBN6168_n_46337), .d(n_11184), .o(n_46370) );
oa22m02 g784550 ( .a(FE_OCP_RBN6864_n_46285), .b(n_11307), .c(FE_OCP_RBN6168_n_46337), .d(n_11282), .o(n_46371) );
oa22m02 g784551 ( .a(FE_OCP_RBN6864_n_46285), .b(n_11252), .c(FE_OCP_RBN6168_n_46337), .d(n_11220), .o(n_46372) );
oa22s02 g784552 ( .a(FE_OCP_RBN6864_n_46285), .b(n_10885), .c(n_46337), .d(n_10799), .o(n_46373) );
oa22f02 g784553 ( .a(FE_OCP_RBN6862_n_46285), .b(n_11356), .c(FE_OCP_RBN6167_n_46337), .d(n_11334), .o(n_46374) );
oa22m02 g784554 ( .a(FE_OCP_RBN6863_n_46285), .b(n_11061), .c(n_46337), .d(n_11036), .o(n_46375) );
oa22m02 g784555 ( .a(FE_OCP_RBN6864_n_46285), .b(n_11278), .c(FE_OCP_RBN6168_n_46337), .d(n_11232), .o(n_46376) );
oa22s02 g784556 ( .a(FE_OCP_RBN6864_n_46285), .b(n_11177), .c(n_46337), .d(n_11151), .o(n_46377) );
oa22f02 g784557 ( .a(FE_OCP_RBN6862_n_46285), .b(n_11297), .c(FE_OCP_RBN6167_n_46337), .d(n_11265), .o(n_46378) );
oa22s02 g784558 ( .a(FE_OCP_RBN6864_n_46285), .b(n_10959), .c(n_46337), .d(n_10928), .o(n_46379) );
oa22s02 g784559 ( .a(FE_OCP_RBN6863_n_46285), .b(n_10680), .c(FE_OCP_RBN6166_n_46337), .d(n_10631), .o(n_46380) );
oa22s02 g784560 ( .a(FE_OCP_RBN6863_n_46285), .b(n_10705), .c(n_46337), .d(FE_OCP_RBN6194_n_10636), .o(n_46381) );
oa22s02 g784561 ( .a(FE_OCP_RBN6863_n_46285), .b(n_10848), .c(FE_OCP_RBN6166_n_46337), .d(n_10814), .o(n_46382) );
oa22s02 g784562 ( .a(FE_OCP_RBN6863_n_46285), .b(n_46988), .c(n_46337), .d(n_10980), .o(n_46383) );
oa22s02 g784563 ( .a(FE_OCP_RBN6864_n_46285), .b(n_10739), .c(n_46337), .d(n_10721), .o(n_46384) );
oa22s02 g784564 ( .a(FE_OCP_RBN6864_n_46285), .b(n_11098), .c(n_46337), .d(n_11055), .o(n_46385) );
oa22f02 g784565 ( .a(FE_OCP_RBN6862_n_46285), .b(n_11411), .c(FE_OCP_RBN6167_n_46337), .d(n_11396), .o(n_46386) );
oa22s02 g784566 ( .a(FE_OCP_RBN6863_n_46285), .b(n_10783), .c(FE_OCP_RBN6166_n_46337), .d(n_10716), .o(n_46387) );
oa22f02 g784567 ( .a(FE_OCP_RBN6862_n_46285), .b(n_11369), .c(FE_OCP_RBN6168_n_46337), .d(n_11338), .o(n_46388) );
no02s10 g784590 ( .a(n_32643), .b(FE_OCPN3542_n_32436), .o(n_46413) );
no02s01 g784591 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_23_), .o(n_46414) );
na02s01 g784592 ( .a(n_12823), .b(n_12892), .o(n_46415) );
na02s01 g784593 ( .a(n_37945), .b(FE_OCP_RBN5563_n_37551), .o(n_46416) );
na02s08 g784594 ( .a(FE_OCP_RBN5683_n_38474), .b(n_38486), .o(n_46417) );
na02m01 g784595 ( .a(n_8493), .b(n_8346), .o(n_46418) );
no02m02 g784596 ( .a(n_14190), .b(FE_OCP_RBN5947_n_14982), .o(n_46419) );
na02m04 g784597 ( .a(n_10465), .b(n_10464), .o(n_46420) );
na02s06 g784598 ( .a(n_16197), .b(FE_OCPN1733_n_14524), .o(n_46421) );
no02f08 g784599 ( .a(n_26920), .b(n_26919), .o(n_46422) );
no02s06 g784600 ( .a(n_11118), .b(FE_OFN4800_n_44498), .o(n_46423) );
no02s08 g784601 ( .a(n_11089), .b(FE_OCPN4845_FE_OFN4779_n_44490), .o(n_46424) );
no02m08 g784602 ( .a(n_11049), .b(FE_OFN756_n_44464), .o(n_44453) );
no02m08 g784603 ( .a(n_16241), .b(n_14805), .o(n_46426) );
no02f06 g784604 ( .a(n_5952), .b(n_5940), .o(n_46427) );
na02s06 g784605 ( .a(n_12406), .b(n_12686), .o(n_46933) );
na02s04 g784606 ( .a(FE_OCP_RBN6871_FE_RN_2289_0), .b(n_26620), .o(n_46934) );
ao12s01 g784607 ( .a(n_42996), .b(n_42985), .c(n_42708), .o(n_46935) );
ao12s02 g784608 ( .a(n_42950), .b(n_42928), .c(n_42673), .o(n_46936) );
ao12s01 g784609 ( .a(n_42930), .b(n_42914), .c(n_42610), .o(n_46937) );
oa12s01 g784610 ( .a(n_42904), .b(n_42881), .c(n_42760), .o(n_46938) );
ao12s01 g784611 ( .a(n_42890), .b(n_42869), .c(n_42616), .o(n_46939) );
ao12s01 g784612 ( .a(n_42874), .b(n_42848), .c(n_42612), .o(n_46940) );
ao12s01 g784613 ( .a(n_42752), .b(n_42734), .c(n_42712), .o(n_46941) );
ao12s01 g784614 ( .a(n_42704), .b(n_42687), .c(n_42681), .o(n_46942) );
ao12s01 g784615 ( .a(n_42634), .b(n_42379), .c(n_42587), .o(n_46943) );
oa12s01 g784616 ( .a(n_42567), .b(n_42552), .c(n_42314), .o(n_46944) );
na02f02 TIMEBOOST_cell_3102 ( .a(FE_RN_90_0), .b(n_24503), .o(TIMEBOOST_net_842) );
ao12s01 g784619 ( .a(n_39533), .b(n_39532), .c(n_39072), .o(n_46948) );
ao12s02 g784620 ( .a(n_39494), .b(n_39408), .c(n_39455), .o(n_46949) );
oa12s02 g784621 ( .a(n_39472), .b(n_39431), .c(n_39391), .o(n_46950) );
oa12s01 g784622 ( .a(n_38479), .b(n_38478), .c(n_38085), .o(n_46951) );
oa12f04 g784623 ( .a(n_37232), .b(n_37377), .c(n_37019), .o(n_46952) );
oa12f02 g784636 ( .a(n_22536), .b(n_22482), .c(n_22347), .o(n_46965) );
oa12f04 g784640 ( .a(n_20854), .b(n_20823), .c(n_20732), .o(n_46969) );
oa12f02 g784643 ( .a(n_16999), .b(n_16753), .c(n_16938), .o(n_46973) );
oa12f02 g784644 ( .a(n_16840), .b(n_16811), .c(n_16785), .o(n_46974) );
oa12f02 g784645 ( .a(n_16787), .b(n_16755), .c(n_16728), .o(n_46975) );
oa12f02 g784646 ( .a(n_16703), .b(n_16640), .c(n_16656), .o(n_46976) );
oa12f02 g784647 ( .a(n_16628), .b(n_16607), .c(n_16585), .o(n_46977) );
oa12s02 g784649 ( .a(n_16559), .b(n_16527), .c(n_16486), .o(n_46979) );
ao12m04 g784650 ( .a(n_15738), .b(n_15696), .c(n_15649), .o(n_46980) );
ao12f04 g784651 ( .a(n_15728), .b(n_15688), .c(n_15727), .o(n_46981) );
no02s06 TIMEBOOST_cell_3159 ( .a(n_30530), .b(TIMEBOOST_net_870), .o(n_30599) );
oa12f04 g784656 ( .a(n_11361), .b(n_11316), .c(n_11187), .o(n_46986) );
ao12m04 g784657 ( .a(n_11080), .b(n_11045), .c(n_10989), .o(n_46987) );
oa12s02 g784658 ( .a(n_10900), .b(n_10813), .c(n_10684), .o(n_46988) );
oa12s02 g784660 ( .a(n_8520), .b(n_8421), .c(n_8466), .o(n_46990) );
ao12s01 g784662 ( .a(n_7490), .b(n_7462), .c(n_7292), .o(n_46992) );
oa12m02 g784664 ( .a(n_6224), .b(n_6178), .c(n_6119), .o(n_46994) );
oa12s02 g784665 ( .a(n_6121), .b(n_6036), .c(n_5889), .o(n_46995) );
oa12m02 g784667 ( .a(n_5928), .b(n_5902), .c(n_5761), .o(n_46997) );
ao12f02 g784668 ( .a(n_5838), .b(n_5793), .c(n_5587), .o(n_46998) );
oa12f02 g784669 ( .a(n_5592), .b(n_5506), .c(n_5559), .o(n_46999) );
ao12m02 g784673 ( .a(n_5161), .b(n_5123), .c(n_4723), .o(n_47003) );
ao12s02 g784674 ( .a(n_5012), .b(n_4933), .c(n_4348), .o(n_47004) );
oa12s02 g784676 ( .a(n_4664), .b(n_4661), .c(n_4267), .o(n_47006) );
oa12m02 g784680 ( .a(n_3949), .b(n_3948), .c(n_3920), .o(n_47010) );
ao12m02 g784682 ( .a(n_3942), .b(n_3894), .c(n_3792), .o(n_47012) );
oa12s02 g784683 ( .a(n_3775), .b(n_3744), .c(n_3613), .o(n_47013) );
oa12s02 g784684 ( .a(n_3683), .b(n_3575), .c(n_3460), .o(n_47014) );
oa12m01 g784685 ( .a(n_3569), .b(n_3557), .c(n_3444), .o(n_47015) );
ao12s02 g784686 ( .a(n_3496), .b(n_3475), .c(n_3248), .o(n_47016) );
oa12s02 g784687 ( .a(n_3493), .b(n_3492), .c(n_2764), .o(n_47017) );
ao12s02 g784688 ( .a(n_3412), .b(FE_OCP_RBN4213_n_3386), .c(n_2695), .o(n_47018) );
ao12s02 g784689 ( .a(n_3360), .b(n_3340), .c(n_3152), .o(n_47019) );
ao12s02 g784690 ( .a(n_3093), .b(n_3092), .c(n_2286), .o(n_47020) );
oa12m02 g784691 ( .a(n_3100), .b(n_2940), .c(n_3049), .o(n_47021) );
oa12m02 g784693 ( .a(n_2915), .b(n_2914), .c(n_2280), .o(n_47023) );
ao12s01 g784694 ( .a(n_2786), .b(n_2722), .c(n_2137), .o(n_47024) );
no02s02 TIMEBOOST_cell_8522 ( .a(n_672), .b(n_666), .o(TIMEBOOST_net_2748) );
oa12f02 g784698 ( .a(FE_OCPN869_n_45003), .b(n_20250), .c(n_20229), .o(n_47174) );
no02f02 g784699 ( .a(n_20229), .b(n_20250), .o(n_47175) );
no02s01 g784702 ( .a(n_7332), .b(n_47179), .o(n_47180) );
na02s01 g784703 ( .a(n_47177), .b(FE_RN_816_0), .o(n_47179) );
in01s01 g784704 ( .a(n_6749), .o(n_47177) );
no02s04 g784706 ( .a(n_11308), .b(FE_OCP_RBN3094_n_10023), .o(n_47182) );
na02s04 g784707 ( .a(n_47183), .b(n_47184), .o(n_47185) );
in01s02 g784708 ( .a(n_11308), .o(n_47183) );
in01s01 g784709 ( .a(FE_OCP_RBN3095_n_10023), .o(n_47184) );
in01s06 g784728 ( .a(n_47212), .o(n_47213) );
no02m10 g784729 ( .a(n_11962), .b(n_11643), .o(n_47212) );
ao22s02 g784753 ( .a(n_7687), .b(n_7310), .c(n_7686), .d(n_7309), .o(n_47235) );
no02s02 g784754 ( .a(n_47235), .b(FE_OCP_RBN6597_n_7708), .o(n_47240) );
no02s02 g784755 ( .a(n_47235), .b(n_7730), .o(n_47241) );
na02s02 g784756 ( .a(n_47235), .b(n_8073), .o(n_47242) );
na02s02 g784757 ( .a(n_8889), .b(FE_OCPN4851_n_47235), .o(n_47243) );
no02m04 g784758 ( .a(n_8889), .b(FE_OCPN4851_n_47235), .o(n_47244) );
na02s06 g784760 ( .a(FE_OFN777_n_18268), .b(n_18368), .o(n_47246) );
na02m03 g784761 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_), .o(n_47247) );
no02s03 g784762 ( .a(FE_OCP_RBN2495_n_18242), .b(delay_add_ln22_unr11_stage5_stallmux_q_21_), .o(n_47248) );
no02m08 g784763 ( .a(n_33594), .b(n_34037), .o(n_47249) );
na02s02 g784764 ( .a(n_12823), .b(n_12834), .o(n_47250) );
no02m06 g784765 ( .a(n_29231), .b(FE_OFN773_n_25834), .o(n_47251) );
na02s02 g784766 ( .a(FE_OCP_RBN5600_n_44875), .b(n_37623), .o(n_47252) );
no02s03 g784768 ( .a(n_44102), .b(FE_OCP_RBN4912_n_33803), .o(n_47254) );
na02s01 g784769 ( .a(FE_OCP_RBN6671_n_34297), .b(n_33584), .o(n_47255) );
no02m06 g784770 ( .a(n_14547), .b(FE_OCP_RBN4200_n_13796), .o(n_47256) );
no02s02 g784771 ( .a(n_20249), .b(FE_OCP_RBN7033_n_18981), .o(n_47257) );
na02s06 g784772 ( .a(FE_OCP_RBN6790_n_20242), .b(FE_OCP_RBN5669_n_19101), .o(n_47258) );
na02f02 g784773 ( .a(n_9410), .b(FE_OCPN1061_n_44460), .o(n_47259) );
no02s04 g784774 ( .a(n_8750), .b(n_9724), .o(n_47260) );
no02s02 g784775 ( .a(n_15103), .b(FE_OCP_RBN2079_n_14149), .o(n_47261) );
no02f04 g784776 ( .a(n_14935), .b(FE_OCP_RBN2834_n_13962), .o(n_47262) );
no02s08 g784778 ( .a(FE_OCP_RBN6075_n_44256), .b(n_35861), .o(n_47264) );
no02s02 g784779 ( .a(FE_OCP_RBN3171_n_44211), .b(n_34946), .o(n_47265) );
no02s06 g784780 ( .a(FE_OCP_RBN4910_n_44222), .b(n_35906), .o(n_47266) );
no02m01 g784781 ( .a(n_35977), .b(FE_OCP_RBN4910_n_44222), .o(n_47267) );
na02m08 g784782 ( .a(n_16241), .b(n_14805), .o(n_47268) );
na02m06 g784783 ( .a(n_11089), .b(n_44511), .o(n_47269) );
na02s02 g784784 ( .a(n_5746), .b(FE_OCP_RBN3066_n_4294), .o(n_47270) );
no02s02 g784785 ( .a(FE_OCP_RBN3391_n_31819), .b(FE_OCP_RBN6038_n_30733), .o(n_47271) );
no02s02 g784786 ( .a(FE_OCP_RBN4472_n_31819), .b(n_30733), .o(n_47272) );
na02s02 g784788 ( .a(FE_OCP_RBN4472_n_31819), .b(FE_OCP_RBN6063_n_30908), .o(n_47274) );
no02s01 g784790 ( .a(FE_OCP_RBN4468_n_44267), .b(FE_OCPN6931_n_22156), .o(n_47278) );
no02s06 g784791 ( .a(FE_OCP_RBN6883_n_11486), .b(FE_OCP_RBN3289_n_10915), .o(n_47279) );
in01f04 g784792 ( .a(n_47332), .o(n_47333) );
no02f04 g784793 ( .a(n_15543), .b(n_15586), .o(n_47332) );
in01f02 g784794 ( .a(n_47334), .o(n_47335) );
no02f02 g784795 ( .a(n_6565), .b(n_6415), .o(n_47334) );
oa12m02 g784796 ( .a(n_44875), .b(n_38269), .c(n_37935), .o(n_47336) );
ao12m04 g784797 ( .a(n_23194), .b(n_23138), .c(n_23047), .o(n_47337) );
oa12f02 g784799 ( .a(n_16372), .b(n_16322), .c(n_16274), .o(n_47340) );
ao12s01 g784800 ( .a(n_3150), .b(n_3149), .c(n_2983), .o(n_47341) );
ms00f80 mux_while_ln12_psv_q_reg_1_ ( .ck(ispd_clk), .d(n_98), .o(mux_while_ln12_psv_q_1_) );
ms00f80 mux_while_ln12_psv_q_reg_2_ ( .ck(ispd_clk), .d(n_173), .o(mux_while_ln12_psv_q_2_) );
ms00f80 mux_while_ln12_psv_q_reg_3_ ( .ck(ispd_clk), .d(n_181), .o(mux_while_ln12_psv_q_3_) );
ms00f80 mux_while_ln12_psv_q_reg_4_ ( .ck(ispd_clk), .d(n_204), .o(mux_while_ln12_psv_q_4_) );
ms00f80 mux_while_ln12_psv_q_reg_5_ ( .ck(ispd_clk), .d(n_213), .o(mux_while_ln12_psv_q_5_) );
ms00f80 mux_while_ln12_psv_q_reg_6_ ( .ck(ispd_clk), .d(n_227), .o(mux_while_ln12_psv_q_6_) );
ms00f80 mux_while_ln12_psv_q_reg_7_ ( .ck(ispd_clk), .d(n_243), .o(mux_while_ln12_psv_q_7_) );
ms00f80 mux_while_ln12_psv_q_reg_8_ ( .ck(ispd_clk), .d(n_265), .o(TIMEBOOST_net_2186) );
ms00f80 sin_out_reg_0_ ( .ck(ispd_clk), .d(n_43155), .o(sin_out_0) );
ms00f80 sin_out_reg_10_ ( .ck(ispd_clk), .d(n_43803), .o(sin_out_10) );
ms00f80 sin_out_reg_11_ ( .ck(ispd_clk), .d(n_43805), .o(sin_out_11) );
ms00f80 sin_out_reg_12_ ( .ck(ispd_clk), .d(n_43802), .o(sin_out_12) );
ms00f80 sin_out_reg_13_ ( .ck(ispd_clk), .d(n_43804), .o(sin_out_13) );
ms00f80 sin_out_reg_14_ ( .ck(ispd_clk), .d(n_43824), .o(sin_out_14) );
ms00f80 sin_out_reg_15_ ( .ck(ispd_clk), .d(n_43813), .o(sin_out_15) );
ms00f80 sin_out_reg_16_ ( .ck(ispd_clk), .d(n_43873), .o(sin_out_16) );
ms00f80 sin_out_reg_17_ ( .ck(ispd_clk), .d(n_43890), .o(sin_out_17) );
ms00f80 sin_out_reg_18_ ( .ck(ispd_clk), .d(n_43889), .o(sin_out_18) );
ms00f80 sin_out_reg_19_ ( .ck(ispd_clk), .d(n_43896), .o(sin_out_19) );
ms00f80 sin_out_reg_1_ ( .ck(ispd_clk), .d(n_43237), .o(sin_out_1) );
ms00f80 sin_out_reg_20_ ( .ck(ispd_clk), .d(n_43888), .o(sin_out_20) );
ms00f80 sin_out_reg_21_ ( .ck(ispd_clk), .d(n_43899), .o(sin_out_21) );
ms00f80 sin_out_reg_22_ ( .ck(ispd_clk), .d(n_43898), .o(sin_out_22) );
ms00f80 sin_out_reg_23_ ( .ck(ispd_clk), .d(n_43903), .o(sin_out_23) );
ms00f80 sin_out_reg_24_ ( .ck(ispd_clk), .d(n_43910), .o(sin_out_24) );
ms00f80 sin_out_reg_25_ ( .ck(ispd_clk), .d(n_43913), .o(sin_out_25) );
ms00f80 sin_out_reg_26_ ( .ck(ispd_clk), .d(n_43915), .o(sin_out_26) );
ms00f80 sin_out_reg_27_ ( .ck(ispd_clk), .d(n_43917), .o(sin_out_27) );
ms00f80 sin_out_reg_28_ ( .ck(ispd_clk), .d(n_43914), .o(sin_out_28) );
ms00f80 sin_out_reg_29_ ( .ck(ispd_clk), .d(n_43920), .o(sin_out_29) );
ms00f80 sin_out_reg_2_ ( .ck(ispd_clk), .d(n_43337), .o(sin_out_2) );
ms00f80 sin_out_reg_30_ ( .ck(ispd_clk), .d(n_43919), .o(sin_out_30) );
ms00f80 sin_out_reg_31_ ( .ck(ispd_clk), .d(n_43916), .o(sin_out_31) );
ms00f80 sin_out_reg_3_ ( .ck(ispd_clk), .d(n_43680), .o(sin_out_3) );
ms00f80 sin_out_reg_4_ ( .ck(ispd_clk), .d(n_43685), .o(sin_out_4) );
ms00f80 sin_out_reg_5_ ( .ck(ispd_clk), .d(n_43703), .o(sin_out_5) );
ms00f80 sin_out_reg_6_ ( .ck(ispd_clk), .d(n_43677), .o(sin_out_6) );
ms00f80 sin_out_reg_7_ ( .ck(ispd_clk), .d(n_43707), .o(sin_out_7) );
ms00f80 sin_out_reg_8_ ( .ck(ispd_clk), .d(n_43746), .o(sin_out_8) );
ms00f80 sin_out_reg_9_ ( .ck(ispd_clk), .d(n_43773), .o(sin_out_9) );
ms00f80 state_cordic_reg_1_ ( .ck(ispd_clk), .d(rst), .o(TIMEBOOST_net_1375) );
no02s02 TIMEBOOST_cell_1564 ( .a(TIMEBOOST_net_396), .b(n_4131), .o(n_4184) );

endmodule
